module aes_cipher_top (clk,
    done,
    ld,
    rst,
    key,
    text_in,
    text_out);
 input clk;
 output done;
 input ld;
 input rst;
 input [127:0] key;
 input [127:0] text_in;
 output [127:0] text_out;

 INV_X1 _17732_ (.A(_01330_),
    .ZN(_03727_));
 BUF_X4 _17733_ (.A(_03727_),
    .Z(_03738_));
 BUF_X4 _17734_ (.A(_03738_),
    .Z(_03749_));
 AND2_X1 _17735_ (.A1(_17140_),
    .A2(_17141_),
    .ZN(_03760_));
 INV_X1 _17736_ (.A(_03760_),
    .ZN(_03771_));
 INV_X1 _17737_ (.A(_17142_),
    .ZN(_03782_));
 OAI21_X1 _17738_ (.A(_03749_),
    .B1(_03771_),
    .B2(_03782_),
    .ZN(_01186_));
 AND2_X1 _17739_ (.A1(_03760_),
    .A2(_17142_),
    .ZN(_03803_));
 INV_X1 _17740_ (.A(_17143_),
    .ZN(_03814_));
 NAND2_X1 _17741_ (.A1(_03803_),
    .A2(_03814_),
    .ZN(_03825_));
 BUF_X4 _17742_ (.A(_01330_),
    .Z(_03836_));
 BUF_X4 _17743_ (.A(_03836_),
    .Z(_03847_));
 NOR2_X1 _17744_ (.A1(_01330_),
    .A2(_17140_),
    .ZN(_01194_));
 INV_X1 _17745_ (.A(_17141_),
    .ZN(_03868_));
 AND2_X1 _17746_ (.A1(_01194_),
    .A2(_03868_),
    .ZN(_03879_));
 INV_X1 _17747_ (.A(_03879_),
    .ZN(_03890_));
 OAI22_X1 _17748_ (.A1(_03825_),
    .A2(_03847_),
    .B1(_03890_),
    .B2(_17142_),
    .ZN(_01187_));
 XNOR2_X1 _17749_ (.A(_03803_),
    .B(_03814_),
    .ZN(_03911_));
 XNOR2_X1 _17750_ (.A(_03760_),
    .B(_03782_),
    .ZN(_03922_));
 BUF_X4 _17751_ (.A(_03727_),
    .Z(_03933_));
 NAND3_X1 _17752_ (.A1(_03933_),
    .A2(_03868_),
    .A3(_17140_),
    .ZN(_03944_));
 OR3_X1 _17753_ (.A1(_03911_),
    .A2(_03922_),
    .A3(_03944_),
    .ZN(_03955_));
 INV_X1 _17754_ (.A(_03922_),
    .ZN(_03966_));
 NAND3_X1 _17755_ (.A1(_03911_),
    .A2(_03966_),
    .A3(_03879_),
    .ZN(_03977_));
 NAND2_X1 _17756_ (.A1(_03955_),
    .A2(_03977_),
    .ZN(_01188_));
 OR4_X1 _17757_ (.A1(_17140_),
    .A2(_03868_),
    .A3(_17142_),
    .A4(_17143_),
    .ZN(_03998_));
 AOI21_X1 _17758_ (.A(_03847_),
    .B1(_03825_),
    .B2(_03998_),
    .ZN(_01189_));
 NAND4_X1 _17759_ (.A1(_03749_),
    .A2(_03814_),
    .A3(_17140_),
    .A4(_17141_),
    .ZN(_04019_));
 NAND2_X1 _17760_ (.A1(_03977_),
    .A2(_04019_),
    .ZN(_01190_));
 NAND2_X1 _17761_ (.A1(_03922_),
    .A2(_03814_),
    .ZN(_04040_));
 OAI21_X1 _17762_ (.A(_03977_),
    .B1(_03890_),
    .B2(_04040_),
    .ZN(_01191_));
 NOR2_X1 _17763_ (.A1(_04040_),
    .A2(_03944_),
    .ZN(_01192_));
 AND4_X1 _17764_ (.A1(_17141_),
    .A2(_03922_),
    .A3(_03814_),
    .A4(_01194_),
    .ZN(_01193_));
 NOR2_X1 _17765_ (.A1(_17140_),
    .A2(_17141_),
    .ZN(_04080_));
 NOR3_X1 _17766_ (.A1(_03760_),
    .A2(_04080_),
    .A3(_03847_),
    .ZN(_01195_));
 AOI21_X1 _17767_ (.A(_01186_),
    .B1(_03782_),
    .B2(_03771_),
    .ZN(_01196_));
 AND2_X1 _17768_ (.A1(_03911_),
    .A2(_03749_),
    .ZN(_01197_));
 BUF_X4 _17769_ (.A(_17144_),
    .Z(_04121_));
 BUF_X4 _17770_ (.A(_04121_),
    .Z(_04132_));
 XOR2_X1 _17771_ (.A(_04132_),
    .B(_17012_),
    .Z(_04143_));
 INV_X32 _17772_ (.A(_16833_),
    .ZN(_04154_));
 AND2_X4 _17773_ (.A1(_04154_),
    .A2(_16832_),
    .ZN(_04165_));
 NOR2_X4 _17774_ (.A1(_16835_),
    .A2(_16834_),
    .ZN(_04176_));
 BUF_X4 _17775_ (.A(_04176_),
    .Z(_04187_));
 AND2_X2 _17776_ (.A1(_04165_),
    .A2(_04187_),
    .ZN(_04198_));
 BUF_X4 _17777_ (.A(_04198_),
    .Z(_04209_));
 INV_X32 _17778_ (.A(_16831_),
    .ZN(_04220_));
 NOR2_X4 _17779_ (.A1(_04220_),
    .A2(_16830_),
    .ZN(_04231_));
 NOR2_X4 _17780_ (.A1(_16829_),
    .A2(_16828_),
    .ZN(_04242_));
 AND2_X2 _17781_ (.A1(_04231_),
    .A2(_04242_),
    .ZN(_04253_));
 NAND2_X1 _17782_ (.A1(_04209_),
    .A2(_04253_),
    .ZN(_04264_));
 BUF_X32 _17783_ (.A(_16829_),
    .Z(_04275_));
 AND2_X4 _17784_ (.A1(_04275_),
    .A2(_16828_),
    .ZN(_04286_));
 AND2_X4 _17785_ (.A1(_04231_),
    .A2(_04286_),
    .ZN(_04297_));
 NAND3_X1 _17786_ (.A1(_04297_),
    .A2(_04187_),
    .A3(_04165_),
    .ZN(_04308_));
 AND2_X1 _17787_ (.A1(_04264_),
    .A2(_04308_),
    .ZN(_04319_));
 NOR2_X4 _17788_ (.A1(_16833_),
    .A2(_16832_),
    .ZN(_04329_));
 AND2_X4 _17789_ (.A1(_04187_),
    .A2(_04329_),
    .ZN(_04340_));
 INV_X32 _17790_ (.A(_16830_),
    .ZN(_04351_));
 NOR2_X4 _17791_ (.A1(_04351_),
    .A2(_16831_),
    .ZN(_04362_));
 INV_X32 _17792_ (.A(_16828_),
    .ZN(_04373_));
 NOR2_X4 _17793_ (.A1(_04373_),
    .A2(_16829_),
    .ZN(_04384_));
 BUF_X8 _17794_ (.A(_04384_),
    .Z(_04395_));
 AND3_X1 _17795_ (.A1(_04340_),
    .A2(_04362_),
    .A3(_04395_),
    .ZN(_04406_));
 AND2_X2 _17796_ (.A1(_04362_),
    .A2(_04275_),
    .ZN(_04417_));
 BUF_X4 _17797_ (.A(_04340_),
    .Z(_04428_));
 AND2_X1 _17798_ (.A1(_04417_),
    .A2(_04428_),
    .ZN(_04439_));
 NOR2_X4 _17799_ (.A1(_16830_),
    .A2(_16831_),
    .ZN(_04450_));
 AND2_X1 _17800_ (.A1(_04450_),
    .A2(_04275_),
    .ZN(_04461_));
 AOI211_X2 _17801_ (.A(_04406_),
    .B(_04439_),
    .C1(_04461_),
    .C2(_04428_),
    .ZN(_04472_));
 BUF_X2 _17802_ (.A(_04209_),
    .Z(_04483_));
 BUF_X8 _17803_ (.A(_04286_),
    .Z(_04494_));
 INV_X4 _17804_ (.A(_04494_),
    .ZN(_04505_));
 AND2_X1 _17805_ (.A1(_04505_),
    .A2(_04362_),
    .ZN(_04516_));
 INV_X1 _17806_ (.A(_04242_),
    .ZN(_04527_));
 AND2_X2 _17807_ (.A1(_04516_),
    .A2(_04527_),
    .ZN(_04538_));
 BUF_X2 _17808_ (.A(_04461_),
    .Z(_04549_));
 OAI21_X1 _17809_ (.A(_04483_),
    .B1(_04538_),
    .B2(_04549_),
    .ZN(_04560_));
 INV_X32 _17810_ (.A(_16829_),
    .ZN(_04571_));
 NOR2_X4 _17811_ (.A1(_04571_),
    .A2(_16828_),
    .ZN(_04581_));
 BUF_X8 _17812_ (.A(_04231_),
    .Z(_04592_));
 AND3_X1 _17813_ (.A1(_04428_),
    .A2(_04581_),
    .A3(_04592_),
    .ZN(_04603_));
 INV_X1 _17814_ (.A(_04603_),
    .ZN(_04614_));
 AND2_X4 _17815_ (.A1(_16830_),
    .A2(_16831_),
    .ZN(_04625_));
 INV_X1 _17816_ (.A(_04625_),
    .ZN(_04636_));
 BUF_X8 _17817_ (.A(_04242_),
    .Z(_04647_));
 NOR2_X2 _17818_ (.A1(_04636_),
    .A2(_04647_),
    .ZN(_04658_));
 BUF_X8 _17819_ (.A(_04505_),
    .Z(_04669_));
 NAND3_X1 _17820_ (.A1(_04658_),
    .A2(_04669_),
    .A3(_04428_),
    .ZN(_04680_));
 NAND2_X1 _17821_ (.A1(_04297_),
    .A2(_04428_),
    .ZN(_04691_));
 NAND3_X1 _17822_ (.A1(_04428_),
    .A2(_04395_),
    .A3(_04592_),
    .ZN(_04702_));
 AND4_X1 _17823_ (.A1(_04614_),
    .A2(_04680_),
    .A3(_04691_),
    .A4(_04702_),
    .ZN(_04713_));
 AND4_X1 _17824_ (.A1(_04319_),
    .A2(_04472_),
    .A3(_04560_),
    .A4(_04713_),
    .ZN(_04724_));
 NOR2_X4 _17825_ (.A1(_04154_),
    .A2(_16832_),
    .ZN(_04735_));
 AND2_X1 _17826_ (.A1(_04735_),
    .A2(_04187_),
    .ZN(_04746_));
 BUF_X4 _17827_ (.A(_04746_),
    .Z(_04757_));
 BUF_X4 _17828_ (.A(_04757_),
    .Z(_04768_));
 BUF_X4 _17829_ (.A(_04450_),
    .Z(_04779_));
 INV_X1 _17830_ (.A(_04779_),
    .ZN(_04790_));
 NOR2_X1 _17831_ (.A1(_04790_),
    .A2(_04494_),
    .ZN(_04801_));
 AND2_X1 _17832_ (.A1(_04768_),
    .A2(_04801_),
    .ZN(_04812_));
 AOI21_X1 _17833_ (.A(_04812_),
    .B1(_04538_),
    .B2(_04768_),
    .ZN(_04823_));
 BUF_X8 _17834_ (.A(_04625_),
    .Z(_04833_));
 AND2_X4 _17835_ (.A1(_04833_),
    .A2(_04647_),
    .ZN(_04844_));
 BUF_X8 _17836_ (.A(_04844_),
    .Z(_04855_));
 AND2_X1 _17837_ (.A1(_04757_),
    .A2(_04855_),
    .ZN(_04866_));
 INV_X1 _17838_ (.A(_04866_),
    .ZN(_04877_));
 AND2_X2 _17839_ (.A1(_04527_),
    .A2(_04592_),
    .ZN(_04888_));
 NAND2_X1 _17840_ (.A1(_04888_),
    .A2(_04768_),
    .ZN(_04899_));
 AND2_X4 _17841_ (.A1(_04625_),
    .A2(_04275_),
    .ZN(_04910_));
 BUF_X2 _17842_ (.A(_04910_),
    .Z(_04921_));
 BUF_X2 _17843_ (.A(_04735_),
    .Z(_04932_));
 NAND3_X1 _17844_ (.A1(_04921_),
    .A2(_04187_),
    .A3(_04932_),
    .ZN(_04943_));
 AND3_X1 _17845_ (.A1(_04877_),
    .A2(_04899_),
    .A3(_04943_),
    .ZN(_04954_));
 AND2_X4 _17846_ (.A1(_04494_),
    .A2(_04833_),
    .ZN(_04965_));
 BUF_X8 _17847_ (.A(_04965_),
    .Z(_04976_));
 AND2_X4 _17848_ (.A1(_16833_),
    .A2(_16832_),
    .ZN(_04987_));
 AND2_X4 _17849_ (.A1(_04987_),
    .A2(_04176_),
    .ZN(_04998_));
 BUF_X8 _17850_ (.A(_04998_),
    .Z(_05009_));
 NAND2_X1 _17851_ (.A1(_04976_),
    .A2(_05009_),
    .ZN(_05018_));
 NAND2_X1 _17852_ (.A1(_04527_),
    .A2(_04779_),
    .ZN(_05028_));
 INV_X1 _17853_ (.A(_05028_),
    .ZN(_05037_));
 AND2_X1 _17854_ (.A1(_04362_),
    .A2(_04581_),
    .ZN(_05047_));
 BUF_X2 _17855_ (.A(_05047_),
    .Z(_05056_));
 OAI21_X1 _17856_ (.A(_05009_),
    .B1(_05037_),
    .B2(_05056_),
    .ZN(_05066_));
 NAND2_X1 _17857_ (.A1(_04253_),
    .A2(_05009_),
    .ZN(_05075_));
 AND2_X2 _17858_ (.A1(_04625_),
    .A2(_04571_),
    .ZN(_05085_));
 NAND2_X1 _17859_ (.A1(_04998_),
    .A2(_05085_),
    .ZN(_05095_));
 AND4_X1 _17860_ (.A1(_05018_),
    .A2(_05066_),
    .A3(_05075_),
    .A4(_05095_),
    .ZN(_05105_));
 AND4_X2 _17861_ (.A1(_04724_),
    .A2(_04823_),
    .A3(_04954_),
    .A4(_05105_),
    .ZN(_05114_));
 INV_X32 _17862_ (.A(_16835_),
    .ZN(_05124_));
 AND2_X4 _17863_ (.A1(_05124_),
    .A2(_16834_),
    .ZN(_05133_));
 AND2_X2 _17864_ (.A1(_05133_),
    .A2(_04735_),
    .ZN(_05143_));
 AND2_X4 _17865_ (.A1(_04581_),
    .A2(_04833_),
    .ZN(_05152_));
 AND2_X2 _17866_ (.A1(_05143_),
    .A2(_05152_),
    .ZN(_05161_));
 AND2_X4 _17867_ (.A1(_04362_),
    .A2(_04571_),
    .ZN(_05170_));
 BUF_X4 _17868_ (.A(_05170_),
    .Z(_05180_));
 NAND2_X4 _17869_ (.A1(_05143_),
    .A2(_05180_),
    .ZN(_05184_));
 AND2_X4 _17870_ (.A1(_04362_),
    .A2(_04286_),
    .ZN(_05188_));
 NAND2_X1 _17871_ (.A1(_05143_),
    .A2(_05188_),
    .ZN(_05190_));
 INV_X1 _17872_ (.A(_05143_),
    .ZN(_05192_));
 INV_X1 _17873_ (.A(_05047_),
    .ZN(_05194_));
 OAI211_X2 _17874_ (.A(_05184_),
    .B(_05190_),
    .C1(_05192_),
    .C2(_05194_),
    .ZN(_05196_));
 BUF_X4 _17875_ (.A(_16828_),
    .Z(_05198_));
 AND2_X4 _17876_ (.A1(_04779_),
    .A2(_05198_),
    .ZN(_05200_));
 BUF_X2 _17877_ (.A(_05133_),
    .Z(_05202_));
 AND3_X1 _17878_ (.A1(_05200_),
    .A2(_05202_),
    .A3(_04932_),
    .ZN(_05204_));
 NAND4_X1 _17879_ (.A1(_05202_),
    .A2(_04592_),
    .A3(_04932_),
    .A4(_04494_),
    .ZN(_05206_));
 NAND2_X2 _17880_ (.A1(_04231_),
    .A2(_04571_),
    .ZN(_05214_));
 OAI21_X1 _17881_ (.A(_05206_),
    .B1(_05192_),
    .B2(_05214_),
    .ZN(_05225_));
 OR4_X2 _17882_ (.A1(_05161_),
    .A2(_05196_),
    .A3(_05204_),
    .A4(_05225_),
    .ZN(_05236_));
 AND2_X2 _17883_ (.A1(_05133_),
    .A2(_04329_),
    .ZN(_05247_));
 OAI21_X1 _17884_ (.A(_05247_),
    .B1(_05152_),
    .B2(_05085_),
    .ZN(_05258_));
 BUF_X4 _17885_ (.A(_04592_),
    .Z(_05269_));
 NAND4_X1 _17886_ (.A1(_05202_),
    .A2(_05269_),
    .A3(_05198_),
    .A4(_04329_),
    .ZN(_05280_));
 AND2_X1 _17887_ (.A1(_05258_),
    .A2(_05280_),
    .ZN(_05291_));
 AND2_X1 _17888_ (.A1(_04450_),
    .A2(_04571_),
    .ZN(_05302_));
 BUF_X2 _17889_ (.A(_05302_),
    .Z(_05313_));
 NAND3_X1 _17890_ (.A1(_05313_),
    .A2(_04329_),
    .A3(_05202_),
    .ZN(_05324_));
 AND2_X2 _17891_ (.A1(_04362_),
    .A2(_04242_),
    .ZN(_05335_));
 INV_X1 _17892_ (.A(_05335_),
    .ZN(_05346_));
 BUF_X4 _17893_ (.A(_05247_),
    .Z(_05357_));
 INV_X1 _17894_ (.A(_05357_),
    .ZN(_05368_));
 OAI211_X2 _17895_ (.A(_05291_),
    .B(_05324_),
    .C1(_05346_),
    .C2(_05368_),
    .ZN(_05379_));
 AND2_X4 _17896_ (.A1(_05133_),
    .A2(_04987_),
    .ZN(_05390_));
 BUF_X4 _17897_ (.A(_04362_),
    .Z(_05401_));
 AND2_X2 _17898_ (.A1(_05401_),
    .A2(_05198_),
    .ZN(_05412_));
 AND2_X1 _17899_ (.A1(_05390_),
    .A2(_05412_),
    .ZN(_05423_));
 INV_X1 _17900_ (.A(_05423_),
    .ZN(_05434_));
 NAND3_X1 _17901_ (.A1(_05390_),
    .A2(_04669_),
    .A3(_04658_),
    .ZN(_05445_));
 BUF_X4 _17902_ (.A(_04297_),
    .Z(_05456_));
 BUF_X2 _17903_ (.A(_04987_),
    .Z(_05467_));
 NAND3_X1 _17904_ (.A1(_05456_),
    .A2(_05202_),
    .A3(_05467_),
    .ZN(_05478_));
 BUF_X4 _17905_ (.A(_05390_),
    .Z(_05489_));
 BUF_X4 _17906_ (.A(_04779_),
    .Z(_05500_));
 BUF_X4 _17907_ (.A(_04571_),
    .Z(_05511_));
 BUF_X4 _17908_ (.A(_05198_),
    .Z(_05522_));
 OAI211_X2 _17909_ (.A(_05489_),
    .B(_05500_),
    .C1(_05511_),
    .C2(_05522_),
    .ZN(_05533_));
 NAND4_X1 _17910_ (.A1(_05434_),
    .A2(_05445_),
    .A3(_05478_),
    .A4(_05533_),
    .ZN(_05544_));
 AND2_X2 _17911_ (.A1(_05133_),
    .A2(_04165_),
    .ZN(_05555_));
 AND2_X4 _17912_ (.A1(_04494_),
    .A2(_04779_),
    .ZN(_05566_));
 AND2_X1 _17913_ (.A1(_05555_),
    .A2(_05566_),
    .ZN(_05577_));
 INV_X1 _17914_ (.A(_05577_),
    .ZN(_05588_));
 BUF_X2 _17915_ (.A(_05555_),
    .Z(_05599_));
 NAND2_X1 _17916_ (.A1(_05599_),
    .A2(_04417_),
    .ZN(_05610_));
 AND2_X1 _17917_ (.A1(_04592_),
    .A2(_05198_),
    .ZN(_05621_));
 OAI21_X2 _17918_ (.A(_05599_),
    .B1(_05621_),
    .B2(_04976_),
    .ZN(_05632_));
 NAND2_X1 _17919_ (.A1(_05599_),
    .A2(_05313_),
    .ZN(_05643_));
 NAND4_X1 _17920_ (.A1(_05588_),
    .A2(_05610_),
    .A3(_05632_),
    .A4(_05643_),
    .ZN(_05654_));
 NOR4_X4 _17921_ (.A1(_05236_),
    .A2(_05379_),
    .A3(_05544_),
    .A4(_05654_),
    .ZN(_05665_));
 NOR2_X4 _17922_ (.A1(_05124_),
    .A2(_16834_),
    .ZN(_05676_));
 AND2_X4 _17923_ (.A1(_04165_),
    .A2(_05676_),
    .ZN(_05687_));
 INV_X1 _17924_ (.A(_05687_),
    .ZN(_05698_));
 AND2_X4 _17925_ (.A1(_04395_),
    .A2(_04779_),
    .ZN(_05709_));
 INV_X1 _17926_ (.A(_05709_),
    .ZN(_05720_));
 INV_X1 _17927_ (.A(_04910_),
    .ZN(_05731_));
 AOI21_X1 _17928_ (.A(_05698_),
    .B1(_05720_),
    .B2(_05731_),
    .ZN(_05742_));
 BUF_X4 _17929_ (.A(_04373_),
    .Z(_05753_));
 BUF_X4 _17930_ (.A(_05753_),
    .Z(_05764_));
 BUF_X4 _17931_ (.A(_05687_),
    .Z(_05775_));
 AND2_X1 _17932_ (.A1(_05775_),
    .A2(_04549_),
    .ZN(_05786_));
 AOI21_X1 _17933_ (.A(_05742_),
    .B1(_05764_),
    .B2(_05786_),
    .ZN(_05797_));
 AND2_X4 _17934_ (.A1(_04735_),
    .A2(_05676_),
    .ZN(_05808_));
 AND2_X1 _17935_ (.A1(_05808_),
    .A2(_05335_),
    .ZN(_05819_));
 INV_X1 _17936_ (.A(_05819_),
    .ZN(_05830_));
 BUF_X4 _17937_ (.A(_05808_),
    .Z(_05841_));
 OAI21_X2 _17938_ (.A(_05841_),
    .B1(_04976_),
    .B2(_05085_),
    .ZN(_05852_));
 BUF_X2 _17939_ (.A(_05676_),
    .Z(_05863_));
 NAND4_X1 _17940_ (.A1(_04395_),
    .A2(_05269_),
    .A3(_04932_),
    .A4(_05863_),
    .ZN(_05874_));
 NAND3_X1 _17941_ (.A1(_05830_),
    .A2(_05852_),
    .A3(_05874_),
    .ZN(_05885_));
 INV_X1 _17942_ (.A(_05401_),
    .ZN(_05896_));
 BUF_X4 _17943_ (.A(_04581_),
    .Z(_05907_));
 NOR2_X1 _17944_ (.A1(_05896_),
    .A2(_05907_),
    .ZN(_05918_));
 AND2_X2 _17945_ (.A1(_05676_),
    .A2(_04987_),
    .ZN(_05929_));
 BUF_X4 _17946_ (.A(_05929_),
    .Z(_05940_));
 AND2_X2 _17947_ (.A1(_05918_),
    .A2(_05940_),
    .ZN(_05951_));
 INV_X1 _17948_ (.A(_05929_),
    .ZN(_05962_));
 INV_X1 _17949_ (.A(_04461_),
    .ZN(_05973_));
 AND2_X4 _17950_ (.A1(_04450_),
    .A2(_04647_),
    .ZN(_05984_));
 INV_X2 _17951_ (.A(_05984_),
    .ZN(_05995_));
 AOI21_X1 _17952_ (.A(_05962_),
    .B1(_05973_),
    .B2(_05995_),
    .ZN(_06006_));
 AND3_X1 _17953_ (.A1(_04855_),
    .A2(_05467_),
    .A3(_05863_),
    .ZN(_06017_));
 NOR4_X1 _17954_ (.A1(_05885_),
    .A2(_05951_),
    .A3(_06006_),
    .A4(_06017_),
    .ZN(_06028_));
 AND2_X1 _17955_ (.A1(_05676_),
    .A2(_04329_),
    .ZN(_06039_));
 BUF_X4 _17956_ (.A(_06039_),
    .Z(_06050_));
 BUF_X4 _17957_ (.A(_06050_),
    .Z(_06061_));
 AND2_X1 _17958_ (.A1(_04779_),
    .A2(_04373_),
    .ZN(_06072_));
 OAI21_X1 _17959_ (.A(_06061_),
    .B1(_05918_),
    .B2(_06072_),
    .ZN(_06083_));
 OAI21_X1 _17960_ (.A(_06061_),
    .B1(_04658_),
    .B2(_05621_),
    .ZN(_06094_));
 AND4_X2 _17961_ (.A1(_05797_),
    .A2(_06028_),
    .A3(_06083_),
    .A4(_06094_),
    .ZN(_06105_));
 AND2_X4 _17962_ (.A1(_16835_),
    .A2(_16834_),
    .ZN(_06116_));
 BUF_X8 _17963_ (.A(_06116_),
    .Z(_06127_));
 AND2_X4 _17964_ (.A1(_06127_),
    .A2(_04329_),
    .ZN(_06138_));
 BUF_X8 _17965_ (.A(_06138_),
    .Z(_06149_));
 AND3_X1 _17966_ (.A1(_06149_),
    .A2(_05907_),
    .A3(_04833_),
    .ZN(_06160_));
 AND2_X1 _17967_ (.A1(_05621_),
    .A2(_06149_),
    .ZN(_06171_));
 AND3_X1 _17968_ (.A1(_06149_),
    .A2(_05753_),
    .A3(_04549_),
    .ZN(_06182_));
 AND2_X2 _17969_ (.A1(_05085_),
    .A2(_06149_),
    .ZN(_06193_));
 OR4_X2 _17970_ (.A1(_06160_),
    .A2(_06171_),
    .A3(_06182_),
    .A4(_06193_),
    .ZN(_06204_));
 AND2_X4 _17971_ (.A1(_04932_),
    .A2(_06127_),
    .ZN(_06215_));
 BUF_X4 _17972_ (.A(_06215_),
    .Z(_06226_));
 INV_X4 _17973_ (.A(_05566_),
    .ZN(_06237_));
 NAND2_X1 _17974_ (.A1(_06237_),
    .A2(_05995_),
    .ZN(_06248_));
 OAI21_X1 _17975_ (.A(_06226_),
    .B1(_06248_),
    .B2(_05180_),
    .ZN(_06259_));
 BUF_X4 _17976_ (.A(_05269_),
    .Z(_06270_));
 NAND4_X1 _17977_ (.A1(_06270_),
    .A2(_04932_),
    .A3(_04647_),
    .A4(_06127_),
    .ZN(_06281_));
 OAI211_X2 _17978_ (.A(_06226_),
    .B(_06270_),
    .C1(_05907_),
    .C2(_04494_),
    .ZN(_06292_));
 BUF_X16 _17979_ (.A(_06215_),
    .Z(_06303_));
 AND2_X1 _17980_ (.A1(_04833_),
    .A2(_05198_),
    .ZN(_06314_));
 AND2_X1 _17981_ (.A1(_06303_),
    .A2(_06314_),
    .ZN(_06325_));
 INV_X1 _17982_ (.A(_06325_),
    .ZN(_06336_));
 NAND4_X1 _17983_ (.A1(_06259_),
    .A2(_06281_),
    .A3(_06292_),
    .A4(_06336_),
    .ZN(_06341_));
 AND2_X4 _17984_ (.A1(_04165_),
    .A2(_06127_),
    .ZN(_06347_));
 INV_X1 _17985_ (.A(_06347_),
    .ZN(_06358_));
 AOI21_X1 _17986_ (.A(_06270_),
    .B1(_04658_),
    .B2(_04669_),
    .ZN(_06369_));
 AND2_X2 _17987_ (.A1(_05401_),
    .A2(_04395_),
    .ZN(_06380_));
 AND2_X2 _17988_ (.A1(_04581_),
    .A2(_04450_),
    .ZN(_06391_));
 NOR2_X1 _17989_ (.A1(_06380_),
    .A2(_06391_),
    .ZN(_06402_));
 AOI21_X1 _17990_ (.A(_06358_),
    .B1(_06369_),
    .B2(_06402_),
    .ZN(_06413_));
 AND2_X1 _17991_ (.A1(_04987_),
    .A2(_06116_),
    .ZN(_06424_));
 BUF_X2 _17992_ (.A(_06424_),
    .Z(_06435_));
 BUF_X4 _17993_ (.A(_06435_),
    .Z(_06446_));
 OAI211_X2 _17994_ (.A(_06446_),
    .B(_16831_),
    .C1(_04351_),
    .C2(_05907_),
    .ZN(_06457_));
 NAND2_X1 _17995_ (.A1(_05335_),
    .A2(_06446_),
    .ZN(_06468_));
 NAND2_X1 _17996_ (.A1(_05709_),
    .A2(_06435_),
    .ZN(_06479_));
 NAND2_X1 _17997_ (.A1(_06446_),
    .A2(_04549_),
    .ZN(_06490_));
 NAND4_X1 _17998_ (.A1(_06457_),
    .A2(_06468_),
    .A3(_06479_),
    .A4(_06490_),
    .ZN(_06501_));
 NOR4_X4 _17999_ (.A1(_06204_),
    .A2(_06341_),
    .A3(_06413_),
    .A4(_06501_),
    .ZN(_06512_));
 NAND4_X4 _18000_ (.A1(_05114_),
    .A2(_05665_),
    .A3(_06105_),
    .A4(_06512_),
    .ZN(_06523_));
 OAI21_X1 _18001_ (.A(_04220_),
    .B1(_04527_),
    .B2(_16830_),
    .ZN(_06534_));
 AND3_X1 _18002_ (.A1(_04187_),
    .A2(_04329_),
    .A3(_04220_),
    .ZN(_06545_));
 AND2_X1 _18003_ (.A1(_06534_),
    .A2(_06545_),
    .ZN(_06556_));
 NOR2_X4 _18004_ (.A1(_06523_),
    .A2(_06556_),
    .ZN(_06567_));
 NOR2_X1 _18005_ (.A1(_16793_),
    .A2(_16792_),
    .ZN(_06578_));
 NOR2_X1 _18006_ (.A1(_16795_),
    .A2(_16794_),
    .ZN(_06589_));
 AND2_X1 _18007_ (.A1(_06578_),
    .A2(_06589_),
    .ZN(_06600_));
 BUF_X4 _18008_ (.A(_06600_),
    .Z(_06611_));
 NOR2_X4 _18009_ (.A1(_16790_),
    .A2(_16791_),
    .ZN(_06622_));
 BUF_X8 _18010_ (.A(_06622_),
    .Z(_06633_));
 BUF_X32 _18011_ (.A(_16789_),
    .Z(_06644_));
 AND2_X2 _18012_ (.A1(_06633_),
    .A2(_06644_),
    .ZN(_06655_));
 AND2_X1 _18013_ (.A1(_06611_),
    .A2(_06655_),
    .ZN(_06666_));
 INV_X32 _18014_ (.A(_16794_),
    .ZN(_06677_));
 AND2_X4 _18015_ (.A1(_06677_),
    .A2(_16795_),
    .ZN(_06688_));
 AND2_X2 _18016_ (.A1(_16793_),
    .A2(_16792_),
    .ZN(_06699_));
 AND2_X2 _18017_ (.A1(_06688_),
    .A2(_06699_),
    .ZN(_06710_));
 INV_X4 _18018_ (.A(_06633_),
    .ZN(_06721_));
 INV_X32 _18019_ (.A(_16788_),
    .ZN(_06732_));
 NOR2_X4 _18020_ (.A1(_06732_),
    .A2(_16789_),
    .ZN(_06743_));
 NOR2_X2 _18021_ (.A1(_06721_),
    .A2(_06743_),
    .ZN(_06754_));
 AND2_X1 _18022_ (.A1(_06710_),
    .A2(_06754_),
    .ZN(_06765_));
 INV_X32 _18023_ (.A(_16790_),
    .ZN(_06776_));
 NOR2_X4 _18024_ (.A1(_06776_),
    .A2(_16791_),
    .ZN(_06787_));
 INV_X4 _18025_ (.A(_16789_),
    .ZN(_06792_));
 AND2_X2 _18026_ (.A1(_06787_),
    .A2(_06792_),
    .ZN(_06798_));
 INV_X16 _18027_ (.A(_16793_),
    .ZN(_06809_));
 NOR2_X1 _18028_ (.A1(_06809_),
    .A2(_16792_),
    .ZN(_06820_));
 AND2_X4 _18029_ (.A1(_16795_),
    .A2(_16794_),
    .ZN(_06831_));
 BUF_X8 _18030_ (.A(_06831_),
    .Z(_06842_));
 AND2_X2 _18031_ (.A1(_06820_),
    .A2(_06842_),
    .ZN(_06853_));
 AND2_X4 _18032_ (.A1(_06798_),
    .A2(_06853_),
    .ZN(_06864_));
 BUF_X32 _18033_ (.A(_16788_),
    .Z(_06875_));
 NOR2_X4 _18034_ (.A1(_06644_),
    .A2(_06875_),
    .ZN(_06886_));
 BUF_X8 _18035_ (.A(_06886_),
    .Z(_06897_));
 AND2_X2 _18036_ (.A1(_06633_),
    .A2(_06897_),
    .ZN(_06908_));
 AND2_X1 _18037_ (.A1(_06908_),
    .A2(_06600_),
    .ZN(_06919_));
 OR4_X4 _18038_ (.A1(_06666_),
    .A2(_06765_),
    .A3(_06864_),
    .A4(_06919_),
    .ZN(_06930_));
 NOR2_X4 _18039_ (.A1(_06677_),
    .A2(_16795_),
    .ZN(_06941_));
 AND2_X2 _18040_ (.A1(_06820_),
    .A2(_06941_),
    .ZN(_06952_));
 BUF_X2 _18041_ (.A(_06952_),
    .Z(_06963_));
 INV_X4 _18042_ (.A(_16791_),
    .ZN(_06974_));
 NOR2_X4 _18043_ (.A1(_06974_),
    .A2(_16790_),
    .ZN(_06985_));
 INV_X1 _18044_ (.A(_06985_),
    .ZN(_06996_));
 NOR2_X4 _18045_ (.A1(_06792_),
    .A2(_06875_),
    .ZN(_07007_));
 BUF_X8 _18046_ (.A(_07007_),
    .Z(_07018_));
 BUF_X4 _18047_ (.A(_06732_),
    .Z(_07029_));
 OAI22_X1 _18048_ (.A1(_06996_),
    .A2(_07018_),
    .B1(_07029_),
    .B2(_06721_),
    .ZN(_07040_));
 BUF_X2 _18049_ (.A(_06787_),
    .Z(_07051_));
 BUF_X4 _18050_ (.A(_07051_),
    .Z(_07062_));
 OAI21_X1 _18051_ (.A(_06963_),
    .B1(_07040_),
    .B2(_07062_),
    .ZN(_07073_));
 AND2_X2 _18052_ (.A1(_06743_),
    .A2(_06985_),
    .ZN(_07084_));
 INV_X1 _18053_ (.A(_07084_),
    .ZN(_07095_));
 AND2_X2 _18054_ (.A1(_06842_),
    .A2(_06578_),
    .ZN(_07106_));
 BUF_X4 _18055_ (.A(_07106_),
    .Z(_07117_));
 INV_X1 _18056_ (.A(_07117_),
    .ZN(_07128_));
 NOR2_X1 _18057_ (.A1(_06996_),
    .A2(_06743_),
    .ZN(_07130_));
 INV_X1 _18058_ (.A(_07130_),
    .ZN(_07139_));
 INV_X1 _18059_ (.A(_06853_),
    .ZN(_07150_));
 OAI221_X1 _18060_ (.A(_07073_),
    .B1(_07095_),
    .B2(_07128_),
    .C1(_07139_),
    .C2(_07150_),
    .ZN(_07161_));
 BUF_X4 _18061_ (.A(_06710_),
    .Z(_07172_));
 AND2_X4 _18062_ (.A1(_16790_),
    .A2(_16791_),
    .ZN(_07183_));
 AND2_X1 _18063_ (.A1(_07183_),
    .A2(_06886_),
    .ZN(_07194_));
 BUF_X4 _18064_ (.A(_07194_),
    .Z(_07205_));
 AND2_X4 _18065_ (.A1(_07183_),
    .A2(_06792_),
    .ZN(_07216_));
 BUF_X4 _18066_ (.A(_07216_),
    .Z(_07227_));
 BUF_X2 _18067_ (.A(_06589_),
    .Z(_07238_));
 AND2_X1 _18068_ (.A1(_06699_),
    .A2(_07238_),
    .ZN(_07249_));
 BUF_X4 _18069_ (.A(_07249_),
    .Z(_07260_));
 AOI22_X1 _18070_ (.A1(_07172_),
    .A2(_07205_),
    .B1(_07227_),
    .B2(_07260_),
    .ZN(_07271_));
 INV_X1 _18071_ (.A(_06787_),
    .ZN(_07282_));
 NOR2_X1 _18072_ (.A1(_07282_),
    .A2(_07018_),
    .ZN(_07293_));
 BUF_X8 _18073_ (.A(_06688_),
    .Z(_07304_));
 AND2_X2 _18074_ (.A1(_07304_),
    .A2(_06578_),
    .ZN(_07315_));
 BUF_X2 _18075_ (.A(_07315_),
    .Z(_07326_));
 NAND2_X4 _18076_ (.A1(_07293_),
    .A2(_07326_),
    .ZN(_07337_));
 INV_X1 _18077_ (.A(_06600_),
    .ZN(_07348_));
 AND2_X2 _18078_ (.A1(_06787_),
    .A2(_06644_),
    .ZN(_07359_));
 INV_X2 _18079_ (.A(_07359_),
    .ZN(_07370_));
 OAI211_X2 _18080_ (.A(_07271_),
    .B(_07337_),
    .C1(_07348_),
    .C2(_07370_),
    .ZN(_07381_));
 AND2_X2 _18081_ (.A1(_06743_),
    .A2(_06633_),
    .ZN(_07392_));
 AND2_X1 _18082_ (.A1(_06831_),
    .A2(_06699_),
    .ZN(_07403_));
 BUF_X4 _18083_ (.A(_07403_),
    .Z(_07414_));
 AND2_X4 _18084_ (.A1(_16789_),
    .A2(_06875_),
    .ZN(_07425_));
 BUF_X8 _18085_ (.A(_07425_),
    .Z(_07436_));
 BUF_X4 _18086_ (.A(_07183_),
    .Z(_07447_));
 AND2_X4 _18087_ (.A1(_07436_),
    .A2(_07447_),
    .ZN(_07458_));
 AOI22_X1 _18088_ (.A1(_07392_),
    .A2(_07414_),
    .B1(_07458_),
    .B2(_07260_),
    .ZN(_07466_));
 AND2_X2 _18089_ (.A1(_07304_),
    .A2(_06820_),
    .ZN(_07477_));
 INV_X1 _18090_ (.A(_07477_),
    .ZN(_07488_));
 AND2_X2 _18091_ (.A1(_06787_),
    .A2(_06897_),
    .ZN(_07499_));
 INV_X4 _18092_ (.A(_07499_),
    .ZN(_07510_));
 AND2_X2 _18093_ (.A1(_06941_),
    .A2(_06699_),
    .ZN(_07521_));
 BUF_X4 _18094_ (.A(_07521_),
    .Z(_07532_));
 INV_X2 _18095_ (.A(_07532_),
    .ZN(_07543_));
 AND2_X1 _18096_ (.A1(_06622_),
    .A2(_06792_),
    .ZN(_07554_));
 BUF_X2 _18097_ (.A(_07554_),
    .Z(_07565_));
 INV_X1 _18098_ (.A(_07565_),
    .ZN(_07576_));
 OAI221_X1 _18099_ (.A(_07466_),
    .B1(_07488_),
    .B2(_07510_),
    .C1(_07543_),
    .C2(_07576_),
    .ZN(_07587_));
 NOR4_X2 _18100_ (.A1(_06930_),
    .A2(_07161_),
    .A3(_07381_),
    .A4(_07587_),
    .ZN(_07598_));
 INV_X1 _18101_ (.A(_07183_),
    .ZN(_07609_));
 NOR2_X4 _18102_ (.A1(_07609_),
    .A2(_07436_),
    .ZN(_07620_));
 AND2_X2 _18103_ (.A1(_07018_),
    .A2(_06633_),
    .ZN(_07631_));
 OAI21_X1 _18104_ (.A(_07117_),
    .B1(_07620_),
    .B2(_07631_),
    .ZN(_07642_));
 BUF_X4 _18105_ (.A(_07260_),
    .Z(_07653_));
 AND2_X1 _18106_ (.A1(_07007_),
    .A2(_06787_),
    .ZN(_07664_));
 BUF_X2 _18107_ (.A(_07664_),
    .Z(_07675_));
 AND2_X1 _18108_ (.A1(_06985_),
    .A2(_06897_),
    .ZN(_07686_));
 OAI21_X1 _18109_ (.A(_07653_),
    .B1(_07675_),
    .B2(_07686_),
    .ZN(_07697_));
 AND2_X2 _18110_ (.A1(_06820_),
    .A2(_07238_),
    .ZN(_07708_));
 BUF_X4 _18111_ (.A(_07708_),
    .Z(_07719_));
 INV_X1 _18112_ (.A(_06886_),
    .ZN(_07730_));
 BUF_X2 _18113_ (.A(_06985_),
    .Z(_07740_));
 AND2_X1 _18114_ (.A1(_07730_),
    .A2(_07740_),
    .ZN(_07751_));
 NOR2_X1 _18115_ (.A1(_06721_),
    .A2(_07436_),
    .ZN(_07762_));
 OAI21_X1 _18116_ (.A(_07719_),
    .B1(_07751_),
    .B2(_07762_),
    .ZN(_07773_));
 AND2_X1 _18117_ (.A1(_06941_),
    .A2(_06578_),
    .ZN(_07784_));
 BUF_X4 _18118_ (.A(_07784_),
    .Z(_07795_));
 OAI21_X1 _18119_ (.A(_07795_),
    .B1(_07499_),
    .B2(_07565_),
    .ZN(_07806_));
 NAND4_X1 _18120_ (.A1(_07642_),
    .A2(_07697_),
    .A3(_07773_),
    .A4(_07806_),
    .ZN(_07817_));
 AND2_X4 _18121_ (.A1(_06985_),
    .A2(_07425_),
    .ZN(_07828_));
 INV_X1 _18122_ (.A(_07828_),
    .ZN(_07839_));
 INV_X1 _18123_ (.A(_07686_),
    .ZN(_07850_));
 NAND2_X1 _18124_ (.A1(_07839_),
    .A2(_07850_),
    .ZN(_07861_));
 AND2_X4 _18125_ (.A1(_06809_),
    .A2(_16792_),
    .ZN(_07872_));
 BUF_X8 _18126_ (.A(_07872_),
    .Z(_07883_));
 AND2_X4 _18127_ (.A1(_07883_),
    .A2(_06589_),
    .ZN(_07894_));
 BUF_X4 _18128_ (.A(_07894_),
    .Z(_07905_));
 AND2_X1 _18129_ (.A1(_07861_),
    .A2(_07905_),
    .ZN(_07916_));
 NOR2_X1 _18130_ (.A1(_07609_),
    .A2(_06897_),
    .ZN(_07927_));
 NAND2_X1 _18131_ (.A1(_07326_),
    .A2(_07927_),
    .ZN(_07938_));
 BUF_X4 _18132_ (.A(_07883_),
    .Z(_07949_));
 BUF_X4 _18133_ (.A(_07304_),
    .Z(_07960_));
 NAND4_X1 _18134_ (.A1(_07949_),
    .A2(_07960_),
    .A3(_06644_),
    .A4(_07447_),
    .ZN(_07971_));
 AND2_X1 _18135_ (.A1(_07872_),
    .A2(_06941_),
    .ZN(_07982_));
 INV_X1 _18136_ (.A(_07982_),
    .ZN(_07992_));
 OAI211_X2 _18137_ (.A(_07938_),
    .B(_07971_),
    .C1(_07992_),
    .C2(_07370_),
    .ZN(_08003_));
 AND2_X1 _18138_ (.A1(_07007_),
    .A2(_07183_),
    .ZN(_08014_));
 BUF_X2 _18139_ (.A(_08014_),
    .Z(_08025_));
 OAI21_X1 _18140_ (.A(_07795_),
    .B1(_08025_),
    .B2(_07227_),
    .ZN(_08036_));
 BUF_X4 _18141_ (.A(_07740_),
    .Z(_08047_));
 BUF_X2 _18142_ (.A(_06941_),
    .Z(_08058_));
 BUF_X4 _18143_ (.A(_06875_),
    .Z(_08069_));
 BUF_X2 _18144_ (.A(_06578_),
    .Z(_08080_));
 NAND4_X1 _18145_ (.A1(_08047_),
    .A2(_08058_),
    .A3(_08069_),
    .A4(_08080_),
    .ZN(_08091_));
 NAND2_X1 _18146_ (.A1(_08036_),
    .A2(_08091_),
    .ZN(_08102_));
 NOR4_X1 _18147_ (.A1(_07817_),
    .A2(_07916_),
    .A3(_08003_),
    .A4(_08102_),
    .ZN(_08113_));
 AND2_X2 _18148_ (.A1(_06787_),
    .A2(_06743_),
    .ZN(_08124_));
 INV_X1 _18149_ (.A(_08124_),
    .ZN(_08135_));
 INV_X1 _18150_ (.A(_07664_),
    .ZN(_08146_));
 NAND2_X1 _18151_ (.A1(_08135_),
    .A2(_08146_),
    .ZN(_08157_));
 NOR2_X1 _18152_ (.A1(_07609_),
    .A2(_06743_),
    .ZN(_08168_));
 OAI21_X1 _18153_ (.A(_07719_),
    .B1(_08157_),
    .B2(_08168_),
    .ZN(_08179_));
 BUF_X2 _18154_ (.A(_07982_),
    .Z(_08190_));
 AND2_X1 _18155_ (.A1(_07740_),
    .A2(_06875_),
    .ZN(_08201_));
 OR2_X1 _18156_ (.A1(_08201_),
    .A2(_07458_),
    .ZN(_08212_));
 NOR2_X2 _18157_ (.A1(_06721_),
    .A2(_07018_),
    .ZN(_08222_));
 OAI21_X1 _18158_ (.A(_08190_),
    .B1(_08212_),
    .B2(_08222_),
    .ZN(_08233_));
 INV_X1 _18159_ (.A(_07436_),
    .ZN(_08244_));
 NAND3_X1 _18160_ (.A1(_07927_),
    .A2(_07532_),
    .A3(_08244_),
    .ZN(_08255_));
 NAND2_X1 _18161_ (.A1(_07828_),
    .A2(_07532_),
    .ZN(_08266_));
 NAND2_X1 _18162_ (.A1(_08255_),
    .A2(_08266_),
    .ZN(_08277_));
 INV_X1 _18163_ (.A(_08277_),
    .ZN(_08288_));
 BUF_X2 _18164_ (.A(_06853_),
    .Z(_08299_));
 AND2_X4 _18165_ (.A1(_07425_),
    .A2(_06633_),
    .ZN(_08310_));
 INV_X1 _18166_ (.A(_08310_),
    .ZN(_08321_));
 INV_X1 _18167_ (.A(_06908_),
    .ZN(_08332_));
 NAND2_X1 _18168_ (.A1(_08321_),
    .A2(_08332_),
    .ZN(_08343_));
 AND2_X1 _18169_ (.A1(_07447_),
    .A2(_06875_),
    .ZN(_08354_));
 OAI21_X1 _18170_ (.A(_08299_),
    .B1(_08343_),
    .B2(_08354_),
    .ZN(_08365_));
 AND4_X1 _18171_ (.A1(_08179_),
    .A2(_08233_),
    .A3(_08288_),
    .A4(_08365_),
    .ZN(_08376_));
 INV_X1 _18172_ (.A(_07007_),
    .ZN(_08386_));
 BUF_X4 _18173_ (.A(_06792_),
    .Z(_08396_));
 OAI22_X1 _18174_ (.A1(_08386_),
    .A2(_07609_),
    .B1(_08396_),
    .B2(_06721_),
    .ZN(_08405_));
 OAI21_X1 _18175_ (.A(_07414_),
    .B1(_08405_),
    .B2(_08047_),
    .ZN(_08415_));
 OAI21_X1 _18176_ (.A(_07905_),
    .B1(_08124_),
    .B2(_07675_),
    .ZN(_08424_));
 INV_X1 _18177_ (.A(_06655_),
    .ZN(_08433_));
 INV_X1 _18178_ (.A(_07894_),
    .ZN(_08443_));
 OAI211_X2 _18179_ (.A(_08415_),
    .B(_08424_),
    .C1(_08433_),
    .C2(_08443_),
    .ZN(_08453_));
 AND2_X1 _18180_ (.A1(_07620_),
    .A2(_07730_),
    .ZN(_08462_));
 INV_X2 _18181_ (.A(_08462_),
    .ZN(_08472_));
 AOI22_X1 _18182_ (.A1(_08047_),
    .A2(_07730_),
    .B1(_07062_),
    .B2(_06743_),
    .ZN(_08481_));
 AOI21_X1 _18183_ (.A(_07348_),
    .B1(_08472_),
    .B2(_08481_),
    .ZN(_08491_));
 AND2_X4 _18184_ (.A1(_06787_),
    .A2(_07436_),
    .ZN(_08500_));
 NAND2_X1 _18185_ (.A1(_07172_),
    .A2(_08500_),
    .ZN(_08510_));
 BUF_X2 _18186_ (.A(_06699_),
    .Z(_08519_));
 NAND3_X1 _18187_ (.A1(_06798_),
    .A2(_07304_),
    .A3(_08519_),
    .ZN(_08528_));
 NOR2_X4 _18188_ (.A1(_06721_),
    .A2(_06897_),
    .ZN(_08532_));
 NAND2_X1 _18189_ (.A1(_08532_),
    .A2(_07653_),
    .ZN(_08533_));
 NAND2_X1 _18190_ (.A1(_07499_),
    .A2(_07414_),
    .ZN(_08534_));
 NAND4_X1 _18191_ (.A1(_08510_),
    .A2(_08528_),
    .A3(_08533_),
    .A4(_08534_),
    .ZN(_08535_));
 NOR3_X1 _18192_ (.A1(_08453_),
    .A2(_08491_),
    .A3(_08535_),
    .ZN(_08536_));
 AND4_X1 _18193_ (.A1(_07598_),
    .A2(_08113_),
    .A3(_08376_),
    .A4(_08536_),
    .ZN(_08537_));
 BUF_X4 _18194_ (.A(_06633_),
    .Z(_08538_));
 AND2_X1 _18195_ (.A1(_08538_),
    .A2(_07029_),
    .ZN(_08539_));
 OAI21_X1 _18196_ (.A(_07326_),
    .B1(_08201_),
    .B2(_08539_),
    .ZN(_08540_));
 INV_X1 _18197_ (.A(_08014_),
    .ZN(_08541_));
 INV_X1 _18198_ (.A(_06952_),
    .ZN(_08542_));
 OAI221_X1 _18199_ (.A(_08540_),
    .B1(_07839_),
    .B2(_07128_),
    .C1(_08541_),
    .C2(_08542_),
    .ZN(_08543_));
 BUF_X4 _18200_ (.A(_07477_),
    .Z(_08544_));
 AND2_X4 _18201_ (.A1(_08544_),
    .A2(_07458_),
    .ZN(_08545_));
 INV_X1 _18202_ (.A(_08545_),
    .ZN(_08546_));
 OAI21_X1 _18203_ (.A(_08544_),
    .B1(_07084_),
    .B2(_07227_),
    .ZN(_08547_));
 NAND2_X1 _18204_ (.A1(_08546_),
    .A2(_08547_),
    .ZN(_08548_));
 AND2_X1 _18205_ (.A1(_07883_),
    .A2(_06842_),
    .ZN(_08549_));
 BUF_X4 _18206_ (.A(_08549_),
    .Z(_08550_));
 INV_X1 _18207_ (.A(_08550_),
    .ZN(_08551_));
 AOI21_X1 _18208_ (.A(_08047_),
    .B1(_07927_),
    .B2(_08244_),
    .ZN(_08552_));
 NOR2_X1 _18209_ (.A1(_08124_),
    .A2(_07631_),
    .ZN(_08553_));
 AOI21_X1 _18210_ (.A(_08551_),
    .B1(_08552_),
    .B2(_08553_),
    .ZN(_08554_));
 NAND4_X1 _18211_ (.A1(_08532_),
    .A2(_07949_),
    .A3(_08244_),
    .A4(_07960_),
    .ZN(_08555_));
 AND2_X2 _18212_ (.A1(_06787_),
    .A2(_06875_),
    .ZN(_08556_));
 NAND2_X1 _18213_ (.A1(_07521_),
    .A2(_08556_),
    .ZN(_08557_));
 OAI211_X2 _18214_ (.A(_08555_),
    .B(_08557_),
    .C1(_07543_),
    .C2(_08321_),
    .ZN(_08558_));
 NOR4_X1 _18215_ (.A1(_08543_),
    .A2(_08548_),
    .A3(_08554_),
    .A4(_08558_),
    .ZN(_08559_));
 AND2_X2 _18216_ (.A1(_08537_),
    .A2(_08559_),
    .ZN(_08560_));
 XOR2_X1 _18217_ (.A(_06567_),
    .B(_08560_),
    .Z(_08561_));
 NOR2_X4 _18218_ (.A1(_16787_),
    .A2(_16786_),
    .ZN(_08562_));
 NOR2_X4 _18219_ (.A1(_16785_),
    .A2(_16784_),
    .ZN(_08563_));
 AND2_X2 _18220_ (.A1(_08562_),
    .A2(_08563_),
    .ZN(_08564_));
 BUF_X4 _18221_ (.A(_08564_),
    .Z(_08565_));
 INV_X32 _18222_ (.A(_16780_),
    .ZN(_08566_));
 NOR2_X4 _18223_ (.A1(_08566_),
    .A2(_16781_),
    .ZN(_08567_));
 INV_X32 _18224_ (.A(_16782_),
    .ZN(_08568_));
 NOR2_X4 _18225_ (.A1(_08568_),
    .A2(_16783_),
    .ZN(_08569_));
 BUF_X8 _18226_ (.A(_08569_),
    .Z(_08570_));
 AND3_X1 _18227_ (.A1(_08565_),
    .A2(_08567_),
    .A3(_08570_),
    .ZN(_08571_));
 AND2_X1 _18228_ (.A1(_08569_),
    .A2(_16781_),
    .ZN(_08572_));
 BUF_X2 _18229_ (.A(_08572_),
    .Z(_08573_));
 AND2_X1 _18230_ (.A1(_08573_),
    .A2(_08565_),
    .ZN(_08574_));
 BUF_X4 _18231_ (.A(_08565_),
    .Z(_08575_));
 NOR2_X4 _18232_ (.A1(_16783_),
    .A2(_16782_),
    .ZN(_08576_));
 AND2_X1 _18233_ (.A1(_08576_),
    .A2(_16781_),
    .ZN(_08577_));
 BUF_X2 _18234_ (.A(_08577_),
    .Z(_08578_));
 AOI211_X4 _18235_ (.A(_08571_),
    .B(_08574_),
    .C1(_08575_),
    .C2(_08578_),
    .ZN(_08579_));
 INV_X32 _18236_ (.A(_16783_),
    .ZN(_08580_));
 NOR2_X4 _18237_ (.A1(_08580_),
    .A2(_16782_),
    .ZN(_08581_));
 BUF_X2 _18238_ (.A(_08581_),
    .Z(_08582_));
 BUF_X4 _18239_ (.A(_08582_),
    .Z(_08583_));
 BUF_X4 _18240_ (.A(_16780_),
    .Z(_08584_));
 BUF_X4 _18241_ (.A(_08584_),
    .Z(_08585_));
 BUF_X4 _18242_ (.A(_16781_),
    .Z(_08586_));
 OAI211_X2 _18243_ (.A(_08575_),
    .B(_08583_),
    .C1(_08585_),
    .C2(_08586_),
    .ZN(_08587_));
 INV_X1 _18244_ (.A(_08564_),
    .ZN(_08588_));
 AND2_X4 _18245_ (.A1(_16783_),
    .A2(_16782_),
    .ZN(_08589_));
 INV_X2 _18246_ (.A(_08589_),
    .ZN(_08590_));
 NOR2_X4 _18247_ (.A1(_16780_),
    .A2(_16781_),
    .ZN(_08591_));
 BUF_X8 _18248_ (.A(_08591_),
    .Z(_08592_));
 NOR2_X1 _18249_ (.A1(_08590_),
    .A2(_08592_),
    .ZN(_08593_));
 AND2_X4 _18250_ (.A1(_16780_),
    .A2(_16781_),
    .ZN(_08594_));
 INV_X1 _18251_ (.A(_08594_),
    .ZN(_08595_));
 AND2_X1 _18252_ (.A1(_08593_),
    .A2(_08595_),
    .ZN(_08596_));
 INV_X1 _18253_ (.A(_08596_),
    .ZN(_08597_));
 OAI211_X2 _18254_ (.A(_08579_),
    .B(_08587_),
    .C1(_08588_),
    .C2(_08597_),
    .ZN(_08598_));
 BUF_X2 _18255_ (.A(_08562_),
    .Z(_08599_));
 INV_X32 _18256_ (.A(_16784_),
    .ZN(_08600_));
 NOR2_X1 _18257_ (.A1(_08600_),
    .A2(_16785_),
    .ZN(_08601_));
 BUF_X2 _18258_ (.A(_08601_),
    .Z(_08602_));
 NAND3_X1 _18259_ (.A1(_08578_),
    .A2(_08599_),
    .A3(_08602_),
    .ZN(_08603_));
 INV_X1 _18260_ (.A(_08591_),
    .ZN(_08604_));
 BUF_X8 _18261_ (.A(_08570_),
    .Z(_08605_));
 AND2_X1 _18262_ (.A1(_08604_),
    .A2(_08605_),
    .ZN(_08606_));
 AND2_X2 _18263_ (.A1(_08601_),
    .A2(_08562_),
    .ZN(_08607_));
 BUF_X4 _18264_ (.A(_08607_),
    .Z(_08608_));
 NAND3_X1 _18265_ (.A1(_08606_),
    .A2(_08608_),
    .A3(_08595_),
    .ZN(_08609_));
 NOR3_X1 _18266_ (.A1(_08567_),
    .A2(_08580_),
    .A3(_16782_),
    .ZN(_08610_));
 INV_X32 _18267_ (.A(_16781_),
    .ZN(_08611_));
 NOR2_X4 _18268_ (.A1(_08611_),
    .A2(_16780_),
    .ZN(_08612_));
 BUF_X8 _18269_ (.A(_08612_),
    .Z(_08613_));
 INV_X1 _18270_ (.A(_08613_),
    .ZN(_08614_));
 AND2_X1 _18271_ (.A1(_08610_),
    .A2(_08614_),
    .ZN(_08615_));
 INV_X1 _18272_ (.A(_08615_),
    .ZN(_08616_));
 INV_X1 _18273_ (.A(_08607_),
    .ZN(_08617_));
 OAI211_X2 _18274_ (.A(_08603_),
    .B(_08609_),
    .C1(_08616_),
    .C2(_08617_),
    .ZN(_08618_));
 AND2_X4 _18275_ (.A1(_08600_),
    .A2(_16785_),
    .ZN(_08619_));
 BUF_X4 _18276_ (.A(_08619_),
    .Z(_08620_));
 AND2_X4 _18277_ (.A1(_08620_),
    .A2(_08599_),
    .ZN(_08621_));
 BUF_X2 _18278_ (.A(_08621_),
    .Z(_08622_));
 INV_X1 _18279_ (.A(_08576_),
    .ZN(_08623_));
 NOR2_X1 _18280_ (.A1(_08623_),
    .A2(_08594_),
    .ZN(_08624_));
 AND2_X4 _18281_ (.A1(_08622_),
    .A2(_08624_),
    .ZN(_08625_));
 INV_X1 _18282_ (.A(_08625_),
    .ZN(_08626_));
 NAND3_X1 _18283_ (.A1(_08622_),
    .A2(_08606_),
    .A3(_08595_),
    .ZN(_08627_));
 AND2_X1 _18284_ (.A1(_08604_),
    .A2(_08581_),
    .ZN(_08628_));
 NAND2_X1 _18285_ (.A1(_08621_),
    .A2(_08628_),
    .ZN(_08629_));
 AND2_X2 _18286_ (.A1(_08589_),
    .A2(_08591_),
    .ZN(_08630_));
 BUF_X4 _18287_ (.A(_08630_),
    .Z(_08631_));
 AND2_X2 _18288_ (.A1(_08589_),
    .A2(_08586_),
    .ZN(_08632_));
 BUF_X4 _18289_ (.A(_08632_),
    .Z(_08633_));
 OAI21_X1 _18290_ (.A(_08622_),
    .B1(_08631_),
    .B2(_08633_),
    .ZN(_08634_));
 NAND4_X1 _18291_ (.A1(_08626_),
    .A2(_08627_),
    .A3(_08629_),
    .A4(_08634_),
    .ZN(_08635_));
 AND2_X4 _18292_ (.A1(_08613_),
    .A2(_08576_),
    .ZN(_08636_));
 BUF_X4 _18293_ (.A(_08636_),
    .Z(_08637_));
 AND2_X4 _18294_ (.A1(_16785_),
    .A2(_16784_),
    .ZN(_08638_));
 AND2_X1 _18295_ (.A1(_08638_),
    .A2(_08599_),
    .ZN(_08639_));
 BUF_X4 _18296_ (.A(_08639_),
    .Z(_08640_));
 AND2_X1 _18297_ (.A1(_08637_),
    .A2(_08640_),
    .ZN(_08641_));
 AND2_X2 _18298_ (.A1(_08576_),
    .A2(_16780_),
    .ZN(_08642_));
 AND2_X1 _18299_ (.A1(_08640_),
    .A2(_08642_),
    .ZN(_08643_));
 NOR2_X1 _18300_ (.A1(_08641_),
    .A2(_08643_),
    .ZN(_08644_));
 BUF_X8 _18301_ (.A(_08640_),
    .Z(_08645_));
 BUF_X4 _18302_ (.A(_08589_),
    .Z(_08646_));
 NAND3_X1 _18303_ (.A1(_08645_),
    .A2(_08614_),
    .A3(_08646_),
    .ZN(_08647_));
 BUF_X2 _18304_ (.A(_08612_),
    .Z(_08648_));
 BUF_X4 _18305_ (.A(_08605_),
    .Z(_08649_));
 BUF_X4 _18306_ (.A(_08638_),
    .Z(_08650_));
 NAND4_X1 _18307_ (.A1(_08648_),
    .A2(_08649_),
    .A3(_08599_),
    .A4(_08650_),
    .ZN(_08651_));
 NAND3_X1 _18308_ (.A1(_08645_),
    .A2(_08583_),
    .A3(_08592_),
    .ZN(_08652_));
 NAND4_X1 _18309_ (.A1(_08644_),
    .A2(_08647_),
    .A3(_08651_),
    .A4(_08652_),
    .ZN(_08653_));
 NOR4_X1 _18310_ (.A1(_08598_),
    .A2(_08618_),
    .A3(_08635_),
    .A4(_08653_),
    .ZN(_08654_));
 INV_X16 _18311_ (.A(_16786_),
    .ZN(_08655_));
 NOR2_X1 _18312_ (.A1(_08655_),
    .A2(_16787_),
    .ZN(_08656_));
 AND2_X2 _18313_ (.A1(_08656_),
    .A2(_08638_),
    .ZN(_08657_));
 BUF_X2 _18314_ (.A(_08657_),
    .Z(_08658_));
 INV_X2 _18315_ (.A(_08658_),
    .ZN(_08659_));
 AND2_X1 _18316_ (.A1(_08581_),
    .A2(_08594_),
    .ZN(_08660_));
 INV_X1 _18317_ (.A(_08660_),
    .ZN(_08661_));
 AND2_X2 _18318_ (.A1(_08613_),
    .A2(_08589_),
    .ZN(_08662_));
 INV_X4 _18319_ (.A(_08662_),
    .ZN(_08663_));
 AOI21_X1 _18320_ (.A(_08659_),
    .B1(_08661_),
    .B2(_08663_),
    .ZN(_08664_));
 AND2_X1 _18321_ (.A1(_08567_),
    .A2(_08589_),
    .ZN(_08665_));
 BUF_X2 _18322_ (.A(_08665_),
    .Z(_08666_));
 AND2_X1 _18323_ (.A1(_08666_),
    .A2(_08658_),
    .ZN(_08667_));
 NOR2_X1 _18324_ (.A1(_08664_),
    .A2(_08667_),
    .ZN(_08668_));
 AND2_X2 _18325_ (.A1(_08594_),
    .A2(_08576_),
    .ZN(_08669_));
 NAND2_X1 _18326_ (.A1(_08658_),
    .A2(_08669_),
    .ZN(_08670_));
 AND2_X2 _18327_ (.A1(_08570_),
    .A2(_16780_),
    .ZN(_08671_));
 NAND2_X1 _18328_ (.A1(_08671_),
    .A2(_08658_),
    .ZN(_08672_));
 AND2_X2 _18329_ (.A1(_08576_),
    .A2(_08611_),
    .ZN(_08673_));
 BUF_X4 _18330_ (.A(_08673_),
    .Z(_08674_));
 BUF_X2 _18331_ (.A(_08656_),
    .Z(_08675_));
 NAND3_X1 _18332_ (.A1(_08674_),
    .A2(_08650_),
    .A3(_08675_),
    .ZN(_08676_));
 NAND4_X1 _18333_ (.A1(_08668_),
    .A2(_08670_),
    .A3(_08672_),
    .A4(_08676_),
    .ZN(_08677_));
 AND2_X1 _18334_ (.A1(_08656_),
    .A2(_08563_),
    .ZN(_08678_));
 BUF_X2 _18335_ (.A(_08678_),
    .Z(_08679_));
 AND2_X1 _18336_ (.A1(_08589_),
    .A2(_08611_),
    .ZN(_08680_));
 BUF_X4 _18337_ (.A(_08680_),
    .Z(_08681_));
 OAI21_X1 _18338_ (.A(_08679_),
    .B1(_08662_),
    .B2(_08681_),
    .ZN(_08682_));
 BUF_X2 _18339_ (.A(_08563_),
    .Z(_08683_));
 NAND4_X1 _18340_ (.A1(_08583_),
    .A2(_08675_),
    .A3(_08584_),
    .A4(_08683_),
    .ZN(_08684_));
 AND2_X1 _18341_ (.A1(_08682_),
    .A2(_08684_),
    .ZN(_08685_));
 AND2_X1 _18342_ (.A1(_08570_),
    .A2(_08592_),
    .ZN(_08686_));
 AND2_X1 _18343_ (.A1(_08686_),
    .A2(_08679_),
    .ZN(_08687_));
 INV_X1 _18344_ (.A(_08687_),
    .ZN(_08688_));
 INV_X1 _18345_ (.A(_08674_),
    .ZN(_08689_));
 INV_X1 _18346_ (.A(_08678_),
    .ZN(_08690_));
 OAI211_X2 _18347_ (.A(_08685_),
    .B(_08688_),
    .C1(_08689_),
    .C2(_08690_),
    .ZN(_08691_));
 AND2_X1 _18348_ (.A1(_08601_),
    .A2(_08656_),
    .ZN(_08692_));
 BUF_X4 _18349_ (.A(_08692_),
    .Z(_08693_));
 BUF_X4 _18350_ (.A(_08693_),
    .Z(_08694_));
 AND2_X2 _18351_ (.A1(_08582_),
    .A2(_08584_),
    .ZN(_08695_));
 AND2_X4 _18352_ (.A1(_08594_),
    .A2(_08589_),
    .ZN(_08696_));
 BUF_X2 _18353_ (.A(_08696_),
    .Z(_08697_));
 OAI21_X1 _18354_ (.A(_08694_),
    .B1(_08695_),
    .B2(_08697_),
    .ZN(_08698_));
 NAND3_X1 _18355_ (.A1(_08674_),
    .A2(_08602_),
    .A3(_08675_),
    .ZN(_08699_));
 NAND2_X1 _18356_ (.A1(_08693_),
    .A2(_08669_),
    .ZN(_08700_));
 NAND2_X1 _18357_ (.A1(_08694_),
    .A2(_08573_),
    .ZN(_08701_));
 NAND4_X1 _18358_ (.A1(_08698_),
    .A2(_08699_),
    .A3(_08700_),
    .A4(_08701_),
    .ZN(_08702_));
 AND2_X2 _18359_ (.A1(_08619_),
    .A2(_08656_),
    .ZN(_08703_));
 BUF_X4 _18360_ (.A(_08703_),
    .Z(_08704_));
 OAI21_X1 _18361_ (.A(_08704_),
    .B1(_08642_),
    .B2(_08649_),
    .ZN(_08705_));
 BUF_X4 _18362_ (.A(_08611_),
    .Z(_08706_));
 NAND4_X1 _18363_ (.A1(_08620_),
    .A2(_08583_),
    .A3(_08675_),
    .A4(_08706_),
    .ZN(_08707_));
 NAND2_X1 _18364_ (.A1(_08704_),
    .A2(_08662_),
    .ZN(_08708_));
 BUF_X2 _18365_ (.A(_08660_),
    .Z(_08709_));
 NAND3_X1 _18366_ (.A1(_08709_),
    .A2(_08675_),
    .A3(_08620_),
    .ZN(_08710_));
 NAND4_X1 _18367_ (.A1(_08705_),
    .A2(_08707_),
    .A3(_08708_),
    .A4(_08710_),
    .ZN(_08711_));
 NOR4_X1 _18368_ (.A1(_08677_),
    .A2(_08691_),
    .A3(_08702_),
    .A4(_08711_),
    .ZN(_08712_));
 AND2_X4 _18369_ (.A1(_08655_),
    .A2(_16787_),
    .ZN(_08713_));
 AND2_X2 _18370_ (.A1(_08713_),
    .A2(_08563_),
    .ZN(_08714_));
 BUF_X4 _18371_ (.A(_08714_),
    .Z(_08715_));
 INV_X1 _18372_ (.A(_08570_),
    .ZN(_08716_));
 NOR2_X1 _18373_ (.A1(_08716_),
    .A2(_08613_),
    .ZN(_08717_));
 AND2_X1 _18374_ (.A1(_08576_),
    .A2(_08566_),
    .ZN(_08718_));
 OAI21_X1 _18375_ (.A(_08715_),
    .B1(_08717_),
    .B2(_08718_),
    .ZN(_08719_));
 AND2_X2 _18376_ (.A1(_08619_),
    .A2(_08713_),
    .ZN(_08720_));
 BUF_X4 _18377_ (.A(_08720_),
    .Z(_08721_));
 OAI21_X1 _18378_ (.A(_08721_),
    .B1(_08697_),
    .B2(_08680_),
    .ZN(_08722_));
 AND2_X1 _18379_ (.A1(_08581_),
    .A2(_08611_),
    .ZN(_08723_));
 BUF_X2 _18380_ (.A(_08723_),
    .Z(_08724_));
 BUF_X2 _18381_ (.A(_08713_),
    .Z(_08725_));
 NAND4_X1 _18382_ (.A1(_08724_),
    .A2(_08584_),
    .A3(_08725_),
    .A4(_08620_),
    .ZN(_08726_));
 AND2_X1 _18383_ (.A1(_08722_),
    .A2(_08726_),
    .ZN(_08727_));
 NAND3_X1 _18384_ (.A1(_08631_),
    .A2(_08725_),
    .A3(_08650_),
    .ZN(_08728_));
 NAND2_X1 _18385_ (.A1(_08720_),
    .A2(_08686_),
    .ZN(_08729_));
 AND2_X2 _18386_ (.A1(_08713_),
    .A2(_08638_),
    .ZN(_08730_));
 BUF_X4 _18387_ (.A(_08730_),
    .Z(_08731_));
 NOR2_X1 _18388_ (.A1(_08623_),
    .A2(_08567_),
    .ZN(_08732_));
 OAI21_X1 _18389_ (.A(_08731_),
    .B1(_08717_),
    .B2(_08732_),
    .ZN(_08733_));
 AND4_X1 _18390_ (.A1(_08727_),
    .A2(_08728_),
    .A3(_08729_),
    .A4(_08733_),
    .ZN(_08734_));
 INV_X1 _18391_ (.A(_08714_),
    .ZN(_08735_));
 INV_X1 _18392_ (.A(_08666_),
    .ZN(_08736_));
 INV_X1 _18393_ (.A(_08632_),
    .ZN(_08737_));
 AOI21_X1 _18394_ (.A(_08735_),
    .B1(_08736_),
    .B2(_08737_),
    .ZN(_08738_));
 AOI21_X1 _18395_ (.A(_08738_),
    .B1(_08695_),
    .B2(_08715_),
    .ZN(_08739_));
 AND2_X4 _18396_ (.A1(_08713_),
    .A2(_08601_),
    .ZN(_08740_));
 BUF_X2 _18397_ (.A(_08740_),
    .Z(_08741_));
 AND3_X1 _18398_ (.A1(_08741_),
    .A2(_08604_),
    .A3(_08624_),
    .ZN(_08742_));
 AOI21_X1 _18399_ (.A(_08742_),
    .B1(_08741_),
    .B2(_08633_),
    .ZN(_08743_));
 AND4_X1 _18400_ (.A1(_08719_),
    .A2(_08734_),
    .A3(_08739_),
    .A4(_08743_),
    .ZN(_08744_));
 AND2_X4 _18401_ (.A1(_16787_),
    .A2(_16786_),
    .ZN(_08745_));
 AND2_X4 _18402_ (.A1(_08602_),
    .A2(_08745_),
    .ZN(_08746_));
 BUF_X4 _18403_ (.A(_08746_),
    .Z(_08747_));
 BUF_X4 _18404_ (.A(_08747_),
    .Z(_08748_));
 AND2_X2 _18405_ (.A1(_08567_),
    .A2(_08569_),
    .ZN(_08749_));
 OR3_X4 _18406_ (.A1(_08666_),
    .A2(_08749_),
    .A3(_08637_),
    .ZN(_08750_));
 AOI21_X1 _18407_ (.A(_08580_),
    .B1(_08614_),
    .B2(_16782_),
    .ZN(_08751_));
 OAI21_X1 _18408_ (.A(_08748_),
    .B1(_08750_),
    .B2(_08751_),
    .ZN(_08752_));
 BUF_X4 _18409_ (.A(_08576_),
    .Z(_08753_));
 BUF_X2 _18410_ (.A(_08745_),
    .Z(_08754_));
 AND4_X1 _18411_ (.A1(_08563_),
    .A2(_08648_),
    .A3(_08753_),
    .A4(_08754_),
    .ZN(_08755_));
 AND2_X4 _18412_ (.A1(_08745_),
    .A2(_08563_),
    .ZN(_08756_));
 INV_X1 _18413_ (.A(_08756_),
    .ZN(_08757_));
 INV_X1 _18414_ (.A(_08680_),
    .ZN(_08758_));
 AOI21_X1 _18415_ (.A(_08757_),
    .B1(_08663_),
    .B2(_08758_),
    .ZN(_08759_));
 BUF_X4 _18416_ (.A(_08756_),
    .Z(_08760_));
 AOI211_X4 _18417_ (.A(_08755_),
    .B(_08759_),
    .C1(_08695_),
    .C2(_08760_),
    .ZN(_08761_));
 INV_X1 _18418_ (.A(_08567_),
    .ZN(_08762_));
 NOR2_X1 _18419_ (.A1(_08623_),
    .A2(_08648_),
    .ZN(_08763_));
 AND4_X1 _18420_ (.A1(_08762_),
    .A2(_08763_),
    .A3(_08754_),
    .A4(_08620_),
    .ZN(_08764_));
 AND2_X2 _18421_ (.A1(_08619_),
    .A2(_08745_),
    .ZN(_08765_));
 BUF_X4 _18422_ (.A(_08765_),
    .Z(_08766_));
 AND2_X2 _18423_ (.A1(_08570_),
    .A2(_08611_),
    .ZN(_08767_));
 AND2_X1 _18424_ (.A1(_08766_),
    .A2(_08767_),
    .ZN(_08768_));
 AND2_X1 _18425_ (.A1(_08766_),
    .A2(_08610_),
    .ZN(_08769_));
 AND2_X2 _18426_ (.A1(_08646_),
    .A2(_16780_),
    .ZN(_08770_));
 AND2_X1 _18427_ (.A1(_08766_),
    .A2(_08770_),
    .ZN(_08771_));
 NOR4_X1 _18428_ (.A1(_08764_),
    .A2(_08768_),
    .A3(_08769_),
    .A4(_08771_),
    .ZN(_08772_));
 AND2_X1 _18429_ (.A1(_08638_),
    .A2(_08745_),
    .ZN(_08773_));
 BUF_X4 _18430_ (.A(_08773_),
    .Z(_08774_));
 AND2_X1 _18431_ (.A1(_08686_),
    .A2(_08774_),
    .ZN(_08775_));
 INV_X1 _18432_ (.A(_08775_),
    .ZN(_08776_));
 OAI211_X2 _18433_ (.A(_08774_),
    .B(_08753_),
    .C1(_08584_),
    .C2(_08586_),
    .ZN(_08777_));
 AND2_X1 _18434_ (.A1(_08581_),
    .A2(_16781_),
    .ZN(_08778_));
 BUF_X2 _18435_ (.A(_08778_),
    .Z(_08779_));
 OAI21_X1 _18436_ (.A(_08774_),
    .B1(_08779_),
    .B2(_08724_),
    .ZN(_08780_));
 NAND3_X1 _18437_ (.A1(_08774_),
    .A2(_08648_),
    .A3(_08646_),
    .ZN(_08781_));
 AND4_X1 _18438_ (.A1(_08776_),
    .A2(_08777_),
    .A3(_08780_),
    .A4(_08781_),
    .ZN(_08782_));
 AND4_X1 _18439_ (.A1(_08752_),
    .A2(_08761_),
    .A3(_08772_),
    .A4(_08782_),
    .ZN(_08783_));
 NAND4_X1 _18440_ (.A1(_08654_),
    .A2(_08712_),
    .A3(_08744_),
    .A4(_08783_),
    .ZN(_08784_));
 AND2_X2 _18441_ (.A1(_08591_),
    .A2(_08576_),
    .ZN(_08785_));
 AND2_X1 _18442_ (.A1(_08564_),
    .A2(_08785_),
    .ZN(_08786_));
 NOR2_X2 _18443_ (.A1(_08784_),
    .A2(_08786_),
    .ZN(_08787_));
 BUF_X4 _18444_ (.A(_08774_),
    .Z(_08788_));
 AND2_X2 _18445_ (.A1(_08581_),
    .A2(_08567_),
    .ZN(_08789_));
 AND2_X1 _18446_ (.A1(_08646_),
    .A2(_08566_),
    .ZN(_08790_));
 OAI21_X1 _18447_ (.A(_08788_),
    .B1(_08789_),
    .B2(_08790_),
    .ZN(_08791_));
 AND2_X2 _18448_ (.A1(_08766_),
    .A2(_08673_),
    .ZN(_08792_));
 NAND3_X1 _18449_ (.A1(_08572_),
    .A2(_08754_),
    .A3(_08619_),
    .ZN(_08793_));
 INV_X1 _18450_ (.A(_08765_),
    .ZN(_08794_));
 INV_X1 _18451_ (.A(_08749_),
    .ZN(_08795_));
 OAI21_X1 _18452_ (.A(_08793_),
    .B1(_08794_),
    .B2(_08795_),
    .ZN(_08796_));
 AOI211_X2 _18453_ (.A(_08792_),
    .B(_08796_),
    .C1(_08637_),
    .C2(_08766_),
    .ZN(_08797_));
 BUF_X4 _18454_ (.A(_08767_),
    .Z(_08798_));
 OAI21_X1 _18455_ (.A(_08788_),
    .B1(_08798_),
    .B2(_08624_),
    .ZN(_08799_));
 NOR2_X1 _18456_ (.A1(_08590_),
    .A2(_08613_),
    .ZN(_08800_));
 OAI211_X2 _18457_ (.A(_08766_),
    .B(_08762_),
    .C1(_08800_),
    .C2(_08583_),
    .ZN(_08801_));
 AND4_X1 _18458_ (.A1(_08791_),
    .A2(_08797_),
    .A3(_08799_),
    .A4(_08801_),
    .ZN(_08802_));
 OAI21_X1 _18459_ (.A(_08760_),
    .B1(_08606_),
    .B2(_08785_),
    .ZN(_08803_));
 AND2_X1 _18460_ (.A1(_08723_),
    .A2(_08756_),
    .ZN(_08804_));
 AND2_X1 _18461_ (.A1(_08665_),
    .A2(_08756_),
    .ZN(_08805_));
 AOI211_X2 _18462_ (.A(_08804_),
    .B(_08805_),
    .C1(_08632_),
    .C2(_08756_),
    .ZN(_08806_));
 OAI21_X1 _18463_ (.A(_08748_),
    .B1(_08800_),
    .B2(_08709_),
    .ZN(_08807_));
 NAND2_X1 _18464_ (.A1(_08637_),
    .A2(_08747_),
    .ZN(_08808_));
 AND2_X4 _18465_ (.A1(_08612_),
    .A2(_08570_),
    .ZN(_08809_));
 BUF_X4 _18466_ (.A(_08809_),
    .Z(_08810_));
 NAND2_X1 _18467_ (.A1(_08810_),
    .A2(_08747_),
    .ZN(_08811_));
 AND2_X1 _18468_ (.A1(_08808_),
    .A2(_08811_),
    .ZN(_08812_));
 AND4_X1 _18469_ (.A1(_08803_),
    .A2(_08806_),
    .A3(_08807_),
    .A4(_08812_),
    .ZN(_08813_));
 OAI21_X1 _18470_ (.A(_08741_),
    .B1(_08573_),
    .B2(_08642_),
    .ZN(_08814_));
 AND2_X2 _18471_ (.A1(_08628_),
    .A2(_08595_),
    .ZN(_08815_));
 OR2_X1 _18472_ (.A1(_08696_),
    .A2(_08630_),
    .ZN(_08816_));
 OAI21_X1 _18473_ (.A(_08741_),
    .B1(_08815_),
    .B2(_08816_),
    .ZN(_08817_));
 AND3_X1 _18474_ (.A1(_08724_),
    .A2(_08683_),
    .A3(_08725_),
    .ZN(_08818_));
 INV_X1 _18475_ (.A(_08818_),
    .ZN(_08819_));
 INV_X1 _18476_ (.A(_08669_),
    .ZN(_08820_));
 INV_X1 _18477_ (.A(_08785_),
    .ZN(_08821_));
 NAND2_X1 _18478_ (.A1(_08820_),
    .A2(_08821_),
    .ZN(_08822_));
 OAI21_X1 _18479_ (.A(_08715_),
    .B1(_08822_),
    .B2(_08749_),
    .ZN(_08823_));
 AND4_X1 _18480_ (.A1(_08814_),
    .A2(_08817_),
    .A3(_08819_),
    .A4(_08823_),
    .ZN(_08824_));
 NOR2_X1 _18481_ (.A1(_08778_),
    .A2(_08662_),
    .ZN(_08825_));
 INV_X1 _18482_ (.A(_08730_),
    .ZN(_08826_));
 NOR2_X1 _18483_ (.A1(_08825_),
    .A2(_08826_),
    .ZN(_08827_));
 INV_X1 _18484_ (.A(_08827_),
    .ZN(_08828_));
 NAND2_X1 _18485_ (.A1(_08721_),
    .A2(_08785_),
    .ZN(_08829_));
 BUF_X2 _18486_ (.A(_08566_),
    .Z(_08830_));
 OAI221_X1 _18487_ (.A(_08721_),
    .B1(_08830_),
    .B2(_08706_),
    .C1(_08583_),
    .C2(_08646_),
    .ZN(_08831_));
 OAI21_X1 _18488_ (.A(_08731_),
    .B1(_08717_),
    .B2(_08674_),
    .ZN(_08832_));
 AND4_X1 _18489_ (.A1(_08828_),
    .A2(_08829_),
    .A3(_08831_),
    .A4(_08832_),
    .ZN(_08833_));
 NAND4_X2 _18490_ (.A1(_08802_),
    .A2(_08813_),
    .A3(_08824_),
    .A4(_08833_),
    .ZN(_08834_));
 AND2_X1 _18491_ (.A1(_08724_),
    .A2(_08658_),
    .ZN(_08835_));
 AND2_X4 _18492_ (.A1(_08581_),
    .A2(_08613_),
    .ZN(_08836_));
 AND2_X1 _18493_ (.A1(_08836_),
    .A2(_08657_),
    .ZN(_08837_));
 NOR2_X1 _18494_ (.A1(_08835_),
    .A2(_08837_),
    .ZN(_08838_));
 INV_X1 _18495_ (.A(_08703_),
    .ZN(_08839_));
 INV_X1 _18496_ (.A(_08789_),
    .ZN(_08840_));
 AOI21_X1 _18497_ (.A(_08839_),
    .B1(_08840_),
    .B2(_08737_),
    .ZN(_08841_));
 AND2_X1 _18498_ (.A1(_08703_),
    .A2(_08578_),
    .ZN(_08842_));
 AND2_X4 _18499_ (.A1(_08570_),
    .A2(_08594_),
    .ZN(_08843_));
 AND2_X1 _18500_ (.A1(_08703_),
    .A2(_08843_),
    .ZN(_08844_));
 AND2_X1 _18501_ (.A1(_08703_),
    .A2(_08673_),
    .ZN(_08845_));
 NOR4_X1 _18502_ (.A1(_08841_),
    .A2(_08842_),
    .A3(_08844_),
    .A4(_08845_),
    .ZN(_08846_));
 AND2_X2 _18503_ (.A1(_08593_),
    .A2(_08657_),
    .ZN(_08847_));
 INV_X1 _18504_ (.A(_08847_),
    .ZN(_08848_));
 AND2_X1 _18505_ (.A1(_08657_),
    .A2(_08642_),
    .ZN(_08849_));
 AND2_X1 _18506_ (.A1(_08843_),
    .A2(_08657_),
    .ZN(_08850_));
 AOI211_X2 _18507_ (.A(_08849_),
    .B(_08850_),
    .C1(_08767_),
    .C2(_08657_),
    .ZN(_08851_));
 AND4_X1 _18508_ (.A1(_08838_),
    .A2(_08846_),
    .A3(_08848_),
    .A4(_08851_),
    .ZN(_08852_));
 NAND2_X1 _18509_ (.A1(_08749_),
    .A2(_08693_),
    .ZN(_08853_));
 INV_X1 _18510_ (.A(_08809_),
    .ZN(_08854_));
 INV_X1 _18511_ (.A(_08693_),
    .ZN(_08855_));
 OAI21_X1 _18512_ (.A(_08853_),
    .B1(_08854_),
    .B2(_08855_),
    .ZN(_08856_));
 AOI21_X1 _18513_ (.A(_08856_),
    .B1(_08694_),
    .B2(_08642_),
    .ZN(_08857_));
 OAI21_X1 _18514_ (.A(_08693_),
    .B1(_08815_),
    .B2(_08697_),
    .ZN(_08858_));
 AND2_X1 _18515_ (.A1(_08567_),
    .A2(_08576_),
    .ZN(_08859_));
 BUF_X4 _18516_ (.A(_08859_),
    .Z(_08860_));
 OAI21_X1 _18517_ (.A(_08679_),
    .B1(_08860_),
    .B2(_08843_),
    .ZN(_08861_));
 OAI21_X1 _18518_ (.A(_08679_),
    .B1(_08779_),
    .B2(_08770_),
    .ZN(_08862_));
 AND4_X1 _18519_ (.A1(_08857_),
    .A2(_08858_),
    .A3(_08861_),
    .A4(_08862_),
    .ZN(_08863_));
 AND3_X1 _18520_ (.A1(_08717_),
    .A2(_08762_),
    .A3(_08607_),
    .ZN(_08864_));
 INV_X1 _18521_ (.A(_08864_),
    .ZN(_08865_));
 NAND3_X1 _18522_ (.A1(_08673_),
    .A2(_08599_),
    .A3(_08602_),
    .ZN(_08866_));
 NAND4_X1 _18523_ (.A1(_08648_),
    .A2(_08602_),
    .A3(_08599_),
    .A4(_08753_),
    .ZN(_08867_));
 NAND3_X1 _18524_ (.A1(_08865_),
    .A2(_08866_),
    .A3(_08867_),
    .ZN(_08868_));
 AOI211_X4 _18525_ (.A(_08590_),
    .B(_08617_),
    .C1(_08830_),
    .C2(_08586_),
    .ZN(_08869_));
 NAND4_X1 _18526_ (.A1(_08565_),
    .A2(_08614_),
    .A3(_08762_),
    .A4(_08605_),
    .ZN(_08870_));
 NAND2_X4 _18527_ (.A1(_08681_),
    .A2(_08575_),
    .ZN(_08871_));
 OAI211_X2 _18528_ (.A(_08870_),
    .B(_08871_),
    .C1(_08663_),
    .C2(_08588_),
    .ZN(_08872_));
 INV_X4 _18529_ (.A(_08778_),
    .ZN(_08873_));
 INV_X1 _18530_ (.A(_08723_),
    .ZN(_08874_));
 AOI21_X1 _18531_ (.A(_08617_),
    .B1(_08873_),
    .B2(_08874_),
    .ZN(_08875_));
 NOR4_X2 _18532_ (.A1(_08868_),
    .A2(_08869_),
    .A3(_08872_),
    .A4(_08875_),
    .ZN(_08876_));
 AND2_X1 _18533_ (.A1(_08671_),
    .A2(_08640_),
    .ZN(_08877_));
 INV_X1 _18534_ (.A(_08877_),
    .ZN(_08878_));
 INV_X1 _18535_ (.A(_08643_),
    .ZN(_08879_));
 OAI21_X1 _18536_ (.A(_08645_),
    .B1(_08779_),
    .B2(_08790_),
    .ZN(_08880_));
 NAND3_X1 _18537_ (.A1(_08878_),
    .A2(_08879_),
    .A3(_08880_),
    .ZN(_08881_));
 AND2_X1 _18538_ (.A1(_08621_),
    .A2(_08573_),
    .ZN(_08882_));
 NAND2_X1 _18539_ (.A1(_08621_),
    .A2(_08666_),
    .ZN(_08883_));
 NAND2_X1 _18540_ (.A1(_08629_),
    .A2(_08883_),
    .ZN(_08884_));
 NOR4_X1 _18541_ (.A1(_08881_),
    .A2(_08625_),
    .A3(_08882_),
    .A4(_08884_),
    .ZN(_08885_));
 NAND4_X1 _18542_ (.A1(_08852_),
    .A2(_08863_),
    .A3(_08876_),
    .A4(_08885_),
    .ZN(_08886_));
 NOR2_X4 _18543_ (.A1(_08834_),
    .A2(_08886_),
    .ZN(_08887_));
 XNOR2_X1 _18544_ (.A(_08787_),
    .B(_08887_),
    .ZN(_08888_));
 XNOR2_X1 _18545_ (.A(_08561_),
    .B(_08888_),
    .ZN(_08889_));
 INV_X32 _18546_ (.A(_16875_),
    .ZN(_08890_));
 AND2_X4 _18547_ (.A1(_08890_),
    .A2(_16874_),
    .ZN(_08891_));
 AND2_X4 _18548_ (.A1(_16873_),
    .A2(_16872_),
    .ZN(_08892_));
 AND2_X2 _18549_ (.A1(_08891_),
    .A2(_08892_),
    .ZN(_08893_));
 INV_X32 _18550_ (.A(_16871_),
    .ZN(_08894_));
 NOR2_X4 _18551_ (.A1(_08894_),
    .A2(_16870_),
    .ZN(_08895_));
 INV_X32 _18552_ (.A(_16869_),
    .ZN(_08896_));
 NOR2_X4 _18553_ (.A1(_08896_),
    .A2(_16868_),
    .ZN(_08897_));
 AND2_X1 _18554_ (.A1(_08895_),
    .A2(_08897_),
    .ZN(_08898_));
 BUF_X2 _18555_ (.A(_08898_),
    .Z(_08899_));
 BUF_X32 _18556_ (.A(_08896_),
    .Z(_08900_));
 AND2_X2 _18557_ (.A1(_08895_),
    .A2(_08900_),
    .ZN(_08901_));
 OAI21_X1 _18558_ (.A(_08893_),
    .B1(_08899_),
    .B2(_08901_),
    .ZN(_08902_));
 INV_X32 _18559_ (.A(_16872_),
    .ZN(_08903_));
 AND2_X2 _18560_ (.A1(_08903_),
    .A2(_16873_),
    .ZN(_08904_));
 BUF_X8 _18561_ (.A(_08891_),
    .Z(_08905_));
 AND2_X2 _18562_ (.A1(_08904_),
    .A2(_08905_),
    .ZN(_08906_));
 INV_X32 _18563_ (.A(_16868_),
    .ZN(_08907_));
 BUF_X32 _18564_ (.A(_16869_),
    .Z(_08908_));
 NOR2_X4 _18565_ (.A1(_08907_),
    .A2(_08908_),
    .ZN(_08909_));
 AND2_X2 _18566_ (.A1(_08895_),
    .A2(_08909_),
    .ZN(_08910_));
 AND2_X4 _18567_ (.A1(_16871_),
    .A2(_16870_),
    .ZN(_08911_));
 AND2_X4 _18568_ (.A1(_08911_),
    .A2(_08908_),
    .ZN(_08912_));
 OAI21_X1 _18569_ (.A(_08906_),
    .B1(_08910_),
    .B2(_08912_),
    .ZN(_08913_));
 INV_X32 _18570_ (.A(_16870_),
    .ZN(_08914_));
 NOR2_X4 _18571_ (.A1(_08914_),
    .A2(_16871_),
    .ZN(_08915_));
 BUF_X4 _18572_ (.A(_08915_),
    .Z(_08916_));
 AND2_X4 _18573_ (.A1(_16868_),
    .A2(_16869_),
    .ZN(_08917_));
 BUF_X16 _18574_ (.A(_08917_),
    .Z(_08918_));
 AND2_X4 _18575_ (.A1(_08916_),
    .A2(_08918_),
    .ZN(_08919_));
 NAND2_X1 _18576_ (.A1(_08906_),
    .A2(_08919_),
    .ZN(_08920_));
 BUF_X4 _18577_ (.A(_08904_),
    .Z(_08921_));
 NOR2_X4 _18578_ (.A1(_16871_),
    .A2(_16870_),
    .ZN(_08922_));
 AND2_X1 _18579_ (.A1(_08922_),
    .A2(_08896_),
    .ZN(_08923_));
 BUF_X4 _18580_ (.A(_08923_),
    .Z(_08924_));
 BUF_X8 _18581_ (.A(_08922_),
    .Z(_08925_));
 AND2_X2 _18582_ (.A1(_08925_),
    .A2(_08908_),
    .ZN(_08926_));
 OAI211_X2 _18583_ (.A(_08921_),
    .B(_08905_),
    .C1(_08924_),
    .C2(_08926_),
    .ZN(_08927_));
 AND3_X1 _18584_ (.A1(_08913_),
    .A2(_08920_),
    .A3(_08927_),
    .ZN(_08928_));
 BUF_X32 _18585_ (.A(_16868_),
    .Z(_08929_));
 NOR2_X4 _18586_ (.A1(_08929_),
    .A2(_08908_),
    .ZN(_08930_));
 INV_X2 _18587_ (.A(_08930_),
    .ZN(_08931_));
 BUF_X2 _18588_ (.A(_08911_),
    .Z(_08932_));
 NAND2_X4 _18589_ (.A1(_08931_),
    .A2(_08932_),
    .ZN(_08933_));
 INV_X1 _18590_ (.A(_08933_),
    .ZN(_08934_));
 AND2_X1 _18591_ (.A1(_08934_),
    .A2(_08893_),
    .ZN(_08935_));
 INV_X1 _18592_ (.A(_08935_),
    .ZN(_08936_));
 AND2_X2 _18593_ (.A1(_08925_),
    .A2(_08929_),
    .ZN(_08937_));
 NAND2_X1 _18594_ (.A1(_08893_),
    .A2(_08937_),
    .ZN(_08938_));
 AND2_X2 _18595_ (.A1(_08915_),
    .A2(_08900_),
    .ZN(_08939_));
 NAND2_X1 _18596_ (.A1(_08893_),
    .A2(_08939_),
    .ZN(_08940_));
 NAND2_X1 _18597_ (.A1(_08893_),
    .A2(_08919_),
    .ZN(_08941_));
 AND3_X1 _18598_ (.A1(_08938_),
    .A2(_08940_),
    .A3(_08941_),
    .ZN(_08942_));
 AND4_X1 _18599_ (.A1(_08902_),
    .A2(_08928_),
    .A3(_08936_),
    .A4(_08942_),
    .ZN(_08943_));
 NOR2_X1 _18600_ (.A1(_16875_),
    .A2(_16874_),
    .ZN(_08944_));
 NOR2_X4 _18601_ (.A1(_16873_),
    .A2(_16872_),
    .ZN(_08945_));
 AND2_X1 _18602_ (.A1(_08944_),
    .A2(_08945_),
    .ZN(_08946_));
 BUF_X4 _18603_ (.A(_08946_),
    .Z(_08947_));
 AND2_X2 _18604_ (.A1(_08915_),
    .A2(_08930_),
    .ZN(_08948_));
 OAI21_X1 _18605_ (.A(_08947_),
    .B1(_08948_),
    .B2(_08919_),
    .ZN(_08949_));
 NOR2_X2 _18606_ (.A1(_08903_),
    .A2(_16873_),
    .ZN(_08950_));
 AND2_X1 _18607_ (.A1(_08950_),
    .A2(_08944_),
    .ZN(_08951_));
 AND2_X1 _18608_ (.A1(_08951_),
    .A2(_08923_),
    .ZN(_08952_));
 BUF_X4 _18609_ (.A(_08951_),
    .Z(_08953_));
 BUF_X8 _18610_ (.A(_08897_),
    .Z(_08954_));
 AND2_X2 _18611_ (.A1(_08954_),
    .A2(_08925_),
    .ZN(_08955_));
 INV_X1 _18612_ (.A(_08897_),
    .ZN(_08956_));
 AND2_X4 _18613_ (.A1(_08956_),
    .A2(_08915_),
    .ZN(_08957_));
 AND2_X1 _18614_ (.A1(_08957_),
    .A2(_08953_),
    .ZN(_08958_));
 INV_X1 _18615_ (.A(_08909_),
    .ZN(_08959_));
 AOI221_X1 _18616_ (.A(_08952_),
    .B1(_08953_),
    .B2(_08955_),
    .C1(_08958_),
    .C2(_08959_),
    .ZN(_08960_));
 BUF_X4 _18617_ (.A(_08932_),
    .Z(_08961_));
 BUF_X4 _18618_ (.A(_08907_),
    .Z(_08962_));
 OAI211_X2 _18619_ (.A(_08947_),
    .B(_08961_),
    .C1(_08962_),
    .C2(_08900_),
    .ZN(_08963_));
 AND2_X4 _18620_ (.A1(_08895_),
    .A2(_08908_),
    .ZN(_08964_));
 OAI21_X1 _18621_ (.A(_08953_),
    .B1(_08901_),
    .B2(_08964_),
    .ZN(_08965_));
 AND2_X1 _18622_ (.A1(_08911_),
    .A2(_08900_),
    .ZN(_08966_));
 NAND2_X1 _18623_ (.A1(_08953_),
    .A2(_08966_),
    .ZN(_08967_));
 AND2_X4 _18624_ (.A1(_08918_),
    .A2(_08911_),
    .ZN(_08968_));
 BUF_X8 _18625_ (.A(_08968_),
    .Z(_08969_));
 NAND2_X1 _18626_ (.A1(_08953_),
    .A2(_08969_),
    .ZN(_08970_));
 AND3_X1 _18627_ (.A1(_08965_),
    .A2(_08967_),
    .A3(_08970_),
    .ZN(_08971_));
 AND4_X1 _18628_ (.A1(_08949_),
    .A2(_08960_),
    .A3(_08963_),
    .A4(_08971_),
    .ZN(_08972_));
 AND2_X2 _18629_ (.A1(_08891_),
    .A2(_08950_),
    .ZN(_08973_));
 AND2_X1 _18630_ (.A1(_08909_),
    .A2(_08915_),
    .ZN(_08974_));
 AND2_X1 _18631_ (.A1(_08954_),
    .A2(_08915_),
    .ZN(_08975_));
 OAI21_X1 _18632_ (.A(_08973_),
    .B1(_08974_),
    .B2(_08975_),
    .ZN(_08976_));
 BUF_X4 _18633_ (.A(_08925_),
    .Z(_08977_));
 NAND4_X1 _18634_ (.A1(_08905_),
    .A2(_08929_),
    .A3(_08950_),
    .A4(_08977_),
    .ZN(_08978_));
 AND2_X1 _18635_ (.A1(_08976_),
    .A2(_08978_),
    .ZN(_08979_));
 NAND2_X1 _18636_ (.A1(_08931_),
    .A2(_08895_),
    .ZN(_08980_));
 NOR2_X2 _18637_ (.A1(_08980_),
    .A2(_08918_),
    .ZN(_08981_));
 OAI21_X1 _18638_ (.A(_08973_),
    .B1(_08981_),
    .B2(_08969_),
    .ZN(_08982_));
 AND2_X2 _18639_ (.A1(_08905_),
    .A2(_08945_),
    .ZN(_08983_));
 AND2_X2 _18640_ (.A1(_08909_),
    .A2(_08925_),
    .ZN(_08984_));
 BUF_X2 _18641_ (.A(_08984_),
    .Z(_08985_));
 OAI21_X1 _18642_ (.A(_08983_),
    .B1(_08919_),
    .B2(_08985_),
    .ZN(_08986_));
 BUF_X2 _18643_ (.A(_08964_),
    .Z(_08987_));
 AND2_X2 _18644_ (.A1(_08932_),
    .A2(_08929_),
    .ZN(_08988_));
 OAI21_X1 _18645_ (.A(_08983_),
    .B1(_08987_),
    .B2(_08988_),
    .ZN(_08989_));
 AND4_X1 _18646_ (.A1(_08979_),
    .A2(_08982_),
    .A3(_08986_),
    .A4(_08989_),
    .ZN(_08990_));
 AND2_X2 _18647_ (.A1(_08904_),
    .A2(_08944_),
    .ZN(_08991_));
 INV_X4 _18648_ (.A(_08991_),
    .ZN(_08992_));
 INV_X2 _18649_ (.A(_08918_),
    .ZN(_08993_));
 NAND2_X1 _18650_ (.A1(_08993_),
    .A2(_08925_),
    .ZN(_08994_));
 NOR2_X1 _18651_ (.A1(_08992_),
    .A2(_08994_),
    .ZN(_08995_));
 INV_X1 _18652_ (.A(_08995_),
    .ZN(_08996_));
 OR2_X1 _18653_ (.A1(_08992_),
    .A2(_08980_),
    .ZN(_08997_));
 AND2_X2 _18654_ (.A1(_08916_),
    .A2(_08908_),
    .ZN(_08998_));
 AND2_X1 _18655_ (.A1(_08991_),
    .A2(_08998_),
    .ZN(_08999_));
 INV_X1 _18656_ (.A(_08999_),
    .ZN(_09000_));
 AND2_X1 _18657_ (.A1(_08909_),
    .A2(_08911_),
    .ZN(_09001_));
 BUF_X4 _18658_ (.A(_09001_),
    .Z(_09002_));
 NAND2_X1 _18659_ (.A1(_08991_),
    .A2(_09002_),
    .ZN(_09003_));
 NAND4_X1 _18660_ (.A1(_08996_),
    .A2(_08997_),
    .A3(_09000_),
    .A4(_09003_),
    .ZN(_09004_));
 AND2_X2 _18661_ (.A1(_08892_),
    .A2(_08944_),
    .ZN(_09005_));
 AND2_X1 _18662_ (.A1(_09005_),
    .A2(_08937_),
    .ZN(_09006_));
 AND3_X1 _18663_ (.A1(_09005_),
    .A2(_08929_),
    .A3(_08916_),
    .ZN(_09007_));
 INV_X1 _18664_ (.A(_09005_),
    .ZN(_09008_));
 INV_X1 _18665_ (.A(_08987_),
    .ZN(_09009_));
 AND2_X1 _18666_ (.A1(_08932_),
    .A2(_08907_),
    .ZN(_09010_));
 INV_X1 _18667_ (.A(_09010_),
    .ZN(_09011_));
 AOI21_X1 _18668_ (.A(_09008_),
    .B1(_09009_),
    .B2(_09011_),
    .ZN(_09012_));
 NOR4_X1 _18669_ (.A1(_09004_),
    .A2(_09006_),
    .A3(_09007_),
    .A4(_09012_),
    .ZN(_09013_));
 AND4_X1 _18670_ (.A1(_08943_),
    .A2(_08972_),
    .A3(_08990_),
    .A4(_09013_),
    .ZN(_09014_));
 AND2_X4 _18671_ (.A1(_16875_),
    .A2(_16874_),
    .ZN(_09015_));
 AND2_X2 _18672_ (.A1(_08904_),
    .A2(_09015_),
    .ZN(_09016_));
 BUF_X4 _18673_ (.A(_08930_),
    .Z(_09017_));
 AND2_X2 _18674_ (.A1(_08911_),
    .A2(_09017_),
    .ZN(_09018_));
 AND2_X2 _18675_ (.A1(_09016_),
    .A2(_09018_),
    .ZN(_09019_));
 INV_X1 _18676_ (.A(_09019_),
    .ZN(_09020_));
 AND3_X1 _18677_ (.A1(_08969_),
    .A2(_08921_),
    .A3(_09015_),
    .ZN(_09021_));
 INV_X1 _18678_ (.A(_09021_),
    .ZN(_09022_));
 INV_X1 _18679_ (.A(_09016_),
    .ZN(_09023_));
 NAND2_X4 _18680_ (.A1(_08959_),
    .A2(_08895_),
    .ZN(_09024_));
 OAI211_X2 _18681_ (.A(_09020_),
    .B(_09022_),
    .C1(_09023_),
    .C2(_09024_),
    .ZN(_09025_));
 BUF_X4 _18682_ (.A(_08974_),
    .Z(_09026_));
 OAI21_X1 _18683_ (.A(_09016_),
    .B1(_09026_),
    .B2(_08998_),
    .ZN(_09027_));
 NAND2_X1 _18684_ (.A1(_09016_),
    .A2(_08924_),
    .ZN(_09028_));
 INV_X1 _18685_ (.A(_08955_),
    .ZN(_09029_));
 OAI211_X2 _18686_ (.A(_09027_),
    .B(_09028_),
    .C1(_09023_),
    .C2(_09029_),
    .ZN(_09030_));
 AND2_X4 _18687_ (.A1(_08892_),
    .A2(_09015_),
    .ZN(_09031_));
 INV_X1 _18688_ (.A(_09031_),
    .ZN(_09032_));
 INV_X1 _18689_ (.A(_08910_),
    .ZN(_09033_));
 AOI21_X1 _18690_ (.A(_09032_),
    .B1(_09033_),
    .B2(_09011_),
    .ZN(_09034_));
 INV_X1 _18691_ (.A(_08939_),
    .ZN(_09035_));
 AOI21_X1 _18692_ (.A(_09032_),
    .B1(_09035_),
    .B2(_08994_),
    .ZN(_09036_));
 NOR4_X1 _18693_ (.A1(_09025_),
    .A2(_09030_),
    .A3(_09034_),
    .A4(_09036_),
    .ZN(_09037_));
 AND2_X4 _18694_ (.A1(_09015_),
    .A2(_08945_),
    .ZN(_09038_));
 BUF_X4 _18695_ (.A(_09038_),
    .Z(_09039_));
 NAND2_X1 _18696_ (.A1(_08901_),
    .A2(_09039_),
    .ZN(_09040_));
 AND2_X2 _18697_ (.A1(_08950_),
    .A2(_09015_),
    .ZN(_09041_));
 NAND2_X1 _18698_ (.A1(_08955_),
    .A2(_09041_),
    .ZN(_09042_));
 NAND2_X1 _18699_ (.A1(_08975_),
    .A2(_09041_),
    .ZN(_09043_));
 AND2_X1 _18700_ (.A1(_09042_),
    .A2(_09043_),
    .ZN(_09044_));
 AND2_X1 _18701_ (.A1(_08895_),
    .A2(_08917_),
    .ZN(_09045_));
 AND2_X1 _18702_ (.A1(_09045_),
    .A2(_09041_),
    .ZN(_09046_));
 INV_X1 _18703_ (.A(_09046_),
    .ZN(_09047_));
 OAI211_X2 _18704_ (.A(_09041_),
    .B(_08932_),
    .C1(_08929_),
    .C2(_08900_),
    .ZN(_09048_));
 AND3_X1 _18705_ (.A1(_09044_),
    .A2(_09047_),
    .A3(_09048_),
    .ZN(_09049_));
 AND3_X1 _18706_ (.A1(_08916_),
    .A2(_08945_),
    .A3(_09015_),
    .ZN(_09050_));
 AND2_X2 _18707_ (.A1(_08925_),
    .A2(_08930_),
    .ZN(_09051_));
 AOI22_X1 _18708_ (.A1(_09050_),
    .A2(_08931_),
    .B1(_09039_),
    .B2(_09051_),
    .ZN(_09052_));
 BUF_X4 _18709_ (.A(_09039_),
    .Z(_09053_));
 BUF_X4 _18710_ (.A(_08929_),
    .Z(_09054_));
 OAI211_X2 _18711_ (.A(_09053_),
    .B(_08961_),
    .C1(_09054_),
    .C2(_08908_),
    .ZN(_09055_));
 AND4_X1 _18712_ (.A1(_09040_),
    .A2(_09049_),
    .A3(_09052_),
    .A4(_09055_),
    .ZN(_09056_));
 NOR2_X2 _18713_ (.A1(_08890_),
    .A2(_16874_),
    .ZN(_09057_));
 AND2_X2 _18714_ (.A1(_08950_),
    .A2(_09057_),
    .ZN(_09058_));
 AND2_X1 _18715_ (.A1(_08981_),
    .A2(_09058_),
    .ZN(_09059_));
 INV_X1 _18716_ (.A(_09059_),
    .ZN(_09060_));
 NOR2_X1 _18717_ (.A1(_08969_),
    .A2(_09018_),
    .ZN(_09061_));
 INV_X1 _18718_ (.A(_09058_),
    .ZN(_09062_));
 OAI21_X1 _18719_ (.A(_09060_),
    .B1(_09061_),
    .B2(_09062_),
    .ZN(_09063_));
 AND2_X2 _18720_ (.A1(_09057_),
    .A2(_08945_),
    .ZN(_09064_));
 AND2_X1 _18721_ (.A1(_08901_),
    .A2(_09064_),
    .ZN(_09065_));
 INV_X1 _18722_ (.A(_08937_),
    .ZN(_09066_));
 INV_X1 _18723_ (.A(_08998_),
    .ZN(_09067_));
 AOI21_X1 _18724_ (.A(_09062_),
    .B1(_09066_),
    .B2(_09067_),
    .ZN(_09068_));
 AND2_X1 _18725_ (.A1(_08917_),
    .A2(_08925_),
    .ZN(_09069_));
 INV_X2 _18726_ (.A(_09069_),
    .ZN(_09070_));
 INV_X4 _18727_ (.A(_09051_),
    .ZN(_09071_));
 NAND2_X4 _18728_ (.A1(_09070_),
    .A2(_09071_),
    .ZN(_09072_));
 NAND2_X1 _18729_ (.A1(_09072_),
    .A2(_09064_),
    .ZN(_09073_));
 BUF_X2 _18730_ (.A(_09064_),
    .Z(_09074_));
 NAND2_X1 _18731_ (.A1(_09026_),
    .A2(_09074_),
    .ZN(_09075_));
 NAND2_X1 _18732_ (.A1(_09073_),
    .A2(_09075_),
    .ZN(_09076_));
 NOR4_X1 _18733_ (.A1(_09063_),
    .A2(_09065_),
    .A3(_09068_),
    .A4(_09076_),
    .ZN(_09077_));
 AND2_X1 _18734_ (.A1(_09057_),
    .A2(_08892_),
    .ZN(_09078_));
 AND2_X2 _18735_ (.A1(_08954_),
    .A2(_08911_),
    .ZN(_09079_));
 AND2_X1 _18736_ (.A1(_09078_),
    .A2(_09079_),
    .ZN(_09080_));
 BUF_X2 _18737_ (.A(_09078_),
    .Z(_09081_));
 AND2_X1 _18738_ (.A1(_09081_),
    .A2(_08964_),
    .ZN(_09082_));
 NOR2_X1 _18739_ (.A1(_09080_),
    .A2(_09082_),
    .ZN(_09083_));
 AND2_X2 _18740_ (.A1(_08904_),
    .A2(_09057_),
    .ZN(_09084_));
 AND2_X1 _18741_ (.A1(_09084_),
    .A2(_09051_),
    .ZN(_09085_));
 INV_X1 _18742_ (.A(_09085_),
    .ZN(_09086_));
 BUF_X4 _18743_ (.A(_08895_),
    .Z(_09087_));
 OAI221_X1 _18744_ (.A(_09084_),
    .B1(_08907_),
    .B2(_08900_),
    .C1(_09087_),
    .C2(_08932_),
    .ZN(_09088_));
 OAI21_X1 _18745_ (.A(_09081_),
    .B1(_08957_),
    .B2(_08924_),
    .ZN(_09089_));
 AND4_X1 _18746_ (.A1(_09083_),
    .A2(_09086_),
    .A3(_09088_),
    .A4(_09089_),
    .ZN(_09090_));
 AND4_X1 _18747_ (.A1(_09037_),
    .A2(_09056_),
    .A3(_09077_),
    .A4(_09090_),
    .ZN(_09091_));
 AND2_X2 _18748_ (.A1(_09014_),
    .A2(_09091_),
    .ZN(_09092_));
 BUF_X4 _18749_ (.A(_09092_),
    .Z(_09093_));
 XNOR2_X1 _18750_ (.A(_08889_),
    .B(_09093_),
    .ZN(_09094_));
 INV_X2 _18751_ (.A(_04121_),
    .ZN(_09095_));
 BUF_X4 _18752_ (.A(_09095_),
    .Z(_09096_));
 XNOR2_X1 _18753_ (.A(_09094_),
    .B(_09096_),
    .ZN(_09097_));
 INV_X2 _18754_ (.A(_01331_),
    .ZN(_09098_));
 BUF_X4 _18755_ (.A(_09098_),
    .Z(_09099_));
 BUF_X4 _18756_ (.A(_09099_),
    .Z(_09100_));
 MUX2_X1 _18757_ (.A(_04143_),
    .B(_09097_),
    .S(_09100_),
    .Z(_00724_));
 BUF_X4 _18758_ (.A(_17155_),
    .Z(_09101_));
 XOR2_X1 _18759_ (.A(_09101_),
    .B(_17051_),
    .Z(_09102_));
 AND2_X4 _18760_ (.A1(_16789_),
    .A2(_16791_),
    .ZN(_09103_));
 NAND2_X4 _18761_ (.A1(_09103_),
    .A2(_06776_),
    .ZN(_09104_));
 INV_X1 _18762_ (.A(_09104_),
    .ZN(_09105_));
 BUF_X4 _18763_ (.A(_09105_),
    .Z(_09106_));
 OAI21_X1 _18764_ (.A(_07905_),
    .B1(_08025_),
    .B2(_09106_),
    .ZN(_09107_));
 NAND4_X1 _18765_ (.A1(_07949_),
    .A2(_07062_),
    .A3(_07029_),
    .A4(_07238_),
    .ZN(_09108_));
 OAI211_X2 _18766_ (.A(_09107_),
    .B(_09108_),
    .C1(_07576_),
    .C2(_08443_),
    .ZN(_09109_));
 INV_X1 _18767_ (.A(_06666_),
    .ZN(_09110_));
 NAND2_X1 _18768_ (.A1(_07227_),
    .A2(_06611_),
    .ZN(_09111_));
 AND2_X1 _18769_ (.A1(_08244_),
    .A2(_07051_),
    .ZN(_09112_));
 NAND2_X1 _18770_ (.A1(_09112_),
    .A2(_06611_),
    .ZN(_09113_));
 NAND2_X1 _18771_ (.A1(_06611_),
    .A2(_09103_),
    .ZN(_09114_));
 NAND4_X1 _18772_ (.A1(_09110_),
    .A2(_09111_),
    .A3(_09113_),
    .A4(_09114_),
    .ZN(_09115_));
 OAI211_X2 _18773_ (.A(_07653_),
    .B(_08047_),
    .C1(_08396_),
    .C2(_08069_),
    .ZN(_09116_));
 OAI211_X2 _18774_ (.A(_07260_),
    .B(_07447_),
    .C1(_08396_),
    .C2(_07029_),
    .ZN(_09117_));
 NAND2_X1 _18775_ (.A1(_08556_),
    .A2(_07653_),
    .ZN(_09118_));
 NAND4_X1 _18776_ (.A1(_09116_),
    .A2(_09117_),
    .A3(_08533_),
    .A4(_09118_),
    .ZN(_09119_));
 INV_X1 _18777_ (.A(_07708_),
    .ZN(_09120_));
 INV_X1 _18778_ (.A(_09112_),
    .ZN(_09121_));
 INV_X1 _18779_ (.A(_06754_),
    .ZN(_09122_));
 AOI21_X1 _18780_ (.A(_09120_),
    .B1(_09121_),
    .B2(_09122_),
    .ZN(_09123_));
 NOR4_X1 _18781_ (.A1(_09109_),
    .A2(_09115_),
    .A3(_09119_),
    .A4(_09123_),
    .ZN(_09124_));
 AND2_X2 _18782_ (.A1(_06743_),
    .A2(_07183_),
    .ZN(_09125_));
 AND2_X1 _18783_ (.A1(_09125_),
    .A2(_07784_),
    .ZN(_09126_));
 NAND4_X1 _18784_ (.A1(_07740_),
    .A2(_06941_),
    .A3(_08396_),
    .A4(_06578_),
    .ZN(_09127_));
 INV_X1 _18785_ (.A(_07784_),
    .ZN(_09128_));
 OAI21_X1 _18786_ (.A(_09127_),
    .B1(_09104_),
    .B2(_09128_),
    .ZN(_09129_));
 AOI211_X4 _18787_ (.A(_09126_),
    .B(_09129_),
    .C1(_08025_),
    .C2(_07784_),
    .ZN(_09130_));
 BUF_X4 _18788_ (.A(_06798_),
    .Z(_09131_));
 OAI21_X1 _18789_ (.A(_07795_),
    .B1(_07675_),
    .B2(_09131_),
    .ZN(_09132_));
 AND2_X2 _18790_ (.A1(_06633_),
    .A2(_06875_),
    .ZN(_09133_));
 INV_X1 _18791_ (.A(_09133_),
    .ZN(_09134_));
 OAI211_X2 _18792_ (.A(_09130_),
    .B(_09132_),
    .C1(_09134_),
    .C2(_09128_),
    .ZN(_09135_));
 NOR2_X2 _18793_ (.A1(_06974_),
    .A2(_06644_),
    .ZN(_09136_));
 AND2_X2 _18794_ (.A1(_09136_),
    .A2(_06776_),
    .ZN(_09137_));
 BUF_X4 _18795_ (.A(_09137_),
    .Z(_09138_));
 AND2_X1 _18796_ (.A1(_08190_),
    .A2(_09138_),
    .ZN(_09139_));
 INV_X4 _18797_ (.A(_08500_),
    .ZN(_09140_));
 AOI21_X1 _18798_ (.A(_07992_),
    .B1(_08332_),
    .B2(_09140_),
    .ZN(_09141_));
 AND2_X2 _18799_ (.A1(_07007_),
    .A2(_06985_),
    .ZN(_09142_));
 AND2_X1 _18800_ (.A1(_07982_),
    .A2(_09142_),
    .ZN(_09143_));
 NOR2_X1 _18801_ (.A1(_07609_),
    .A2(_07007_),
    .ZN(_09144_));
 INV_X1 _18802_ (.A(_06743_),
    .ZN(_09145_));
 AND3_X1 _18803_ (.A1(_07982_),
    .A2(_09144_),
    .A3(_09145_),
    .ZN(_09146_));
 OR4_X1 _18804_ (.A1(_09139_),
    .A2(_09141_),
    .A3(_09143_),
    .A4(_09146_),
    .ZN(_09147_));
 OAI21_X1 _18805_ (.A(_06963_),
    .B1(_08025_),
    .B2(_09106_),
    .ZN(_09148_));
 NAND2_X1 _18806_ (.A1(_06963_),
    .A2(_08532_),
    .ZN(_09149_));
 NAND4_X1 _18807_ (.A1(_07062_),
    .A2(_06820_),
    .A3(_08058_),
    .A4(_07029_),
    .ZN(_09150_));
 NAND3_X1 _18808_ (.A1(_09148_),
    .A2(_09149_),
    .A3(_09150_),
    .ZN(_09151_));
 AND2_X1 _18809_ (.A1(_07927_),
    .A2(_07521_),
    .ZN(_09152_));
 NOR3_X2 _18810_ (.A1(_07436_),
    .A2(_16790_),
    .A3(_06974_),
    .ZN(_09153_));
 AND3_X1 _18811_ (.A1(_07521_),
    .A2(_07730_),
    .A3(_09153_),
    .ZN(_09154_));
 AND2_X1 _18812_ (.A1(_07521_),
    .A2(_09133_),
    .ZN(_09155_));
 AND4_X1 _18813_ (.A1(_07051_),
    .A2(_08058_),
    .A3(_06897_),
    .A4(_08519_),
    .ZN(_09156_));
 OR4_X1 _18814_ (.A1(_09152_),
    .A2(_09154_),
    .A3(_09155_),
    .A4(_09156_),
    .ZN(_09157_));
 NOR4_X1 _18815_ (.A1(_09135_),
    .A2(_09147_),
    .A3(_09151_),
    .A4(_09157_),
    .ZN(_09158_));
 OAI21_X4 _18816_ (.A(_06853_),
    .B1(_07458_),
    .B2(_07194_),
    .ZN(_09159_));
 NAND2_X1 _18817_ (.A1(_09138_),
    .A2(_06853_),
    .ZN(_09160_));
 INV_X1 _18818_ (.A(_09142_),
    .ZN(_09161_));
 OAI211_X2 _18819_ (.A(_09159_),
    .B(_09160_),
    .C1(_09161_),
    .C2(_07150_),
    .ZN(_09162_));
 INV_X2 _18820_ (.A(_07403_),
    .ZN(_09163_));
 AOI211_X4 _18821_ (.A(_07282_),
    .B(_09163_),
    .C1(_06644_),
    .C2(_06875_),
    .ZN(_09164_));
 AND2_X4 _18822_ (.A1(_09103_),
    .A2(_16790_),
    .ZN(_09165_));
 BUF_X4 _18823_ (.A(_09165_),
    .Z(_09166_));
 INV_X1 _18824_ (.A(_09166_),
    .ZN(_09167_));
 AOI21_X1 _18825_ (.A(_09163_),
    .B1(_07839_),
    .B2(_09167_),
    .ZN(_09168_));
 AND2_X1 _18826_ (.A1(_07675_),
    .A2(_06853_),
    .ZN(_09169_));
 OR4_X1 _18827_ (.A1(_09162_),
    .A2(_09164_),
    .A3(_09168_),
    .A4(_09169_),
    .ZN(_09170_));
 NAND3_X1 _18828_ (.A1(_08124_),
    .A2(_07949_),
    .A3(_06842_),
    .ZN(_09171_));
 NAND3_X1 _18829_ (.A1(_07359_),
    .A2(_07949_),
    .A3(_06842_),
    .ZN(_09172_));
 OAI211_X2 _18830_ (.A(_09171_),
    .B(_09172_),
    .C1(_08551_),
    .C2(_09134_),
    .ZN(_09173_));
 OAI21_X1 _18831_ (.A(_08550_),
    .B1(_07458_),
    .B2(_07205_),
    .ZN(_09174_));
 OAI21_X1 _18832_ (.A(_09174_),
    .B1(_08551_),
    .B2(_09161_),
    .ZN(_09175_));
 OAI21_X1 _18833_ (.A(_07117_),
    .B1(_08343_),
    .B2(_08556_),
    .ZN(_09176_));
 AND2_X1 _18834_ (.A1(_07828_),
    .A2(_07106_),
    .ZN(_09177_));
 INV_X1 _18835_ (.A(_09177_),
    .ZN(_09178_));
 AND2_X1 _18836_ (.A1(_07205_),
    .A2(_07106_),
    .ZN(_09179_));
 INV_X1 _18837_ (.A(_09179_),
    .ZN(_09180_));
 NAND2_X1 _18838_ (.A1(_07106_),
    .A2(_09166_),
    .ZN(_09181_));
 NAND4_X1 _18839_ (.A1(_09176_),
    .A2(_09178_),
    .A3(_09180_),
    .A4(_09181_),
    .ZN(_09182_));
 NOR4_X1 _18840_ (.A1(_09170_),
    .A2(_09173_),
    .A3(_09175_),
    .A4(_09182_),
    .ZN(_09183_));
 NAND4_X1 _18841_ (.A1(_07960_),
    .A2(_08538_),
    .A3(_07018_),
    .A4(_08080_),
    .ZN(_09184_));
 AND2_X2 _18842_ (.A1(_07337_),
    .A2(_09184_),
    .ZN(_09185_));
 NAND2_X1 _18843_ (.A1(_07326_),
    .A2(_07458_),
    .ZN(_09186_));
 INV_X1 _18844_ (.A(_07315_),
    .ZN(_09187_));
 AND2_X2 _18845_ (.A1(_09153_),
    .A2(_07730_),
    .ZN(_09188_));
 INV_X1 _18846_ (.A(_09188_),
    .ZN(_09189_));
 OAI211_X2 _18847_ (.A(_09185_),
    .B(_09186_),
    .C1(_09187_),
    .C2(_09189_),
    .ZN(_09190_));
 AND2_X1 _18848_ (.A1(_07872_),
    .A2(_06688_),
    .ZN(_09191_));
 BUF_X2 _18849_ (.A(_09191_),
    .Z(_09192_));
 NAND2_X1 _18850_ (.A1(_09192_),
    .A2(_09131_),
    .ZN(_09193_));
 NAND3_X1 _18851_ (.A1(_07631_),
    .A2(_07883_),
    .A3(_07960_),
    .ZN(_09194_));
 NAND2_X1 _18852_ (.A1(_09193_),
    .A2(_09194_),
    .ZN(_09195_));
 AND2_X1 _18853_ (.A1(_09192_),
    .A2(_07447_),
    .ZN(_09196_));
 AND2_X1 _18854_ (.A1(_09191_),
    .A2(_09138_),
    .ZN(_09197_));
 OR3_X1 _18855_ (.A1(_09195_),
    .A2(_09196_),
    .A3(_09197_),
    .ZN(_09198_));
 NOR2_X1 _18856_ (.A1(_06996_),
    .A2(_07018_),
    .ZN(_09199_));
 AND2_X1 _18857_ (.A1(_09199_),
    .A2(_07477_),
    .ZN(_09200_));
 INV_X1 _18858_ (.A(_09200_),
    .ZN(_09201_));
 NAND2_X1 _18859_ (.A1(_07477_),
    .A2(_08124_),
    .ZN(_09202_));
 NAND2_X1 _18860_ (.A1(_08544_),
    .A2(_07392_),
    .ZN(_09203_));
 NAND2_X1 _18861_ (.A1(_08544_),
    .A2(_06655_),
    .ZN(_09204_));
 NAND4_X1 _18862_ (.A1(_09201_),
    .A2(_09202_),
    .A3(_09203_),
    .A4(_09204_),
    .ZN(_09205_));
 OAI21_X1 _18863_ (.A(_07172_),
    .B1(_09125_),
    .B2(_08025_),
    .ZN(_09206_));
 OAI21_X1 _18864_ (.A(_07172_),
    .B1(_07675_),
    .B2(_08539_),
    .ZN(_09207_));
 NAND4_X1 _18865_ (.A1(_07960_),
    .A2(_08069_),
    .A3(_08047_),
    .A4(_08519_),
    .ZN(_09208_));
 NAND3_X1 _18866_ (.A1(_09206_),
    .A2(_09207_),
    .A3(_09208_),
    .ZN(_09209_));
 NOR4_X1 _18867_ (.A1(_09190_),
    .A2(_09198_),
    .A3(_09205_),
    .A4(_09209_),
    .ZN(_09210_));
 AND4_X1 _18868_ (.A1(_09124_),
    .A2(_09158_),
    .A3(_09183_),
    .A4(_09210_),
    .ZN(_09211_));
 INV_X1 _18869_ (.A(_06919_),
    .ZN(_09212_));
 AND2_X2 _18870_ (.A1(_09211_),
    .A2(_09212_),
    .ZN(_09213_));
 AND2_X1 _18871_ (.A1(_08720_),
    .A2(_08577_),
    .ZN(_09214_));
 AND2_X1 _18872_ (.A1(_08720_),
    .A2(_08859_),
    .ZN(_09215_));
 AOI211_X4 _18873_ (.A(_09214_),
    .B(_09215_),
    .C1(_08749_),
    .C2(_08721_),
    .ZN(_09216_));
 OAI21_X1 _18874_ (.A(_08731_),
    .B1(_08596_),
    .B2(_08695_),
    .ZN(_09217_));
 INV_X1 _18875_ (.A(_08582_),
    .ZN(_09218_));
 NOR2_X1 _18876_ (.A1(_09218_),
    .A2(_08648_),
    .ZN(_09219_));
 NAND2_X1 _18877_ (.A1(_09219_),
    .A2(_08721_),
    .ZN(_09220_));
 OAI21_X1 _18878_ (.A(_08731_),
    .B1(_08810_),
    .B2(_08718_),
    .ZN(_09221_));
 NAND4_X1 _18879_ (.A1(_09216_),
    .A2(_09217_),
    .A3(_09220_),
    .A4(_09221_),
    .ZN(_09222_));
 NAND2_X1 _18880_ (.A1(_08717_),
    .A2(_08715_),
    .ZN(_09223_));
 NAND4_X1 _18881_ (.A1(_08725_),
    .A2(_08683_),
    .A3(_08648_),
    .A4(_08753_),
    .ZN(_09224_));
 NAND2_X1 _18882_ (.A1(_09223_),
    .A2(_09224_),
    .ZN(_09225_));
 NAND2_X1 _18883_ (.A1(_08715_),
    .A2(_08697_),
    .ZN(_09226_));
 INV_X1 _18884_ (.A(_08815_),
    .ZN(_09227_));
 OAI21_X1 _18885_ (.A(_09226_),
    .B1(_09227_),
    .B2(_08735_),
    .ZN(_09228_));
 OAI21_X1 _18886_ (.A(_08741_),
    .B1(_08637_),
    .B2(_08798_),
    .ZN(_09229_));
 NAND2_X1 _18887_ (.A1(_08740_),
    .A2(_08723_),
    .ZN(_09230_));
 INV_X4 _18888_ (.A(_08740_),
    .ZN(_09231_));
 OAI211_X2 _18889_ (.A(_09229_),
    .B(_09230_),
    .C1(_08590_),
    .C2(_09231_),
    .ZN(_09232_));
 NOR4_X1 _18890_ (.A1(_09222_),
    .A2(_09225_),
    .A3(_09228_),
    .A4(_09232_),
    .ZN(_09233_));
 INV_X1 _18891_ (.A(_08767_),
    .ZN(_09234_));
 AOI21_X1 _18892_ (.A(_08588_),
    .B1(_08854_),
    .B2(_09234_),
    .ZN(_09235_));
 AOI211_X4 _18893_ (.A(_08580_),
    .B(_08588_),
    .C1(_08611_),
    .C2(_08568_),
    .ZN(_09236_));
 AOI211_X4 _18894_ (.A(_09235_),
    .B(_09236_),
    .C1(_08575_),
    .C2(_08578_),
    .ZN(_09237_));
 AND2_X1 _18895_ (.A1(_08662_),
    .A2(_08607_),
    .ZN(_09238_));
 AND2_X1 _18896_ (.A1(_08570_),
    .A2(_08566_),
    .ZN(_09239_));
 INV_X1 _18897_ (.A(_09239_),
    .ZN(_09240_));
 OAI21_X1 _18898_ (.A(_08866_),
    .B1(_08617_),
    .B2(_09240_),
    .ZN(_09241_));
 AOI211_X4 _18899_ (.A(_09238_),
    .B(_09241_),
    .C1(_08779_),
    .C2(_08607_),
    .ZN(_09242_));
 AND2_X1 _18900_ (.A1(_08595_),
    .A2(_08605_),
    .ZN(_09243_));
 OAI21_X1 _18901_ (.A(_08622_),
    .B1(_09243_),
    .B2(_08732_),
    .ZN(_09244_));
 OAI211_X2 _18902_ (.A(_08645_),
    .B(_08583_),
    .C1(_08585_),
    .C2(_08706_),
    .ZN(_09245_));
 OAI211_X2 _18903_ (.A(_08640_),
    .B(_08646_),
    .C1(_08830_),
    .C2(_08706_),
    .ZN(_09246_));
 AND4_X1 _18904_ (.A1(_08644_),
    .A2(_08878_),
    .A3(_09245_),
    .A4(_09246_),
    .ZN(_09247_));
 AND4_X1 _18905_ (.A1(_09237_),
    .A2(_09242_),
    .A3(_09244_),
    .A4(_09247_),
    .ZN(_09248_));
 AND4_X1 _18906_ (.A1(_08582_),
    .A2(_08613_),
    .A3(_08602_),
    .A4(_08745_),
    .ZN(_09249_));
 AND3_X1 _18907_ (.A1(_08630_),
    .A2(_08602_),
    .A3(_08754_),
    .ZN(_09250_));
 AOI211_X4 _18908_ (.A(_09249_),
    .B(_09250_),
    .C1(_08697_),
    .C2(_08747_),
    .ZN(_09251_));
 NAND4_X1 _18909_ (.A1(_08602_),
    .A2(_08585_),
    .A3(_08754_),
    .A4(_08753_),
    .ZN(_09252_));
 OAI211_X2 _18910_ (.A(_08748_),
    .B(_08649_),
    .C1(_08585_),
    .C2(_08586_),
    .ZN(_09253_));
 AND3_X1 _18911_ (.A1(_09251_),
    .A2(_09252_),
    .A3(_09253_),
    .ZN(_09254_));
 NAND2_X1 _18912_ (.A1(_08709_),
    .A2(_08760_),
    .ZN(_09255_));
 OAI21_X1 _18913_ (.A(_08760_),
    .B1(_08822_),
    .B2(_08671_),
    .ZN(_09256_));
 NAND2_X1 _18914_ (.A1(_08756_),
    .A2(_08632_),
    .ZN(_09257_));
 NAND2_X1 _18915_ (.A1(_08631_),
    .A2(_08760_),
    .ZN(_09258_));
 AND4_X1 _18916_ (.A1(_09255_),
    .A2(_09256_),
    .A3(_09257_),
    .A4(_09258_),
    .ZN(_09259_));
 AND2_X1 _18917_ (.A1(_08766_),
    .A2(_08810_),
    .ZN(_09260_));
 INV_X1 _18918_ (.A(_08836_),
    .ZN(_09261_));
 AOI21_X1 _18919_ (.A(_08794_),
    .B1(_09261_),
    .B2(_08874_),
    .ZN(_09262_));
 AOI211_X4 _18920_ (.A(_09260_),
    .B(_09262_),
    .C1(_08766_),
    .C2(_08816_),
    .ZN(_09263_));
 AND4_X1 _18921_ (.A1(_08582_),
    .A2(_08594_),
    .A3(_08650_),
    .A4(_08754_),
    .ZN(_09264_));
 NAND2_X1 _18922_ (.A1(_08767_),
    .A2(_08774_),
    .ZN(_09265_));
 INV_X1 _18923_ (.A(_08774_),
    .ZN(_09266_));
 OAI21_X1 _18924_ (.A(_09265_),
    .B1(_08854_),
    .B2(_09266_),
    .ZN(_09267_));
 AOI211_X4 _18925_ (.A(_09264_),
    .B(_09267_),
    .C1(_08633_),
    .C2(_08774_),
    .ZN(_09268_));
 AND4_X1 _18926_ (.A1(_09254_),
    .A2(_09259_),
    .A3(_09263_),
    .A4(_09268_),
    .ZN(_09269_));
 AND2_X1 _18927_ (.A1(_09243_),
    .A2(_08679_),
    .ZN(_09270_));
 AOI21_X1 _18928_ (.A(_08690_),
    .B1(_08873_),
    .B2(_08874_),
    .ZN(_09271_));
 AOI21_X1 _18929_ (.A(_08690_),
    .B1(_08736_),
    .B2(_08663_),
    .ZN(_09272_));
 AND4_X1 _18930_ (.A1(_08584_),
    .A2(_08675_),
    .A3(_08683_),
    .A4(_08753_),
    .ZN(_09273_));
 OR4_X2 _18931_ (.A1(_09270_),
    .A2(_09271_),
    .A3(_09272_),
    .A4(_09273_),
    .ZN(_09274_));
 OAI21_X1 _18932_ (.A(_08694_),
    .B1(_08836_),
    .B2(_08724_),
    .ZN(_09275_));
 OAI21_X1 _18933_ (.A(_08694_),
    .B1(_08843_),
    .B2(_08785_),
    .ZN(_09276_));
 OAI21_X1 _18934_ (.A(_08694_),
    .B1(_08697_),
    .B2(_08631_),
    .ZN(_09277_));
 NAND3_X1 _18935_ (.A1(_09275_),
    .A2(_09276_),
    .A3(_09277_),
    .ZN(_09278_));
 OAI21_X1 _18936_ (.A(_08753_),
    .B1(_16780_),
    .B2(_08586_),
    .ZN(_09279_));
 INV_X1 _18937_ (.A(_09279_),
    .ZN(_09280_));
 OAI21_X1 _18938_ (.A(_08704_),
    .B1(_09239_),
    .B2(_09280_),
    .ZN(_09281_));
 OAI211_X2 _18939_ (.A(_09281_),
    .B(_08708_),
    .C1(_08873_),
    .C2(_08839_),
    .ZN(_09282_));
 OAI21_X1 _18940_ (.A(_08658_),
    .B1(_08686_),
    .B2(_08642_),
    .ZN(_09283_));
 OAI211_X2 _18941_ (.A(_08848_),
    .B(_09283_),
    .C1(_09227_),
    .C2(_08659_),
    .ZN(_09284_));
 NOR4_X1 _18942_ (.A1(_09274_),
    .A2(_09278_),
    .A3(_09282_),
    .A4(_09284_),
    .ZN(_09285_));
 NAND4_X1 _18943_ (.A1(_09233_),
    .A2(_09248_),
    .A3(_09269_),
    .A4(_09285_),
    .ZN(_09286_));
 NOR2_X2 _18944_ (.A1(_09286_),
    .A2(_08786_),
    .ZN(_09287_));
 XNOR2_X2 _18945_ (.A(_09213_),
    .B(_09287_),
    .ZN(_09288_));
 XNOR2_X1 _18946_ (.A(_09288_),
    .B(_08888_),
    .ZN(_09289_));
 AND2_X1 _18947_ (.A1(_09016_),
    .A2(_08898_),
    .ZN(_09290_));
 AND2_X1 _18948_ (.A1(_09016_),
    .A2(_09045_),
    .ZN(_09291_));
 OR2_X2 _18949_ (.A1(_09290_),
    .A2(_09291_),
    .ZN(_09292_));
 AND2_X1 _18950_ (.A1(_08895_),
    .A2(_09017_),
    .ZN(_09293_));
 AOI221_X1 _18951_ (.A(_09292_),
    .B1(_09293_),
    .B2(_09016_),
    .C1(_08957_),
    .C2(_09081_),
    .ZN(_09294_));
 NAND2_X1 _18952_ (.A1(_09084_),
    .A2(_08948_),
    .ZN(_09295_));
 AND2_X1 _18953_ (.A1(_08925_),
    .A2(_08907_),
    .ZN(_09296_));
 AND3_X1 _18954_ (.A1(_09296_),
    .A2(_08892_),
    .A3(_08891_),
    .ZN(_09297_));
 INV_X1 _18955_ (.A(_09297_),
    .ZN(_09298_));
 OAI21_X1 _18956_ (.A(_09295_),
    .B1(_09298_),
    .B2(_08908_),
    .ZN(_09299_));
 AOI221_X1 _18957_ (.A(_09299_),
    .B1(_09081_),
    .B2(_09018_),
    .C1(_09053_),
    .C2(_08955_),
    .ZN(_09300_));
 AND4_X1 _18958_ (.A1(_08997_),
    .A2(_09294_),
    .A3(_08996_),
    .A4(_09300_),
    .ZN(_09301_));
 INV_X1 _18959_ (.A(_08948_),
    .ZN(_09302_));
 INV_X1 _18960_ (.A(_08953_),
    .ZN(_09303_));
 OAI221_X1 _18961_ (.A(_09042_),
    .B1(_09302_),
    .B2(_09032_),
    .C1(_09303_),
    .C2(_09029_),
    .ZN(_09304_));
 BUF_X4 _18962_ (.A(_08947_),
    .Z(_09305_));
 AND2_X1 _18963_ (.A1(_08998_),
    .A2(_09305_),
    .ZN(_09306_));
 AND2_X1 _18964_ (.A1(_08987_),
    .A2(_09305_),
    .ZN(_09307_));
 NAND2_X1 _18965_ (.A1(_08993_),
    .A2(_08916_),
    .ZN(_09308_));
 INV_X1 _18966_ (.A(_09308_),
    .ZN(_09309_));
 BUF_X4 _18967_ (.A(_08953_),
    .Z(_09310_));
 AND3_X1 _18968_ (.A1(_09309_),
    .A2(_09310_),
    .A3(_08931_),
    .ZN(_09311_));
 NOR4_X1 _18969_ (.A1(_09304_),
    .A2(_09306_),
    .A3(_09307_),
    .A4(_09311_),
    .ZN(_09312_));
 NAND3_X1 _18970_ (.A1(_08934_),
    .A2(_08993_),
    .A3(_09305_),
    .ZN(_09313_));
 NAND2_X1 _18971_ (.A1(_09305_),
    .A2(_08926_),
    .ZN(_09314_));
 NAND2_X1 _18972_ (.A1(_09026_),
    .A2(_09305_),
    .ZN(_09315_));
 AND4_X1 _18973_ (.A1(_08938_),
    .A2(_09313_),
    .A3(_09314_),
    .A4(_09315_),
    .ZN(_09316_));
 AND2_X1 _18974_ (.A1(_08953_),
    .A2(_09293_),
    .ZN(_09317_));
 BUF_X2 _18975_ (.A(_09045_),
    .Z(_09318_));
 AND2_X1 _18976_ (.A1(_08953_),
    .A2(_09318_),
    .ZN(_09319_));
 NOR2_X1 _18977_ (.A1(_09317_),
    .A2(_09319_),
    .ZN(_09320_));
 AND2_X1 _18978_ (.A1(_09005_),
    .A2(_08966_),
    .ZN(_09321_));
 AND2_X1 _18979_ (.A1(_08991_),
    .A2(_08912_),
    .ZN(_09322_));
 NOR2_X1 _18980_ (.A1(_09308_),
    .A2(_09017_),
    .ZN(_09323_));
 AOI211_X4 _18981_ (.A(_09321_),
    .B(_09322_),
    .C1(_08991_),
    .C2(_09323_),
    .ZN(_09324_));
 AND2_X2 _18982_ (.A1(_08916_),
    .A2(_08929_),
    .ZN(_09325_));
 BUF_X2 _18983_ (.A(_08893_),
    .Z(_09326_));
 BUF_X2 _18984_ (.A(_08973_),
    .Z(_09327_));
 AOI22_X1 _18985_ (.A1(_09325_),
    .A2(_09326_),
    .B1(_09327_),
    .B2(_08998_),
    .ZN(_09328_));
 BUF_X4 _18986_ (.A(_08983_),
    .Z(_09329_));
 BUF_X2 _18987_ (.A(_09058_),
    .Z(_09330_));
 BUF_X4 _18988_ (.A(_08912_),
    .Z(_09331_));
 AOI22_X1 _18989_ (.A1(_09329_),
    .A2(_08924_),
    .B1(_09330_),
    .B2(_09331_),
    .ZN(_09332_));
 AND4_X1 _18990_ (.A1(_09320_),
    .A2(_09324_),
    .A3(_09328_),
    .A4(_09332_),
    .ZN(_09333_));
 NAND4_X1 _18991_ (.A1(_09301_),
    .A2(_09312_),
    .A3(_09316_),
    .A4(_09333_),
    .ZN(_09334_));
 AND2_X1 _18992_ (.A1(_08957_),
    .A2(_09074_),
    .ZN(_09335_));
 AND3_X1 _18993_ (.A1(_08934_),
    .A2(_08893_),
    .A3(_08993_),
    .ZN(_09336_));
 AND3_X1 _18994_ (.A1(_09318_),
    .A2(_08892_),
    .A3(_08905_),
    .ZN(_09337_));
 OR3_X1 _18995_ (.A1(_09335_),
    .A2(_09336_),
    .A3(_09337_),
    .ZN(_09338_));
 BUF_X2 _18996_ (.A(_09084_),
    .Z(_09339_));
 BUF_X4 _18997_ (.A(_08966_),
    .Z(_09340_));
 OAI21_X1 _18998_ (.A(_09339_),
    .B1(_08969_),
    .B2(_09340_),
    .ZN(_09341_));
 NAND3_X1 _18999_ (.A1(_08910_),
    .A2(_09057_),
    .A3(_08921_),
    .ZN(_09342_));
 AND2_X1 _19000_ (.A1(_09341_),
    .A2(_09342_),
    .ZN(_09343_));
 AND2_X2 _19001_ (.A1(_09087_),
    .A2(_08929_),
    .ZN(_09344_));
 OAI21_X1 _19002_ (.A(_09074_),
    .B1(_09344_),
    .B2(_09296_),
    .ZN(_09345_));
 BUF_X4 _19003_ (.A(_09041_),
    .Z(_09346_));
 NOR2_X1 _19004_ (.A1(_08933_),
    .A2(_08918_),
    .ZN(_09347_));
 OAI21_X1 _19005_ (.A(_09346_),
    .B1(_09347_),
    .B2(_09026_),
    .ZN(_09348_));
 INV_X2 _19006_ (.A(_09081_),
    .ZN(_09349_));
 NAND2_X1 _19007_ (.A1(_08959_),
    .A2(_08977_),
    .ZN(_09350_));
 NOR2_X2 _19008_ (.A1(_09349_),
    .A2(_09350_),
    .ZN(_09351_));
 INV_X1 _19009_ (.A(_09351_),
    .ZN(_09352_));
 NAND4_X1 _19010_ (.A1(_09343_),
    .A2(_09345_),
    .A3(_09348_),
    .A4(_09352_),
    .ZN(_09353_));
 BUF_X8 _19011_ (.A(_08906_),
    .Z(_09354_));
 BUF_X4 _19012_ (.A(_08916_),
    .Z(_09355_));
 OAI21_X1 _19013_ (.A(_09354_),
    .B1(_08937_),
    .B2(_09355_),
    .ZN(_09356_));
 INV_X1 _19014_ (.A(_09064_),
    .ZN(_09357_));
 OAI21_X1 _19015_ (.A(_09356_),
    .B1(_09357_),
    .B2(_08933_),
    .ZN(_09358_));
 NAND2_X1 _19016_ (.A1(_08931_),
    .A2(_08977_),
    .ZN(_09359_));
 NOR2_X1 _19017_ (.A1(_09008_),
    .A2(_09359_),
    .ZN(_09360_));
 INV_X1 _19018_ (.A(_09360_),
    .ZN(_09361_));
 OAI21_X1 _19019_ (.A(_09327_),
    .B1(_09344_),
    .B2(_08969_),
    .ZN(_09362_));
 NAND3_X1 _19020_ (.A1(_09327_),
    .A2(_08977_),
    .A3(_08956_),
    .ZN(_09363_));
 NOR3_X1 _19021_ (.A1(_08954_),
    .A2(_08894_),
    .A3(_16870_),
    .ZN(_09364_));
 NAND3_X1 _19022_ (.A1(_09364_),
    .A2(_08921_),
    .A3(_08905_),
    .ZN(_09365_));
 NAND4_X1 _19023_ (.A1(_09361_),
    .A2(_09362_),
    .A3(_09363_),
    .A4(_09365_),
    .ZN(_09366_));
 NOR4_X1 _19024_ (.A1(_09338_),
    .A2(_09353_),
    .A3(_09358_),
    .A4(_09366_),
    .ZN(_09367_));
 NAND2_X1 _19025_ (.A1(_08906_),
    .A2(_09079_),
    .ZN(_09368_));
 NAND2_X1 _19026_ (.A1(_09293_),
    .A2(_09005_),
    .ZN(_09369_));
 AND2_X1 _19027_ (.A1(_09368_),
    .A2(_09369_),
    .ZN(_09370_));
 INV_X1 _19028_ (.A(_08968_),
    .ZN(_09371_));
 INV_X1 _19029_ (.A(_09329_),
    .ZN(_09372_));
 OAI221_X1 _19030_ (.A(_09370_),
    .B1(_09008_),
    .B2(_09371_),
    .C1(_09302_),
    .C2(_09372_),
    .ZN(_09373_));
 BUF_X4 _19031_ (.A(_09069_),
    .Z(_09374_));
 AND2_X1 _19032_ (.A1(_08953_),
    .A2(_09374_),
    .ZN(_09375_));
 INV_X1 _19033_ (.A(_09375_),
    .ZN(_09376_));
 BUF_X4 _19034_ (.A(_09005_),
    .Z(_09377_));
 BUF_X2 _19035_ (.A(_08975_),
    .Z(_09378_));
 AOI22_X1 _19036_ (.A1(_09377_),
    .A2(_09378_),
    .B1(_08910_),
    .B2(_08947_),
    .ZN(_09379_));
 INV_X1 _19037_ (.A(_09018_),
    .ZN(_09380_));
 OAI211_X2 _19038_ (.A(_09376_),
    .B(_09379_),
    .C1(_08992_),
    .C2(_09380_),
    .ZN(_09381_));
 BUF_X4 _19039_ (.A(_09031_),
    .Z(_09382_));
 AND2_X1 _19040_ (.A1(_08984_),
    .A2(_09382_),
    .ZN(_09383_));
 NAND2_X1 _19041_ (.A1(_09079_),
    .A2(_09382_),
    .ZN(_09384_));
 INV_X2 _19042_ (.A(_09079_),
    .ZN(_09385_));
 INV_X1 _19043_ (.A(_09039_),
    .ZN(_09386_));
 OAI21_X1 _19044_ (.A(_09384_),
    .B1(_09385_),
    .B2(_09386_),
    .ZN(_09387_));
 NOR4_X1 _19045_ (.A1(_09373_),
    .A2(_09381_),
    .A3(_09383_),
    .A4(_09387_),
    .ZN(_09388_));
 OAI21_X1 _19046_ (.A(_08983_),
    .B1(_09079_),
    .B2(_09340_),
    .ZN(_09389_));
 NAND4_X1 _19047_ (.A1(_08905_),
    .A2(_08929_),
    .A3(_09087_),
    .A4(_08945_),
    .ZN(_09390_));
 NAND2_X1 _19048_ (.A1(_09389_),
    .A2(_09390_),
    .ZN(_09391_));
 BUF_X4 _19049_ (.A(_09016_),
    .Z(_09392_));
 OAI21_X1 _19050_ (.A(_09392_),
    .B1(_09072_),
    .B2(_08988_),
    .ZN(_09393_));
 BUF_X4 _19051_ (.A(_08939_),
    .Z(_09394_));
 NAND2_X1 _19052_ (.A1(_09392_),
    .A2(_09394_),
    .ZN(_09395_));
 NAND2_X1 _19053_ (.A1(_09393_),
    .A2(_09395_),
    .ZN(_09396_));
 BUF_X4 _19054_ (.A(_09382_),
    .Z(_09397_));
 NOR2_X1 _19055_ (.A1(_08900_),
    .A2(_16870_),
    .ZN(_09398_));
 AOI211_X2 _19056_ (.A(_09391_),
    .B(_09396_),
    .C1(_09397_),
    .C2(_09398_),
    .ZN(_09399_));
 INV_X1 _19057_ (.A(_09359_),
    .ZN(_09400_));
 NAND3_X1 _19058_ (.A1(_09400_),
    .A2(_08993_),
    .A3(_09330_),
    .ZN(_09401_));
 AND2_X1 _19059_ (.A1(_08966_),
    .A2(_09039_),
    .ZN(_09402_));
 AOI221_X1 _19060_ (.A(_09402_),
    .B1(_08964_),
    .B2(_09346_),
    .C1(_09053_),
    .C2(_09344_),
    .ZN(_09403_));
 BUF_X2 _19061_ (.A(_08901_),
    .Z(_09404_));
 BUF_X4 _19062_ (.A(_09346_),
    .Z(_09405_));
 NAND2_X1 _19063_ (.A1(_09404_),
    .A2(_09405_),
    .ZN(_09406_));
 OAI21_X1 _19064_ (.A(_08894_),
    .B1(_08931_),
    .B2(_16870_),
    .ZN(_09407_));
 AND3_X1 _19065_ (.A1(_08944_),
    .A2(_08945_),
    .A3(_08894_),
    .ZN(_09408_));
 AOI22_X1 _19066_ (.A1(_09407_),
    .A2(_09408_),
    .B1(_09404_),
    .B2(_09382_),
    .ZN(_09409_));
 AND4_X1 _19067_ (.A1(_09401_),
    .A2(_09403_),
    .A3(_09406_),
    .A4(_09409_),
    .ZN(_09410_));
 NAND4_X1 _19068_ (.A1(_09367_),
    .A2(_09388_),
    .A3(_09399_),
    .A4(_09410_),
    .ZN(_09411_));
 NOR2_X4 _19069_ (.A1(_09334_),
    .A2(_09411_),
    .ZN(_09412_));
 XOR2_X2 _19070_ (.A(_09412_),
    .B(_09093_),
    .Z(_09413_));
 NAND2_X1 _19071_ (.A1(_05918_),
    .A2(_06061_),
    .ZN(_09414_));
 NAND4_X1 _19072_ (.A1(_05907_),
    .A2(_05863_),
    .A3(_05500_),
    .A4(_04329_),
    .ZN(_09415_));
 AND2_X1 _19073_ (.A1(_09414_),
    .A2(_09415_),
    .ZN(_09416_));
 AND2_X4 _19074_ (.A1(_04395_),
    .A2(_04625_),
    .ZN(_09417_));
 AND2_X1 _19075_ (.A1(_09417_),
    .A2(_05929_),
    .ZN(_09418_));
 AND2_X1 _19076_ (.A1(_05152_),
    .A2(_05929_),
    .ZN(_09419_));
 AND4_X1 _19077_ (.A1(_05198_),
    .A2(_04592_),
    .A3(_05676_),
    .A4(_05467_),
    .ZN(_09420_));
 OR3_X2 _19078_ (.A1(_09418_),
    .A2(_09419_),
    .A3(_09420_),
    .ZN(_09421_));
 INV_X1 _19079_ (.A(_05214_),
    .ZN(_09422_));
 AND2_X1 _19080_ (.A1(_09422_),
    .A2(_05841_),
    .ZN(_09423_));
 AND2_X1 _19081_ (.A1(_05841_),
    .A2(_04297_),
    .ZN(_09424_));
 NOR2_X1 _19082_ (.A1(_09423_),
    .A2(_09424_),
    .ZN(_09425_));
 INV_X1 _19083_ (.A(_09425_),
    .ZN(_09426_));
 NAND4_X1 _19084_ (.A1(_05863_),
    .A2(_05753_),
    .A3(_05467_),
    .A4(_05500_),
    .ZN(_09427_));
 OAI21_X1 _19085_ (.A(_09427_),
    .B1(_05194_),
    .B2(_05962_),
    .ZN(_09428_));
 NAND2_X1 _19086_ (.A1(_06380_),
    .A2(_05841_),
    .ZN(_09429_));
 NAND2_X1 _19087_ (.A1(_05808_),
    .A2(_05709_),
    .ZN(_09430_));
 NAND2_X1 _19088_ (.A1(_05841_),
    .A2(_04549_),
    .ZN(_09431_));
 NAND3_X1 _19089_ (.A1(_09429_),
    .A2(_09430_),
    .A3(_09431_),
    .ZN(_09432_));
 NOR4_X1 _19090_ (.A1(_09421_),
    .A2(_09426_),
    .A3(_09428_),
    .A4(_09432_),
    .ZN(_09433_));
 AND2_X4 _19091_ (.A1(_04888_),
    .A2(_04669_),
    .ZN(_09434_));
 OAI21_X1 _19092_ (.A(_06061_),
    .B1(_09434_),
    .B2(_04976_),
    .ZN(_09435_));
 AND2_X2 _19093_ (.A1(_05775_),
    .A2(_09422_),
    .ZN(_09436_));
 NAND2_X2 _19094_ (.A1(_05775_),
    .A2(_05180_),
    .ZN(_09437_));
 BUF_X4 _19095_ (.A(_04165_),
    .Z(_09438_));
 NAND3_X1 _19096_ (.A1(_06391_),
    .A2(_09438_),
    .A3(_05676_),
    .ZN(_09439_));
 NAND2_X1 _19097_ (.A1(_09437_),
    .A2(_09439_),
    .ZN(_09440_));
 BUF_X4 _19098_ (.A(_04833_),
    .Z(_09441_));
 AOI211_X4 _19099_ (.A(_09436_),
    .B(_09440_),
    .C1(_09441_),
    .C2(_05775_),
    .ZN(_09442_));
 AND4_X1 _19100_ (.A1(_09416_),
    .A2(_09433_),
    .A3(_09435_),
    .A4(_09442_),
    .ZN(_09443_));
 BUF_X4 _19101_ (.A(_04428_),
    .Z(_09444_));
 NAND2_X1 _19102_ (.A1(_09444_),
    .A2(_04549_),
    .ZN(_09445_));
 AND2_X1 _19103_ (.A1(_04614_),
    .A2(_04691_),
    .ZN(_09446_));
 OAI21_X1 _19104_ (.A(_09444_),
    .B1(_05085_),
    .B2(_04921_),
    .ZN(_09447_));
 AND3_X1 _19105_ (.A1(_04428_),
    .A2(_05401_),
    .A3(_04647_),
    .ZN(_09448_));
 AND3_X1 _19106_ (.A1(_04428_),
    .A2(_05401_),
    .A3(_05907_),
    .ZN(_09449_));
 NOR3_X1 _19107_ (.A1(_04406_),
    .A2(_09448_),
    .A3(_09449_),
    .ZN(_09450_));
 AND4_X1 _19108_ (.A1(_09445_),
    .A2(_09446_),
    .A3(_09447_),
    .A4(_09450_),
    .ZN(_09451_));
 AND2_X1 _19109_ (.A1(_05401_),
    .A2(_04373_),
    .ZN(_09452_));
 AND2_X1 _19110_ (.A1(_04483_),
    .A2(_09452_),
    .ZN(_09453_));
 AND2_X4 _19111_ (.A1(_04592_),
    .A2(_04275_),
    .ZN(_09454_));
 AND2_X1 _19112_ (.A1(_04209_),
    .A2(_09454_),
    .ZN(_09455_));
 AND2_X1 _19113_ (.A1(_04209_),
    .A2(_05152_),
    .ZN(_09456_));
 AND2_X1 _19114_ (.A1(_04198_),
    .A2(_05302_),
    .ZN(_09457_));
 NOR4_X1 _19115_ (.A1(_09453_),
    .A2(_09455_),
    .A3(_09456_),
    .A4(_09457_),
    .ZN(_09458_));
 AND2_X1 _19116_ (.A1(_04516_),
    .A2(_04757_),
    .ZN(_09459_));
 AND2_X1 _19117_ (.A1(_06391_),
    .A2(_04757_),
    .ZN(_09460_));
 AND2_X1 _19118_ (.A1(_04757_),
    .A2(_05566_),
    .ZN(_09461_));
 AND3_X1 _19119_ (.A1(_05984_),
    .A2(_04187_),
    .A3(_04932_),
    .ZN(_09462_));
 NOR4_X1 _19120_ (.A1(_09459_),
    .A2(_09460_),
    .A3(_09461_),
    .A4(_09462_),
    .ZN(_09463_));
 BUF_X4 _19121_ (.A(_05009_),
    .Z(_09464_));
 NAND2_X1 _19122_ (.A1(_05037_),
    .A2(_09464_),
    .ZN(_09465_));
 OAI211_X2 _19123_ (.A(_05009_),
    .B(_06270_),
    .C1(_05511_),
    .C2(_05522_),
    .ZN(_09466_));
 OAI211_X2 _19124_ (.A(_05009_),
    .B(_04833_),
    .C1(_05511_),
    .C2(_05753_),
    .ZN(_09467_));
 BUF_X4 _19125_ (.A(_05401_),
    .Z(_09468_));
 NAND3_X1 _19126_ (.A1(_05009_),
    .A2(_05522_),
    .A3(_09468_),
    .ZN(_09469_));
 AND4_X1 _19127_ (.A1(_09465_),
    .A2(_09466_),
    .A3(_09467_),
    .A4(_09469_),
    .ZN(_09470_));
 AND4_X1 _19128_ (.A1(_09451_),
    .A2(_09458_),
    .A3(_09463_),
    .A4(_09470_),
    .ZN(_09471_));
 AND2_X1 _19129_ (.A1(_04581_),
    .A2(_04592_),
    .ZN(_09472_));
 BUF_X2 _19130_ (.A(_09472_),
    .Z(_09473_));
 AND2_X1 _19131_ (.A1(_09473_),
    .A2(_06303_),
    .ZN(_09474_));
 INV_X4 _19132_ (.A(_04965_),
    .ZN(_09475_));
 INV_X1 _19133_ (.A(_04844_),
    .ZN(_09476_));
 NAND2_X2 _19134_ (.A1(_09475_),
    .A2(_09476_),
    .ZN(_09477_));
 AND2_X2 _19135_ (.A1(_09477_),
    .A2(_06303_),
    .ZN(_09478_));
 AND2_X1 _19136_ (.A1(_09422_),
    .A2(_06215_),
    .ZN(_09479_));
 AND2_X1 _19137_ (.A1(_05047_),
    .A2(_06215_),
    .ZN(_09480_));
 OR4_X2 _19138_ (.A1(_09474_),
    .A2(_09478_),
    .A3(_09479_),
    .A4(_09480_),
    .ZN(_09481_));
 BUF_X2 _19139_ (.A(_06138_),
    .Z(_09482_));
 OAI21_X1 _19140_ (.A(_09482_),
    .B1(_06248_),
    .B2(_05412_),
    .ZN(_09483_));
 NAND2_X1 _19141_ (.A1(_04855_),
    .A2(_09482_),
    .ZN(_09484_));
 AND2_X2 _19142_ (.A1(_05456_),
    .A2(_06149_),
    .ZN(_09485_));
 INV_X1 _19143_ (.A(_09485_),
    .ZN(_09486_));
 AND2_X1 _19144_ (.A1(_04921_),
    .A2(_09482_),
    .ZN(_09487_));
 INV_X1 _19145_ (.A(_09487_),
    .ZN(_09488_));
 NAND4_X1 _19146_ (.A1(_09483_),
    .A2(_09484_),
    .A3(_09486_),
    .A4(_09488_),
    .ZN(_09489_));
 NAND2_X1 _19147_ (.A1(_06347_),
    .A2(_09472_),
    .ZN(_09490_));
 BUF_X4 _19148_ (.A(_06347_),
    .Z(_09491_));
 NAND2_X1 _19149_ (.A1(_09491_),
    .A2(_04976_),
    .ZN(_09492_));
 NAND2_X1 _19150_ (.A1(_09491_),
    .A2(_04855_),
    .ZN(_09493_));
 AND3_X1 _19151_ (.A1(_09490_),
    .A2(_09492_),
    .A3(_09493_),
    .ZN(_09494_));
 OAI21_X1 _19152_ (.A(_09491_),
    .B1(_06380_),
    .B2(_04417_),
    .ZN(_09495_));
 INV_X1 _19153_ (.A(_05200_),
    .ZN(_09496_));
 OAI211_X2 _19154_ (.A(_09494_),
    .B(_09495_),
    .C1(_09496_),
    .C2(_06358_),
    .ZN(_09497_));
 AND2_X1 _19155_ (.A1(_05170_),
    .A2(_06424_),
    .ZN(_09498_));
 INV_X1 _19156_ (.A(_09498_),
    .ZN(_09499_));
 OAI21_X1 _19157_ (.A(_06446_),
    .B1(_05456_),
    .B2(_04921_),
    .ZN(_09500_));
 INV_X1 _19158_ (.A(_06446_),
    .ZN(_09501_));
 OAI211_X2 _19159_ (.A(_09499_),
    .B(_09500_),
    .C1(_05194_),
    .C2(_09501_),
    .ZN(_09502_));
 NOR4_X2 _19160_ (.A1(_09481_),
    .A2(_09489_),
    .A3(_09497_),
    .A4(_09502_),
    .ZN(_09503_));
 NAND2_X1 _19161_ (.A1(_04516_),
    .A2(_05357_),
    .ZN(_09504_));
 BUF_X8 _19162_ (.A(_09454_),
    .Z(_09505_));
 OAI21_X1 _19163_ (.A(_05247_),
    .B1(_09422_),
    .B2(_09505_),
    .ZN(_09506_));
 BUF_X8 _19164_ (.A(_09417_),
    .Z(_09507_));
 OAI21_X1 _19165_ (.A(_05247_),
    .B1(_09507_),
    .B2(_05152_),
    .ZN(_09508_));
 NAND4_X1 _19166_ (.A1(_05202_),
    .A2(_05522_),
    .A3(_05500_),
    .A4(_04329_),
    .ZN(_09509_));
 AND4_X1 _19167_ (.A1(_09504_),
    .A2(_09506_),
    .A3(_09508_),
    .A4(_09509_),
    .ZN(_09510_));
 AND2_X1 _19168_ (.A1(_05390_),
    .A2(_04658_),
    .ZN(_09511_));
 INV_X1 _19169_ (.A(_05390_),
    .ZN(_09512_));
 AOI21_X1 _19170_ (.A(_09512_),
    .B1(_09496_),
    .B2(_05346_),
    .ZN(_09513_));
 AOI211_X4 _19171_ (.A(_09511_),
    .B(_09513_),
    .C1(_05489_),
    .C2(_09434_),
    .ZN(_09514_));
 INV_X1 _19172_ (.A(_05555_),
    .ZN(_09515_));
 INV_X1 _19173_ (.A(_05188_),
    .ZN(_09516_));
 AOI21_X1 _19174_ (.A(_09515_),
    .B1(_09516_),
    .B2(_05995_),
    .ZN(_09517_));
 AOI21_X1 _19175_ (.A(_09515_),
    .B1(_09476_),
    .B2(_09475_),
    .ZN(_09518_));
 AND2_X1 _19176_ (.A1(_05555_),
    .A2(_09422_),
    .ZN(_09519_));
 AND2_X1 _19177_ (.A1(_05599_),
    .A2(_09473_),
    .ZN(_09520_));
 NOR4_X1 _19178_ (.A1(_09517_),
    .A2(_09518_),
    .A3(_09519_),
    .A4(_09520_),
    .ZN(_09521_));
 AND2_X1 _19179_ (.A1(_05037_),
    .A2(_05143_),
    .ZN(_09522_));
 AND4_X1 _19180_ (.A1(_05753_),
    .A2(_05202_),
    .A3(_05401_),
    .A4(_04932_),
    .ZN(_09523_));
 AND4_X1 _19181_ (.A1(_04275_),
    .A2(_05202_),
    .A3(_05269_),
    .A4(_04932_),
    .ZN(_09524_));
 NOR4_X1 _19182_ (.A1(_09522_),
    .A2(_05161_),
    .A3(_09523_),
    .A4(_09524_),
    .ZN(_09525_));
 AND4_X1 _19183_ (.A1(_09510_),
    .A2(_09514_),
    .A3(_09521_),
    .A4(_09525_),
    .ZN(_09526_));
 NAND4_X1 _19184_ (.A1(_09443_),
    .A2(_09471_),
    .A3(_09503_),
    .A4(_09526_),
    .ZN(_09527_));
 NOR2_X2 _19185_ (.A1(_09527_),
    .A2(_06556_),
    .ZN(_09528_));
 XNOR2_X1 _19186_ (.A(_09413_),
    .B(_09528_),
    .ZN(_09529_));
 XNOR2_X1 _19187_ (.A(_09289_),
    .B(_09529_),
    .ZN(_09530_));
 INV_X2 _19188_ (.A(_17155_),
    .ZN(_09531_));
 BUF_X8 _19189_ (.A(_09531_),
    .Z(_09532_));
 XNOR2_X1 _19190_ (.A(_09530_),
    .B(_09532_),
    .ZN(_09533_));
 MUX2_X1 _19191_ (.A(_09102_),
    .B(_09533_),
    .S(_09100_),
    .Z(_00725_));
 XOR2_X1 _19192_ (.A(_17166_),
    .B(_17062_),
    .Z(_09534_));
 NAND3_X1 _19193_ (.A1(_07392_),
    .A2(_07949_),
    .A3(_06842_),
    .ZN(_09535_));
 OAI211_X2 _19194_ (.A(_09172_),
    .B(_09535_),
    .C1(_08551_),
    .C2(_08433_),
    .ZN(_09536_));
 NAND2_X1 _19195_ (.A1(_08550_),
    .A2(_09166_),
    .ZN(_09537_));
 INV_X1 _19196_ (.A(_07205_),
    .ZN(_09538_));
 OAI21_X1 _19197_ (.A(_09537_),
    .B1(_08551_),
    .B2(_09538_),
    .ZN(_09539_));
 AND4_X1 _19198_ (.A1(_07949_),
    .A2(_09153_),
    .A3(_06842_),
    .A4(_07730_),
    .ZN(_09540_));
 NOR3_X1 _19199_ (.A1(_09536_),
    .A2(_09539_),
    .A3(_09540_),
    .ZN(_09541_));
 OAI21_X1 _19200_ (.A(_09202_),
    .B1(_07488_),
    .B2(_07370_),
    .ZN(_09542_));
 AOI21_X2 _19201_ (.A(_07488_),
    .B1(_08472_),
    .B2(_09161_),
    .ZN(_09543_));
 NAND2_X1 _19202_ (.A1(_06710_),
    .A2(_06754_),
    .ZN(_09544_));
 INV_X2 _19203_ (.A(_06710_),
    .ZN(_09545_));
 OAI211_X2 _19204_ (.A(_08528_),
    .B(_09544_),
    .C1(_08146_),
    .C2(_09545_),
    .ZN(_09546_));
 NAND3_X1 _19205_ (.A1(_09137_),
    .A2(_07304_),
    .A3(_08519_),
    .ZN(_09547_));
 NAND4_X1 _19206_ (.A1(_07304_),
    .A2(_07018_),
    .A3(_07740_),
    .A4(_06699_),
    .ZN(_09548_));
 AND2_X1 _19207_ (.A1(_07183_),
    .A2(_06732_),
    .ZN(_09549_));
 INV_X1 _19208_ (.A(_09549_),
    .ZN(_09550_));
 OAI211_X2 _19209_ (.A(_09547_),
    .B(_09548_),
    .C1(_09545_),
    .C2(_09550_),
    .ZN(_09551_));
 OR4_X2 _19210_ (.A1(_09542_),
    .A2(_09543_),
    .A3(_09546_),
    .A4(_09551_),
    .ZN(_09552_));
 AND3_X1 _19211_ (.A1(_09138_),
    .A2(_07960_),
    .A3(_06578_),
    .ZN(_09553_));
 AND2_X1 _19212_ (.A1(_07315_),
    .A2(_09105_),
    .ZN(_09554_));
 AND2_X2 _19213_ (.A1(_07315_),
    .A2(_07227_),
    .ZN(_09555_));
 OR3_X1 _19214_ (.A1(_09553_),
    .A2(_09554_),
    .A3(_09555_),
    .ZN(_09556_));
 NAND2_X1 _19215_ (.A1(_07315_),
    .A2(_08310_),
    .ZN(_09557_));
 NAND4_X1 _19216_ (.A1(_07960_),
    .A2(_08396_),
    .A3(_06633_),
    .A4(_08080_),
    .ZN(_09558_));
 OAI211_X2 _19217_ (.A(_09557_),
    .B(_09558_),
    .C1(_09187_),
    .C2(_07282_),
    .ZN(_09559_));
 AND2_X1 _19218_ (.A1(_09191_),
    .A2(_07216_),
    .ZN(_09560_));
 AND2_X1 _19219_ (.A1(_09191_),
    .A2(_06655_),
    .ZN(_09561_));
 AND3_X4 _19220_ (.A1(_07828_),
    .A2(_07883_),
    .A3(_07304_),
    .ZN(_09562_));
 OR4_X2 _19221_ (.A1(_09560_),
    .A2(_09197_),
    .A3(_09561_),
    .A4(_09562_),
    .ZN(_09563_));
 NOR4_X2 _19222_ (.A1(_09552_),
    .A2(_09556_),
    .A3(_09559_),
    .A4(_09563_),
    .ZN(_09564_));
 OAI21_X1 _19223_ (.A(_07414_),
    .B1(_08343_),
    .B2(_09131_),
    .ZN(_09565_));
 NAND2_X1 _19224_ (.A1(_09106_),
    .A2(_07414_),
    .ZN(_09566_));
 INV_X1 _19225_ (.A(_08354_),
    .ZN(_09567_));
 OAI211_X2 _19226_ (.A(_09565_),
    .B(_09566_),
    .C1(_09163_),
    .C2(_09567_),
    .ZN(_09568_));
 AND2_X1 _19227_ (.A1(_07359_),
    .A2(_08299_),
    .ZN(_09569_));
 AND3_X1 _19228_ (.A1(_06853_),
    .A2(_07730_),
    .A3(_09153_),
    .ZN(_09570_));
 INV_X1 _19229_ (.A(_07458_),
    .ZN(_09571_));
 INV_X1 _19230_ (.A(_07227_),
    .ZN(_09572_));
 AOI21_X1 _19231_ (.A(_07150_),
    .B1(_09571_),
    .B2(_09572_),
    .ZN(_09573_));
 NOR4_X1 _19232_ (.A1(_09568_),
    .A2(_09569_),
    .A3(_09570_),
    .A4(_09573_),
    .ZN(_09574_));
 OAI211_X2 _19233_ (.A(_07117_),
    .B(_08047_),
    .C1(_06644_),
    .C2(_08069_),
    .ZN(_09575_));
 NAND2_X1 _19234_ (.A1(_09125_),
    .A2(_07106_),
    .ZN(_09576_));
 OAI21_X1 _19235_ (.A(_07117_),
    .B1(_06655_),
    .B2(_07062_),
    .ZN(_09577_));
 AND3_X1 _19236_ (.A1(_09575_),
    .A2(_09576_),
    .A3(_09577_),
    .ZN(_09578_));
 AND4_X2 _19237_ (.A1(_09541_),
    .A2(_09564_),
    .A3(_09574_),
    .A4(_09578_),
    .ZN(_09579_));
 AOI21_X1 _19238_ (.A(_07992_),
    .B1(_08135_),
    .B2(_08321_),
    .ZN(_09580_));
 AOI211_X4 _19239_ (.A(_09143_),
    .B(_09580_),
    .C1(_08190_),
    .C2(_08354_),
    .ZN(_09581_));
 INV_X1 _19240_ (.A(_09125_),
    .ZN(_09582_));
 AOI21_X1 _19241_ (.A(_08542_),
    .B1(_09582_),
    .B2(_08541_),
    .ZN(_09583_));
 INV_X1 _19242_ (.A(_08556_),
    .ZN(_09584_));
 INV_X1 _19243_ (.A(_07392_),
    .ZN(_09585_));
 AOI21_X1 _19244_ (.A(_08542_),
    .B1(_09584_),
    .B2(_09585_),
    .ZN(_09586_));
 AOI211_X4 _19245_ (.A(_09583_),
    .B(_09586_),
    .C1(_06952_),
    .C2(_07861_),
    .ZN(_09587_));
 OAI21_X1 _19246_ (.A(_07795_),
    .B1(_08124_),
    .B2(_07631_),
    .ZN(_09588_));
 OAI21_X1 _19247_ (.A(_07795_),
    .B1(_09142_),
    .B2(_09166_),
    .ZN(_09589_));
 AND2_X1 _19248_ (.A1(_09588_),
    .A2(_09589_),
    .ZN(_09590_));
 AND2_X1 _19249_ (.A1(_07521_),
    .A2(_08310_),
    .ZN(_09591_));
 INV_X1 _19250_ (.A(_09591_),
    .ZN(_09592_));
 NAND2_X1 _19251_ (.A1(_09125_),
    .A2(_07521_),
    .ZN(_09593_));
 NAND2_X1 _19252_ (.A1(_09138_),
    .A2(_07532_),
    .ZN(_09594_));
 AND4_X1 _19253_ (.A1(_09592_),
    .A2(_08557_),
    .A3(_09593_),
    .A4(_09594_),
    .ZN(_09595_));
 NAND4_X1 _19254_ (.A1(_09581_),
    .A2(_09587_),
    .A3(_09590_),
    .A4(_09595_),
    .ZN(_09596_));
 OAI21_X1 _19255_ (.A(_07653_),
    .B1(_07686_),
    .B2(_08354_),
    .ZN(_09597_));
 NAND4_X1 _19256_ (.A1(_08519_),
    .A2(_08538_),
    .A3(_07238_),
    .A4(_08396_),
    .ZN(_09598_));
 NAND4_X1 _19257_ (.A1(_07653_),
    .A2(_07062_),
    .A3(_07730_),
    .A4(_08244_),
    .ZN(_09599_));
 NAND3_X1 _19258_ (.A1(_09597_),
    .A2(_09598_),
    .A3(_09599_),
    .ZN(_09600_));
 NAND2_X1 _19259_ (.A1(_09144_),
    .A2(_06611_),
    .ZN(_09601_));
 NAND4_X1 _19260_ (.A1(_07018_),
    .A2(_07740_),
    .A3(_08080_),
    .A4(_07238_),
    .ZN(_09602_));
 NAND2_X1 _19261_ (.A1(_09601_),
    .A2(_09602_),
    .ZN(_09603_));
 OAI21_X1 _19262_ (.A(_07894_),
    .B1(_09138_),
    .B2(_07828_),
    .ZN(_09604_));
 OAI21_X1 _19263_ (.A(_09604_),
    .B1(_09572_),
    .B2(_08443_),
    .ZN(_09605_));
 AOI21_X1 _19264_ (.A(_08443_),
    .B1(_08321_),
    .B2(_08146_),
    .ZN(_09606_));
 NAND2_X1 _19265_ (.A1(_08532_),
    .A2(_06600_),
    .ZN(_09607_));
 OAI22_X1 _19266_ (.A1(_09607_),
    .A2(_07436_),
    .B1(_07370_),
    .B2(_07348_),
    .ZN(_09608_));
 OR4_X2 _19267_ (.A1(_09603_),
    .A2(_09605_),
    .A3(_09606_),
    .A4(_09608_),
    .ZN(_09609_));
 OAI21_X1 _19268_ (.A(_07719_),
    .B1(_07359_),
    .B2(_09131_),
    .ZN(_09610_));
 OAI211_X2 _19269_ (.A(_07719_),
    .B(_08047_),
    .C1(_08396_),
    .C2(_07029_),
    .ZN(_09611_));
 NAND2_X1 _19270_ (.A1(_07719_),
    .A2(_08222_),
    .ZN(_09612_));
 NAND4_X1 _19271_ (.A1(_06820_),
    .A2(_07436_),
    .A3(_07447_),
    .A4(_07238_),
    .ZN(_09613_));
 NAND4_X1 _19272_ (.A1(_09610_),
    .A2(_09611_),
    .A3(_09612_),
    .A4(_09613_),
    .ZN(_09614_));
 NOR4_X4 _19273_ (.A1(_09596_),
    .A2(_09600_),
    .A3(_09609_),
    .A4(_09614_),
    .ZN(_09615_));
 NAND2_X4 _19274_ (.A1(_09579_),
    .A2(_09615_),
    .ZN(_09616_));
 OAI21_X1 _19275_ (.A(_08715_),
    .B1(_08573_),
    .B2(_08798_),
    .ZN(_09617_));
 AND2_X1 _19276_ (.A1(_08740_),
    .A2(_08577_),
    .ZN(_09618_));
 OAI21_X1 _19277_ (.A(_09230_),
    .B1(_09231_),
    .B2(_08661_),
    .ZN(_09619_));
 AOI211_X2 _19278_ (.A(_09618_),
    .B(_09619_),
    .C1(_08741_),
    .C2(_08680_),
    .ZN(_09620_));
 OAI21_X1 _19279_ (.A(_08714_),
    .B1(_08669_),
    .B2(_08673_),
    .ZN(_09621_));
 OAI211_X2 _19280_ (.A(_08715_),
    .B(_16783_),
    .C1(_08706_),
    .C2(_08568_),
    .ZN(_09622_));
 AND4_X1 _19281_ (.A1(_09617_),
    .A2(_09620_),
    .A3(_09621_),
    .A4(_09622_),
    .ZN(_09623_));
 OAI21_X1 _19282_ (.A(_08721_),
    .B1(_08749_),
    .B2(_08573_),
    .ZN(_09624_));
 AND2_X1 _19283_ (.A1(_08730_),
    .A2(_08732_),
    .ZN(_09625_));
 AND2_X1 _19284_ (.A1(_08730_),
    .A2(_08809_),
    .ZN(_09626_));
 AOI211_X2 _19285_ (.A(_09625_),
    .B(_09626_),
    .C1(_08767_),
    .C2(_08730_),
    .ZN(_09627_));
 OAI21_X1 _19286_ (.A(_08721_),
    .B1(_08596_),
    .B2(_08836_),
    .ZN(_09628_));
 AND4_X1 _19287_ (.A1(_08581_),
    .A2(_08713_),
    .A3(_08613_),
    .A4(_08638_),
    .ZN(_09629_));
 AND3_X1 _19288_ (.A1(_08723_),
    .A2(_08713_),
    .A3(_08638_),
    .ZN(_09630_));
 AOI211_X4 _19289_ (.A(_09629_),
    .B(_09630_),
    .C1(_08731_),
    .C2(_08790_),
    .ZN(_09631_));
 AND4_X1 _19290_ (.A1(_09624_),
    .A2(_09627_),
    .A3(_09628_),
    .A4(_09631_),
    .ZN(_09632_));
 BUF_X4 _19291_ (.A(_08766_),
    .Z(_09633_));
 OAI21_X1 _19292_ (.A(_09633_),
    .B1(_08815_),
    .B2(_08800_),
    .ZN(_09634_));
 OAI21_X1 _19293_ (.A(_08788_),
    .B1(_08779_),
    .B2(_08770_),
    .ZN(_09635_));
 OAI21_X1 _19294_ (.A(_08788_),
    .B1(_08822_),
    .B2(_08798_),
    .ZN(_09636_));
 AND4_X1 _19295_ (.A1(_08793_),
    .A2(_09634_),
    .A3(_09635_),
    .A4(_09636_),
    .ZN(_09637_));
 AOI21_X2 _19296_ (.A(_08757_),
    .B1(_08840_),
    .B2(_08873_),
    .ZN(_09638_));
 OR2_X4 _19297_ (.A1(_09638_),
    .A2(_08805_),
    .ZN(_09639_));
 AND2_X1 _19298_ (.A1(_08756_),
    .A2(_08578_),
    .ZN(_09640_));
 INV_X1 _19299_ (.A(_08573_),
    .ZN(_09641_));
 AOI21_X1 _19300_ (.A(_08757_),
    .B1(_09641_),
    .B2(_09234_),
    .ZN(_09642_));
 OAI21_X1 _19301_ (.A(_08747_),
    .B1(_08860_),
    .B2(_08578_),
    .ZN(_09643_));
 NAND3_X1 _19302_ (.A1(_08628_),
    .A2(_08747_),
    .A3(_08595_),
    .ZN(_09644_));
 OAI21_X1 _19303_ (.A(_08747_),
    .B1(_08631_),
    .B2(_08632_),
    .ZN(_09645_));
 NAND2_X1 _19304_ (.A1(_08747_),
    .A2(_08573_),
    .ZN(_09646_));
 NAND4_X1 _19305_ (.A1(_09643_),
    .A2(_09644_),
    .A3(_09645_),
    .A4(_09646_),
    .ZN(_09647_));
 NOR4_X1 _19306_ (.A1(_09639_),
    .A2(_09640_),
    .A3(_09642_),
    .A4(_09647_),
    .ZN(_09648_));
 NAND4_X1 _19307_ (.A1(_09623_),
    .A2(_09632_),
    .A3(_09637_),
    .A4(_09648_),
    .ZN(_09649_));
 INV_X1 _19308_ (.A(_08621_),
    .ZN(_09650_));
 AOI21_X1 _19309_ (.A(_09650_),
    .B1(_09641_),
    .B2(_09234_),
    .ZN(_09651_));
 NAND2_X1 _19310_ (.A1(_08621_),
    .A2(_08724_),
    .ZN(_09652_));
 OAI21_X1 _19311_ (.A(_09652_),
    .B1(_09650_),
    .B2(_09261_),
    .ZN(_09653_));
 AND2_X1 _19312_ (.A1(_08621_),
    .A2(_08697_),
    .ZN(_09654_));
 AND2_X2 _19313_ (.A1(_08621_),
    .A2(_08763_),
    .ZN(_09655_));
 NOR4_X2 _19314_ (.A1(_09651_),
    .A2(_09653_),
    .A3(_09654_),
    .A4(_09655_),
    .ZN(_09656_));
 AND2_X1 _19315_ (.A1(_08606_),
    .A2(_08595_),
    .ZN(_09657_));
 OAI21_X1 _19316_ (.A(_08645_),
    .B1(_09657_),
    .B2(_08674_),
    .ZN(_09658_));
 NAND4_X1 _19317_ (.A1(_08646_),
    .A2(_08650_),
    .A3(_08585_),
    .A4(_08599_),
    .ZN(_09659_));
 AND4_X2 _19318_ (.A1(_08652_),
    .A2(_09656_),
    .A3(_09658_),
    .A4(_09659_),
    .ZN(_09660_));
 NAND3_X1 _19319_ (.A1(_08681_),
    .A2(_08599_),
    .A3(_08602_),
    .ZN(_09661_));
 NAND2_X1 _19320_ (.A1(_08800_),
    .A2(_08565_),
    .ZN(_09662_));
 NAND4_X1 _19321_ (.A1(_08582_),
    .A2(_08648_),
    .A3(_08599_),
    .A4(_08563_),
    .ZN(_09663_));
 AND2_X1 _19322_ (.A1(_09662_),
    .A2(_09663_),
    .ZN(_09664_));
 INV_X1 _19323_ (.A(_09664_),
    .ZN(_09665_));
 AND3_X1 _19324_ (.A1(_08624_),
    .A2(_08565_),
    .A3(_08604_),
    .ZN(_09666_));
 NOR3_X1 _19325_ (.A1(_09665_),
    .A2(_08574_),
    .A3(_09666_),
    .ZN(_09667_));
 OAI21_X1 _19326_ (.A(_08608_),
    .B1(_08810_),
    .B2(_08669_),
    .ZN(_09668_));
 OAI211_X2 _19327_ (.A(_08608_),
    .B(_08583_),
    .C1(_08585_),
    .C2(_08706_),
    .ZN(_09669_));
 AND4_X1 _19328_ (.A1(_09661_),
    .A2(_09667_),
    .A3(_09668_),
    .A4(_09669_),
    .ZN(_09670_));
 NAND2_X1 _19329_ (.A1(_08704_),
    .A2(_08860_),
    .ZN(_09671_));
 INV_X1 _19330_ (.A(_08844_),
    .ZN(_09672_));
 OAI211_X2 _19331_ (.A(_09671_),
    .B(_09672_),
    .C1(_08839_),
    .C2(_08795_),
    .ZN(_09673_));
 AOI21_X1 _19332_ (.A(_08839_),
    .B1(_08616_),
    .B2(_08597_),
    .ZN(_09674_));
 NAND2_X1 _19333_ (.A1(_08672_),
    .A2(_08670_),
    .ZN(_09675_));
 AOI21_X1 _19334_ (.A(_08659_),
    .B1(_08736_),
    .B2(_08874_),
    .ZN(_09676_));
 NOR4_X1 _19335_ (.A1(_09673_),
    .A2(_09674_),
    .A3(_09675_),
    .A4(_09676_),
    .ZN(_09677_));
 OAI21_X1 _19336_ (.A(_08679_),
    .B1(_08749_),
    .B2(_08637_),
    .ZN(_09678_));
 OAI21_X1 _19337_ (.A(_08679_),
    .B1(_08836_),
    .B2(_08633_),
    .ZN(_09679_));
 OAI21_X1 _19338_ (.A(_08694_),
    .B1(_08749_),
    .B2(_08669_),
    .ZN(_09680_));
 OAI21_X1 _19339_ (.A(_08693_),
    .B1(_08836_),
    .B2(_08770_),
    .ZN(_09681_));
 AND4_X1 _19340_ (.A1(_09678_),
    .A2(_09679_),
    .A3(_09680_),
    .A4(_09681_),
    .ZN(_09682_));
 NAND4_X2 _19341_ (.A1(_09660_),
    .A2(_09670_),
    .A3(_09677_),
    .A4(_09682_),
    .ZN(_09683_));
 NOR2_X2 _19342_ (.A1(_09649_),
    .A2(_09683_),
    .ZN(_09684_));
 XNOR2_X2 _19343_ (.A(_09616_),
    .B(_09684_),
    .ZN(_09685_));
 OAI221_X1 _19344_ (.A(_05190_),
    .B1(_05192_),
    .B2(_05720_),
    .C1(_05753_),
    .C2(_05184_),
    .ZN(_09686_));
 AND2_X1 _19345_ (.A1(_05143_),
    .A2(_09417_),
    .ZN(_09687_));
 OR2_X4 _19346_ (.A1(_05161_),
    .A2(_09687_),
    .ZN(_09688_));
 OR2_X2 _19347_ (.A1(_04297_),
    .A2(_04253_),
    .ZN(_09689_));
 AND2_X1 _19348_ (.A1(_09689_),
    .A2(_05143_),
    .ZN(_09690_));
 NOR3_X2 _19349_ (.A1(_09686_),
    .A2(_09688_),
    .A3(_09690_),
    .ZN(_09691_));
 BUF_X4 _19350_ (.A(_05566_),
    .Z(_09692_));
 NAND2_X1 _19351_ (.A1(_05489_),
    .A2(_09692_),
    .ZN(_09693_));
 OAI21_X1 _19352_ (.A(_05489_),
    .B1(_09422_),
    .B2(_09507_),
    .ZN(_09694_));
 AND4_X1 _19353_ (.A1(_05434_),
    .A2(_09691_),
    .A3(_09693_),
    .A4(_09694_),
    .ZN(_09695_));
 OAI21_X1 _19354_ (.A(_05357_),
    .B1(_06380_),
    .B2(_06391_),
    .ZN(_09696_));
 OAI21_X1 _19355_ (.A(_05599_),
    .B1(_06380_),
    .B2(_05566_),
    .ZN(_09697_));
 OAI21_X1 _19356_ (.A(_05599_),
    .B1(_09473_),
    .B2(_06314_),
    .ZN(_09698_));
 OAI21_X1 _19357_ (.A(_05247_),
    .B1(_09473_),
    .B2(_04921_),
    .ZN(_09699_));
 AND4_X1 _19358_ (.A1(_09696_),
    .A2(_09697_),
    .A3(_09698_),
    .A4(_09699_),
    .ZN(_09700_));
 NOR2_X1 _19359_ (.A1(_04636_),
    .A2(_04581_),
    .ZN(_09701_));
 AND2_X1 _19360_ (.A1(_09701_),
    .A2(_04428_),
    .ZN(_09702_));
 OR2_X1 _19361_ (.A1(_09702_),
    .A2(_04603_),
    .ZN(_09703_));
 OAI21_X1 _19362_ (.A(_04209_),
    .B1(_05056_),
    .B2(_05566_),
    .ZN(_09704_));
 NAND2_X1 _19363_ (.A1(_04209_),
    .A2(_05085_),
    .ZN(_09705_));
 NAND2_X1 _19364_ (.A1(_04209_),
    .A2(_09422_),
    .ZN(_09706_));
 NAND4_X1 _19365_ (.A1(_09704_),
    .A2(_09705_),
    .A3(_09706_),
    .A4(_04308_),
    .ZN(_09707_));
 AND3_X1 _19366_ (.A1(_04801_),
    .A2(_04527_),
    .A3(_09444_),
    .ZN(_09708_));
 NOR4_X1 _19367_ (.A1(_09703_),
    .A2(_09707_),
    .A3(_04439_),
    .A4(_09708_),
    .ZN(_09709_));
 OAI21_X1 _19368_ (.A(_09464_),
    .B1(_04538_),
    .B2(_05313_),
    .ZN(_09710_));
 OAI211_X2 _19369_ (.A(_04757_),
    .B(_05269_),
    .C1(_05511_),
    .C2(_05753_),
    .ZN(_09711_));
 NAND4_X1 _19370_ (.A1(_04932_),
    .A2(_04494_),
    .A3(_04833_),
    .A4(_04187_),
    .ZN(_09712_));
 AND2_X1 _19371_ (.A1(_09711_),
    .A2(_09712_),
    .ZN(_09713_));
 OAI21_X1 _19372_ (.A(_09464_),
    .B1(_04253_),
    .B2(_06314_),
    .ZN(_09714_));
 NAND2_X1 _19373_ (.A1(_04757_),
    .A2(_05180_),
    .ZN(_09715_));
 NAND2_X1 _19374_ (.A1(_04757_),
    .A2(_04417_),
    .ZN(_09716_));
 NOR2_X1 _19375_ (.A1(_04790_),
    .A2(_05907_),
    .ZN(_09717_));
 NAND2_X1 _19376_ (.A1(_04746_),
    .A2(_09717_),
    .ZN(_09718_));
 AND3_X1 _19377_ (.A1(_09715_),
    .A2(_09716_),
    .A3(_09718_),
    .ZN(_09719_));
 AND4_X1 _19378_ (.A1(_09710_),
    .A2(_09713_),
    .A3(_09714_),
    .A4(_09719_),
    .ZN(_09720_));
 NAND4_X4 _19379_ (.A1(_09695_),
    .A2(_09700_),
    .A3(_09709_),
    .A4(_09720_),
    .ZN(_09721_));
 NAND2_X1 _19380_ (.A1(_06050_),
    .A2(_09717_),
    .ZN(_09722_));
 AND2_X1 _19381_ (.A1(_05775_),
    .A2(_05085_),
    .ZN(_09723_));
 AND3_X1 _19382_ (.A1(_04297_),
    .A2(_04165_),
    .A3(_05676_),
    .ZN(_09724_));
 NOR4_X1 _19383_ (.A1(_05786_),
    .A2(_09723_),
    .A3(_09436_),
    .A4(_09724_),
    .ZN(_09725_));
 OAI21_X1 _19384_ (.A(_06050_),
    .B1(_04417_),
    .B2(_05180_),
    .ZN(_09726_));
 OAI211_X2 _19385_ (.A(_06050_),
    .B(_16831_),
    .C1(_05511_),
    .C2(_04351_),
    .ZN(_09727_));
 AND4_X1 _19386_ (.A1(_09722_),
    .A2(_09725_),
    .A3(_09726_),
    .A4(_09727_),
    .ZN(_09728_));
 OAI21_X1 _19387_ (.A(_06435_),
    .B1(_09473_),
    .B2(_05456_),
    .ZN(_09729_));
 NAND4_X1 _19388_ (.A1(_04833_),
    .A2(_05467_),
    .A3(_06127_),
    .A4(_05522_),
    .ZN(_09730_));
 OAI21_X1 _19389_ (.A(_06435_),
    .B1(_05566_),
    .B2(_05984_),
    .ZN(_09731_));
 NAND4_X1 _19390_ (.A1(_09499_),
    .A2(_09729_),
    .A3(_09730_),
    .A4(_09731_),
    .ZN(_09732_));
 AND3_X1 _19391_ (.A1(_04888_),
    .A2(_04669_),
    .A3(_06303_),
    .ZN(_09733_));
 AND2_X1 _19392_ (.A1(_04417_),
    .A2(_06303_),
    .ZN(_09734_));
 AND2_X1 _19393_ (.A1(_09701_),
    .A2(_06303_),
    .ZN(_09735_));
 NOR4_X1 _19394_ (.A1(_09732_),
    .A2(_09733_),
    .A3(_09734_),
    .A4(_09735_),
    .ZN(_09736_));
 NAND3_X1 _19395_ (.A1(_04417_),
    .A2(_09438_),
    .A3(_06127_),
    .ZN(_09737_));
 NAND2_X1 _19396_ (.A1(_09491_),
    .A2(_05313_),
    .ZN(_09738_));
 OAI221_X1 _19397_ (.A(_09737_),
    .B1(_06358_),
    .B2(_05973_),
    .C1(_05764_),
    .C2(_09738_),
    .ZN(_09739_));
 OR2_X1 _19398_ (.A1(_04888_),
    .A2(_09507_),
    .ZN(_09740_));
 AND2_X1 _19399_ (.A1(_09740_),
    .A2(_09482_),
    .ZN(_09741_));
 NAND2_X1 _19400_ (.A1(_06347_),
    .A2(_04921_),
    .ZN(_09742_));
 AND2_X2 _19401_ (.A1(_04384_),
    .A2(_04231_),
    .ZN(_09743_));
 NAND3_X1 _19402_ (.A1(_09743_),
    .A2(_09438_),
    .A3(_06127_),
    .ZN(_09744_));
 NAND4_X1 _19403_ (.A1(_09490_),
    .A2(_09493_),
    .A3(_09742_),
    .A4(_09744_),
    .ZN(_09745_));
 OAI211_X2 _19404_ (.A(_06149_),
    .B(_05401_),
    .C1(_04395_),
    .C2(_04647_),
    .ZN(_09746_));
 NAND3_X1 _19405_ (.A1(_06138_),
    .A2(_04275_),
    .A3(_05401_),
    .ZN(_09747_));
 INV_X8 _19406_ (.A(_06149_),
    .ZN(_09748_));
 OAI211_X2 _19407_ (.A(_09746_),
    .B(_09747_),
    .C1(_05973_),
    .C2(_09748_),
    .ZN(_09749_));
 NOR4_X1 _19408_ (.A1(_09739_),
    .A2(_09741_),
    .A3(_09745_),
    .A4(_09749_),
    .ZN(_09750_));
 AND2_X1 _19409_ (.A1(_04658_),
    .A2(_04669_),
    .ZN(_09751_));
 OAI21_X1 _19410_ (.A(_05841_),
    .B1(_09751_),
    .B2(_09473_),
    .ZN(_09752_));
 NAND2_X1 _19411_ (.A1(_05047_),
    .A2(_05808_),
    .ZN(_09753_));
 AND2_X1 _19412_ (.A1(_05808_),
    .A2(_05188_),
    .ZN(_09754_));
 INV_X1 _19413_ (.A(_09754_),
    .ZN(_09755_));
 NAND4_X1 _19414_ (.A1(_09752_),
    .A2(_09429_),
    .A3(_09753_),
    .A4(_09755_),
    .ZN(_09756_));
 AOI211_X4 _19415_ (.A(_05896_),
    .B(_05962_),
    .C1(_04275_),
    .C2(_05198_),
    .ZN(_09757_));
 OAI21_X4 _19416_ (.A(_05940_),
    .B1(_05152_),
    .B2(_04855_),
    .ZN(_09758_));
 NAND4_X1 _19417_ (.A1(_05907_),
    .A2(_05269_),
    .A3(_05863_),
    .A4(_05467_),
    .ZN(_09759_));
 OAI211_X2 _19418_ (.A(_09758_),
    .B(_09759_),
    .C1(_05962_),
    .C2(_05214_),
    .ZN(_09760_));
 NOR4_X1 _19419_ (.A1(_09756_),
    .A2(_09757_),
    .A3(_06006_),
    .A4(_09760_),
    .ZN(_09761_));
 NAND4_X2 _19420_ (.A1(_09728_),
    .A2(_09736_),
    .A3(_09750_),
    .A4(_09761_),
    .ZN(_09762_));
 NOR2_X4 _19421_ (.A1(_09721_),
    .A2(_09762_),
    .ZN(_09763_));
 XNOR2_X1 _19422_ (.A(_09685_),
    .B(_09763_),
    .ZN(_09764_));
 AND2_X1 _19423_ (.A1(_09309_),
    .A2(_08991_),
    .ZN(_09765_));
 AND3_X1 _19424_ (.A1(_08946_),
    .A2(_08916_),
    .A3(_08993_),
    .ZN(_09766_));
 NOR2_X1 _19425_ (.A1(_09765_),
    .A2(_09766_),
    .ZN(_09767_));
 AND2_X1 _19426_ (.A1(_09355_),
    .A2(_08907_),
    .ZN(_09768_));
 OAI21_X1 _19427_ (.A(_09354_),
    .B1(_08987_),
    .B2(_09768_),
    .ZN(_09769_));
 NAND3_X1 _19428_ (.A1(_09330_),
    .A2(_08962_),
    .A3(_08926_),
    .ZN(_09770_));
 NAND2_X1 _19429_ (.A1(_08906_),
    .A2(_09400_),
    .ZN(_09771_));
 NAND4_X1 _19430_ (.A1(_09767_),
    .A2(_09769_),
    .A3(_09770_),
    .A4(_09771_),
    .ZN(_09772_));
 NAND2_X1 _19431_ (.A1(_09026_),
    .A2(_09346_),
    .ZN(_09773_));
 NAND2_X1 _19432_ (.A1(_08998_),
    .A2(_09346_),
    .ZN(_09774_));
 NAND3_X1 _19433_ (.A1(_08937_),
    .A2(_08950_),
    .A3(_09015_),
    .ZN(_09775_));
 NAND3_X1 _19434_ (.A1(_09773_),
    .A2(_09774_),
    .A3(_09775_),
    .ZN(_09776_));
 AND2_X1 _19435_ (.A1(_09084_),
    .A2(_08926_),
    .ZN(_09777_));
 AND2_X1 _19436_ (.A1(_09392_),
    .A2(_08901_),
    .ZN(_09778_));
 OR3_X1 _19437_ (.A1(_09776_),
    .A2(_09777_),
    .A3(_09778_),
    .ZN(_09779_));
 NOR4_X2 _19438_ (.A1(_09772_),
    .A2(_09779_),
    .A3(_08935_),
    .A4(_09360_),
    .ZN(_09780_));
 NAND2_X1 _19439_ (.A1(_09079_),
    .A2(_09310_),
    .ZN(_09781_));
 AND3_X1 _19440_ (.A1(_09378_),
    .A2(_08921_),
    .A3(_09015_),
    .ZN(_09782_));
 AND2_X1 _19441_ (.A1(_09339_),
    .A2(_08985_),
    .ZN(_09783_));
 BUF_X4 _19442_ (.A(_08908_),
    .Z(_09784_));
 AND3_X1 _19443_ (.A1(_09344_),
    .A2(_09784_),
    .A3(_09039_),
    .ZN(_09785_));
 NOR4_X1 _19444_ (.A1(_09290_),
    .A2(_09782_),
    .A3(_09783_),
    .A4(_09785_),
    .ZN(_09786_));
 NAND2_X1 _19445_ (.A1(_09309_),
    .A2(_09329_),
    .ZN(_09787_));
 AND3_X1 _19446_ (.A1(_08987_),
    .A2(_09346_),
    .A3(_08962_),
    .ZN(_09788_));
 BUF_X4 _19447_ (.A(_08991_),
    .Z(_09789_));
 AOI21_X1 _19448_ (.A(_09788_),
    .B1(_09789_),
    .B2(_09374_),
    .ZN(_09790_));
 AND4_X1 _19449_ (.A1(_09781_),
    .A2(_09786_),
    .A3(_09787_),
    .A4(_09790_),
    .ZN(_09791_));
 AND4_X1 _19450_ (.A1(_08977_),
    .A2(_08954_),
    .A3(_09057_),
    .A4(_08945_),
    .ZN(_09792_));
 NOR2_X1 _19451_ (.A1(_09335_),
    .A2(_09792_),
    .ZN(_09793_));
 INV_X1 _19452_ (.A(_08919_),
    .ZN(_09794_));
 NAND4_X1 _19453_ (.A1(_09794_),
    .A2(_09371_),
    .A3(_09380_),
    .A4(_09071_),
    .ZN(_09795_));
 NAND2_X1 _19454_ (.A1(_09795_),
    .A2(_09327_),
    .ZN(_09796_));
 BUF_X4 _19455_ (.A(_09081_),
    .Z(_09797_));
 OAI21_X1 _19456_ (.A(_09797_),
    .B1(_09347_),
    .B2(_09344_),
    .ZN(_09798_));
 OAI21_X1 _19457_ (.A(_09074_),
    .B1(_08981_),
    .B2(_08969_),
    .ZN(_09799_));
 AND4_X1 _19458_ (.A1(_09793_),
    .A2(_09796_),
    .A3(_09798_),
    .A4(_09799_),
    .ZN(_09800_));
 OAI21_X1 _19459_ (.A(_09326_),
    .B1(_08981_),
    .B2(_08948_),
    .ZN(_09801_));
 AND2_X1 _19460_ (.A1(_09327_),
    .A2(_08899_),
    .ZN(_09802_));
 AND3_X1 _19461_ (.A1(_09026_),
    .A2(_09057_),
    .A3(_08921_),
    .ZN(_09803_));
 AND2_X1 _19462_ (.A1(_09378_),
    .A2(_09081_),
    .ZN(_09804_));
 NOR3_X1 _19463_ (.A1(_09802_),
    .A2(_09803_),
    .A3(_09804_),
    .ZN(_09805_));
 OAI21_X1 _19464_ (.A(_09329_),
    .B1(_09347_),
    .B2(_08937_),
    .ZN(_09806_));
 OAI21_X1 _19465_ (.A(_09053_),
    .B1(_09072_),
    .B2(_09325_),
    .ZN(_09807_));
 AND4_X1 _19466_ (.A1(_09801_),
    .A2(_09805_),
    .A3(_09806_),
    .A4(_09807_),
    .ZN(_09808_));
 NAND4_X1 _19467_ (.A1(_09780_),
    .A2(_09791_),
    .A3(_09800_),
    .A4(_09808_),
    .ZN(_09809_));
 AND2_X1 _19468_ (.A1(_08983_),
    .A2(_09087_),
    .ZN(_09810_));
 AND2_X4 _19469_ (.A1(_09394_),
    .A2(_09382_),
    .ZN(_09811_));
 OR4_X2 _19470_ (.A1(_08952_),
    .A2(_09810_),
    .A3(_09811_),
    .A4(_09007_),
    .ZN(_09812_));
 AND2_X4 _19471_ (.A1(_09039_),
    .A2(_09331_),
    .ZN(_09813_));
 AND2_X1 _19472_ (.A1(_08947_),
    .A2(_08932_),
    .ZN(_09814_));
 OAI21_X1 _19473_ (.A(_08938_),
    .B1(_09303_),
    .B2(_09009_),
    .ZN(_09815_));
 NOR4_X2 _19474_ (.A1(_09812_),
    .A2(_09813_),
    .A3(_09814_),
    .A4(_09815_),
    .ZN(_09816_));
 AND2_X1 _19475_ (.A1(_09378_),
    .A2(_09382_),
    .ZN(_09817_));
 AND2_X1 _19476_ (.A1(_09053_),
    .A2(_09018_),
    .ZN(_09818_));
 NOR2_X1 _19477_ (.A1(_09817_),
    .A2(_09818_),
    .ZN(_09819_));
 OAI21_X1 _19478_ (.A(_09377_),
    .B1(_09079_),
    .B2(_09344_),
    .ZN(_09820_));
 NAND4_X1 _19479_ (.A1(_09397_),
    .A2(_09054_),
    .A3(_16871_),
    .A4(_09398_),
    .ZN(_09821_));
 AND4_X1 _19480_ (.A1(_09370_),
    .A2(_09819_),
    .A3(_09820_),
    .A4(_09821_),
    .ZN(_09822_));
 INV_X1 _19481_ (.A(_09405_),
    .ZN(_09823_));
 OR2_X1 _19482_ (.A1(_09061_),
    .A2(_09823_),
    .ZN(_09824_));
 AND2_X1 _19483_ (.A1(_09407_),
    .A2(_09408_),
    .ZN(_09825_));
 NOR3_X1 _19484_ (.A1(_09019_),
    .A2(_09825_),
    .A3(_09021_),
    .ZN(_09826_));
 AOI22_X1 _19485_ (.A1(_09789_),
    .A2(_09296_),
    .B1(_09330_),
    .B2(_09394_),
    .ZN(_09827_));
 AOI22_X1 _19486_ (.A1(_08961_),
    .A2(_09330_),
    .B1(_09397_),
    .B2(_09331_),
    .ZN(_09828_));
 AND4_X1 _19487_ (.A1(_09824_),
    .A2(_09826_),
    .A3(_09827_),
    .A4(_09828_),
    .ZN(_09829_));
 AOI22_X1 _19488_ (.A1(_09327_),
    .A2(_09404_),
    .B1(_09797_),
    .B2(_09296_),
    .ZN(_09830_));
 AOI22_X1 _19489_ (.A1(_09310_),
    .A2(_09768_),
    .B1(_09330_),
    .B2(_09404_),
    .ZN(_09831_));
 BUF_X4 _19490_ (.A(_09087_),
    .Z(_09832_));
 OAI211_X2 _19491_ (.A(_09305_),
    .B(_09784_),
    .C1(_08977_),
    .C2(_09832_),
    .ZN(_09833_));
 AOI22_X1 _19492_ (.A1(_09339_),
    .A2(_09364_),
    .B1(_09377_),
    .B2(_09340_),
    .ZN(_09834_));
 AND4_X1 _19493_ (.A1(_09830_),
    .A2(_09831_),
    .A3(_09833_),
    .A4(_09834_),
    .ZN(_09835_));
 NAND4_X2 _19494_ (.A1(_09816_),
    .A2(_09822_),
    .A3(_09829_),
    .A4(_09835_),
    .ZN(_09836_));
 NOR2_X4 _19495_ (.A1(_09809_),
    .A2(_09836_),
    .ZN(_09837_));
 INV_X1 _19496_ (.A(_09837_),
    .ZN(_09838_));
 XNOR2_X1 _19497_ (.A(_09287_),
    .B(_09838_),
    .ZN(_09839_));
 XNOR2_X1 _19498_ (.A(_09764_),
    .B(_09839_),
    .ZN(_09840_));
 XNOR2_X1 _19499_ (.A(_09840_),
    .B(_17166_),
    .ZN(_09841_));
 MUX2_X1 _19500_ (.A(_09534_),
    .B(_09841_),
    .S(_09100_),
    .Z(_00726_));
 XOR2_X1 _19501_ (.A(_17169_),
    .B(_17073_),
    .Z(_09842_));
 NAND2_X1 _19502_ (.A1(_08956_),
    .A2(_08925_),
    .ZN(_09843_));
 NOR2_X1 _19503_ (.A1(_09357_),
    .A2(_09843_),
    .ZN(_09844_));
 AND2_X1 _19504_ (.A1(_09064_),
    .A2(_08964_),
    .ZN(_09845_));
 OR2_X1 _19505_ (.A1(_09065_),
    .A2(_09845_),
    .ZN(_09846_));
 AND2_X2 _19506_ (.A1(_09074_),
    .A2(_09340_),
    .ZN(_09847_));
 AOI21_X1 _19507_ (.A(_09357_),
    .B1(_09035_),
    .B2(_09067_),
    .ZN(_09848_));
 OR4_X4 _19508_ (.A1(_09844_),
    .A2(_09846_),
    .A3(_09847_),
    .A4(_09848_),
    .ZN(_09849_));
 AND2_X1 _19509_ (.A1(_09330_),
    .A2(_09340_),
    .ZN(_09850_));
 AND2_X1 _19510_ (.A1(_09058_),
    .A2(_08926_),
    .ZN(_09851_));
 AND2_X1 _19511_ (.A1(_09058_),
    .A2(_09404_),
    .ZN(_09852_));
 AND2_X1 _19512_ (.A1(_09058_),
    .A2(_09318_),
    .ZN(_09853_));
 OR2_X1 _19513_ (.A1(_09852_),
    .A2(_09853_),
    .ZN(_09854_));
 NOR4_X4 _19514_ (.A1(_09849_),
    .A2(_09850_),
    .A3(_09851_),
    .A4(_09854_),
    .ZN(_09855_));
 OAI21_X1 _19515_ (.A(_09397_),
    .B1(_08899_),
    .B2(_09318_),
    .ZN(_09856_));
 AND2_X1 _19516_ (.A1(_08981_),
    .A2(_09392_),
    .ZN(_09857_));
 AND2_X1 _19517_ (.A1(_09392_),
    .A2(_08998_),
    .ZN(_09858_));
 AND2_X1 _19518_ (.A1(_09016_),
    .A2(_08988_),
    .ZN(_09859_));
 NOR4_X1 _19519_ (.A1(_09857_),
    .A2(_09858_),
    .A3(_09859_),
    .A4(_09019_),
    .ZN(_09860_));
 NAND4_X1 _19520_ (.A1(_08892_),
    .A2(_08961_),
    .A3(_09015_),
    .A4(_09054_),
    .ZN(_09861_));
 OAI21_X1 _19521_ (.A(_09397_),
    .B1(_09072_),
    .B2(_09394_),
    .ZN(_09862_));
 AND4_X1 _19522_ (.A1(_09856_),
    .A2(_09860_),
    .A3(_09861_),
    .A4(_09862_),
    .ZN(_09863_));
 OAI211_X2 _19523_ (.A(_09405_),
    .B(_09832_),
    .C1(_08909_),
    .C2(_08954_),
    .ZN(_09864_));
 OAI21_X1 _19524_ (.A(_09405_),
    .B1(_08985_),
    .B2(_08926_),
    .ZN(_09865_));
 OAI21_X1 _19525_ (.A(_09405_),
    .B1(_09018_),
    .B2(_09331_),
    .ZN(_09866_));
 NAND4_X1 _19526_ (.A1(_09864_),
    .A2(_09865_),
    .A3(_09866_),
    .A4(_09774_),
    .ZN(_09867_));
 OAI211_X2 _19527_ (.A(_09054_),
    .B(_09053_),
    .C1(_09340_),
    .C2(_09832_),
    .ZN(_09868_));
 NAND2_X1 _19528_ (.A1(_08899_),
    .A2(_09053_),
    .ZN(_09869_));
 NAND2_X1 _19529_ (.A1(_09868_),
    .A2(_09869_),
    .ZN(_09870_));
 AND2_X1 _19530_ (.A1(_09053_),
    .A2(_08926_),
    .ZN(_09871_));
 NOR4_X1 _19531_ (.A1(_09867_),
    .A2(_09870_),
    .A3(_09050_),
    .A4(_09871_),
    .ZN(_09872_));
 INV_X1 _19532_ (.A(_09080_),
    .ZN(_09873_));
 OAI211_X2 _19533_ (.A(_09797_),
    .B(_09832_),
    .C1(_08962_),
    .C2(_08900_),
    .ZN(_09874_));
 OAI211_X2 _19534_ (.A(_09873_),
    .B(_09874_),
    .C1(_09349_),
    .C2(_09380_),
    .ZN(_09875_));
 OAI21_X1 _19535_ (.A(_09339_),
    .B1(_09347_),
    .B2(_08899_),
    .ZN(_09876_));
 OAI211_X2 _19536_ (.A(_09339_),
    .B(_09355_),
    .C1(_09054_),
    .C2(_09784_),
    .ZN(_09877_));
 NAND2_X1 _19537_ (.A1(_09876_),
    .A2(_09877_),
    .ZN(_09878_));
 NAND2_X1 _19538_ (.A1(_09378_),
    .A2(_09797_),
    .ZN(_09879_));
 OAI21_X1 _19539_ (.A(_09879_),
    .B1(_09035_),
    .B2(_09349_),
    .ZN(_09880_));
 NOR4_X1 _19540_ (.A1(_09875_),
    .A2(_09878_),
    .A3(_09351_),
    .A4(_09880_),
    .ZN(_09881_));
 NAND4_X1 _19541_ (.A1(_09855_),
    .A2(_09863_),
    .A3(_09872_),
    .A4(_09881_),
    .ZN(_09882_));
 NOR2_X4 _19542_ (.A1(_08992_),
    .A2(_09843_),
    .ZN(_09883_));
 AOI211_X2 _19543_ (.A(_08999_),
    .B(_09883_),
    .C1(_09394_),
    .C2(_09789_),
    .ZN(_09884_));
 AND4_X1 _19544_ (.A1(_08944_),
    .A2(_08904_),
    .A3(_09087_),
    .A4(_08954_),
    .ZN(_09885_));
 AND4_X1 _19545_ (.A1(_08944_),
    .A2(_08921_),
    .A3(_08918_),
    .A4(_08932_),
    .ZN(_09886_));
 AOI211_X4 _19546_ (.A(_09885_),
    .B(_09886_),
    .C1(_09404_),
    .C2(_08991_),
    .ZN(_09887_));
 OAI21_X1 _19547_ (.A(_09377_),
    .B1(_09323_),
    .B2(_08924_),
    .ZN(_09888_));
 OAI21_X1 _19548_ (.A(_09377_),
    .B1(_09293_),
    .B2(_08988_),
    .ZN(_09889_));
 AND4_X1 _19549_ (.A1(_09884_),
    .A2(_09887_),
    .A3(_09888_),
    .A4(_09889_),
    .ZN(_09890_));
 NAND2_X1 _19550_ (.A1(_09378_),
    .A2(_09310_),
    .ZN(_09891_));
 OAI211_X2 _19551_ (.A(_09310_),
    .B(_09832_),
    .C1(_09054_),
    .C2(_08900_),
    .ZN(_09892_));
 NAND4_X1 _19552_ (.A1(_09376_),
    .A2(_08967_),
    .A3(_09891_),
    .A4(_09892_),
    .ZN(_09893_));
 NAND2_X1 _19553_ (.A1(_09814_),
    .A2(_08956_),
    .ZN(_09894_));
 NAND3_X1 _19554_ (.A1(_08947_),
    .A2(_09087_),
    .A3(_08954_),
    .ZN(_09895_));
 NAND2_X1 _19555_ (.A1(_09894_),
    .A2(_09895_),
    .ZN(_09896_));
 INV_X1 _19556_ (.A(_08947_),
    .ZN(_09897_));
 NOR3_X1 _19557_ (.A1(_09897_),
    .A2(_08994_),
    .A3(_09017_),
    .ZN(_09898_));
 NOR4_X1 _19558_ (.A1(_09893_),
    .A2(_09896_),
    .A3(_09306_),
    .A4(_09898_),
    .ZN(_09899_));
 NOR2_X1 _19559_ (.A1(_09024_),
    .A2(_08954_),
    .ZN(_09900_));
 OAI21_X1 _19560_ (.A(_09354_),
    .B1(_09900_),
    .B2(_09347_),
    .ZN(_09901_));
 NAND2_X1 _19561_ (.A1(_09354_),
    .A2(_08985_),
    .ZN(_09902_));
 NAND2_X1 _19562_ (.A1(_09354_),
    .A2(_09026_),
    .ZN(_09903_));
 AND3_X1 _19563_ (.A1(_08920_),
    .A2(_09902_),
    .A3(_09903_),
    .ZN(_09904_));
 OAI21_X1 _19564_ (.A(_09326_),
    .B1(_09002_),
    .B2(_09404_),
    .ZN(_09905_));
 OAI21_X1 _19565_ (.A(_09326_),
    .B1(_09325_),
    .B2(_09374_),
    .ZN(_09906_));
 AND4_X1 _19566_ (.A1(_09901_),
    .A2(_09904_),
    .A3(_09905_),
    .A4(_09906_),
    .ZN(_09907_));
 OAI21_X1 _19567_ (.A(_09329_),
    .B1(_09026_),
    .B2(_08955_),
    .ZN(_09908_));
 OAI21_X1 _19568_ (.A(_09329_),
    .B1(_08899_),
    .B2(_09331_),
    .ZN(_09909_));
 OAI21_X1 _19569_ (.A(_09327_),
    .B1(_09026_),
    .B2(_09374_),
    .ZN(_09910_));
 OAI21_X1 _19570_ (.A(_09327_),
    .B1(_08899_),
    .B2(_08988_),
    .ZN(_09911_));
 AND4_X1 _19571_ (.A1(_09908_),
    .A2(_09909_),
    .A3(_09910_),
    .A4(_09911_),
    .ZN(_09912_));
 NAND4_X1 _19572_ (.A1(_09890_),
    .A2(_09899_),
    .A3(_09907_),
    .A4(_09912_),
    .ZN(_09913_));
 NOR2_X4 _19573_ (.A1(_09882_),
    .A2(_09913_),
    .ZN(_09914_));
 XOR2_X1 _19574_ (.A(_09914_),
    .B(_09093_),
    .Z(_09915_));
 OAI21_X1 _19575_ (.A(_08714_),
    .B1(_08596_),
    .B2(_08778_),
    .ZN(_09916_));
 NAND4_X1 _19576_ (.A1(_08725_),
    .A2(_08683_),
    .A3(_08649_),
    .A4(_08592_),
    .ZN(_09917_));
 AND3_X1 _19577_ (.A1(_09916_),
    .A2(_09621_),
    .A3(_09917_),
    .ZN(_09918_));
 NAND2_X1 _19578_ (.A1(_08720_),
    .A2(_08843_),
    .ZN(_09919_));
 AND2_X1 _19579_ (.A1(_08729_),
    .A2(_09919_),
    .ZN(_09920_));
 INV_X1 _19580_ (.A(_09920_),
    .ZN(_09921_));
 AND2_X1 _19581_ (.A1(_08721_),
    .A2(_08697_),
    .ZN(_09922_));
 AND2_X1 _19582_ (.A1(_08720_),
    .A2(_08836_),
    .ZN(_09923_));
 NOR4_X2 _19583_ (.A1(_09921_),
    .A2(_09922_),
    .A3(_09923_),
    .A4(_09214_),
    .ZN(_09924_));
 AOI21_X1 _19584_ (.A(_08826_),
    .B1(_08736_),
    .B2(_08737_),
    .ZN(_09925_));
 NAND4_X1 _19585_ (.A1(_08725_),
    .A2(_08584_),
    .A3(_08650_),
    .A4(_08753_),
    .ZN(_09926_));
 NAND4_X1 _19586_ (.A1(_08713_),
    .A2(_08592_),
    .A3(_08605_),
    .A4(_08650_),
    .ZN(_09927_));
 OAI211_X2 _19587_ (.A(_09926_),
    .B(_09927_),
    .C1(_08826_),
    .C2(_09641_),
    .ZN(_09928_));
 AND3_X1 _19588_ (.A1(_08730_),
    .A2(_08614_),
    .A3(_08610_),
    .ZN(_09929_));
 NOR3_X1 _19589_ (.A1(_09925_),
    .A2(_09928_),
    .A3(_09929_),
    .ZN(_09930_));
 AND2_X1 _19590_ (.A1(_08815_),
    .A2(_08741_),
    .ZN(_09931_));
 AND2_X2 _19591_ (.A1(_08740_),
    .A2(_08589_),
    .ZN(_09932_));
 AND3_X1 _19592_ (.A1(_08671_),
    .A2(_08602_),
    .A3(_08713_),
    .ZN(_09933_));
 NOR4_X1 _19593_ (.A1(_09931_),
    .A2(_09932_),
    .A3(_09618_),
    .A4(_09933_),
    .ZN(_09934_));
 AND4_X1 _19594_ (.A1(_09918_),
    .A2(_09924_),
    .A3(_09930_),
    .A4(_09934_),
    .ZN(_09935_));
 OAI211_X2 _19595_ (.A(_08788_),
    .B(_08583_),
    .C1(_08585_),
    .C2(_08586_),
    .ZN(_09936_));
 OAI211_X2 _19596_ (.A(_08788_),
    .B(_08649_),
    .C1(_08594_),
    .C2(_08592_),
    .ZN(_09937_));
 OAI21_X1 _19597_ (.A(_08788_),
    .B1(_08785_),
    .B2(_08578_),
    .ZN(_09938_));
 AND4_X1 _19598_ (.A1(_08781_),
    .A2(_09936_),
    .A3(_09937_),
    .A4(_09938_),
    .ZN(_09939_));
 OAI21_X1 _19599_ (.A(_09633_),
    .B1(_08637_),
    .B2(_08860_),
    .ZN(_09940_));
 OAI21_X1 _19600_ (.A(_09633_),
    .B1(_08810_),
    .B2(_08798_),
    .ZN(_09941_));
 OAI21_X1 _19601_ (.A(_09633_),
    .B1(_08709_),
    .B2(_08724_),
    .ZN(_09942_));
 OAI21_X1 _19602_ (.A(_08766_),
    .B1(_08631_),
    .B2(_08633_),
    .ZN(_09943_));
 AND4_X1 _19603_ (.A1(_09940_),
    .A2(_09941_),
    .A3(_09942_),
    .A4(_09943_),
    .ZN(_09944_));
 NAND2_X1 _19604_ (.A1(_08760_),
    .A2(_08673_),
    .ZN(_09945_));
 NAND4_X1 _19605_ (.A1(_08594_),
    .A2(_08754_),
    .A3(_08683_),
    .A4(_08753_),
    .ZN(_09946_));
 NAND4_X1 _19606_ (.A1(_08605_),
    .A2(_08683_),
    .A3(_08754_),
    .A4(_08592_),
    .ZN(_09947_));
 AND3_X1 _19607_ (.A1(_09945_),
    .A2(_09946_),
    .A3(_09947_),
    .ZN(_09948_));
 AND4_X1 _19608_ (.A1(_08614_),
    .A2(_08746_),
    .A3(_08762_),
    .A4(_08605_),
    .ZN(_09949_));
 AOI21_X1 _19609_ (.A(_09949_),
    .B1(_08860_),
    .B2(_08748_),
    .ZN(_09950_));
 OAI21_X1 _19610_ (.A(_09257_),
    .B1(_08758_),
    .B2(_08757_),
    .ZN(_09951_));
 AND2_X1 _19611_ (.A1(_08709_),
    .A2(_08756_),
    .ZN(_09952_));
 NOR3_X1 _19612_ (.A1(_09951_),
    .A2(_09952_),
    .A3(_08804_),
    .ZN(_09953_));
 OAI21_X1 _19613_ (.A(_08748_),
    .B1(_08709_),
    .B2(_08633_),
    .ZN(_09954_));
 AND4_X1 _19614_ (.A1(_09948_),
    .A2(_09950_),
    .A3(_09953_),
    .A4(_09954_),
    .ZN(_09955_));
 NAND4_X1 _19615_ (.A1(_09935_),
    .A2(_09939_),
    .A3(_09944_),
    .A4(_09955_),
    .ZN(_09956_));
 AND3_X1 _19616_ (.A1(_08565_),
    .A2(_08648_),
    .A3(_08605_),
    .ZN(_09957_));
 AOI211_X2 _19617_ (.A(_08571_),
    .B(_09957_),
    .C1(_08575_),
    .C2(_08642_),
    .ZN(_09958_));
 AND2_X1 _19618_ (.A1(_08630_),
    .A2(_08565_),
    .ZN(_09959_));
 AND3_X1 _19619_ (.A1(_08565_),
    .A2(_08648_),
    .A3(_08646_),
    .ZN(_09960_));
 AOI211_X2 _19620_ (.A(_09959_),
    .B(_09960_),
    .C1(_08565_),
    .C2(_08660_),
    .ZN(_09961_));
 OAI21_X1 _19621_ (.A(_08608_),
    .B1(_08798_),
    .B2(_08732_),
    .ZN(_09962_));
 OAI21_X1 _19622_ (.A(_08608_),
    .B1(_08615_),
    .B2(_08631_),
    .ZN(_09963_));
 AND4_X4 _19623_ (.A1(_09958_),
    .A2(_09961_),
    .A3(_09962_),
    .A4(_09963_),
    .ZN(_09964_));
 NAND2_X1 _19624_ (.A1(_08704_),
    .A2(_08695_),
    .ZN(_09965_));
 AND2_X1 _19625_ (.A1(_08582_),
    .A2(_08830_),
    .ZN(_09966_));
 OAI21_X1 _19626_ (.A(_08658_),
    .B1(_08666_),
    .B2(_09966_),
    .ZN(_09967_));
 NAND3_X1 _19627_ (.A1(_08606_),
    .A2(_08658_),
    .A3(_08595_),
    .ZN(_09968_));
 AND3_X1 _19628_ (.A1(_09967_),
    .A2(_08670_),
    .A3(_09968_),
    .ZN(_09969_));
 OAI21_X1 _19629_ (.A(_08704_),
    .B1(_08749_),
    .B2(_09280_),
    .ZN(_09970_));
 OAI21_X1 _19630_ (.A(_08704_),
    .B1(_08666_),
    .B2(_08633_),
    .ZN(_09971_));
 AND4_X1 _19631_ (.A1(_09965_),
    .A2(_09969_),
    .A3(_09970_),
    .A4(_09971_),
    .ZN(_09972_));
 AOI211_X4 _19632_ (.A(_08623_),
    .B(_08690_),
    .C1(_08584_),
    .C2(_08706_),
    .ZN(_09973_));
 OAI21_X1 _19633_ (.A(_08693_),
    .B1(_08779_),
    .B2(_08724_),
    .ZN(_09974_));
 OAI21_X1 _19634_ (.A(_08693_),
    .B1(_08680_),
    .B2(_08632_),
    .ZN(_09975_));
 NAND2_X1 _19635_ (.A1(_08693_),
    .A2(_08671_),
    .ZN(_09976_));
 NAND4_X1 _19636_ (.A1(_09974_),
    .A2(_08700_),
    .A3(_09975_),
    .A4(_09976_),
    .ZN(_09977_));
 NAND4_X1 _19637_ (.A1(_08675_),
    .A2(_08830_),
    .A3(_08646_),
    .A4(_08683_),
    .ZN(_09978_));
 OAI21_X1 _19638_ (.A(_09978_),
    .B1(_08840_),
    .B2(_08690_),
    .ZN(_09979_));
 NOR4_X1 _19639_ (.A1(_09973_),
    .A2(_09977_),
    .A3(_09270_),
    .A4(_09979_),
    .ZN(_09980_));
 OAI21_X1 _19640_ (.A(_08622_),
    .B1(_08860_),
    .B2(_08671_),
    .ZN(_09981_));
 NAND3_X1 _19641_ (.A1(_08717_),
    .A2(_08762_),
    .A3(_08645_),
    .ZN(_09982_));
 NAND2_X1 _19642_ (.A1(_08645_),
    .A2(_08631_),
    .ZN(_09983_));
 AND4_X1 _19643_ (.A1(_08883_),
    .A2(_09981_),
    .A3(_09982_),
    .A4(_09983_),
    .ZN(_09984_));
 NAND4_X1 _19644_ (.A1(_09964_),
    .A2(_09972_),
    .A3(_09980_),
    .A4(_09984_),
    .ZN(_09985_));
 NOR2_X4 _19645_ (.A1(_09956_),
    .A2(_09985_),
    .ZN(_09986_));
 NAND2_X1 _19646_ (.A1(_07084_),
    .A2(_07403_),
    .ZN(_09987_));
 OAI211_X2 _19647_ (.A(_09987_),
    .B(_09566_),
    .C1(_08541_),
    .C2(_09163_),
    .ZN(_09988_));
 OAI21_X1 _19648_ (.A(_08534_),
    .B1(_09140_),
    .B2(_09163_),
    .ZN(_09989_));
 AOI21_X1 _19649_ (.A(_09163_),
    .B1(_08332_),
    .B2(_08433_),
    .ZN(_09990_));
 NOR3_X1 _19650_ (.A1(_09988_),
    .A2(_09989_),
    .A3(_09990_),
    .ZN(_09991_));
 AND3_X1 _19651_ (.A1(_09125_),
    .A2(_07960_),
    .A3(_08519_),
    .ZN(_09992_));
 AND3_X1 _19652_ (.A1(_09199_),
    .A2(_09145_),
    .A3(_06710_),
    .ZN(_09993_));
 AOI211_X2 _19653_ (.A(_09992_),
    .B(_09993_),
    .C1(_09166_),
    .C2(_07172_),
    .ZN(_09994_));
 OAI211_X2 _19654_ (.A(_09557_),
    .B(_09558_),
    .C1(_09187_),
    .C2(_07510_),
    .ZN(_09995_));
 AND3_X1 _19655_ (.A1(_07326_),
    .A2(_08244_),
    .A3(_07927_),
    .ZN(_09996_));
 NOR3_X1 _19656_ (.A1(_09995_),
    .A2(_09554_),
    .A3(_09996_),
    .ZN(_09997_));
 AND4_X1 _19657_ (.A1(_07051_),
    .A2(_07304_),
    .A3(_06897_),
    .A4(_08519_),
    .ZN(_09998_));
 AND4_X1 _19658_ (.A1(_06644_),
    .A2(_07304_),
    .A3(_07051_),
    .A4(_08519_),
    .ZN(_09999_));
 AOI211_X4 _19659_ (.A(_09998_),
    .B(_09999_),
    .C1(_07172_),
    .C2(_09133_),
    .ZN(_10000_));
 AND4_X1 _19660_ (.A1(_09991_),
    .A2(_09994_),
    .A3(_09997_),
    .A4(_10000_),
    .ZN(_10001_));
 NAND3_X1 _19661_ (.A1(_07293_),
    .A2(_09145_),
    .A3(_07653_),
    .ZN(_10002_));
 NAND2_X4 _19662_ (.A1(_09140_),
    .A2(_07510_),
    .ZN(_10003_));
 AND2_X2 _19663_ (.A1(_10003_),
    .A2(_07477_),
    .ZN(_10004_));
 INV_X1 _19664_ (.A(_10004_),
    .ZN(_10005_));
 OAI21_X1 _19665_ (.A(_07905_),
    .B1(_06754_),
    .B2(_07205_),
    .ZN(_10006_));
 OAI21_X1 _19666_ (.A(_08556_),
    .B1(_09192_),
    .B2(_07719_),
    .ZN(_10007_));
 AND4_X1 _19667_ (.A1(_10002_),
    .A2(_10005_),
    .A3(_10006_),
    .A4(_10007_),
    .ZN(_10008_));
 NAND4_X1 _19668_ (.A1(_08244_),
    .A2(_07062_),
    .A3(_08080_),
    .A4(_08058_),
    .ZN(_10009_));
 NAND4_X1 _19669_ (.A1(_09204_),
    .A2(_09160_),
    .A3(_09149_),
    .A4(_10009_),
    .ZN(_10010_));
 NAND2_X1 _19670_ (.A1(_08190_),
    .A2(_07447_),
    .ZN(_10011_));
 OAI21_X1 _19671_ (.A(_10011_),
    .B1(_09585_),
    .B2(_09120_),
    .ZN(_10012_));
 AND2_X1 _19672_ (.A1(_07631_),
    .A2(_08299_),
    .ZN(_10013_));
 AND2_X1 _19673_ (.A1(_08550_),
    .A2(_07828_),
    .ZN(_10014_));
 NOR4_X1 _19674_ (.A1(_10010_),
    .A2(_10012_),
    .A3(_10013_),
    .A4(_10014_),
    .ZN(_10015_));
 NAND2_X1 _19675_ (.A1(_07205_),
    .A2(_06611_),
    .ZN(_10016_));
 NAND4_X1 _19676_ (.A1(_08047_),
    .A2(_07436_),
    .A3(_08080_),
    .A4(_07238_),
    .ZN(_10017_));
 OAI211_X2 _19677_ (.A(_10016_),
    .B(_10017_),
    .C1(_08541_),
    .C2(_07348_),
    .ZN(_10018_));
 AOI21_X1 _19678_ (.A(_07348_),
    .B1(_08135_),
    .B2(_08146_),
    .ZN(_10019_));
 AND4_X1 _19679_ (.A1(_08069_),
    .A2(_08538_),
    .A3(_08080_),
    .A4(_07238_),
    .ZN(_10020_));
 NOR3_X1 _19680_ (.A1(_10018_),
    .A2(_10019_),
    .A3(_10020_),
    .ZN(_10021_));
 NAND2_X1 _19681_ (.A1(_07905_),
    .A2(_09131_),
    .ZN(_10022_));
 NAND2_X1 _19682_ (.A1(_08190_),
    .A2(_09106_),
    .ZN(_10023_));
 AND2_X1 _19683_ (.A1(_10022_),
    .A2(_10023_),
    .ZN(_10024_));
 AND2_X1 _19684_ (.A1(_09188_),
    .A2(_09192_),
    .ZN(_10025_));
 INV_X1 _19685_ (.A(_10025_),
    .ZN(_10026_));
 AND3_X4 _19686_ (.A1(_08556_),
    .A2(_07883_),
    .A3(_08058_),
    .ZN(_10027_));
 NOR2_X1 _19687_ (.A1(_09561_),
    .A2(_10027_),
    .ZN(_10028_));
 AND4_X1 _19688_ (.A1(_10021_),
    .A2(_10024_),
    .A3(_10026_),
    .A4(_10028_),
    .ZN(_10029_));
 NAND4_X1 _19689_ (.A1(_10001_),
    .A2(_10008_),
    .A3(_10015_),
    .A4(_10029_),
    .ZN(_10030_));
 OR2_X1 _19690_ (.A1(_07916_),
    .A2(_08545_),
    .ZN(_10031_));
 AND2_X1 _19691_ (.A1(_06952_),
    .A2(_08025_),
    .ZN(_10032_));
 NOR2_X1 _19692_ (.A1(_10032_),
    .A2(_09177_),
    .ZN(_10033_));
 INV_X1 _19693_ (.A(_10033_),
    .ZN(_10034_));
 NOR4_X1 _19694_ (.A1(_10031_),
    .A2(_10034_),
    .A3(_06864_),
    .A4(_09196_),
    .ZN(_10035_));
 OAI21_X1 _19695_ (.A(_09550_),
    .B1(_09145_),
    .B2(_06996_),
    .ZN(_10036_));
 OAI21_X1 _19696_ (.A(_07795_),
    .B1(_10036_),
    .B2(_06754_),
    .ZN(_10037_));
 AND2_X1 _19697_ (.A1(_07740_),
    .A2(_07029_),
    .ZN(_10038_));
 INV_X1 _19698_ (.A(_10038_),
    .ZN(_10039_));
 NAND3_X1 _19699_ (.A1(_08135_),
    .A2(_08146_),
    .A3(_10039_),
    .ZN(_10040_));
 NAND2_X1 _19700_ (.A1(_10040_),
    .A2(_07532_),
    .ZN(_10041_));
 OAI22_X1 _19701_ (.A1(_08386_),
    .A2(_07282_),
    .B1(_09145_),
    .B2(_06721_),
    .ZN(_10042_));
 OAI21_X1 _19702_ (.A(_08299_),
    .B1(_10042_),
    .B2(_08168_),
    .ZN(_10043_));
 AND3_X1 _19703_ (.A1(_10037_),
    .A2(_10041_),
    .A3(_10043_),
    .ZN(_10044_));
 AND2_X1 _19704_ (.A1(_07982_),
    .A2(_08310_),
    .ZN(_10045_));
 INV_X1 _19705_ (.A(_10045_),
    .ZN(_10046_));
 INV_X1 _19706_ (.A(_09139_),
    .ZN(_10047_));
 NAND2_X1 _19707_ (.A1(_09138_),
    .A2(_07106_),
    .ZN(_10048_));
 NAND4_X1 _19708_ (.A1(_10046_),
    .A2(_10047_),
    .A3(_09593_),
    .A4(_10048_),
    .ZN(_10049_));
 AND2_X1 _19709_ (.A1(_08069_),
    .A2(_16791_),
    .ZN(_10050_));
 AND2_X1 _19710_ (.A1(_06963_),
    .A2(_10050_),
    .ZN(_10051_));
 OAI21_X1 _19711_ (.A(_09537_),
    .B1(_08135_),
    .B2(_08542_),
    .ZN(_10052_));
 NOR4_X1 _19712_ (.A1(_10049_),
    .A2(_09591_),
    .A3(_10051_),
    .A4(_10052_),
    .ZN(_10053_));
 OAI21_X1 _19713_ (.A(_08550_),
    .B1(_10003_),
    .B2(_07392_),
    .ZN(_10054_));
 OR2_X1 _19714_ (.A1(_07499_),
    .A2(_08222_),
    .ZN(_10055_));
 OAI21_X1 _19715_ (.A(_07117_),
    .B1(_10055_),
    .B2(_07447_),
    .ZN(_10056_));
 AND2_X1 _19716_ (.A1(_08544_),
    .A2(_09142_),
    .ZN(_10057_));
 AND2_X1 _19717_ (.A1(_09125_),
    .A2(_07708_),
    .ZN(_10058_));
 NOR2_X1 _19718_ (.A1(_10057_),
    .A2(_10058_),
    .ZN(_10059_));
 NAND2_X1 _19719_ (.A1(_07828_),
    .A2(_06853_),
    .ZN(_10060_));
 NAND2_X1 _19720_ (.A1(_07205_),
    .A2(_07260_),
    .ZN(_10061_));
 AND2_X1 _19721_ (.A1(_10060_),
    .A2(_10061_),
    .ZN(_10062_));
 AND4_X1 _19722_ (.A1(_10054_),
    .A2(_10056_),
    .A3(_10059_),
    .A4(_10062_),
    .ZN(_10063_));
 NAND4_X1 _19723_ (.A1(_10035_),
    .A2(_10044_),
    .A3(_10053_),
    .A4(_10063_),
    .ZN(_10064_));
 NOR2_X2 _19724_ (.A1(_10030_),
    .A2(_10064_),
    .ZN(_10065_));
 XOR2_X1 _19725_ (.A(_09986_),
    .B(_10065_),
    .Z(_10066_));
 XNOR2_X1 _19726_ (.A(_09915_),
    .B(_10066_),
    .ZN(_10067_));
 XNOR2_X1 _19727_ (.A(_09684_),
    .B(_08887_),
    .ZN(_10068_));
 OAI21_X1 _19728_ (.A(_05555_),
    .B1(_05152_),
    .B2(_04976_),
    .ZN(_10069_));
 INV_X1 _19729_ (.A(_05085_),
    .ZN(_10070_));
 OAI21_X1 _19730_ (.A(_10069_),
    .B1(_10070_),
    .B2(_09515_),
    .ZN(_10071_));
 NAND2_X1 _19731_ (.A1(_05555_),
    .A2(_05412_),
    .ZN(_10072_));
 OAI21_X1 _19732_ (.A(_10072_),
    .B1(_09515_),
    .B2(_06237_),
    .ZN(_10073_));
 AND2_X1 _19733_ (.A1(_05555_),
    .A2(_09505_),
    .ZN(_10074_));
 NOR4_X2 _19734_ (.A1(_10071_),
    .A2(_10073_),
    .A3(_09519_),
    .A4(_10074_),
    .ZN(_10075_));
 BUF_X4 _19735_ (.A(_04275_),
    .Z(_10076_));
 OAI211_X2 _19736_ (.A(_05357_),
    .B(_05500_),
    .C1(_10076_),
    .C2(_05764_),
    .ZN(_10077_));
 AND2_X2 _19737_ (.A1(_04625_),
    .A2(_04373_),
    .ZN(_10078_));
 OAI21_X1 _19738_ (.A(_05357_),
    .B1(_09743_),
    .B2(_10078_),
    .ZN(_10079_));
 AND4_X1 _19739_ (.A1(_09504_),
    .A2(_10075_),
    .A3(_10077_),
    .A4(_10079_),
    .ZN(_10080_));
 AND2_X1 _19740_ (.A1(_04592_),
    .A2(_05753_),
    .ZN(_10081_));
 OAI21_X1 _19741_ (.A(_05489_),
    .B1(_09507_),
    .B2(_10081_),
    .ZN(_10082_));
 INV_X1 _19742_ (.A(_09687_),
    .ZN(_10083_));
 NAND2_X1 _19743_ (.A1(_05143_),
    .A2(_05621_),
    .ZN(_10084_));
 BUF_X4 _19744_ (.A(_05143_),
    .Z(_10085_));
 NAND2_X1 _19745_ (.A1(_10085_),
    .A2(_04921_),
    .ZN(_10086_));
 AND3_X1 _19746_ (.A1(_10083_),
    .A2(_10084_),
    .A3(_10086_),
    .ZN(_10087_));
 OAI21_X1 _19747_ (.A(_05489_),
    .B1(_04538_),
    .B2(_09692_),
    .ZN(_10088_));
 OAI21_X1 _19748_ (.A(_10085_),
    .B1(_05037_),
    .B2(_06380_),
    .ZN(_10089_));
 AND4_X1 _19749_ (.A1(_10082_),
    .A2(_10087_),
    .A3(_10088_),
    .A4(_10089_),
    .ZN(_10090_));
 NAND2_X1 _19750_ (.A1(_04483_),
    .A2(_04855_),
    .ZN(_10091_));
 AND3_X1 _19751_ (.A1(_04461_),
    .A2(_04187_),
    .A3(_04165_),
    .ZN(_10092_));
 AND4_X1 _19752_ (.A1(_04779_),
    .A2(_04165_),
    .A3(_04647_),
    .A4(_04187_),
    .ZN(_10093_));
 NOR2_X1 _19753_ (.A1(_10092_),
    .A2(_10093_),
    .ZN(_10094_));
 NAND2_X1 _19754_ (.A1(_04483_),
    .A2(_05180_),
    .ZN(_10095_));
 AND4_X1 _19755_ (.A1(_04319_),
    .A2(_10091_),
    .A3(_10094_),
    .A4(_10095_),
    .ZN(_10096_));
 OAI21_X1 _19756_ (.A(_09444_),
    .B1(_04538_),
    .B2(_05200_),
    .ZN(_10097_));
 OAI211_X2 _19757_ (.A(_09444_),
    .B(_09441_),
    .C1(_05907_),
    .C2(_04647_),
    .ZN(_10098_));
 AND4_X1 _19758_ (.A1(_04691_),
    .A2(_10096_),
    .A3(_10097_),
    .A4(_10098_),
    .ZN(_10099_));
 AND2_X1 _19759_ (.A1(_09507_),
    .A2(_04757_),
    .ZN(_10100_));
 INV_X1 _19760_ (.A(_10100_),
    .ZN(_10101_));
 OAI21_X1 _19761_ (.A(_09464_),
    .B1(_05188_),
    .B2(_05335_),
    .ZN(_10102_));
 OAI21_X1 _19762_ (.A(_04768_),
    .B1(_05709_),
    .B2(_05412_),
    .ZN(_10103_));
 NAND2_X1 _19763_ (.A1(_04855_),
    .A2(_09464_),
    .ZN(_10104_));
 AND4_X1 _19764_ (.A1(_10101_),
    .A2(_10102_),
    .A3(_10103_),
    .A4(_10104_),
    .ZN(_10105_));
 NAND4_X4 _19765_ (.A1(_10080_),
    .A2(_10090_),
    .A3(_10099_),
    .A4(_10105_),
    .ZN(_10106_));
 NAND4_X1 _19766_ (.A1(_05863_),
    .A2(_05522_),
    .A3(_05467_),
    .A4(_05500_),
    .ZN(_10107_));
 NAND2_X1 _19767_ (.A1(_05841_),
    .A2(_04976_),
    .ZN(_10108_));
 NOR2_X1 _19768_ (.A1(_05819_),
    .A2(_09754_),
    .ZN(_10109_));
 AND2_X1 _19769_ (.A1(_09472_),
    .A2(_05808_),
    .ZN(_10110_));
 INV_X1 _19770_ (.A(_10110_),
    .ZN(_10111_));
 AND4_X1 _19771_ (.A1(_10108_),
    .A2(_10109_),
    .A3(_09431_),
    .A4(_10111_),
    .ZN(_10112_));
 OAI211_X2 _19772_ (.A(_05940_),
    .B(_09468_),
    .C1(_10076_),
    .C2(_05764_),
    .ZN(_10113_));
 AND4_X1 _19773_ (.A1(_04275_),
    .A2(_05676_),
    .A3(_04833_),
    .A4(_05467_),
    .ZN(_10114_));
 AOI211_X4 _19774_ (.A(_10114_),
    .B(_09418_),
    .C1(_05940_),
    .C2(_09689_),
    .ZN(_10115_));
 AND4_X1 _19775_ (.A1(_10107_),
    .A2(_10112_),
    .A3(_10113_),
    .A4(_10115_),
    .ZN(_10116_));
 AND2_X1 _19776_ (.A1(_05152_),
    .A2(_06435_),
    .ZN(_10117_));
 AND2_X1 _19777_ (.A1(_09473_),
    .A2(_06435_),
    .ZN(_10118_));
 AND2_X2 _19778_ (.A1(_09743_),
    .A2(_06424_),
    .ZN(_10119_));
 AND3_X1 _19779_ (.A1(_06424_),
    .A2(_04494_),
    .A3(_05269_),
    .ZN(_10120_));
 NOR4_X1 _19780_ (.A1(_10117_),
    .A2(_10118_),
    .A3(_10119_),
    .A4(_10120_),
    .ZN(_10121_));
 OAI21_X1 _19781_ (.A(_06446_),
    .B1(_05984_),
    .B2(_04549_),
    .ZN(_10122_));
 OAI211_X2 _19782_ (.A(_06446_),
    .B(_09468_),
    .C1(_04494_),
    .C2(_04647_),
    .ZN(_10123_));
 OAI21_X1 _19783_ (.A(_06303_),
    .B1(_05056_),
    .B2(_05180_),
    .ZN(_10124_));
 OAI211_X2 _19784_ (.A(_06303_),
    .B(_05269_),
    .C1(_05511_),
    .C2(_05198_),
    .ZN(_10125_));
 OAI211_X2 _19785_ (.A(_06215_),
    .B(_04779_),
    .C1(_05907_),
    .C2(_04395_),
    .ZN(_10126_));
 OAI21_X1 _19786_ (.A(_06303_),
    .B1(_04855_),
    .B2(_04921_),
    .ZN(_10127_));
 AND4_X1 _19787_ (.A1(_10124_),
    .A2(_10125_),
    .A3(_10126_),
    .A4(_10127_),
    .ZN(_10128_));
 AND4_X1 _19788_ (.A1(_10121_),
    .A2(_10122_),
    .A3(_10123_),
    .A4(_10128_),
    .ZN(_10129_));
 NAND2_X1 _19789_ (.A1(_09516_),
    .A2(_05346_),
    .ZN(_10130_));
 OAI21_X1 _19790_ (.A(_09491_),
    .B1(_10130_),
    .B2(_05709_),
    .ZN(_10131_));
 AND2_X2 _19791_ (.A1(_06347_),
    .A2(_05456_),
    .ZN(_10132_));
 INV_X1 _19792_ (.A(_10132_),
    .ZN(_10133_));
 NAND3_X1 _19793_ (.A1(_10131_),
    .A2(_10133_),
    .A3(_09742_),
    .ZN(_10134_));
 OAI21_X1 _19794_ (.A(_09482_),
    .B1(_09692_),
    .B2(_05313_),
    .ZN(_10135_));
 NAND2_X1 _19795_ (.A1(_05335_),
    .A2(_09482_),
    .ZN(_10136_));
 NAND2_X1 _19796_ (.A1(_10135_),
    .A2(_10136_),
    .ZN(_10137_));
 AOI21_X1 _19797_ (.A(_09748_),
    .B1(_10070_),
    .B2(_05731_),
    .ZN(_10138_));
 NOR2_X1 _19798_ (.A1(_09748_),
    .A2(_05214_),
    .ZN(_10139_));
 OR2_X1 _19799_ (.A1(_10139_),
    .A2(_09485_),
    .ZN(_10140_));
 NOR4_X2 _19800_ (.A1(_10134_),
    .A2(_10137_),
    .A3(_10138_),
    .A4(_10140_),
    .ZN(_10141_));
 OAI21_X1 _19801_ (.A(_06061_),
    .B1(_05335_),
    .B2(_09717_),
    .ZN(_10142_));
 OAI21_X1 _19802_ (.A(_05775_),
    .B1(_09434_),
    .B2(_09441_),
    .ZN(_10143_));
 OAI21_X1 _19803_ (.A(_06061_),
    .B1(_09751_),
    .B2(_09505_),
    .ZN(_10144_));
 OAI21_X1 _19804_ (.A(_05775_),
    .B1(_05412_),
    .B2(_04549_),
    .ZN(_10145_));
 AND4_X1 _19805_ (.A1(_10142_),
    .A2(_10143_),
    .A3(_10144_),
    .A4(_10145_),
    .ZN(_10146_));
 NAND4_X2 _19806_ (.A1(_10116_),
    .A2(_10129_),
    .A3(_10141_),
    .A4(_10146_),
    .ZN(_10147_));
 NOR2_X4 _19807_ (.A1(_10106_),
    .A2(_10147_),
    .ZN(_10148_));
 XNOR2_X1 _19808_ (.A(_10068_),
    .B(_10148_),
    .ZN(_10149_));
 XNOR2_X1 _19809_ (.A(_10067_),
    .B(_10149_),
    .ZN(_10150_));
 XNOR2_X1 _19810_ (.A(_10150_),
    .B(_17169_),
    .ZN(_10151_));
 MUX2_X1 _19811_ (.A(_09842_),
    .B(_10151_),
    .S(_09100_),
    .Z(_00727_));
 XOR2_X1 _19812_ (.A(_17170_),
    .B(_17084_),
    .Z(_10152_));
 XNOR2_X1 _19813_ (.A(_09986_),
    .B(_08887_),
    .ZN(_10153_));
 AND2_X1 _19814_ (.A1(_04483_),
    .A2(_09692_),
    .ZN(_10154_));
 INV_X1 _19815_ (.A(_10154_),
    .ZN(_10155_));
 AND2_X1 _19816_ (.A1(_04209_),
    .A2(_09743_),
    .ZN(_10156_));
 AOI211_X2 _19817_ (.A(_09456_),
    .B(_10156_),
    .C1(_04483_),
    .C2(_04855_),
    .ZN(_10157_));
 NAND2_X1 _19818_ (.A1(_05918_),
    .A2(_04483_),
    .ZN(_10158_));
 INV_X1 _19819_ (.A(_09444_),
    .ZN(_10159_));
 NOR2_X1 _19820_ (.A1(_10159_),
    .A2(_05028_),
    .ZN(_10160_));
 AND3_X1 _19821_ (.A1(_09444_),
    .A2(_04647_),
    .A3(_05269_),
    .ZN(_10161_));
 NOR4_X1 _19822_ (.A1(_10160_),
    .A2(_09702_),
    .A3(_09448_),
    .A4(_10161_),
    .ZN(_10162_));
 AND4_X1 _19823_ (.A1(_10155_),
    .A2(_10157_),
    .A3(_10158_),
    .A4(_10162_),
    .ZN(_10163_));
 AND2_X1 _19824_ (.A1(_05143_),
    .A2(_05056_),
    .ZN(_10164_));
 INV_X1 _19825_ (.A(_10164_),
    .ZN(_10165_));
 OAI21_X1 _19826_ (.A(_10085_),
    .B1(_09692_),
    .B2(_05984_),
    .ZN(_10166_));
 OAI211_X2 _19827_ (.A(_10085_),
    .B(_09441_),
    .C1(_05511_),
    .C2(_05764_),
    .ZN(_10167_));
 NAND4_X1 _19828_ (.A1(_10165_),
    .A2(_10084_),
    .A3(_10166_),
    .A4(_10167_),
    .ZN(_10168_));
 AOI21_X1 _19829_ (.A(_09512_),
    .B1(_10070_),
    .B2(_05731_),
    .ZN(_10169_));
 AND3_X2 _19830_ (.A1(_05489_),
    .A2(_04669_),
    .A3(_05269_),
    .ZN(_10170_));
 NAND2_X1 _19831_ (.A1(_05390_),
    .A2(_04417_),
    .ZN(_10171_));
 NAND2_X1 _19832_ (.A1(_05390_),
    .A2(_05180_),
    .ZN(_10172_));
 OAI211_X2 _19833_ (.A(_10171_),
    .B(_10172_),
    .C1(_09512_),
    .C2(_05995_),
    .ZN(_10173_));
 NOR4_X1 _19834_ (.A1(_10168_),
    .A2(_10169_),
    .A3(_10170_),
    .A4(_10173_),
    .ZN(_10174_));
 OAI211_X2 _19835_ (.A(_05610_),
    .B(_05643_),
    .C1(_10072_),
    .C2(_10076_),
    .ZN(_10175_));
 OAI21_X1 _19836_ (.A(_05357_),
    .B1(_05056_),
    .B2(_05335_),
    .ZN(_10176_));
 NAND3_X1 _19837_ (.A1(_09692_),
    .A2(_04329_),
    .A3(_05202_),
    .ZN(_10177_));
 NAND3_X1 _19838_ (.A1(_09506_),
    .A2(_10176_),
    .A3(_10177_),
    .ZN(_10178_));
 AND2_X1 _19839_ (.A1(_05599_),
    .A2(_05152_),
    .ZN(_10179_));
 NOR4_X1 _19840_ (.A1(_10175_),
    .A2(_10178_),
    .A3(_10074_),
    .A4(_10179_),
    .ZN(_10180_));
 NAND2_X1 _19841_ (.A1(_05918_),
    .A2(_09464_),
    .ZN(_10181_));
 OAI21_X1 _19842_ (.A(_04768_),
    .B1(_09689_),
    .B2(_09441_),
    .ZN(_10182_));
 OAI211_X2 _19843_ (.A(_04768_),
    .B(_04669_),
    .C1(_09468_),
    .C2(_05500_),
    .ZN(_10183_));
 OAI21_X1 _19844_ (.A(_09464_),
    .B1(_09743_),
    .B2(_04921_),
    .ZN(_10184_));
 AND4_X1 _19845_ (.A1(_10181_),
    .A2(_10182_),
    .A3(_10183_),
    .A4(_10184_),
    .ZN(_10185_));
 NAND4_X2 _19846_ (.A1(_10163_),
    .A2(_10174_),
    .A3(_10180_),
    .A4(_10185_),
    .ZN(_10186_));
 AND2_X1 _19847_ (.A1(_05335_),
    .A2(_06424_),
    .ZN(_10187_));
 AOI211_X4 _19848_ (.A(_10187_),
    .B(_10119_),
    .C1(_09441_),
    .C2(_06435_),
    .ZN(_10188_));
 INV_X1 _19849_ (.A(_09479_),
    .ZN(_10189_));
 OAI21_X1 _19850_ (.A(_06226_),
    .B1(_05037_),
    .B2(_05412_),
    .ZN(_10190_));
 AND4_X1 _19851_ (.A1(_06336_),
    .A2(_10188_),
    .A3(_10189_),
    .A4(_10190_),
    .ZN(_10191_));
 NAND4_X1 _19852_ (.A1(_09490_),
    .A2(_09744_),
    .A3(_10133_),
    .A4(_09742_),
    .ZN(_10192_));
 AND2_X1 _19853_ (.A1(_09452_),
    .A2(_06149_),
    .ZN(_10193_));
 AND2_X1 _19854_ (.A1(_06149_),
    .A2(_05313_),
    .ZN(_10194_));
 OR2_X1 _19855_ (.A1(_10193_),
    .A2(_10194_),
    .ZN(_10195_));
 NAND3_X1 _19856_ (.A1(_06391_),
    .A2(_09438_),
    .A3(_06127_),
    .ZN(_10196_));
 OAI211_X2 _19857_ (.A(_10196_),
    .B(_09738_),
    .C1(_05194_),
    .C2(_06358_),
    .ZN(_10197_));
 NOR4_X1 _19858_ (.A1(_10192_),
    .A2(_09741_),
    .A3(_10195_),
    .A4(_10197_),
    .ZN(_10198_));
 OAI21_X1 _19859_ (.A(_06061_),
    .B1(_04658_),
    .B2(_09505_),
    .ZN(_10199_));
 OAI21_X1 _19860_ (.A(_05775_),
    .B1(_05056_),
    .B2(_09692_),
    .ZN(_10200_));
 OAI21_X1 _19861_ (.A(_05775_),
    .B1(_09701_),
    .B2(_09505_),
    .ZN(_10201_));
 AND4_X1 _19862_ (.A1(_09416_),
    .A2(_10199_),
    .A3(_10200_),
    .A4(_10201_),
    .ZN(_10202_));
 INV_X2 _19863_ (.A(_09434_),
    .ZN(_10203_));
 INV_X1 _19864_ (.A(_09507_),
    .ZN(_10204_));
 AOI21_X1 _19865_ (.A(_05962_),
    .B1(_10203_),
    .B2(_10204_),
    .ZN(_10205_));
 NAND2_X1 _19866_ (.A1(_05841_),
    .A2(_06391_),
    .ZN(_10206_));
 NAND3_X1 _19867_ (.A1(_09755_),
    .A2(_09430_),
    .A3(_10206_),
    .ZN(_10207_));
 NAND2_X1 _19868_ (.A1(_05852_),
    .A2(_05874_),
    .ZN(_10208_));
 NOR2_X1 _19869_ (.A1(_06402_),
    .A2(_05962_),
    .ZN(_10209_));
 NOR4_X1 _19870_ (.A1(_10205_),
    .A2(_10207_),
    .A3(_10208_),
    .A4(_10209_),
    .ZN(_10210_));
 NAND4_X1 _19871_ (.A1(_10191_),
    .A2(_10198_),
    .A3(_10202_),
    .A4(_10210_),
    .ZN(_10211_));
 NOR2_X4 _19872_ (.A1(_10186_),
    .A2(_10211_),
    .ZN(_10212_));
 XNOR2_X1 _19873_ (.A(_10153_),
    .B(_10212_),
    .ZN(_10213_));
 AND4_X1 _19874_ (.A1(_08830_),
    .A2(_08605_),
    .A3(_08563_),
    .A4(_08754_),
    .ZN(_10214_));
 AOI211_X2 _19875_ (.A(_10214_),
    .B(_09639_),
    .C1(_08760_),
    .C2(_08673_),
    .ZN(_10215_));
 AND2_X1 _19876_ (.A1(_08586_),
    .A2(_16783_),
    .ZN(_10216_));
 OAI21_X1 _19877_ (.A(_08748_),
    .B1(_08695_),
    .B2(_10216_),
    .ZN(_10217_));
 OAI21_X1 _19878_ (.A(_08748_),
    .B1(_08637_),
    .B2(_08674_),
    .ZN(_10218_));
 AND4_X2 _19879_ (.A1(_08811_),
    .A2(_10215_),
    .A3(_10217_),
    .A4(_10218_),
    .ZN(_10219_));
 AOI21_X1 _19880_ (.A(_09266_),
    .B1(_08758_),
    .B2(_08737_),
    .ZN(_10220_));
 AOI211_X2 _19881_ (.A(_08775_),
    .B(_10220_),
    .C1(_08789_),
    .C2(_08774_),
    .ZN(_10221_));
 OAI21_X1 _19882_ (.A(_09633_),
    .B1(_08860_),
    .B2(_08578_),
    .ZN(_10222_));
 NAND4_X1 _19883_ (.A1(_08620_),
    .A2(_08585_),
    .A3(_08649_),
    .A4(_08754_),
    .ZN(_10223_));
 OAI21_X1 _19884_ (.A(_09633_),
    .B1(_08724_),
    .B2(_08770_),
    .ZN(_10224_));
 AND4_X1 _19885_ (.A1(_10221_),
    .A2(_10222_),
    .A3(_10223_),
    .A4(_10224_),
    .ZN(_10225_));
 OAI21_X1 _19886_ (.A(_08741_),
    .B1(_08800_),
    .B2(_08779_),
    .ZN(_10226_));
 OAI21_X1 _19887_ (.A(_08741_),
    .B1(_08810_),
    .B2(_08669_),
    .ZN(_10227_));
 NAND2_X1 _19888_ (.A1(_10226_),
    .A2(_10227_),
    .ZN(_10228_));
 AND2_X1 _19889_ (.A1(_08715_),
    .A2(_08779_),
    .ZN(_10229_));
 NOR4_X1 _19890_ (.A1(_08738_),
    .A2(_10228_),
    .A3(_09225_),
    .A4(_10229_),
    .ZN(_10230_));
 OAI21_X1 _19891_ (.A(_08731_),
    .B1(_08750_),
    .B2(_08815_),
    .ZN(_10231_));
 OAI21_X1 _19892_ (.A(_08721_),
    .B1(_08637_),
    .B2(_08860_),
    .ZN(_10232_));
 AND4_X1 _19893_ (.A1(_08727_),
    .A2(_10231_),
    .A3(_09919_),
    .A4(_10232_),
    .ZN(_10233_));
 NAND4_X1 _19894_ (.A1(_10219_),
    .A2(_10225_),
    .A3(_10230_),
    .A4(_10233_),
    .ZN(_10234_));
 AND2_X2 _19895_ (.A1(_08703_),
    .A2(_08810_),
    .ZN(_10235_));
 INV_X1 _19896_ (.A(_10235_),
    .ZN(_10236_));
 NAND4_X1 _19897_ (.A1(_08763_),
    .A2(_08762_),
    .A3(_08675_),
    .A4(_08620_),
    .ZN(_10237_));
 OAI21_X1 _19898_ (.A(_08704_),
    .B1(_08662_),
    .B2(_08681_),
    .ZN(_10238_));
 AND4_X1 _19899_ (.A1(_09965_),
    .A2(_10236_),
    .A3(_10237_),
    .A4(_10238_),
    .ZN(_10239_));
 AND4_X1 _19900_ (.A1(_08592_),
    .A2(_08656_),
    .A3(_08753_),
    .A4(_08638_),
    .ZN(_10240_));
 AND2_X1 _19901_ (.A1(_08573_),
    .A2(_08657_),
    .ZN(_10241_));
 AOI211_X2 _19902_ (.A(_10240_),
    .B(_10241_),
    .C1(_08767_),
    .C2(_08658_),
    .ZN(_10242_));
 OAI21_X1 _19903_ (.A(_08658_),
    .B1(_08681_),
    .B2(_08633_),
    .ZN(_10243_));
 AND4_X1 _19904_ (.A1(_08838_),
    .A2(_10239_),
    .A3(_10242_),
    .A4(_10243_),
    .ZN(_10244_));
 NAND2_X1 _19905_ (.A1(_08810_),
    .A2(_08679_),
    .ZN(_10245_));
 OAI211_X2 _19906_ (.A(_08688_),
    .B(_10245_),
    .C1(_08820_),
    .C2(_08690_),
    .ZN(_10246_));
 NAND3_X1 _19907_ (.A1(_08853_),
    .A2(_08701_),
    .A3(_08699_),
    .ZN(_10247_));
 AOI21_X1 _19908_ (.A(_08855_),
    .B1(_08873_),
    .B2(_08663_),
    .ZN(_10248_));
 NOR4_X1 _19909_ (.A1(_10246_),
    .A2(_10247_),
    .A3(_10248_),
    .A4(_09271_),
    .ZN(_10249_));
 OAI211_X2 _19910_ (.A(_08608_),
    .B(_08649_),
    .C1(_08585_),
    .C2(_08706_),
    .ZN(_10250_));
 OAI21_X1 _19911_ (.A(_08608_),
    .B1(_08662_),
    .B2(_08631_),
    .ZN(_10251_));
 NAND2_X1 _19912_ (.A1(_08607_),
    .A2(_08669_),
    .ZN(_10252_));
 NAND2_X1 _19913_ (.A1(_08789_),
    .A2(_08608_),
    .ZN(_10253_));
 NAND4_X1 _19914_ (.A1(_10250_),
    .A2(_10251_),
    .A3(_10252_),
    .A4(_10253_),
    .ZN(_10254_));
 NAND2_X1 _19915_ (.A1(_09280_),
    .A2(_08575_),
    .ZN(_10255_));
 INV_X1 _19916_ (.A(_10255_),
    .ZN(_10256_));
 AND3_X1 _19917_ (.A1(_08575_),
    .A2(_08592_),
    .A3(_08649_),
    .ZN(_10257_));
 AND2_X1 _19918_ (.A1(_08582_),
    .A2(_08592_),
    .ZN(_10258_));
 NAND2_X1 _19919_ (.A1(_10258_),
    .A2(_08575_),
    .ZN(_10259_));
 NAND2_X1 _19920_ (.A1(_09662_),
    .A2(_10259_),
    .ZN(_10260_));
 NOR4_X1 _19921_ (.A1(_10254_),
    .A2(_10256_),
    .A3(_10257_),
    .A4(_10260_),
    .ZN(_10261_));
 NAND3_X1 _19922_ (.A1(_08622_),
    .A2(_08614_),
    .A3(_08610_),
    .ZN(_10262_));
 OAI21_X1 _19923_ (.A(_08645_),
    .B1(_08789_),
    .B2(_08632_),
    .ZN(_10263_));
 OAI211_X2 _19924_ (.A(_08640_),
    .B(_08649_),
    .C1(_08584_),
    .C2(_08706_),
    .ZN(_10264_));
 AND2_X1 _19925_ (.A1(_10263_),
    .A2(_10264_),
    .ZN(_10265_));
 OAI21_X1 _19926_ (.A(_08622_),
    .B1(_09243_),
    .B2(_08624_),
    .ZN(_10266_));
 OAI21_X1 _19927_ (.A(_08622_),
    .B1(_08681_),
    .B2(_08633_),
    .ZN(_10267_));
 AND4_X1 _19928_ (.A1(_10262_),
    .A2(_10265_),
    .A3(_10266_),
    .A4(_10267_),
    .ZN(_10268_));
 NAND4_X1 _19929_ (.A1(_10244_),
    .A2(_10249_),
    .A3(_10261_),
    .A4(_10268_),
    .ZN(_10269_));
 NOR2_X2 _19930_ (.A1(_10234_),
    .A2(_10269_),
    .ZN(_10270_));
 OAI221_X1 _19931_ (.A(_09203_),
    .B1(_07488_),
    .B2(_09140_),
    .C1(_08069_),
    .C2(_09204_),
    .ZN(_10271_));
 AOI21_X1 _19932_ (.A(_09545_),
    .B1(_09189_),
    .B2(_09582_),
    .ZN(_10272_));
 NOR2_X1 _19933_ (.A1(_08553_),
    .A2(_09545_),
    .ZN(_10273_));
 NOR4_X1 _19934_ (.A1(_10271_),
    .A2(_08548_),
    .A3(_10272_),
    .A4(_10273_),
    .ZN(_10274_));
 OAI21_X1 _19935_ (.A(_08299_),
    .B1(_08556_),
    .B2(_08532_),
    .ZN(_10275_));
 OAI21_X1 _19936_ (.A(_08299_),
    .B1(_09138_),
    .B2(_08354_),
    .ZN(_10276_));
 OAI211_X2 _19937_ (.A(_07414_),
    .B(_16791_),
    .C1(_16790_),
    .C2(_06743_),
    .ZN(_10277_));
 AND4_X1 _19938_ (.A1(_08534_),
    .A2(_10275_),
    .A3(_10276_),
    .A4(_10277_),
    .ZN(_10278_));
 AND2_X1 _19939_ (.A1(_09575_),
    .A2(_09576_),
    .ZN(_10279_));
 NAND3_X1 _19940_ (.A1(_07675_),
    .A2(_07883_),
    .A3(_06842_),
    .ZN(_10280_));
 NAND3_X1 _19941_ (.A1(_07631_),
    .A2(_07883_),
    .A3(_06842_),
    .ZN(_10281_));
 NAND2_X1 _19942_ (.A1(_10280_),
    .A2(_10281_),
    .ZN(_10282_));
 AND2_X4 _19943_ (.A1(_08550_),
    .A2(_07565_),
    .ZN(_10283_));
 NOR2_X1 _19944_ (.A1(_10282_),
    .A2(_10283_),
    .ZN(_10284_));
 AND2_X1 _19945_ (.A1(_07062_),
    .A2(_07029_),
    .ZN(_10285_));
 OAI21_X1 _19946_ (.A(_07117_),
    .B1(_10285_),
    .B2(_07565_),
    .ZN(_10286_));
 OAI21_X1 _19947_ (.A(_08550_),
    .B1(_07751_),
    .B2(_09166_),
    .ZN(_10287_));
 AND4_X1 _19948_ (.A1(_10279_),
    .A2(_10284_),
    .A3(_10286_),
    .A4(_10287_),
    .ZN(_10288_));
 OAI21_X1 _19949_ (.A(_07326_),
    .B1(_07927_),
    .B2(_09106_),
    .ZN(_10289_));
 OAI21_X1 _19950_ (.A(_09192_),
    .B1(_07675_),
    .B2(_08310_),
    .ZN(_10290_));
 OAI21_X1 _19951_ (.A(_09192_),
    .B1(_09144_),
    .B2(_09106_),
    .ZN(_10291_));
 AND4_X1 _19952_ (.A1(_09185_),
    .A2(_10289_),
    .A3(_10290_),
    .A4(_10291_),
    .ZN(_10292_));
 NAND4_X1 _19953_ (.A1(_10274_),
    .A2(_10278_),
    .A3(_10288_),
    .A4(_10292_),
    .ZN(_10293_));
 NAND2_X4 _19954_ (.A1(_07905_),
    .A2(_08310_),
    .ZN(_10294_));
 OAI21_X1 _19955_ (.A(_07894_),
    .B1(_08500_),
    .B2(_09131_),
    .ZN(_10295_));
 OAI21_X1 _19956_ (.A(_07894_),
    .B1(_08025_),
    .B2(_07205_),
    .ZN(_10296_));
 NAND3_X1 _19957_ (.A1(_07084_),
    .A2(_07949_),
    .A3(_07238_),
    .ZN(_10297_));
 AND4_X1 _19958_ (.A1(_10294_),
    .A2(_10295_),
    .A3(_10296_),
    .A4(_10297_),
    .ZN(_10298_));
 NAND2_X1 _19959_ (.A1(_07686_),
    .A2(_06611_),
    .ZN(_10299_));
 OAI21_X1 _19960_ (.A(_06611_),
    .B1(_07499_),
    .B2(_08532_),
    .ZN(_10300_));
 AND4_X1 _19961_ (.A1(_09601_),
    .A2(_10298_),
    .A3(_10299_),
    .A4(_10300_),
    .ZN(_10301_));
 OAI21_X1 _19962_ (.A(_06963_),
    .B1(_08025_),
    .B2(_07227_),
    .ZN(_10302_));
 NAND3_X1 _19963_ (.A1(_06952_),
    .A2(_08222_),
    .A3(_09145_),
    .ZN(_10303_));
 NAND2_X1 _19964_ (.A1(_06963_),
    .A2(_07675_),
    .ZN(_10304_));
 NAND2_X1 _19965_ (.A1(_06963_),
    .A2(_08201_),
    .ZN(_10305_));
 NAND4_X1 _19966_ (.A1(_10302_),
    .A2(_10303_),
    .A3(_10304_),
    .A4(_10305_),
    .ZN(_10306_));
 NAND2_X1 _19967_ (.A1(_07532_),
    .A2(_09131_),
    .ZN(_10307_));
 NAND4_X1 _19968_ (.A1(_08058_),
    .A2(_08538_),
    .A3(_08519_),
    .A4(_06897_),
    .ZN(_10308_));
 OAI211_X2 _19969_ (.A(_10307_),
    .B(_10308_),
    .C1(_07543_),
    .C2(_07370_),
    .ZN(_10309_));
 AOI21_X1 _19970_ (.A(_07543_),
    .B1(_09167_),
    .B2(_09572_),
    .ZN(_10310_));
 AND2_X4 _19971_ (.A1(_07521_),
    .A2(_09153_),
    .ZN(_10311_));
 NOR4_X1 _19972_ (.A1(_10306_),
    .A2(_10309_),
    .A3(_10310_),
    .A4(_10311_),
    .ZN(_10312_));
 NAND2_X1 _19973_ (.A1(_08190_),
    .A2(_08124_),
    .ZN(_10313_));
 NAND2_X1 _19974_ (.A1(_08190_),
    .A2(_07565_),
    .ZN(_10314_));
 OAI211_X2 _19975_ (.A(_10313_),
    .B(_10314_),
    .C1(_07370_),
    .C2(_07992_),
    .ZN(_10315_));
 NAND2_X1 _19976_ (.A1(_07675_),
    .A2(_07795_),
    .ZN(_10316_));
 NAND4_X1 _19977_ (.A1(_08058_),
    .A2(_08538_),
    .A3(_07436_),
    .A4(_08080_),
    .ZN(_10317_));
 OAI211_X2 _19978_ (.A(_10316_),
    .B(_10317_),
    .C1(_07510_),
    .C2(_09128_),
    .ZN(_10318_));
 OAI21_X1 _19979_ (.A(_10023_),
    .B1(_07992_),
    .B2(_08541_),
    .ZN(_10319_));
 NOR4_X1 _19980_ (.A1(_10315_),
    .A2(_10318_),
    .A3(_10319_),
    .A4(_09129_),
    .ZN(_10320_));
 OAI21_X1 _19981_ (.A(_07719_),
    .B1(_07861_),
    .B2(_07447_),
    .ZN(_10321_));
 OAI211_X2 _19982_ (.A(_07653_),
    .B(_07062_),
    .C1(_08396_),
    .C2(_08069_),
    .ZN(_10322_));
 OAI21_X1 _19983_ (.A(_07653_),
    .B1(_07084_),
    .B2(_09166_),
    .ZN(_10323_));
 OAI211_X2 _19984_ (.A(_07719_),
    .B(_08244_),
    .C1(_08538_),
    .C2(_07062_),
    .ZN(_10324_));
 AND4_X1 _19985_ (.A1(_10321_),
    .A2(_10322_),
    .A3(_10323_),
    .A4(_10324_),
    .ZN(_10325_));
 NAND4_X1 _19986_ (.A1(_10301_),
    .A2(_10312_),
    .A3(_10320_),
    .A4(_10325_),
    .ZN(_10326_));
 NOR2_X2 _19987_ (.A1(_10293_),
    .A2(_10326_),
    .ZN(_10327_));
 XOR2_X2 _19988_ (.A(_10270_),
    .B(_10327_),
    .Z(_10328_));
 XNOR2_X1 _19989_ (.A(_10213_),
    .B(_10328_),
    .ZN(_10329_));
 NAND2_X1 _19990_ (.A1(_08973_),
    .A2(_09325_),
    .ZN(_10330_));
 INV_X1 _19991_ (.A(_08973_),
    .ZN(_10331_));
 AOI21_X1 _19992_ (.A(_10331_),
    .B1(_09385_),
    .B2(_09371_),
    .ZN(_10332_));
 AOI21_X1 _19993_ (.A(_10332_),
    .B1(_09340_),
    .B2(_08973_),
    .ZN(_10333_));
 NAND2_X1 _19994_ (.A1(_08973_),
    .A2(_09374_),
    .ZN(_10334_));
 OAI21_X1 _19995_ (.A(_08973_),
    .B1(_08901_),
    .B2(_08987_),
    .ZN(_10335_));
 AND4_X1 _19996_ (.A1(_10330_),
    .A2(_10333_),
    .A3(_10334_),
    .A4(_10335_),
    .ZN(_10336_));
 OAI211_X2 _19997_ (.A(_09329_),
    .B(_08977_),
    .C1(_08962_),
    .C2(_09784_),
    .ZN(_10337_));
 OAI21_X1 _19998_ (.A(_09329_),
    .B1(_08910_),
    .B2(_09010_),
    .ZN(_10338_));
 AND4_X2 _19999_ (.A1(_09787_),
    .A2(_10336_),
    .A3(_10337_),
    .A4(_10338_),
    .ZN(_10339_));
 NAND2_X1 _20000_ (.A1(_09354_),
    .A2(_09344_),
    .ZN(_10340_));
 OAI211_X2 _20001_ (.A(_08921_),
    .B(_08905_),
    .C1(_09002_),
    .C2(_09331_),
    .ZN(_10341_));
 AND4_X1 _20002_ (.A1(_10340_),
    .A2(_10341_),
    .A3(_09771_),
    .A4(_09903_),
    .ZN(_10342_));
 AND2_X1 _20003_ (.A1(_09087_),
    .A2(_08907_),
    .ZN(_10343_));
 OAI21_X1 _20004_ (.A(_09326_),
    .B1(_09002_),
    .B2(_10343_),
    .ZN(_10344_));
 OAI21_X1 _20005_ (.A(_09326_),
    .B1(_09323_),
    .B2(_09374_),
    .ZN(_10345_));
 AND3_X1 _20006_ (.A1(_10342_),
    .A2(_10344_),
    .A3(_10345_),
    .ZN(_10346_));
 NAND2_X1 _20007_ (.A1(_09310_),
    .A2(_09394_),
    .ZN(_10347_));
 NAND3_X1 _20008_ (.A1(_09018_),
    .A2(_08950_),
    .A3(_08944_),
    .ZN(_10348_));
 OR2_X1 _20009_ (.A1(_09303_),
    .A2(_09350_),
    .ZN(_10349_));
 NAND4_X1 _20010_ (.A1(_09320_),
    .A2(_10347_),
    .A3(_10348_),
    .A4(_10349_),
    .ZN(_10350_));
 AND3_X1 _20011_ (.A1(_09305_),
    .A2(_09832_),
    .A3(_08918_),
    .ZN(_10351_));
 INV_X1 _20012_ (.A(_09323_),
    .ZN(_10352_));
 AOI21_X1 _20013_ (.A(_09897_),
    .B1(_10352_),
    .B2(_09066_),
    .ZN(_10353_));
 AOI21_X1 _20014_ (.A(_09897_),
    .B1(_09385_),
    .B2(_09380_),
    .ZN(_10354_));
 NOR4_X1 _20015_ (.A1(_10350_),
    .A2(_10351_),
    .A3(_10353_),
    .A4(_10354_),
    .ZN(_10355_));
 OAI21_X1 _20016_ (.A(_09789_),
    .B1(_08985_),
    .B2(_09325_),
    .ZN(_10356_));
 OAI21_X1 _20017_ (.A(_09377_),
    .B1(_08948_),
    .B2(_08919_),
    .ZN(_10357_));
 NAND2_X1 _20018_ (.A1(_09018_),
    .A2(_09377_),
    .ZN(_10358_));
 AND4_X1 _20019_ (.A1(_09003_),
    .A2(_10356_),
    .A3(_10357_),
    .A4(_10358_),
    .ZN(_10359_));
 NAND4_X1 _20020_ (.A1(_10339_),
    .A2(_10346_),
    .A3(_10355_),
    .A4(_10359_),
    .ZN(_10360_));
 NAND4_X1 _20021_ (.A1(_09057_),
    .A2(_09054_),
    .A3(_08892_),
    .A4(_08977_),
    .ZN(_10361_));
 AND2_X1 _20022_ (.A1(_09084_),
    .A2(_08919_),
    .ZN(_10362_));
 INV_X1 _20023_ (.A(_10362_),
    .ZN(_10363_));
 NAND2_X1 _20024_ (.A1(_10363_),
    .A2(_09295_),
    .ZN(_10364_));
 AND2_X1 _20025_ (.A1(_09084_),
    .A2(_08899_),
    .ZN(_10365_));
 AND2_X4 _20026_ (.A1(_09084_),
    .A2(_08969_),
    .ZN(_10366_));
 NOR4_X1 _20027_ (.A1(_10364_),
    .A2(_10365_),
    .A3(_10366_),
    .A4(_09777_),
    .ZN(_10367_));
 OAI211_X2 _20028_ (.A(_09797_),
    .B(_09355_),
    .C1(_08962_),
    .C2(_09784_),
    .ZN(_10368_));
 AND4_X1 _20029_ (.A1(_08908_),
    .A2(_09057_),
    .A3(_08892_),
    .A4(_08932_),
    .ZN(_10369_));
 AND2_X1 _20030_ (.A1(_09078_),
    .A2(_09002_),
    .ZN(_10370_));
 AOI211_X2 _20031_ (.A(_10369_),
    .B(_10370_),
    .C1(_09081_),
    .C2(_09900_),
    .ZN(_10371_));
 AND4_X1 _20032_ (.A1(_10361_),
    .A2(_10367_),
    .A3(_10368_),
    .A4(_10371_),
    .ZN(_10372_));
 OAI211_X2 _20033_ (.A(_09382_),
    .B(_09087_),
    .C1(_09054_),
    .C2(_09784_),
    .ZN(_10373_));
 OAI211_X2 _20034_ (.A(_09382_),
    .B(_08916_),
    .C1(_09017_),
    .C2(_08918_),
    .ZN(_10374_));
 OAI21_X1 _20035_ (.A(_09382_),
    .B1(_09051_),
    .B2(_08926_),
    .ZN(_10375_));
 AND4_X1 _20036_ (.A1(_09384_),
    .A2(_10373_),
    .A3(_10374_),
    .A4(_10375_),
    .ZN(_10376_));
 AND2_X4 _20037_ (.A1(_09039_),
    .A2(_08923_),
    .ZN(_10377_));
 INV_X4 _20038_ (.A(_10377_),
    .ZN(_10378_));
 NAND3_X1 _20039_ (.A1(_09039_),
    .A2(_09017_),
    .A3(_08916_),
    .ZN(_10379_));
 OAI211_X2 _20040_ (.A(_10378_),
    .B(_10379_),
    .C1(_09070_),
    .C2(_09386_),
    .ZN(_10380_));
 NAND2_X1 _20041_ (.A1(_09318_),
    .A2(_09039_),
    .ZN(_10381_));
 NAND2_X1 _20042_ (.A1(_09040_),
    .A2(_10381_),
    .ZN(_10382_));
 NOR4_X1 _20043_ (.A1(_10380_),
    .A2(_10382_),
    .A3(_09402_),
    .A4(_09813_),
    .ZN(_10383_));
 OAI21_X1 _20044_ (.A(_09392_),
    .B1(_08985_),
    .B2(_08955_),
    .ZN(_10384_));
 OAI21_X1 _20045_ (.A(_09392_),
    .B1(_09378_),
    .B2(_09394_),
    .ZN(_10385_));
 OAI21_X1 _20046_ (.A(_09392_),
    .B1(_09318_),
    .B2(_08901_),
    .ZN(_10386_));
 OAI21_X1 _20047_ (.A(_09016_),
    .B1(_09018_),
    .B2(_09331_),
    .ZN(_10387_));
 AND4_X1 _20048_ (.A1(_10384_),
    .A2(_10385_),
    .A3(_10386_),
    .A4(_10387_),
    .ZN(_10388_));
 OAI21_X1 _20049_ (.A(_09346_),
    .B1(_08948_),
    .B2(_08919_),
    .ZN(_10389_));
 NAND2_X1 _20050_ (.A1(_09346_),
    .A2(_09331_),
    .ZN(_10390_));
 NAND2_X1 _20051_ (.A1(_08985_),
    .A2(_09346_),
    .ZN(_10391_));
 AND4_X1 _20052_ (.A1(_09047_),
    .A2(_10389_),
    .A3(_10390_),
    .A4(_10391_),
    .ZN(_10392_));
 AND4_X1 _20053_ (.A1(_10376_),
    .A2(_10383_),
    .A3(_10388_),
    .A4(_10392_),
    .ZN(_10393_));
 AND2_X1 _20054_ (.A1(_09347_),
    .A2(_09074_),
    .ZN(_10394_));
 AND2_X1 _20055_ (.A1(_08948_),
    .A2(_09074_),
    .ZN(_10395_));
 NOR4_X1 _20056_ (.A1(_10394_),
    .A2(_09844_),
    .A3(_09845_),
    .A4(_10395_),
    .ZN(_10396_));
 AND2_X1 _20057_ (.A1(_09058_),
    .A2(_08932_),
    .ZN(_10397_));
 AND2_X1 _20058_ (.A1(_09330_),
    .A2(_09325_),
    .ZN(_10398_));
 NOR4_X1 _20059_ (.A1(_09059_),
    .A2(_10397_),
    .A3(_09851_),
    .A4(_10398_),
    .ZN(_10399_));
 NAND4_X2 _20060_ (.A1(_10372_),
    .A2(_10393_),
    .A3(_10396_),
    .A4(_10399_),
    .ZN(_10400_));
 NOR2_X4 _20061_ (.A1(_10360_),
    .A2(_10400_),
    .ZN(_10401_));
 XOR2_X1 _20062_ (.A(_10401_),
    .B(_09093_),
    .Z(_10402_));
 XNOR2_X1 _20063_ (.A(_10329_),
    .B(_10402_),
    .ZN(_10403_));
 XNOR2_X1 _20064_ (.A(_10403_),
    .B(_17170_),
    .ZN(_10404_));
 MUX2_X1 _20065_ (.A(_10152_),
    .B(_10404_),
    .S(_09100_),
    .Z(_00728_));
 XOR2_X1 _20066_ (.A(_17171_),
    .B(_17095_),
    .Z(_10405_));
 NOR4_X1 _20067_ (.A1(_10160_),
    .A2(_04406_),
    .A3(_09448_),
    .A4(_09449_),
    .ZN(_10406_));
 INV_X1 _20068_ (.A(_09459_),
    .ZN(_10407_));
 AND2_X4 _20069_ (.A1(_06391_),
    .A2(_05009_),
    .ZN(_10408_));
 INV_X1 _20070_ (.A(_04998_),
    .ZN(_10409_));
 OAI21_X1 _20071_ (.A(_05095_),
    .B1(_05731_),
    .B2(_10409_),
    .ZN(_10410_));
 AOI211_X2 _20072_ (.A(_10408_),
    .B(_10410_),
    .C1(_04297_),
    .C2(_05009_),
    .ZN(_10411_));
 OAI21_X1 _20073_ (.A(_04757_),
    .B1(_10078_),
    .B2(_06270_),
    .ZN(_10412_));
 AND4_X1 _20074_ (.A1(_10407_),
    .A2(_10411_),
    .A3(_09718_),
    .A4(_10412_),
    .ZN(_10413_));
 OAI221_X1 _20075_ (.A(_09444_),
    .B1(_10076_),
    .B2(_05764_),
    .C1(_06270_),
    .C2(_09441_),
    .ZN(_10414_));
 OAI21_X1 _20076_ (.A(_04483_),
    .B1(_10130_),
    .B2(_05566_),
    .ZN(_10415_));
 INV_X1 _20077_ (.A(_09455_),
    .ZN(_10416_));
 NAND3_X1 _20078_ (.A1(_04483_),
    .A2(_04669_),
    .A3(_04658_),
    .ZN(_10417_));
 AND4_X1 _20079_ (.A1(_04264_),
    .A2(_10415_),
    .A3(_10416_),
    .A4(_10417_),
    .ZN(_10418_));
 AND4_X2 _20080_ (.A1(_10406_),
    .A2(_10413_),
    .A3(_10414_),
    .A4(_10418_),
    .ZN(_10419_));
 OAI21_X1 _20081_ (.A(_05390_),
    .B1(_09422_),
    .B2(_05456_),
    .ZN(_10420_));
 NAND2_X1 _20082_ (.A1(_05489_),
    .A2(_05709_),
    .ZN(_10421_));
 NAND4_X1 _20083_ (.A1(_10420_),
    .A2(_05445_),
    .A3(_10421_),
    .A4(_10171_),
    .ZN(_10422_));
 NAND2_X1 _20084_ (.A1(_10085_),
    .A2(_06314_),
    .ZN(_10423_));
 NAND2_X1 _20085_ (.A1(_10084_),
    .A2(_10423_),
    .ZN(_10424_));
 NOR4_X1 _20086_ (.A1(_10422_),
    .A2(_10424_),
    .A3(_10164_),
    .A4(_09522_),
    .ZN(_10425_));
 OAI21_X1 _20087_ (.A(_05599_),
    .B1(_05056_),
    .B2(_05180_),
    .ZN(_10426_));
 OAI21_X1 _20088_ (.A(_05599_),
    .B1(_04253_),
    .B2(_09505_),
    .ZN(_10427_));
 AND3_X1 _20089_ (.A1(_05588_),
    .A2(_10426_),
    .A3(_10427_),
    .ZN(_10428_));
 OAI21_X1 _20090_ (.A(_05357_),
    .B1(_06391_),
    .B2(_05412_),
    .ZN(_10429_));
 AND4_X1 _20091_ (.A1(_05291_),
    .A2(_10425_),
    .A3(_10428_),
    .A4(_10429_),
    .ZN(_10430_));
 AND2_X2 _20092_ (.A1(_05808_),
    .A2(_05984_),
    .ZN(_10431_));
 INV_X2 _20093_ (.A(_10431_),
    .ZN(_10432_));
 NAND4_X1 _20094_ (.A1(_10432_),
    .A2(_09430_),
    .A3(_09753_),
    .A4(_10206_),
    .ZN(_10433_));
 AND2_X1 _20095_ (.A1(_05841_),
    .A2(_04910_),
    .ZN(_10434_));
 OR4_X2 _20096_ (.A1(_09424_),
    .A2(_10433_),
    .A3(_10110_),
    .A4(_10434_),
    .ZN(_10435_));
 NAND2_X1 _20097_ (.A1(_06061_),
    .A2(_09692_),
    .ZN(_10436_));
 OAI211_X2 _20098_ (.A(_06061_),
    .B(_06270_),
    .C1(_10076_),
    .C2(_05522_),
    .ZN(_10437_));
 INV_X1 _20099_ (.A(_09477_),
    .ZN(_10438_));
 INV_X1 _20100_ (.A(_06050_),
    .ZN(_10439_));
 OAI211_X2 _20101_ (.A(_10436_),
    .B(_10437_),
    .C1(_10438_),
    .C2(_10439_),
    .ZN(_10440_));
 AOI21_X1 _20102_ (.A(_06006_),
    .B1(_05188_),
    .B2(_05940_),
    .ZN(_10441_));
 OAI211_X2 _20103_ (.A(_05940_),
    .B(_06270_),
    .C1(_10076_),
    .C2(_05764_),
    .ZN(_10442_));
 OAI211_X2 _20104_ (.A(_05940_),
    .B(_09441_),
    .C1(_05511_),
    .C2(_05764_),
    .ZN(_10443_));
 NAND3_X1 _20105_ (.A1(_10441_),
    .A2(_10442_),
    .A3(_10443_),
    .ZN(_10444_));
 NAND3_X1 _20106_ (.A1(_05984_),
    .A2(_09438_),
    .A3(_05863_),
    .ZN(_10445_));
 OAI211_X2 _20107_ (.A(_09437_),
    .B(_10445_),
    .C1(_10203_),
    .C2(_05698_),
    .ZN(_10446_));
 NOR4_X4 _20108_ (.A1(_10435_),
    .A2(_10440_),
    .A3(_10444_),
    .A4(_10446_),
    .ZN(_10447_));
 AND2_X1 _20109_ (.A1(_09491_),
    .A2(_05047_),
    .ZN(_10448_));
 INV_X1 _20110_ (.A(_10448_),
    .ZN(_10449_));
 NAND2_X1 _20111_ (.A1(_09491_),
    .A2(_04549_),
    .ZN(_10450_));
 OAI21_X1 _20112_ (.A(_09491_),
    .B1(_09422_),
    .B2(_05456_),
    .ZN(_10451_));
 NAND4_X1 _20113_ (.A1(_10449_),
    .A2(_09738_),
    .A3(_10450_),
    .A4(_10451_),
    .ZN(_10452_));
 AND2_X1 _20114_ (.A1(_05188_),
    .A2(_06435_),
    .ZN(_10453_));
 INV_X1 _20115_ (.A(_10453_),
    .ZN(_10454_));
 OAI21_X1 _20116_ (.A(_06446_),
    .B1(_09473_),
    .B2(_10078_),
    .ZN(_10455_));
 NAND4_X1 _20117_ (.A1(_09499_),
    .A2(_10454_),
    .A3(_06479_),
    .A4(_10455_),
    .ZN(_10456_));
 OAI21_X1 _20118_ (.A(_09482_),
    .B1(_09507_),
    .B2(_10081_),
    .ZN(_10457_));
 NAND4_X1 _20119_ (.A1(_09482_),
    .A2(_09468_),
    .A3(_04669_),
    .A4(_04527_),
    .ZN(_10458_));
 OAI211_X2 _20120_ (.A(_10457_),
    .B(_10458_),
    .C1(_04790_),
    .C2(_09748_),
    .ZN(_10459_));
 OAI21_X1 _20121_ (.A(_06226_),
    .B1(_05456_),
    .B2(_05152_),
    .ZN(_10460_));
 OAI21_X1 _20122_ (.A(_06226_),
    .B1(_05335_),
    .B2(_05313_),
    .ZN(_10461_));
 NAND2_X1 _20123_ (.A1(_10460_),
    .A2(_10461_),
    .ZN(_10462_));
 NOR4_X1 _20124_ (.A1(_10452_),
    .A2(_10456_),
    .A3(_10459_),
    .A4(_10462_),
    .ZN(_10463_));
 NAND4_X1 _20125_ (.A1(_10419_),
    .A2(_10430_),
    .A3(_10447_),
    .A4(_10463_),
    .ZN(_10464_));
 NOR2_X2 _20126_ (.A1(_10464_),
    .A2(_06556_),
    .ZN(_10465_));
 XNOR2_X1 _20127_ (.A(_10465_),
    .B(_10270_),
    .ZN(_10466_));
 OAI21_X1 _20128_ (.A(_07117_),
    .B1(_10040_),
    .B2(_08538_),
    .ZN(_10467_));
 AND3_X1 _20129_ (.A1(_07664_),
    .A2(_07883_),
    .A3(_06941_),
    .ZN(_10468_));
 AOI211_X2 _20130_ (.A(_10468_),
    .B(_10045_),
    .C1(_06798_),
    .C2(_08190_),
    .ZN(_10469_));
 NAND4_X1 _20131_ (.A1(_07949_),
    .A2(_08047_),
    .A3(_08058_),
    .A4(_06897_),
    .ZN(_10470_));
 NAND2_X1 _20132_ (.A1(_09571_),
    .A2(_09538_),
    .ZN(_10471_));
 OAI21_X1 _20133_ (.A(_07326_),
    .B1(_10471_),
    .B2(_07751_),
    .ZN(_10472_));
 AND4_X1 _20134_ (.A1(_10023_),
    .A2(_10469_),
    .A3(_10470_),
    .A4(_10472_),
    .ZN(_10473_));
 AND4_X1 _20135_ (.A1(_07018_),
    .A2(_07304_),
    .A3(_07051_),
    .A4(_06820_),
    .ZN(_10474_));
 AND2_X1 _20136_ (.A1(_07477_),
    .A2(_07631_),
    .ZN(_10475_));
 AOI211_X2 _20137_ (.A(_10474_),
    .B(_10475_),
    .C1(_08544_),
    .C2(_07565_),
    .ZN(_10476_));
 OAI21_X1 _20138_ (.A(_08544_),
    .B1(_09106_),
    .B2(_09166_),
    .ZN(_10477_));
 AND4_X2 _20139_ (.A1(_10467_),
    .A2(_10473_),
    .A3(_10476_),
    .A4(_10477_),
    .ZN(_10478_));
 INV_X1 _20140_ (.A(_07260_),
    .ZN(_10479_));
 AOI21_X1 _20141_ (.A(_10479_),
    .B1(_09167_),
    .B2(_09572_),
    .ZN(_10480_));
 AND2_X1 _20142_ (.A1(_07828_),
    .A2(_07260_),
    .ZN(_10481_));
 AND4_X1 _20143_ (.A1(_08538_),
    .A2(_07018_),
    .A3(_08519_),
    .A4(_07238_),
    .ZN(_10482_));
 NOR3_X1 _20144_ (.A1(_10480_),
    .A2(_10481_),
    .A3(_10482_),
    .ZN(_10483_));
 OAI21_X1 _20145_ (.A(_07795_),
    .B1(_07631_),
    .B2(_08556_),
    .ZN(_10484_));
 NOR2_X1 _20146_ (.A1(_08025_),
    .A2(_09105_),
    .ZN(_10485_));
 NOR2_X1 _20147_ (.A1(_10485_),
    .A2(_09545_),
    .ZN(_10486_));
 INV_X1 _20148_ (.A(_10486_),
    .ZN(_10487_));
 NAND4_X1 _20149_ (.A1(_10483_),
    .A2(_09212_),
    .A3(_10484_),
    .A4(_10487_),
    .ZN(_10488_));
 AOI21_X1 _20150_ (.A(_09120_),
    .B1(_09550_),
    .B2(_06996_),
    .ZN(_10489_));
 OAI211_X2 _20151_ (.A(_09149_),
    .B(_09612_),
    .C1(_09121_),
    .C2(_09120_),
    .ZN(_10490_));
 NOR4_X1 _20152_ (.A1(_10488_),
    .A2(_10051_),
    .A3(_10489_),
    .A4(_10490_),
    .ZN(_10491_));
 NAND2_X1 _20153_ (.A1(_10003_),
    .A2(_07894_),
    .ZN(_10492_));
 AOI22_X1 _20154_ (.A1(_07172_),
    .A2(_07227_),
    .B1(_07414_),
    .B2(_09549_),
    .ZN(_10493_));
 OAI211_X2 _20155_ (.A(_10492_),
    .B(_10493_),
    .C1(_07543_),
    .C2(_07370_),
    .ZN(_10494_));
 AOI21_X1 _20156_ (.A(_08443_),
    .B1(_08472_),
    .B2(_07139_),
    .ZN(_10495_));
 NOR3_X1 _20157_ (.A1(_10494_),
    .A2(_08102_),
    .A3(_10495_),
    .ZN(_10496_));
 OAI211_X2 _20158_ (.A(_10304_),
    .B(_09557_),
    .C1(_09545_),
    .C2(_07850_),
    .ZN(_10497_));
 NAND3_X1 _20159_ (.A1(_09113_),
    .A2(_09544_),
    .A3(_09607_),
    .ZN(_10498_));
 NOR4_X1 _20160_ (.A1(_10497_),
    .A2(_10498_),
    .A3(_08277_),
    .A4(_10014_),
    .ZN(_10499_));
 NAND4_X1 _20161_ (.A1(_10478_),
    .A2(_10491_),
    .A3(_10496_),
    .A4(_10499_),
    .ZN(_10500_));
 INV_X1 _20162_ (.A(_10283_),
    .ZN(_10501_));
 AND4_X1 _20163_ (.A1(_09193_),
    .A2(_10026_),
    .A3(_09594_),
    .A4(_10501_),
    .ZN(_10502_));
 NAND2_X1 _20164_ (.A1(_10294_),
    .A2(_10299_),
    .ZN(_10503_));
 AOI221_X4 _20165_ (.A(_10503_),
    .B1(_07205_),
    .B2(_06611_),
    .C1(_06908_),
    .C2(_09192_),
    .ZN(_10504_));
 OAI21_X1 _20166_ (.A(_07392_),
    .B1(_07532_),
    .B2(_07414_),
    .ZN(_10505_));
 AND4_X1 _20167_ (.A1(_08510_),
    .A2(_10505_),
    .A3(_09114_),
    .A4(_09576_),
    .ZN(_10506_));
 OAI21_X1 _20168_ (.A(_08299_),
    .B1(_07499_),
    .B2(_07565_),
    .ZN(_10507_));
 OAI22_X1 _20169_ (.A1(_08386_),
    .A2(_07282_),
    .B1(_06996_),
    .B2(_06644_),
    .ZN(_10508_));
 OAI21_X1 _20170_ (.A(_08550_),
    .B1(_10508_),
    .B2(_06655_),
    .ZN(_10509_));
 OAI21_X1 _20171_ (.A(_08299_),
    .B1(_08025_),
    .B2(_07828_),
    .ZN(_10510_));
 OAI21_X1 _20172_ (.A(_07414_),
    .B1(_07293_),
    .B2(_09142_),
    .ZN(_10511_));
 AND4_X1 _20173_ (.A1(_10507_),
    .A2(_10509_),
    .A3(_10510_),
    .A4(_10511_),
    .ZN(_10512_));
 NAND4_X1 _20174_ (.A1(_10502_),
    .A2(_10504_),
    .A3(_10506_),
    .A4(_10512_),
    .ZN(_10513_));
 NOR2_X4 _20175_ (.A1(_10500_),
    .A2(_10513_),
    .ZN(_10514_));
 AND4_X1 _20176_ (.A1(_08595_),
    .A2(_08756_),
    .A3(_08604_),
    .A4(_08605_),
    .ZN(_10515_));
 AOI211_X4 _20177_ (.A(_09640_),
    .B(_10515_),
    .C1(_08760_),
    .C2(_08674_),
    .ZN(_10516_));
 INV_X1 _20178_ (.A(_08786_),
    .ZN(_10517_));
 OAI21_X1 _20179_ (.A(_08678_),
    .B1(_08636_),
    .B2(_08671_),
    .ZN(_10518_));
 OAI211_X2 _20180_ (.A(_10517_),
    .B(_10518_),
    .C1(_09279_),
    .C2(_08839_),
    .ZN(_10519_));
 AOI211_X2 _20181_ (.A(_09655_),
    .B(_10519_),
    .C1(_08646_),
    .C2(_08645_),
    .ZN(_10520_));
 OAI21_X1 _20182_ (.A(_08760_),
    .B1(_08666_),
    .B2(_09966_),
    .ZN(_10521_));
 AND4_X1 _20183_ (.A1(_08613_),
    .A2(_08713_),
    .A3(_08619_),
    .A4(_08570_),
    .ZN(_10522_));
 AOI221_X4 _20184_ (.A(_10522_),
    .B1(_08673_),
    .B2(_08720_),
    .C1(_09214_),
    .C2(_08830_),
    .ZN(_10523_));
 NAND2_X1 _20185_ (.A1(_08721_),
    .A2(_08633_),
    .ZN(_10524_));
 NAND4_X1 _20186_ (.A1(_08725_),
    .A2(_08620_),
    .A3(_08586_),
    .A4(_08583_),
    .ZN(_10525_));
 AND3_X1 _20187_ (.A1(_10523_),
    .A2(_10524_),
    .A3(_10525_),
    .ZN(_10526_));
 AND4_X1 _20188_ (.A1(_10516_),
    .A2(_10520_),
    .A3(_10521_),
    .A4(_10526_),
    .ZN(_10527_));
 AND2_X1 _20189_ (.A1(_08622_),
    .A2(_08779_),
    .ZN(_10528_));
 AND2_X1 _20190_ (.A1(_08788_),
    .A2(_08790_),
    .ZN(_10529_));
 NOR4_X1 _20191_ (.A1(_08864_),
    .A2(_10528_),
    .A3(_08835_),
    .A4(_10529_),
    .ZN(_10530_));
 AOI221_X4 _20192_ (.A(_09931_),
    .B1(_08695_),
    .B2(_08704_),
    .C1(_08748_),
    .C2(_08578_),
    .ZN(_10531_));
 OAI21_X1 _20193_ (.A(_09652_),
    .B1(_09641_),
    .B2(_08659_),
    .ZN(_10532_));
 AOI221_X4 _20194_ (.A(_10532_),
    .B1(_08575_),
    .B2(_10216_),
    .C1(_08741_),
    .C2(_08798_),
    .ZN(_10533_));
 NAND4_X1 _20195_ (.A1(_10527_),
    .A2(_10530_),
    .A3(_10531_),
    .A4(_10533_),
    .ZN(_10534_));
 OAI211_X2 _20196_ (.A(_10259_),
    .B(_10252_),
    .C1(_09231_),
    .C2(_08821_),
    .ZN(_10535_));
 NOR4_X1 _20197_ (.A1(_10535_),
    .A2(_08664_),
    .A3(_10256_),
    .A4(_08667_),
    .ZN(_10536_));
 NOR3_X1 _20198_ (.A1(_16784_),
    .A2(_16787_),
    .A3(_16786_),
    .ZN(_10537_));
 AOI211_X4 _20199_ (.A(_09625_),
    .B(_08827_),
    .C1(_09243_),
    .C2(_10537_),
    .ZN(_10538_));
 NAND3_X1 _20200_ (.A1(_10258_),
    .A2(_08725_),
    .A3(_08650_),
    .ZN(_10539_));
 NAND3_X1 _20201_ (.A1(_08669_),
    .A2(_08683_),
    .A3(_08725_),
    .ZN(_10540_));
 NAND2_X1 _20202_ (.A1(_10539_),
    .A2(_10540_),
    .ZN(_10541_));
 AND2_X1 _20203_ (.A1(_08709_),
    .A2(_08640_),
    .ZN(_10542_));
 AND3_X1 _20204_ (.A1(_08681_),
    .A2(_08575_),
    .A3(_08830_),
    .ZN(_10543_));
 NOR4_X1 _20205_ (.A1(_10541_),
    .A2(_10235_),
    .A3(_10542_),
    .A4(_10543_),
    .ZN(_10544_));
 NAND2_X1 _20206_ (.A1(_08731_),
    .A2(_08843_),
    .ZN(_10545_));
 AOI22_X1 _20207_ (.A1(_08622_),
    .A2(_08790_),
    .B1(_08637_),
    .B2(_08640_),
    .ZN(_10546_));
 NAND3_X1 _20208_ (.A1(_08860_),
    .A2(_16786_),
    .A3(_08650_),
    .ZN(_10547_));
 OAI21_X1 _20209_ (.A(_08747_),
    .B1(_08810_),
    .B2(_08709_),
    .ZN(_10548_));
 AND4_X1 _20210_ (.A1(_10545_),
    .A2(_10546_),
    .A3(_10547_),
    .A4(_10548_),
    .ZN(_10549_));
 AND4_X1 _20211_ (.A1(_10536_),
    .A2(_10538_),
    .A3(_10544_),
    .A4(_10549_),
    .ZN(_10550_));
 OAI21_X1 _20212_ (.A(_08788_),
    .B1(_08717_),
    .B2(_08836_),
    .ZN(_10551_));
 OAI21_X1 _20213_ (.A(_08694_),
    .B1(_08810_),
    .B2(_08798_),
    .ZN(_10552_));
 OAI21_X1 _20214_ (.A(_08694_),
    .B1(_10258_),
    .B2(_08779_),
    .ZN(_10553_));
 AND4_X1 _20215_ (.A1(_08700_),
    .A2(_10551_),
    .A3(_10552_),
    .A4(_10553_),
    .ZN(_10554_));
 OAI21_X1 _20216_ (.A(_08715_),
    .B1(_08816_),
    .B2(_08628_),
    .ZN(_10555_));
 OAI21_X1 _20217_ (.A(_09633_),
    .B1(_08686_),
    .B2(_08674_),
    .ZN(_10556_));
 OAI21_X1 _20218_ (.A(_09633_),
    .B1(_08709_),
    .B2(_08662_),
    .ZN(_10557_));
 AND3_X1 _20219_ (.A1(_10555_),
    .A2(_10556_),
    .A3(_10557_),
    .ZN(_10558_));
 OAI21_X1 _20220_ (.A(_08608_),
    .B1(_08596_),
    .B2(_08610_),
    .ZN(_10559_));
 OAI21_X1 _20221_ (.A(_08748_),
    .B1(_08724_),
    .B2(_08674_),
    .ZN(_10560_));
 AOI22_X1 _20222_ (.A1(_08704_),
    .A2(_08770_),
    .B1(_08731_),
    .B2(_08681_),
    .ZN(_10561_));
 AND4_X1 _20223_ (.A1(_08685_),
    .A2(_10559_),
    .A3(_10560_),
    .A4(_10561_),
    .ZN(_10562_));
 NAND4_X1 _20224_ (.A1(_10550_),
    .A2(_10554_),
    .A3(_10558_),
    .A4(_10562_),
    .ZN(_10563_));
 NOR2_X4 _20225_ (.A1(_10534_),
    .A2(_10563_),
    .ZN(_10564_));
 XNOR2_X2 _20226_ (.A(_10514_),
    .B(_10564_),
    .ZN(_10565_));
 XNOR2_X1 _20227_ (.A(_10466_),
    .B(_10565_),
    .ZN(_10566_));
 AND2_X1 _20228_ (.A1(_08893_),
    .A2(_09051_),
    .ZN(_10567_));
 AND2_X1 _20229_ (.A1(_08893_),
    .A2(_08998_),
    .ZN(_10568_));
 AOI211_X4 _20230_ (.A(_10567_),
    .B(_10568_),
    .C1(_09394_),
    .C2(_09326_),
    .ZN(_10569_));
 NAND2_X1 _20231_ (.A1(_09326_),
    .A2(_08961_),
    .ZN(_10570_));
 NAND2_X1 _20232_ (.A1(_09072_),
    .A2(_09354_),
    .ZN(_10571_));
 NAND2_X1 _20233_ (.A1(_09354_),
    .A2(_09378_),
    .ZN(_10572_));
 OAI211_X2 _20234_ (.A(_08906_),
    .B(_08961_),
    .C1(_08962_),
    .C2(_08900_),
    .ZN(_10573_));
 AND4_X1 _20235_ (.A1(_10340_),
    .A2(_10571_),
    .A3(_10572_),
    .A4(_10573_),
    .ZN(_10574_));
 AND4_X1 _20236_ (.A1(_08902_),
    .A2(_10569_),
    .A3(_10570_),
    .A4(_10574_),
    .ZN(_10575_));
 NAND2_X1 _20237_ (.A1(_09327_),
    .A2(_08924_),
    .ZN(_10576_));
 OAI221_X1 _20238_ (.A(_10576_),
    .B1(_10331_),
    .B2(_09067_),
    .C1(_09784_),
    .C2(_10330_),
    .ZN(_10577_));
 INV_X1 _20239_ (.A(_09768_),
    .ZN(_10578_));
 AOI21_X1 _20240_ (.A(_09372_),
    .B1(_09070_),
    .B2(_10578_),
    .ZN(_10579_));
 AOI21_X1 _20241_ (.A(_10331_),
    .B1(_09009_),
    .B2(_09385_),
    .ZN(_10580_));
 NOR4_X1 _20242_ (.A1(_10577_),
    .A2(_09810_),
    .A3(_10579_),
    .A4(_10580_),
    .ZN(_10581_));
 NAND3_X1 _20243_ (.A1(_09305_),
    .A2(_09017_),
    .A3(_09355_),
    .ZN(_10582_));
 NAND3_X1 _20244_ (.A1(_09305_),
    .A2(_09832_),
    .A3(_09017_),
    .ZN(_10583_));
 NAND2_X1 _20245_ (.A1(_09400_),
    .A2(_09305_),
    .ZN(_10584_));
 NAND4_X1 _20246_ (.A1(_09894_),
    .A2(_10582_),
    .A3(_10583_),
    .A4(_10584_),
    .ZN(_10585_));
 AOI21_X1 _20247_ (.A(_09303_),
    .B1(_09033_),
    .B2(_09011_),
    .ZN(_10586_));
 NOR4_X1 _20248_ (.A1(_10585_),
    .A2(_08958_),
    .A3(_09375_),
    .A4(_10586_),
    .ZN(_10587_));
 NAND3_X1 _20249_ (.A1(_09789_),
    .A2(_08959_),
    .A3(_09364_),
    .ZN(_10588_));
 AND2_X1 _20250_ (.A1(_09005_),
    .A2(_08912_),
    .ZN(_10589_));
 AND2_X1 _20251_ (.A1(_08910_),
    .A2(_09005_),
    .ZN(_10590_));
 AOI211_X4 _20252_ (.A(_10589_),
    .B(_10590_),
    .C1(_09377_),
    .C2(_08957_),
    .ZN(_10591_));
 OAI211_X2 _20253_ (.A(_09789_),
    .B(_08993_),
    .C1(_08977_),
    .C2(_09355_),
    .ZN(_10592_));
 OAI21_X1 _20254_ (.A(_09789_),
    .B1(_09340_),
    .B2(_09331_),
    .ZN(_10593_));
 AND4_X1 _20255_ (.A1(_10588_),
    .A2(_10591_),
    .A3(_10592_),
    .A4(_10593_),
    .ZN(_10594_));
 NAND4_X1 _20256_ (.A1(_10575_),
    .A2(_10581_),
    .A3(_10587_),
    .A4(_10594_),
    .ZN(_10595_));
 AOI221_X2 _20257_ (.A(_10362_),
    .B1(_09339_),
    .B2(_08984_),
    .C1(_08962_),
    .C2(_09777_),
    .ZN(_10596_));
 OAI21_X1 _20258_ (.A(_09797_),
    .B1(_09026_),
    .B2(_08955_),
    .ZN(_10597_));
 OAI21_X1 _20259_ (.A(_09797_),
    .B1(_08981_),
    .B2(_09002_),
    .ZN(_10598_));
 AND4_X1 _20260_ (.A1(_09343_),
    .A2(_10596_),
    .A3(_10597_),
    .A4(_10598_),
    .ZN(_10599_));
 OAI211_X2 _20261_ (.A(_09405_),
    .B(_09832_),
    .C1(_09054_),
    .C2(_09784_),
    .ZN(_10600_));
 OAI21_X1 _20262_ (.A(_09405_),
    .B1(_08955_),
    .B2(_08924_),
    .ZN(_10601_));
 NAND4_X1 _20263_ (.A1(_10600_),
    .A2(_10601_),
    .A3(_09043_),
    .A4(_10390_),
    .ZN(_10602_));
 AND2_X1 _20264_ (.A1(_09768_),
    .A2(_09053_),
    .ZN(_10603_));
 NOR4_X1 _20265_ (.A1(_10602_),
    .A2(_09870_),
    .A3(_10377_),
    .A4(_10603_),
    .ZN(_10604_));
 INV_X1 _20266_ (.A(_09325_),
    .ZN(_10605_));
 AOI21_X1 _20267_ (.A(_09023_),
    .B1(_10605_),
    .B2(_09359_),
    .ZN(_10606_));
 NAND3_X1 _20268_ (.A1(_09397_),
    .A2(_09832_),
    .A3(_08909_),
    .ZN(_10607_));
 NAND2_X1 _20269_ (.A1(_09397_),
    .A2(_08961_),
    .ZN(_10608_));
 OAI211_X2 _20270_ (.A(_10607_),
    .B(_10608_),
    .C1(_09302_),
    .C2(_09032_),
    .ZN(_10609_));
 NOR4_X1 _20271_ (.A1(_10606_),
    .A2(_10609_),
    .A3(_09859_),
    .A4(_09778_),
    .ZN(_10610_));
 AOI22_X1 _20272_ (.A1(_10397_),
    .A2(_08956_),
    .B1(_08987_),
    .B2(_09330_),
    .ZN(_10611_));
 OAI21_X1 _20273_ (.A(_09074_),
    .B1(_08934_),
    .B2(_08987_),
    .ZN(_10612_));
 OAI21_X1 _20274_ (.A(_09330_),
    .B1(_09378_),
    .B2(_09374_),
    .ZN(_10613_));
 AND4_X1 _20275_ (.A1(_09793_),
    .A2(_10611_),
    .A3(_10612_),
    .A4(_10613_),
    .ZN(_10614_));
 NAND4_X1 _20276_ (.A1(_10599_),
    .A2(_10604_),
    .A3(_10610_),
    .A4(_10614_),
    .ZN(_10615_));
 NOR2_X4 _20277_ (.A1(_10595_),
    .A2(_10615_),
    .ZN(_10616_));
 XNOR2_X1 _20278_ (.A(_10566_),
    .B(_10616_),
    .ZN(_10617_));
 XNOR2_X1 _20279_ (.A(_10617_),
    .B(_17171_),
    .ZN(_10618_));
 MUX2_X1 _20280_ (.A(_10405_),
    .B(_10618_),
    .S(_09100_),
    .Z(_00729_));
 XOR2_X1 _20281_ (.A(_17172_),
    .B(_17106_),
    .Z(_10619_));
 AOI21_X1 _20282_ (.A(_08826_),
    .B1(_08820_),
    .B2(_08689_),
    .ZN(_10620_));
 AOI21_X1 _20283_ (.A(_10620_),
    .B1(_08731_),
    .B2(_09657_),
    .ZN(_10621_));
 OAI21_X1 _20284_ (.A(_08715_),
    .B1(_08822_),
    .B2(_09239_),
    .ZN(_10622_));
 AOI211_X2 _20285_ (.A(_08623_),
    .B(_09231_),
    .C1(_16780_),
    .C2(_08611_),
    .ZN(_10623_));
 AOI221_X1 _20286_ (.A(_10623_),
    .B1(_08614_),
    .B2(_09932_),
    .C1(_08740_),
    .C2(_08723_),
    .ZN(_10624_));
 NAND4_X1 _20287_ (.A1(_08725_),
    .A2(_08830_),
    .A3(_08582_),
    .A4(_08683_),
    .ZN(_10625_));
 OAI21_X1 _20288_ (.A(_08714_),
    .B1(_08697_),
    .B2(_08681_),
    .ZN(_10626_));
 AND4_X1 _20289_ (.A1(_10622_),
    .A2(_10624_),
    .A3(_10625_),
    .A4(_10626_),
    .ZN(_10627_));
 OAI211_X2 _20290_ (.A(_08731_),
    .B(_16783_),
    .C1(_08706_),
    .C2(_08568_),
    .ZN(_10628_));
 AND4_X1 _20291_ (.A1(_10524_),
    .A2(_09920_),
    .A3(_08829_),
    .A4(_09220_),
    .ZN(_10629_));
 AND4_X1 _20292_ (.A1(_10621_),
    .A2(_10627_),
    .A3(_10628_),
    .A4(_10629_),
    .ZN(_10630_));
 AOI221_X1 _20293_ (.A(_08845_),
    .B1(_08767_),
    .B2(_08703_),
    .C1(_08584_),
    .C2(_08842_),
    .ZN(_10631_));
 NAND3_X1 _20294_ (.A1(_08631_),
    .A2(_08675_),
    .A3(_08620_),
    .ZN(_10632_));
 NAND4_X1 _20295_ (.A1(_10631_),
    .A2(_08707_),
    .A3(_08710_),
    .A4(_10632_),
    .ZN(_10633_));
 AND3_X1 _20296_ (.A1(_08606_),
    .A2(_08595_),
    .A3(_08679_),
    .ZN(_10634_));
 AND2_X1 _20297_ (.A1(_08666_),
    .A2(_08679_),
    .ZN(_10635_));
 AND4_X1 _20298_ (.A1(_08830_),
    .A2(_08582_),
    .A3(_08675_),
    .A4(_08563_),
    .ZN(_10636_));
 OR3_X1 _20299_ (.A1(_10634_),
    .A2(_10635_),
    .A3(_10636_),
    .ZN(_10637_));
 OAI21_X1 _20300_ (.A(_08694_),
    .B1(_08671_),
    .B2(_08763_),
    .ZN(_10638_));
 OAI211_X2 _20301_ (.A(_10638_),
    .B(_09975_),
    .C1(_08855_),
    .C2(_08874_),
    .ZN(_10639_));
 AND3_X1 _20302_ (.A1(_08718_),
    .A2(_08650_),
    .A3(_08656_),
    .ZN(_10640_));
 OR4_X4 _20303_ (.A1(_08850_),
    .A2(_08837_),
    .A3(_08847_),
    .A4(_10640_),
    .ZN(_10641_));
 NOR4_X2 _20304_ (.A1(_10633_),
    .A2(_10637_),
    .A3(_10639_),
    .A4(_10641_),
    .ZN(_10642_));
 OAI21_X1 _20305_ (.A(_08608_),
    .B1(_08573_),
    .B2(_08798_),
    .ZN(_10643_));
 OAI21_X1 _20306_ (.A(_08607_),
    .B1(_08789_),
    .B2(_08632_),
    .ZN(_10644_));
 OAI21_X1 _20307_ (.A(_08607_),
    .B1(_08785_),
    .B2(_08578_),
    .ZN(_10645_));
 AND3_X1 _20308_ (.A1(_10643_),
    .A2(_10644_),
    .A3(_10645_),
    .ZN(_10646_));
 AND2_X1 _20309_ (.A1(_08621_),
    .A2(_08681_),
    .ZN(_10647_));
 AND3_X1 _20310_ (.A1(_08859_),
    .A2(_08599_),
    .A3(_08620_),
    .ZN(_10648_));
 NOR4_X1 _20311_ (.A1(_10528_),
    .A2(_08882_),
    .A3(_10647_),
    .A4(_10648_),
    .ZN(_10649_));
 AOI21_X1 _20312_ (.A(_08588_),
    .B1(_09279_),
    .B2(_08716_),
    .ZN(_10650_));
 NOR2_X1 _20313_ (.A1(_09665_),
    .A2(_10650_),
    .ZN(_10651_));
 AND2_X1 _20314_ (.A1(_08697_),
    .A2(_08645_),
    .ZN(_10652_));
 AND2_X1 _20315_ (.A1(_08640_),
    .A2(_08630_),
    .ZN(_10653_));
 NOR4_X1 _20316_ (.A1(_10652_),
    .A2(_10542_),
    .A3(_10653_),
    .A4(_08643_),
    .ZN(_10654_));
 AND4_X1 _20317_ (.A1(_10646_),
    .A2(_10649_),
    .A3(_10651_),
    .A4(_10654_),
    .ZN(_10655_));
 OAI21_X1 _20318_ (.A(_08788_),
    .B1(_10258_),
    .B2(_08666_),
    .ZN(_10656_));
 OAI211_X2 _20319_ (.A(_08774_),
    .B(_08649_),
    .C1(_08585_),
    .C2(_08586_),
    .ZN(_10657_));
 AND2_X1 _20320_ (.A1(_10656_),
    .A2(_10657_),
    .ZN(_10658_));
 OAI21_X1 _20321_ (.A(_08748_),
    .B1(_08822_),
    .B2(_09239_),
    .ZN(_10659_));
 AND4_X1 _20322_ (.A1(_08563_),
    .A2(_08581_),
    .A3(_08613_),
    .A4(_08745_),
    .ZN(_10660_));
 AOI211_X2 _20323_ (.A(_10660_),
    .B(_08804_),
    .C1(_08630_),
    .C2(_08756_),
    .ZN(_10661_));
 OAI21_X1 _20324_ (.A(_08747_),
    .B1(_08666_),
    .B2(_09966_),
    .ZN(_10662_));
 OAI21_X1 _20325_ (.A(_08760_),
    .B1(_08860_),
    .B2(_08843_),
    .ZN(_10663_));
 AND4_X1 _20326_ (.A1(_10659_),
    .A2(_10661_),
    .A3(_10662_),
    .A4(_10663_),
    .ZN(_10664_));
 OAI21_X1 _20327_ (.A(_09633_),
    .B1(_08798_),
    .B2(_08674_),
    .ZN(_10665_));
 OAI21_X1 _20328_ (.A(_09633_),
    .B1(_08800_),
    .B2(_08709_),
    .ZN(_10666_));
 AND4_X2 _20329_ (.A1(_10658_),
    .A2(_10664_),
    .A3(_10665_),
    .A4(_10666_),
    .ZN(_10667_));
 NAND4_X1 _20330_ (.A1(_10630_),
    .A2(_10642_),
    .A3(_10655_),
    .A4(_10667_),
    .ZN(_10668_));
 NOR2_X2 _20331_ (.A1(_10668_),
    .A2(_08786_),
    .ZN(_10669_));
 OAI21_X1 _20332_ (.A(_08550_),
    .B1(_08343_),
    .B2(_10285_),
    .ZN(_10670_));
 OR3_X1 _20333_ (.A1(_09561_),
    .A2(_09555_),
    .A3(_10027_),
    .ZN(_10671_));
 AND2_X1 _20334_ (.A1(_07708_),
    .A2(_07227_),
    .ZN(_10672_));
 OAI211_X2 _20335_ (.A(_10303_),
    .B(_10048_),
    .C1(_07370_),
    .C2(_09120_),
    .ZN(_10673_));
 NOR4_X2 _20336_ (.A1(_10671_),
    .A2(_10672_),
    .A3(_10004_),
    .A4(_10673_),
    .ZN(_10674_));
 OAI21_X1 _20337_ (.A(_08550_),
    .B1(_09125_),
    .B2(_10038_),
    .ZN(_10675_));
 AND4_X1 _20338_ (.A1(_07051_),
    .A2(_07795_),
    .A3(_07730_),
    .A4(_08244_),
    .ZN(_10676_));
 AND4_X1 _20339_ (.A1(_07029_),
    .A2(_07740_),
    .A3(_08058_),
    .A4(_08080_),
    .ZN(_10677_));
 NOR4_X1 _20340_ (.A1(_10676_),
    .A2(_09603_),
    .A3(_09126_),
    .A4(_10677_),
    .ZN(_10678_));
 AND4_X2 _20341_ (.A1(_10670_),
    .A2(_10674_),
    .A3(_10675_),
    .A4(_10678_),
    .ZN(_10679_));
 AND2_X1 _20342_ (.A1(_07719_),
    .A2(_09106_),
    .ZN(_10680_));
 NOR4_X1 _20343_ (.A1(_09139_),
    .A2(_09197_),
    .A3(_06864_),
    .A4(_10680_),
    .ZN(_10681_));
 NAND2_X1 _20344_ (.A1(_09140_),
    .A2(_09585_),
    .ZN(_10682_));
 OAI21_X1 _20345_ (.A(_07117_),
    .B1(_10682_),
    .B2(_09142_),
    .ZN(_10683_));
 OAI21_X1 _20346_ (.A(_07532_),
    .B1(_08500_),
    .B2(_08539_),
    .ZN(_10684_));
 OAI21_X1 _20347_ (.A(_06963_),
    .B1(_09131_),
    .B2(_07205_),
    .ZN(_10685_));
 AND3_X1 _20348_ (.A1(_10683_),
    .A2(_10684_),
    .A3(_10685_),
    .ZN(_10686_));
 OAI21_X1 _20349_ (.A(_07326_),
    .B1(_10285_),
    .B2(_10038_),
    .ZN(_10687_));
 OAI21_X1 _20350_ (.A(_09144_),
    .B1(_09192_),
    .B2(_08299_),
    .ZN(_10688_));
 AND4_X1 _20351_ (.A1(_09201_),
    .A2(_10011_),
    .A3(_10687_),
    .A4(_10688_),
    .ZN(_10689_));
 NAND4_X2 _20352_ (.A1(_10679_),
    .A2(_10681_),
    .A3(_10686_),
    .A4(_10689_),
    .ZN(_10690_));
 AOI21_X1 _20353_ (.A(_09545_),
    .B1(_08321_),
    .B2(_07576_),
    .ZN(_10691_));
 AOI21_X1 _20354_ (.A(_10691_),
    .B1(_07172_),
    .B2(_08157_),
    .ZN(_10692_));
 OAI211_X2 _20355_ (.A(_07172_),
    .B(_16791_),
    .C1(_08396_),
    .C2(_06776_),
    .ZN(_10693_));
 OAI21_X1 _20356_ (.A(_07905_),
    .B1(_07359_),
    .B2(_09131_),
    .ZN(_10694_));
 OAI21_X1 _20357_ (.A(_07905_),
    .B1(_07084_),
    .B2(_09166_),
    .ZN(_10695_));
 OAI21_X1 _20358_ (.A(_07905_),
    .B1(_06908_),
    .B2(_06655_),
    .ZN(_10696_));
 AND3_X1 _20359_ (.A1(_10694_),
    .A2(_10695_),
    .A3(_10696_),
    .ZN(_10697_));
 AND4_X1 _20360_ (.A1(_09212_),
    .A2(_10692_),
    .A3(_10693_),
    .A4(_10697_),
    .ZN(_10698_));
 AOI21_X1 _20361_ (.A(_09571_),
    .B1(_09187_),
    .B2(_10479_),
    .ZN(_10699_));
 AND2_X1 _20362_ (.A1(_06963_),
    .A2(_07392_),
    .ZN(_10700_));
 AND2_X1 _20363_ (.A1(_07392_),
    .A2(_07719_),
    .ZN(_10701_));
 NOR4_X1 _20364_ (.A1(_10699_),
    .A2(_10700_),
    .A3(_10701_),
    .A4(_10481_),
    .ZN(_10702_));
 AOI22_X1 _20365_ (.A1(_06908_),
    .A2(_09192_),
    .B1(_08190_),
    .B2(_08222_),
    .ZN(_10703_));
 AND3_X1 _20366_ (.A1(_09180_),
    .A2(_10061_),
    .A3(_10060_),
    .ZN(_10704_));
 AOI22_X1 _20367_ (.A1(_06963_),
    .A2(_09199_),
    .B1(_07927_),
    .B2(_07532_),
    .ZN(_10705_));
 AOI22_X1 _20368_ (.A1(_08544_),
    .A2(_06908_),
    .B1(_09142_),
    .B2(_07532_),
    .ZN(_10706_));
 AND4_X1 _20369_ (.A1(_10703_),
    .A2(_10704_),
    .A3(_10705_),
    .A4(_10706_),
    .ZN(_10707_));
 AOI22_X1 _20370_ (.A1(_08544_),
    .A2(_09166_),
    .B1(_07653_),
    .B2(_09133_),
    .ZN(_10708_));
 NAND2_X1 _20371_ (.A1(_08299_),
    .A2(_07565_),
    .ZN(_10709_));
 NAND3_X1 _20372_ (.A1(_07326_),
    .A2(_08222_),
    .A3(_09145_),
    .ZN(_10710_));
 NAND3_X1 _20373_ (.A1(_10708_),
    .A2(_10709_),
    .A3(_10710_),
    .ZN(_10711_));
 AOI21_X1 _20374_ (.A(_09163_),
    .B1(_08135_),
    .B2(_07370_),
    .ZN(_10712_));
 AOI21_X1 _20375_ (.A(_09163_),
    .B1(_09582_),
    .B2(_07850_),
    .ZN(_10713_));
 OAI21_X1 _20376_ (.A(_09607_),
    .B1(_07282_),
    .B2(_07348_),
    .ZN(_10714_));
 NOR4_X1 _20377_ (.A1(_10711_),
    .A2(_10712_),
    .A3(_10713_),
    .A4(_10714_),
    .ZN(_10715_));
 NAND4_X1 _20378_ (.A1(_10698_),
    .A2(_10702_),
    .A3(_10707_),
    .A4(_10715_),
    .ZN(_10716_));
 NOR2_X4 _20379_ (.A1(_10690_),
    .A2(_10716_),
    .ZN(_10717_));
 XOR2_X2 _20380_ (.A(_10669_),
    .B(_10717_),
    .Z(_10718_));
 AND2_X1 _20381_ (.A1(_10085_),
    .A2(_04855_),
    .ZN(_10719_));
 INV_X1 _20382_ (.A(_10719_),
    .ZN(_10720_));
 INV_X1 _20383_ (.A(_10434_),
    .ZN(_10721_));
 AND4_X1 _20384_ (.A1(_10072_),
    .A2(_10720_),
    .A3(_10721_),
    .A4(_10094_),
    .ZN(_10722_));
 NAND2_X1 _20385_ (.A1(_05709_),
    .A2(_04768_),
    .ZN(_10723_));
 OAI21_X1 _20386_ (.A(_10723_),
    .B1(_05214_),
    .B2(_09748_),
    .ZN(_10724_));
 AND2_X1 _20387_ (.A1(_05456_),
    .A2(_06303_),
    .ZN(_10725_));
 NOR4_X1 _20388_ (.A1(_10724_),
    .A2(_10071_),
    .A3(_10725_),
    .A4(_09519_),
    .ZN(_10726_));
 NAND2_X2 _20389_ (.A1(_04209_),
    .A2(_04976_),
    .ZN(_10727_));
 NAND2_X1 _20390_ (.A1(_05489_),
    .A2(_05188_),
    .ZN(_10728_));
 NAND2_X1 _20391_ (.A1(_09473_),
    .A2(_09482_),
    .ZN(_10729_));
 AND4_X1 _20392_ (.A1(_09716_),
    .A2(_10727_),
    .A3(_10728_),
    .A4(_10729_),
    .ZN(_10730_));
 AOI22_X1 _20393_ (.A1(_05489_),
    .A2(_09473_),
    .B1(_05200_),
    .B2(_09464_),
    .ZN(_10731_));
 NAND2_X1 _20394_ (.A1(_10085_),
    .A2(_05313_),
    .ZN(_10732_));
 AND3_X1 _20395_ (.A1(_10731_),
    .A2(_10732_),
    .A3(_10158_),
    .ZN(_10733_));
 AND4_X1 _20396_ (.A1(_10722_),
    .A2(_10726_),
    .A3(_10730_),
    .A4(_10733_),
    .ZN(_10734_));
 OAI22_X1 _20397_ (.A1(_05698_),
    .A2(_05214_),
    .B1(_10439_),
    .B2(_09475_),
    .ZN(_10735_));
 AOI221_X4 _20398_ (.A(_10735_),
    .B1(_05390_),
    .B2(_06072_),
    .C1(_06226_),
    .C2(_05180_),
    .ZN(_10736_));
 AND2_X1 _20399_ (.A1(_05056_),
    .A2(_06435_),
    .ZN(_10737_));
 AND2_X1 _20400_ (.A1(_05456_),
    .A2(_05009_),
    .ZN(_10738_));
 NOR4_X1 _20401_ (.A1(_09511_),
    .A2(_09456_),
    .A3(_10737_),
    .A4(_10738_),
    .ZN(_10739_));
 AND2_X1 _20402_ (.A1(_04483_),
    .A2(_05056_),
    .ZN(_10740_));
 AND2_X1 _20403_ (.A1(_06050_),
    .A2(_05085_),
    .ZN(_10741_));
 NOR4_X1 _20404_ (.A1(_05786_),
    .A2(_10740_),
    .A3(_09735_),
    .A4(_10741_),
    .ZN(_10742_));
 AND3_X1 _20405_ (.A1(_04877_),
    .A2(_05184_),
    .A3(_05018_),
    .ZN(_10743_));
 AND4_X1 _20406_ (.A1(_10736_),
    .A2(_10739_),
    .A3(_10742_),
    .A4(_10743_),
    .ZN(_10744_));
 AND2_X1 _20407_ (.A1(_10432_),
    .A2(_10445_),
    .ZN(_10745_));
 INV_X1 _20408_ (.A(_10156_),
    .ZN(_10746_));
 NAND2_X1 _20409_ (.A1(_05775_),
    .A2(_09701_),
    .ZN(_10747_));
 AOI21_X1 _20410_ (.A(_10453_),
    .B1(_06226_),
    .B2(_05313_),
    .ZN(_10748_));
 NAND4_X1 _20411_ (.A1(_10745_),
    .A2(_10746_),
    .A3(_10747_),
    .A4(_10748_),
    .ZN(_10749_));
 NAND4_X1 _20412_ (.A1(_05830_),
    .A2(_09755_),
    .A3(_10101_),
    .A4(_10104_),
    .ZN(_10750_));
 NOR4_X1 _20413_ (.A1(_10749_),
    .A2(_10750_),
    .A3(_09426_),
    .A4(_09703_),
    .ZN(_10751_));
 OAI221_X1 _20414_ (.A(_05643_),
    .B1(_09515_),
    .B2(_06237_),
    .C1(_10084_),
    .C2(_10076_),
    .ZN(_10752_));
 AOI22_X1 _20415_ (.A1(_05357_),
    .A2(_10081_),
    .B1(_04768_),
    .B2(_09505_),
    .ZN(_10753_));
 NAND2_X1 _20416_ (.A1(_10085_),
    .A2(_09692_),
    .ZN(_10754_));
 OAI211_X2 _20417_ (.A(_10753_),
    .B(_10754_),
    .C1(_10204_),
    .C2(_05368_),
    .ZN(_10755_));
 NOR4_X1 _20418_ (.A1(_10752_),
    .A2(_09690_),
    .A3(_06545_),
    .A4(_10755_),
    .ZN(_10756_));
 NAND4_X1 _20419_ (.A1(_10734_),
    .A2(_10744_),
    .A3(_10751_),
    .A4(_10756_),
    .ZN(_10757_));
 NAND2_X1 _20420_ (.A1(_06380_),
    .A2(_06446_),
    .ZN(_10758_));
 AND2_X1 _20421_ (.A1(_04844_),
    .A2(_06138_),
    .ZN(_10759_));
 AOI221_X2 _20422_ (.A(_10759_),
    .B1(_06248_),
    .B2(_06050_),
    .C1(_04538_),
    .C2(_05247_),
    .ZN(_10760_));
 OAI21_X1 _20423_ (.A(_06061_),
    .B1(_09452_),
    .B2(_10081_),
    .ZN(_10761_));
 OAI21_X1 _20424_ (.A(_09482_),
    .B1(_05709_),
    .B2(_05188_),
    .ZN(_10762_));
 OAI21_X1 _20425_ (.A(_06446_),
    .B1(_04253_),
    .B2(_09507_),
    .ZN(_10763_));
 AND2_X1 _20426_ (.A1(_10762_),
    .A2(_10763_),
    .ZN(_10764_));
 AND4_X1 _20427_ (.A1(_10758_),
    .A2(_10760_),
    .A3(_10761_),
    .A4(_10764_),
    .ZN(_10765_));
 AND3_X1 _20428_ (.A1(_05302_),
    .A2(_05467_),
    .A3(_05676_),
    .ZN(_10766_));
 AND4_X1 _20429_ (.A1(_05500_),
    .A2(_05863_),
    .A3(_04494_),
    .A4(_05467_),
    .ZN(_10767_));
 AOI211_X4 _20430_ (.A(_10766_),
    .B(_10767_),
    .C1(_04538_),
    .C2(_05940_),
    .ZN(_10768_));
 AND2_X1 _20431_ (.A1(_09422_),
    .A2(_05940_),
    .ZN(_10769_));
 AND2_X4 _20432_ (.A1(_05940_),
    .A2(_09505_),
    .ZN(_10770_));
 NOR4_X1 _20433_ (.A1(_09418_),
    .A2(_10769_),
    .A3(_10770_),
    .A4(_06017_),
    .ZN(_10771_));
 OAI21_X1 _20434_ (.A(_09491_),
    .B1(_09507_),
    .B2(_10081_),
    .ZN(_10772_));
 OAI211_X2 _20435_ (.A(_09438_),
    .B(_06127_),
    .C1(_09692_),
    .C2(_05984_),
    .ZN(_10773_));
 NAND4_X1 _20436_ (.A1(_09438_),
    .A2(_05764_),
    .A3(_09468_),
    .A4(_06127_),
    .ZN(_10774_));
 AND3_X1 _20437_ (.A1(_10772_),
    .A2(_10773_),
    .A3(_10774_),
    .ZN(_10775_));
 NAND4_X1 _20438_ (.A1(_10765_),
    .A2(_10768_),
    .A3(_10771_),
    .A4(_10775_),
    .ZN(_10776_));
 NOR2_X4 _20439_ (.A1(_10757_),
    .A2(_10776_),
    .ZN(_10777_));
 XNOR2_X1 _20440_ (.A(_10564_),
    .B(_10777_),
    .ZN(_10778_));
 XNOR2_X1 _20441_ (.A(_10718_),
    .B(_10778_),
    .ZN(_10779_));
 OAI211_X2 _20442_ (.A(_09083_),
    .B(_10584_),
    .C1(_09897_),
    .C2(_09024_),
    .ZN(_10780_));
 AND3_X1 _20443_ (.A1(_09378_),
    .A2(_09057_),
    .A3(_08921_),
    .ZN(_10781_));
 AND2_X1 _20444_ (.A1(_09293_),
    .A2(_09081_),
    .ZN(_10782_));
 NOR2_X1 _20445_ (.A1(_10781_),
    .A2(_10782_),
    .ZN(_10783_));
 NAND2_X1 _20446_ (.A1(_09339_),
    .A2(_09318_),
    .ZN(_10784_));
 OAI211_X2 _20447_ (.A(_10783_),
    .B(_10784_),
    .C1(_09357_),
    .C2(_09070_),
    .ZN(_10785_));
 NAND3_X1 _20448_ (.A1(_09767_),
    .A2(_09352_),
    .A3(_09771_),
    .ZN(_10786_));
 OR2_X1 _20449_ (.A1(_09336_),
    .A2(_09337_),
    .ZN(_10787_));
 NOR4_X1 _20450_ (.A1(_10780_),
    .A2(_10785_),
    .A3(_10786_),
    .A4(_10787_),
    .ZN(_10788_));
 AND2_X1 _20451_ (.A1(_08899_),
    .A2(_09382_),
    .ZN(_10789_));
 AND2_X1 _20452_ (.A1(_08955_),
    .A2(_09005_),
    .ZN(_10790_));
 OR4_X1 _20453_ (.A1(_09383_),
    .A2(_10365_),
    .A3(_10789_),
    .A4(_10790_),
    .ZN(_10791_));
 AND3_X1 _20454_ (.A1(_08947_),
    .A2(_09017_),
    .A3(_08961_),
    .ZN(_10792_));
 OAI221_X1 _20455_ (.A(_10572_),
    .B1(_09794_),
    .B2(_09032_),
    .C1(_09071_),
    .C2(_09062_),
    .ZN(_10793_));
 AOI22_X1 _20456_ (.A1(_09392_),
    .A2(_08948_),
    .B1(_09318_),
    .B2(_09005_),
    .ZN(_10794_));
 OAI211_X2 _20457_ (.A(_09376_),
    .B(_10794_),
    .C1(_09349_),
    .C2(_09794_),
    .ZN(_10795_));
 NOR4_X1 _20458_ (.A1(_10791_),
    .A2(_10792_),
    .A3(_10793_),
    .A4(_10795_),
    .ZN(_10796_));
 INV_X1 _20459_ (.A(_10343_),
    .ZN(_10797_));
 AOI21_X1 _20460_ (.A(_09386_),
    .B1(_10352_),
    .B2(_10797_),
    .ZN(_10798_));
 AOI21_X1 _20461_ (.A(_09372_),
    .B1(_10605_),
    .B2(_09029_),
    .ZN(_10799_));
 AND3_X1 _20462_ (.A1(_09339_),
    .A2(_08977_),
    .A3(_08993_),
    .ZN(_10800_));
 NOR4_X1 _20463_ (.A1(_10798_),
    .A2(_10799_),
    .A3(_09883_),
    .A4(_10800_),
    .ZN(_10801_));
 INV_X1 _20464_ (.A(_09825_),
    .ZN(_10802_));
 OAI21_X1 _20465_ (.A(_09789_),
    .B1(_09832_),
    .B2(_09010_),
    .ZN(_10803_));
 NAND3_X1 _20466_ (.A1(_10802_),
    .A2(_10334_),
    .A3(_10803_),
    .ZN(_10804_));
 NAND2_X1 _20467_ (.A1(_09405_),
    .A2(_08926_),
    .ZN(_10805_));
 NAND3_X1 _20468_ (.A1(_10378_),
    .A2(_10340_),
    .A3(_10805_),
    .ZN(_10806_));
 AOI21_X1 _20469_ (.A(_10331_),
    .B1(_09024_),
    .B2(_09308_),
    .ZN(_10807_));
 AOI21_X1 _20470_ (.A(_09357_),
    .B1(_09061_),
    .B2(_08980_),
    .ZN(_10808_));
 NOR4_X1 _20471_ (.A1(_10804_),
    .A2(_10806_),
    .A3(_10807_),
    .A4(_10808_),
    .ZN(_10809_));
 AND4_X1 _20472_ (.A1(_10788_),
    .A2(_10796_),
    .A3(_10801_),
    .A4(_10809_),
    .ZN(_10810_));
 AND2_X1 _20473_ (.A1(_08906_),
    .A2(_08988_),
    .ZN(_10811_));
 AND2_X1 _20474_ (.A1(_09346_),
    .A2(_08924_),
    .ZN(_10812_));
 OR4_X1 _20475_ (.A1(_10589_),
    .A2(_10811_),
    .A3(_10568_),
    .A4(_10812_),
    .ZN(_10813_));
 AND2_X1 _20476_ (.A1(_09339_),
    .A2(_09331_),
    .ZN(_10814_));
 AND2_X1 _20477_ (.A1(_09081_),
    .A2(_09340_),
    .ZN(_10815_));
 INV_X1 _20478_ (.A(_10815_),
    .ZN(_10816_));
 OAI21_X1 _20479_ (.A(_09392_),
    .B1(_09079_),
    .B2(_09318_),
    .ZN(_10817_));
 NAND2_X1 _20480_ (.A1(_10816_),
    .A2(_10817_),
    .ZN(_10818_));
 OAI211_X2 _20481_ (.A(_09310_),
    .B(_09087_),
    .C1(_08962_),
    .C2(_09784_),
    .ZN(_10819_));
 NAND4_X1 _20482_ (.A1(_09310_),
    .A2(_08931_),
    .A3(_08993_),
    .A4(_08961_),
    .ZN(_10820_));
 NAND4_X1 _20483_ (.A1(_09389_),
    .A2(_10819_),
    .A3(_09390_),
    .A4(_10820_),
    .ZN(_10821_));
 NOR4_X1 _20484_ (.A1(_10813_),
    .A2(_10814_),
    .A3(_10818_),
    .A4(_10821_),
    .ZN(_10822_));
 INV_X1 _20485_ (.A(_09002_),
    .ZN(_10823_));
 OAI21_X1 _20486_ (.A(_09043_),
    .B1(_10823_),
    .B2(_09386_),
    .ZN(_10824_));
 NAND2_X1 _20487_ (.A1(_08893_),
    .A2(_08985_),
    .ZN(_10825_));
 NAND2_X1 _20488_ (.A1(_09047_),
    .A2(_10825_),
    .ZN(_10826_));
 AOI211_X4 _20489_ (.A(_10824_),
    .B(_10826_),
    .C1(_08959_),
    .C2(_08958_),
    .ZN(_10827_));
 NAND2_X1 _20490_ (.A1(_09079_),
    .A2(_08947_),
    .ZN(_10828_));
 NAND2_X1 _20491_ (.A1(_08969_),
    .A2(_08947_),
    .ZN(_10829_));
 AND2_X1 _20492_ (.A1(_10828_),
    .A2(_10829_),
    .ZN(_10830_));
 NAND2_X1 _20493_ (.A1(_09326_),
    .A2(_09404_),
    .ZN(_10831_));
 OAI21_X1 _20494_ (.A(_09397_),
    .B1(_09394_),
    .B2(_09010_),
    .ZN(_10832_));
 AND4_X1 _20495_ (.A1(_09028_),
    .A2(_10830_),
    .A3(_10831_),
    .A4(_10832_),
    .ZN(_10833_));
 OAI21_X1 _20496_ (.A(_09406_),
    .B1(_09062_),
    .B2(_09035_),
    .ZN(_10834_));
 NOR4_X1 _20497_ (.A1(_10834_),
    .A2(_09059_),
    .A3(_09321_),
    .A4(_09871_),
    .ZN(_10835_));
 AND4_X1 _20498_ (.A1(_10822_),
    .A2(_10827_),
    .A3(_10833_),
    .A4(_10835_),
    .ZN(_10836_));
 NAND2_X1 _20499_ (.A1(_10810_),
    .A2(_10836_),
    .ZN(_10837_));
 XNOR2_X1 _20500_ (.A(_10779_),
    .B(_10837_),
    .ZN(_10838_));
 XNOR2_X1 _20501_ (.A(_10838_),
    .B(_17172_),
    .ZN(_10839_));
 MUX2_X1 _20502_ (.A(_10619_),
    .B(_10839_),
    .S(_09100_),
    .Z(_00730_));
 OAI21_X1 _20503_ (.A(_06611_),
    .B1(_10003_),
    .B2(_07620_),
    .ZN(_10840_));
 OAI21_X1 _20504_ (.A(_08190_),
    .B1(_09188_),
    .B2(_07458_),
    .ZN(_10841_));
 NAND4_X1 _20505_ (.A1(_07883_),
    .A2(_08058_),
    .A3(_06875_),
    .A4(_06633_),
    .ZN(_10842_));
 OAI21_X1 _20506_ (.A(_07982_),
    .B1(_08124_),
    .B2(_07675_),
    .ZN(_10843_));
 AND3_X1 _20507_ (.A1(_10841_),
    .A2(_10842_),
    .A3(_10843_),
    .ZN(_10844_));
 AOI21_X1 _20508_ (.A(_08542_),
    .B1(_07576_),
    .B2(_08433_),
    .ZN(_10845_));
 AOI21_X1 _20509_ (.A(_08542_),
    .B1(_09167_),
    .B2(_07095_),
    .ZN(_10846_));
 AOI211_X2 _20510_ (.A(_10845_),
    .B(_10846_),
    .C1(_06952_),
    .C2(_08500_),
    .ZN(_10847_));
 AOI21_X1 _20511_ (.A(_09128_),
    .B1(_09567_),
    .B2(_09104_),
    .ZN(_10848_));
 AOI21_X1 _20512_ (.A(_10848_),
    .B1(_07795_),
    .B2(_10682_),
    .ZN(_10849_));
 AND3_X1 _20513_ (.A1(_07521_),
    .A2(_08386_),
    .A3(_07051_),
    .ZN(_10850_));
 NOR4_X1 _20514_ (.A1(_09152_),
    .A2(_10850_),
    .A3(_09155_),
    .A4(_10311_),
    .ZN(_10851_));
 AND4_X1 _20515_ (.A1(_10844_),
    .A2(_10847_),
    .A3(_10849_),
    .A4(_10851_),
    .ZN(_10852_));
 OAI21_X1 _20516_ (.A(_07905_),
    .B1(_07631_),
    .B2(_07565_),
    .ZN(_10853_));
 OAI21_X1 _20517_ (.A(_07894_),
    .B1(_09138_),
    .B2(_09106_),
    .ZN(_10854_));
 OAI21_X1 _20518_ (.A(_07894_),
    .B1(_07458_),
    .B2(_07227_),
    .ZN(_10855_));
 AND4_X1 _20519_ (.A1(_10492_),
    .A2(_10853_),
    .A3(_10854_),
    .A4(_10855_),
    .ZN(_10856_));
 OAI21_X1 _20520_ (.A(_07260_),
    .B1(_09106_),
    .B2(_09549_),
    .ZN(_10857_));
 OAI21_X1 _20521_ (.A(_07708_),
    .B1(_07751_),
    .B2(_09125_),
    .ZN(_10858_));
 OAI21_X1 _20522_ (.A(_07708_),
    .B1(_07359_),
    .B2(_07762_),
    .ZN(_10859_));
 OAI211_X2 _20523_ (.A(_07260_),
    .B(_08069_),
    .C1(_08538_),
    .C2(_07051_),
    .ZN(_10860_));
 AND4_X1 _20524_ (.A1(_10857_),
    .A2(_10858_),
    .A3(_10859_),
    .A4(_10860_),
    .ZN(_10861_));
 AND4_X2 _20525_ (.A1(_10840_),
    .A2(_10852_),
    .A3(_10856_),
    .A4(_10861_),
    .ZN(_10862_));
 AOI211_X4 _20526_ (.A(_06721_),
    .B(_07150_),
    .C1(_06644_),
    .C2(_08069_),
    .ZN(_10863_));
 OAI21_X1 _20527_ (.A(_07414_),
    .B1(_09131_),
    .B2(_07762_),
    .ZN(_10864_));
 OAI211_X2 _20528_ (.A(_10864_),
    .B(_09987_),
    .C1(_09163_),
    .C2(_09550_),
    .ZN(_10865_));
 NAND4_X1 _20529_ (.A1(_07740_),
    .A2(_06820_),
    .A3(_06842_),
    .A4(_06897_),
    .ZN(_10866_));
 OAI211_X2 _20530_ (.A(_09159_),
    .B(_10866_),
    .C1(_09104_),
    .C2(_07150_),
    .ZN(_10867_));
 AND2_X1 _20531_ (.A1(_07730_),
    .A2(_07051_),
    .ZN(_10868_));
 AND2_X1 _20532_ (.A1(_10868_),
    .A2(_06853_),
    .ZN(_10869_));
 NOR4_X2 _20533_ (.A1(_10863_),
    .A2(_10865_),
    .A3(_10867_),
    .A4(_10869_),
    .ZN(_10870_));
 NAND2_X1 _20534_ (.A1(_08544_),
    .A2(_06908_),
    .ZN(_10871_));
 OAI221_X1 _20535_ (.A(_07477_),
    .B1(_08396_),
    .B2(_07029_),
    .C1(_07740_),
    .C2(_07447_),
    .ZN(_10872_));
 OAI21_X1 _20536_ (.A(_07172_),
    .B1(_07293_),
    .B2(_07565_),
    .ZN(_10873_));
 AND4_X1 _20537_ (.A1(_10487_),
    .A2(_10871_),
    .A3(_10872_),
    .A4(_10873_),
    .ZN(_10874_));
 NAND3_X1 _20538_ (.A1(_09138_),
    .A2(_07960_),
    .A3(_08080_),
    .ZN(_10875_));
 OAI21_X1 _20539_ (.A(_09192_),
    .B1(_10471_),
    .B2(_09188_),
    .ZN(_10876_));
 OAI211_X2 _20540_ (.A(_07949_),
    .B(_07960_),
    .C1(_07359_),
    .C2(_09133_),
    .ZN(_10877_));
 OAI21_X1 _20541_ (.A(_07326_),
    .B1(_08343_),
    .B2(_08124_),
    .ZN(_10878_));
 AND4_X1 _20542_ (.A1(_10875_),
    .A2(_10876_),
    .A3(_10877_),
    .A4(_10878_),
    .ZN(_10879_));
 INV_X1 _20543_ (.A(_10282_),
    .ZN(_10880_));
 AND3_X1 _20544_ (.A1(_09576_),
    .A2(_10048_),
    .A3(_09181_),
    .ZN(_10881_));
 OAI21_X1 _20545_ (.A(_07117_),
    .B1(_10868_),
    .B2(_06908_),
    .ZN(_10882_));
 OAI21_X1 _20546_ (.A(_08549_),
    .B1(_09144_),
    .B2(_07828_),
    .ZN(_10883_));
 AND4_X1 _20547_ (.A1(_10880_),
    .A2(_10881_),
    .A3(_10882_),
    .A4(_10883_),
    .ZN(_10884_));
 AND4_X1 _20548_ (.A1(_10870_),
    .A2(_10874_),
    .A3(_10879_),
    .A4(_10884_),
    .ZN(_10885_));
 AND2_X4 _20549_ (.A1(_10862_),
    .A2(_10885_),
    .ZN(_10886_));
 AND2_X1 _20550_ (.A1(_06424_),
    .A2(_10078_),
    .ZN(_10887_));
 OR2_X2 _20551_ (.A1(_10119_),
    .A2(_10887_),
    .ZN(_10888_));
 AOI211_X2 _20552_ (.A(_09498_),
    .B(_10888_),
    .C1(_04801_),
    .C2(_06435_),
    .ZN(_10889_));
 OAI21_X1 _20553_ (.A(_06226_),
    .B1(_06391_),
    .B2(_05313_),
    .ZN(_10890_));
 OAI211_X2 _20554_ (.A(_06226_),
    .B(_09468_),
    .C1(_10076_),
    .C2(_05522_),
    .ZN(_10891_));
 OAI221_X1 _20555_ (.A(_06226_),
    .B1(_10076_),
    .B2(_05753_),
    .C1(_09701_),
    .C2(_06270_),
    .ZN(_10892_));
 AND4_X2 _20556_ (.A1(_10889_),
    .A2(_10890_),
    .A3(_10891_),
    .A4(_10892_),
    .ZN(_10893_));
 OAI21_X1 _20557_ (.A(_09491_),
    .B1(_04976_),
    .B2(_05085_),
    .ZN(_10894_));
 NAND4_X1 _20558_ (.A1(_10449_),
    .A2(_10196_),
    .A3(_10133_),
    .A4(_10894_),
    .ZN(_10895_));
 NAND3_X1 _20559_ (.A1(_06149_),
    .A2(_09468_),
    .A3(_04395_),
    .ZN(_10896_));
 OAI211_X2 _20560_ (.A(_10896_),
    .B(_09747_),
    .C1(_05995_),
    .C2(_09748_),
    .ZN(_10897_));
 AOI21_X1 _20561_ (.A(_09748_),
    .B1(_10204_),
    .B2(_05731_),
    .ZN(_10898_));
 NOR4_X1 _20562_ (.A1(_10895_),
    .A2(_10139_),
    .A3(_10897_),
    .A4(_10898_),
    .ZN(_10899_));
 NOR4_X1 _20563_ (.A1(_05951_),
    .A2(_09419_),
    .A3(_10770_),
    .A4(_10766_),
    .ZN(_10900_));
 OAI221_X1 _20564_ (.A(_05841_),
    .B1(_05511_),
    .B2(_05753_),
    .C1(_06270_),
    .C2(_09441_),
    .ZN(_10901_));
 AND3_X2 _20565_ (.A1(_10900_),
    .A2(_10432_),
    .A3(_10901_),
    .ZN(_10902_));
 AOI21_X1 _20566_ (.A(_05698_),
    .B1(_10203_),
    .B2(_10438_),
    .ZN(_10903_));
 NAND2_X1 _20567_ (.A1(_06380_),
    .A2(_06050_),
    .ZN(_10904_));
 OAI221_X1 _20568_ (.A(_10904_),
    .B1(_10439_),
    .B2(_05214_),
    .C1(_04395_),
    .C2(_09722_),
    .ZN(_10905_));
 AND4_X1 _20569_ (.A1(_10076_),
    .A2(_09438_),
    .A3(_09468_),
    .A4(_05863_),
    .ZN(_10906_));
 AND4_X1 _20570_ (.A1(_05522_),
    .A2(_09438_),
    .A3(_05863_),
    .A4(_05500_),
    .ZN(_10907_));
 NOR4_X1 _20571_ (.A1(_10903_),
    .A2(_10905_),
    .A3(_10906_),
    .A4(_10907_),
    .ZN(_10908_));
 NAND4_X1 _20572_ (.A1(_10893_),
    .A2(_10899_),
    .A3(_10902_),
    .A4(_10908_),
    .ZN(_10909_));
 OAI21_X1 _20573_ (.A(_09444_),
    .B1(_05188_),
    .B2(_05335_),
    .ZN(_10910_));
 AND2_X1 _20574_ (.A1(_04198_),
    .A2(_06391_),
    .ZN(_10911_));
 AOI211_X2 _20575_ (.A(_09457_),
    .B(_10911_),
    .C1(_04209_),
    .C2(_10130_),
    .ZN(_10912_));
 OAI211_X2 _20576_ (.A(_09444_),
    .B(_09441_),
    .C1(_05511_),
    .C2(_05764_),
    .ZN(_10913_));
 AND4_X2 _20577_ (.A1(_10416_),
    .A2(_09705_),
    .A3(_09706_),
    .A4(_10727_),
    .ZN(_10914_));
 AND4_X2 _20578_ (.A1(_10910_),
    .A2(_10912_),
    .A3(_10913_),
    .A4(_10914_),
    .ZN(_10915_));
 OAI21_X1 _20579_ (.A(_10085_),
    .B1(_09743_),
    .B2(_04921_),
    .ZN(_10916_));
 NAND2_X1 _20580_ (.A1(_10085_),
    .A2(_04549_),
    .ZN(_10917_));
 NAND4_X1 _20581_ (.A1(_10916_),
    .A2(_10917_),
    .A3(_10732_),
    .A4(_05190_),
    .ZN(_10918_));
 OAI211_X2 _20582_ (.A(_10172_),
    .B(_10728_),
    .C1(_09512_),
    .C2(_09496_),
    .ZN(_10919_));
 NOR4_X1 _20583_ (.A1(_10918_),
    .A2(_10919_),
    .A3(_09511_),
    .A4(_10170_),
    .ZN(_10920_));
 OAI21_X1 _20584_ (.A(_05555_),
    .B1(_05056_),
    .B2(_06380_),
    .ZN(_10921_));
 NAND4_X1 _20585_ (.A1(_05202_),
    .A2(_09438_),
    .A3(_05198_),
    .A4(_04779_),
    .ZN(_10922_));
 AND2_X1 _20586_ (.A1(_10921_),
    .A2(_10922_),
    .ZN(_10923_));
 OAI21_X1 _20587_ (.A(_05599_),
    .B1(_09434_),
    .B2(_04976_),
    .ZN(_10924_));
 OAI21_X1 _20588_ (.A(_05357_),
    .B1(_05709_),
    .B2(_05188_),
    .ZN(_10925_));
 OAI21_X1 _20589_ (.A(_05357_),
    .B1(_09505_),
    .B2(_06314_),
    .ZN(_10926_));
 AND4_X1 _20590_ (.A1(_10923_),
    .A2(_10924_),
    .A3(_10925_),
    .A4(_10926_),
    .ZN(_10927_));
 OAI21_X1 _20591_ (.A(_09464_),
    .B1(_09505_),
    .B2(_10078_),
    .ZN(_10928_));
 OAI21_X1 _20592_ (.A(_04768_),
    .B1(_04888_),
    .B2(_09507_),
    .ZN(_10929_));
 OAI21_X1 _20593_ (.A(_04768_),
    .B1(_04417_),
    .B2(_04801_),
    .ZN(_10930_));
 OAI211_X2 _20594_ (.A(_09464_),
    .B(_05522_),
    .C1(_09468_),
    .C2(_05500_),
    .ZN(_10931_));
 AND4_X1 _20595_ (.A1(_10928_),
    .A2(_10929_),
    .A3(_10930_),
    .A4(_10931_),
    .ZN(_10932_));
 NAND4_X2 _20596_ (.A1(_10915_),
    .A2(_10920_),
    .A3(_10927_),
    .A4(_10932_),
    .ZN(_10933_));
 NOR2_X4 _20597_ (.A1(_10909_),
    .A2(_10933_),
    .ZN(_10934_));
 XOR2_X2 _20598_ (.A(_10886_),
    .B(_10934_),
    .Z(_10935_));
 AND2_X1 _20599_ (.A1(_09339_),
    .A2(_09364_),
    .ZN(_10936_));
 OR4_X1 _20600_ (.A1(_09085_),
    .A2(_10364_),
    .A3(_10814_),
    .A4(_10936_),
    .ZN(_10937_));
 AND2_X1 _20601_ (.A1(_09074_),
    .A2(_08969_),
    .ZN(_10938_));
 AOI211_X2 _20602_ (.A(_10938_),
    .B(_09847_),
    .C1(_09074_),
    .C2(_10343_),
    .ZN(_10939_));
 OAI211_X2 _20603_ (.A(_10939_),
    .B(_09073_),
    .C1(_09357_),
    .C2(_10578_),
    .ZN(_10940_));
 AND2_X1 _20604_ (.A1(_10397_),
    .A2(_08956_),
    .ZN(_10941_));
 AND2_X1 _20605_ (.A1(_09058_),
    .A2(_09051_),
    .ZN(_10942_));
 OR4_X1 _20606_ (.A1(_09852_),
    .A2(_10941_),
    .A3(_09851_),
    .A4(_10942_),
    .ZN(_10943_));
 OAI21_X1 _20607_ (.A(_09797_),
    .B1(_09374_),
    .B2(_08924_),
    .ZN(_10944_));
 NAND4_X1 _20608_ (.A1(_09797_),
    .A2(_08931_),
    .A3(_09355_),
    .A4(_08993_),
    .ZN(_10945_));
 OAI21_X1 _20609_ (.A(_09797_),
    .B1(_09404_),
    .B2(_08987_),
    .ZN(_10946_));
 NAND4_X1 _20610_ (.A1(_10816_),
    .A2(_10944_),
    .A3(_10945_),
    .A4(_10946_),
    .ZN(_10947_));
 NOR4_X1 _20611_ (.A1(_10937_),
    .A2(_10940_),
    .A3(_10943_),
    .A4(_10947_),
    .ZN(_10948_));
 AND3_X1 _20612_ (.A1(_09002_),
    .A2(_08945_),
    .A3(_08905_),
    .ZN(_10949_));
 AND3_X1 _20613_ (.A1(_09309_),
    .A2(_08931_),
    .A3(_09329_),
    .ZN(_10950_));
 AOI211_X4 _20614_ (.A(_10949_),
    .B(_10950_),
    .C1(_10343_),
    .C2(_09329_),
    .ZN(_10951_));
 NAND2_X1 _20615_ (.A1(_09327_),
    .A2(_09404_),
    .ZN(_10952_));
 AND4_X1 _20616_ (.A1(_10330_),
    .A2(_10333_),
    .A3(_09363_),
    .A4(_10952_),
    .ZN(_10953_));
 NAND2_X1 _20617_ (.A1(_09354_),
    .A2(_09394_),
    .ZN(_10954_));
 AND2_X1 _20618_ (.A1(_09354_),
    .A2(_09018_),
    .ZN(_10955_));
 INV_X1 _20619_ (.A(_10955_),
    .ZN(_10956_));
 OAI211_X2 _20620_ (.A(_08921_),
    .B(_08905_),
    .C1(_09374_),
    .C2(_08924_),
    .ZN(_10957_));
 AND4_X1 _20621_ (.A1(_10954_),
    .A2(_10956_),
    .A3(_09365_),
    .A4(_10957_),
    .ZN(_10958_));
 AND2_X1 _20622_ (.A1(_09326_),
    .A2(_08899_),
    .ZN(_10959_));
 INV_X1 _20623_ (.A(_10959_),
    .ZN(_10960_));
 AND4_X1 _20624_ (.A1(_10960_),
    .A2(_08936_),
    .A3(_08941_),
    .A4(_09298_),
    .ZN(_10961_));
 AND4_X1 _20625_ (.A1(_10951_),
    .A2(_10953_),
    .A3(_10958_),
    .A4(_10961_),
    .ZN(_10962_));
 NAND2_X1 _20626_ (.A1(_08910_),
    .A2(_09310_),
    .ZN(_10963_));
 AND3_X1 _20627_ (.A1(_10963_),
    .A2(_09781_),
    .A3(_08970_),
    .ZN(_10964_));
 OAI211_X2 _20628_ (.A(_09310_),
    .B(_09355_),
    .C1(_08954_),
    .C2(_08918_),
    .ZN(_10965_));
 NAND4_X1 _20629_ (.A1(_10964_),
    .A2(_10347_),
    .A3(_10349_),
    .A4(_10965_),
    .ZN(_10966_));
 OAI211_X2 _20630_ (.A(_09894_),
    .B(_09895_),
    .C1(_09897_),
    .C2(_09407_),
    .ZN(_10967_));
 OAI21_X1 _20631_ (.A(_09789_),
    .B1(_08987_),
    .B2(_09340_),
    .ZN(_10968_));
 NAND2_X1 _20632_ (.A1(_09789_),
    .A2(_08985_),
    .ZN(_10969_));
 OAI211_X2 _20633_ (.A(_10968_),
    .B(_10969_),
    .C1(_09067_),
    .C2(_08992_),
    .ZN(_10970_));
 OAI211_X2 _20634_ (.A(_09377_),
    .B(_08961_),
    .C1(_09017_),
    .C2(_08918_),
    .ZN(_10971_));
 NAND2_X1 _20635_ (.A1(_09318_),
    .A2(_09377_),
    .ZN(_10972_));
 OAI211_X2 _20636_ (.A(_10971_),
    .B(_10972_),
    .C1(_09066_),
    .C2(_09008_),
    .ZN(_10973_));
 NOR4_X1 _20637_ (.A1(_10966_),
    .A2(_10967_),
    .A3(_10970_),
    .A4(_10973_),
    .ZN(_10974_));
 OAI21_X1 _20638_ (.A(_09405_),
    .B1(_09002_),
    .B2(_10343_),
    .ZN(_10975_));
 OAI21_X1 _20639_ (.A(_09405_),
    .B1(_09374_),
    .B2(_09051_),
    .ZN(_10976_));
 NAND4_X1 _20640_ (.A1(_08950_),
    .A2(_09355_),
    .A3(_08962_),
    .A4(_09015_),
    .ZN(_10977_));
 AND3_X1 _20641_ (.A1(_10975_),
    .A2(_10976_),
    .A3(_10977_),
    .ZN(_10978_));
 NAND2_X1 _20642_ (.A1(_09028_),
    .A2(_09395_),
    .ZN(_10979_));
 NOR4_X1 _20643_ (.A1(_10979_),
    .A2(_09859_),
    .A3(_09019_),
    .A4(_09291_),
    .ZN(_10980_));
 INV_X1 _20644_ (.A(_09818_),
    .ZN(_10981_));
 OAI21_X1 _20645_ (.A(_09053_),
    .B1(_08919_),
    .B2(_08985_),
    .ZN(_10982_));
 AND4_X1 _20646_ (.A1(_10981_),
    .A2(_10982_),
    .A3(_09040_),
    .A4(_09869_),
    .ZN(_10983_));
 OAI21_X1 _20647_ (.A(_09397_),
    .B1(_09002_),
    .B2(_09293_),
    .ZN(_10984_));
 OAI211_X2 _20648_ (.A(_09397_),
    .B(_09355_),
    .C1(_09054_),
    .C2(_09784_),
    .ZN(_10985_));
 AND2_X1 _20649_ (.A1(_10984_),
    .A2(_10985_),
    .ZN(_10986_));
 AND4_X1 _20650_ (.A1(_10978_),
    .A2(_10980_),
    .A3(_10983_),
    .A4(_10986_),
    .ZN(_10987_));
 NAND4_X1 _20651_ (.A1(_10948_),
    .A2(_10962_),
    .A3(_10974_),
    .A4(_10987_),
    .ZN(_10988_));
 NOR2_X4 _20652_ (.A1(_10988_),
    .A2(_09825_),
    .ZN(_10989_));
 XOR2_X1 _20653_ (.A(_10935_),
    .B(_10989_),
    .Z(_10990_));
 XNOR2_X1 _20654_ (.A(_10669_),
    .B(_08887_),
    .ZN(_10991_));
 OAI21_X1 _20655_ (.A(_09098_),
    .B1(_10990_),
    .B2(_10991_),
    .ZN(_10992_));
 AOI21_X1 _20656_ (.A(_10992_),
    .B1(_10991_),
    .B2(_10990_),
    .ZN(_10993_));
 AND2_X1 _20657_ (.A1(_01331_),
    .A2(_17117_),
    .ZN(_10994_));
 NOR2_X1 _20658_ (.A1(_10993_),
    .A2(_10994_),
    .ZN(_10995_));
 XNOR2_X1 _20659_ (.A(_10995_),
    .B(_17173_),
    .ZN(_00731_));
 BUF_X4 _20660_ (.A(_17174_),
    .Z(_10996_));
 BUF_X4 _20661_ (.A(_10996_),
    .Z(_10997_));
 XOR2_X1 _20662_ (.A(_17128_),
    .B(_10997_),
    .Z(_10998_));
 XOR2_X1 _20663_ (.A(_08787_),
    .B(_08560_),
    .Z(_10999_));
 XNOR2_X1 _20664_ (.A(_10934_),
    .B(_01049_),
    .ZN(_11000_));
 XNOR2_X1 _20665_ (.A(_10999_),
    .B(_11000_),
    .ZN(_11001_));
 XOR2_X1 _20666_ (.A(_11001_),
    .B(_09413_),
    .Z(_11002_));
 MUX2_X1 _20667_ (.A(_10998_),
    .B(_11002_),
    .S(_09100_),
    .Z(_00692_));
 BUF_X4 _20668_ (.A(_17175_),
    .Z(_11003_));
 BUF_X4 _20669_ (.A(_11003_),
    .Z(_11004_));
 XOR2_X1 _20670_ (.A(_11004_),
    .B(_17139_),
    .Z(_11005_));
 XOR2_X2 _20671_ (.A(_06567_),
    .B(_10934_),
    .Z(_11006_));
 XNOR2_X2 _20672_ (.A(_09288_),
    .B(_11006_),
    .ZN(_11007_));
 XNOR2_X1 _20673_ (.A(_09413_),
    .B(_09838_),
    .ZN(_11008_));
 XNOR2_X2 _20674_ (.A(_11007_),
    .B(_11008_),
    .ZN(_11009_));
 INV_X1 _20675_ (.A(_17175_),
    .ZN(_11010_));
 BUF_X4 _20676_ (.A(_11010_),
    .Z(_11011_));
 XNOR2_X1 _20677_ (.A(_11009_),
    .B(_11011_),
    .ZN(_11012_));
 MUX2_X1 _20678_ (.A(_11005_),
    .B(_11012_),
    .S(_09100_),
    .Z(_00693_));
 XOR2_X1 _20679_ (.A(_17145_),
    .B(_17023_),
    .Z(_11013_));
 XNOR2_X2 _20680_ (.A(_09528_),
    .B(_09837_),
    .ZN(_11014_));
 XOR2_X1 _20681_ (.A(_09685_),
    .B(_11014_),
    .Z(_11015_));
 XNOR2_X1 _20682_ (.A(_11015_),
    .B(_09914_),
    .ZN(_11016_));
 XNOR2_X1 _20683_ (.A(_11016_),
    .B(_17145_),
    .ZN(_11017_));
 MUX2_X1 _20684_ (.A(_11013_),
    .B(_11017_),
    .S(_09100_),
    .Z(_00694_));
 XOR2_X1 _20685_ (.A(_17146_),
    .B(_17034_),
    .Z(_11018_));
 XNOR2_X1 _20686_ (.A(_10934_),
    .B(_09763_),
    .ZN(_11019_));
 XNOR2_X1 _20687_ (.A(_11019_),
    .B(_10401_),
    .ZN(_11020_));
 XNOR2_X1 _20688_ (.A(_10067_),
    .B(_11020_),
    .ZN(_11021_));
 XNOR2_X1 _20689_ (.A(_11021_),
    .B(_17146_),
    .ZN(_11022_));
 BUF_X4 _20690_ (.A(_09099_),
    .Z(_11023_));
 MUX2_X1 _20691_ (.A(_11018_),
    .B(_11022_),
    .S(_11023_),
    .Z(_00695_));
 XOR2_X1 _20692_ (.A(_17147_),
    .B(_17043_),
    .Z(_11024_));
 XOR2_X2 _20693_ (.A(_10934_),
    .B(_10148_),
    .Z(_11025_));
 XNOR2_X1 _20694_ (.A(_10328_),
    .B(_11025_),
    .ZN(_11026_));
 XNOR2_X1 _20695_ (.A(_10402_),
    .B(_10616_),
    .ZN(_11027_));
 XNOR2_X1 _20696_ (.A(_11026_),
    .B(_11027_),
    .ZN(_11028_));
 INV_X1 _20697_ (.A(_17147_),
    .ZN(_11029_));
 XNOR2_X1 _20698_ (.A(_11028_),
    .B(_11029_),
    .ZN(_11030_));
 MUX2_X1 _20699_ (.A(_11024_),
    .B(_11030_),
    .S(_11023_),
    .Z(_00696_));
 XOR2_X1 _20700_ (.A(_17148_),
    .B(_17044_),
    .Z(_11031_));
 XNOR2_X1 _20701_ (.A(_10616_),
    .B(_10212_),
    .ZN(_11032_));
 XNOR2_X1 _20702_ (.A(_11032_),
    .B(_10837_),
    .ZN(_11033_));
 XNOR2_X1 _20703_ (.A(_11033_),
    .B(_10565_),
    .ZN(_11034_));
 INV_X1 _20704_ (.A(_17148_),
    .ZN(_11035_));
 XNOR2_X1 _20705_ (.A(_11034_),
    .B(_11035_),
    .ZN(_11036_));
 MUX2_X1 _20706_ (.A(_11031_),
    .B(_11036_),
    .S(_11023_),
    .Z(_00697_));
 XOR2_X1 _20707_ (.A(_17149_),
    .B(_17045_),
    .Z(_11037_));
 XOR2_X1 _20708_ (.A(_10465_),
    .B(_10837_),
    .Z(_11038_));
 XNOR2_X1 _20709_ (.A(_10718_),
    .B(_11038_),
    .ZN(_11039_));
 XNOR2_X1 _20710_ (.A(_11039_),
    .B(_10989_),
    .ZN(_11040_));
 INV_X1 _20711_ (.A(_17149_),
    .ZN(_11041_));
 XNOR2_X1 _20712_ (.A(_11040_),
    .B(_11041_),
    .ZN(_11042_));
 MUX2_X1 _20713_ (.A(_11037_),
    .B(_11042_),
    .S(_11023_),
    .Z(_00698_));
 XOR2_X1 _20714_ (.A(_17150_),
    .B(_17046_),
    .Z(_11043_));
 XNOR2_X1 _20715_ (.A(_10777_),
    .B(_08887_),
    .ZN(_11044_));
 XNOR2_X1 _20716_ (.A(_11044_),
    .B(_10886_),
    .ZN(_11045_));
 XNOR2_X1 _20717_ (.A(_10989_),
    .B(_09093_),
    .ZN(_11046_));
 XNOR2_X1 _20718_ (.A(_11045_),
    .B(_11046_),
    .ZN(_11047_));
 XNOR2_X1 _20719_ (.A(_11047_),
    .B(_17150_),
    .ZN(_11048_));
 MUX2_X1 _20720_ (.A(_11043_),
    .B(_11048_),
    .S(_11023_),
    .Z(_00699_));
 BUF_X4 _20721_ (.A(_17151_),
    .Z(_11049_));
 BUF_X4 _20722_ (.A(_11049_),
    .Z(_11050_));
 XOR2_X1 _20723_ (.A(_17047_),
    .B(_11050_),
    .Z(_11051_));
 XOR2_X1 _20724_ (.A(_06567_),
    .B(_01050_),
    .Z(_11052_));
 XNOR2_X1 _20725_ (.A(_10935_),
    .B(_11052_),
    .ZN(_11053_));
 XOR2_X1 _20726_ (.A(_09412_),
    .B(_08787_),
    .Z(_11054_));
 XNOR2_X1 _20727_ (.A(_11053_),
    .B(_11054_),
    .ZN(_11055_));
 MUX2_X1 _20728_ (.A(_11051_),
    .B(_11055_),
    .S(_11023_),
    .Z(_00660_));
 BUF_X4 _20729_ (.A(_17152_),
    .Z(_11056_));
 XOR2_X1 _20730_ (.A(_17048_),
    .B(_11056_),
    .Z(_11057_));
 XNOR2_X1 _20731_ (.A(_11006_),
    .B(_11014_),
    .ZN(_11058_));
 XNOR2_X1 _20732_ (.A(_10886_),
    .B(_08560_),
    .ZN(_11059_));
 XNOR2_X1 _20733_ (.A(_09287_),
    .B(_01051_),
    .ZN(_11060_));
 XNOR2_X1 _20734_ (.A(_11059_),
    .B(_11060_),
    .ZN(_11061_));
 XNOR2_X1 _20735_ (.A(_11058_),
    .B(_11061_),
    .ZN(_11062_));
 MUX2_X1 _20736_ (.A(_11057_),
    .B(_11062_),
    .S(_11023_),
    .Z(_00661_));
 XOR2_X1 _20737_ (.A(_17153_),
    .B(_17049_),
    .Z(_11063_));
 XOR2_X1 _20738_ (.A(_09763_),
    .B(_09684_),
    .Z(_11064_));
 XNOR2_X1 _20739_ (.A(_11064_),
    .B(_09914_),
    .ZN(_11065_));
 XNOR2_X1 _20740_ (.A(_09213_),
    .B(_09528_),
    .ZN(_11066_));
 XNOR2_X1 _20741_ (.A(_11065_),
    .B(_11066_),
    .ZN(_11067_));
 INV_X32 _20742_ (.A(_17153_),
    .ZN(_11068_));
 XNOR2_X1 _20743_ (.A(_11067_),
    .B(_11068_),
    .ZN(_11069_));
 MUX2_X1 _20744_ (.A(_11063_),
    .B(_11069_),
    .S(_11023_),
    .Z(_00662_));
 XOR2_X1 _20745_ (.A(_17154_),
    .B(_17050_),
    .Z(_11070_));
 XNOR2_X2 _20746_ (.A(_09616_),
    .B(_10886_),
    .ZN(_11071_));
 XNOR2_X1 _20747_ (.A(_11071_),
    .B(_09986_),
    .ZN(_11072_));
 XNOR2_X2 _20748_ (.A(_11019_),
    .B(_10148_),
    .ZN(_11073_));
 XNOR2_X2 _20749_ (.A(_11072_),
    .B(_11073_),
    .ZN(_11074_));
 XNOR2_X1 _20750_ (.A(_11074_),
    .B(_10401_),
    .ZN(_11075_));
 INV_X1 _20751_ (.A(_17154_),
    .ZN(_11076_));
 XNOR2_X1 _20752_ (.A(_11075_),
    .B(_11076_),
    .ZN(_11077_));
 MUX2_X1 _20753_ (.A(_11070_),
    .B(_11077_),
    .S(_11023_),
    .Z(_00663_));
 XOR2_X1 _20754_ (.A(_17156_),
    .B(_17052_),
    .Z(_11078_));
 XOR2_X1 _20755_ (.A(_10270_),
    .B(_10212_),
    .Z(_11079_));
 XNOR2_X1 _20756_ (.A(_11079_),
    .B(_10616_),
    .ZN(_11080_));
 XNOR2_X1 _20757_ (.A(_10886_),
    .B(_10065_),
    .ZN(_11081_));
 XNOR2_X1 _20758_ (.A(_11025_),
    .B(_11081_),
    .ZN(_11082_));
 XNOR2_X1 _20759_ (.A(_11080_),
    .B(_11082_),
    .ZN(_11083_));
 XNOR2_X1 _20760_ (.A(_11083_),
    .B(_17156_),
    .ZN(_11084_));
 MUX2_X1 _20761_ (.A(_11078_),
    .B(_11084_),
    .S(_11023_),
    .Z(_00664_));
 XOR2_X1 _20762_ (.A(_17053_),
    .B(_17157_),
    .Z(_11085_));
 XNOR2_X1 _20763_ (.A(_10837_),
    .B(_10212_),
    .ZN(_11086_));
 XNOR2_X1 _20764_ (.A(_11086_),
    .B(_10564_),
    .ZN(_11087_));
 XNOR2_X1 _20765_ (.A(_10327_),
    .B(_01052_),
    .ZN(_11088_));
 XNOR2_X1 _20766_ (.A(_10465_),
    .B(_11088_),
    .ZN(_11089_));
 XNOR2_X1 _20767_ (.A(_11087_),
    .B(_11089_),
    .ZN(_11090_));
 BUF_X4 _20768_ (.A(_09099_),
    .Z(_11091_));
 MUX2_X1 _20769_ (.A(_11085_),
    .B(_11090_),
    .S(_11091_),
    .Z(_00665_));
 XOR2_X1 _20770_ (.A(_17054_),
    .B(_17158_),
    .Z(_11092_));
 XOR2_X1 _20771_ (.A(_10669_),
    .B(_10465_),
    .Z(_11093_));
 XNOR2_X1 _20772_ (.A(_11093_),
    .B(_10989_),
    .ZN(_11094_));
 XNOR2_X1 _20773_ (.A(_10514_),
    .B(_01053_),
    .ZN(_11095_));
 XNOR2_X1 _20774_ (.A(_11095_),
    .B(_10777_),
    .ZN(_11096_));
 XNOR2_X1 _20775_ (.A(_11094_),
    .B(_11096_),
    .ZN(_11097_));
 MUX2_X1 _20776_ (.A(_11092_),
    .B(_11097_),
    .S(_11091_),
    .Z(_00666_));
 XOR2_X1 _20777_ (.A(_17159_),
    .B(_17055_),
    .Z(_11098_));
 XNOR2_X1 _20778_ (.A(_10717_),
    .B(_10934_),
    .ZN(_11099_));
 XNOR2_X1 _20779_ (.A(_11099_),
    .B(_11044_),
    .ZN(_11100_));
 XNOR2_X1 _20780_ (.A(_11100_),
    .B(_09093_),
    .ZN(_11101_));
 XNOR2_X1 _20781_ (.A(_11101_),
    .B(_17159_),
    .ZN(_11102_));
 MUX2_X1 _20782_ (.A(_11098_),
    .B(_11102_),
    .S(_11091_),
    .Z(_00667_));
 BUF_X32 _20783_ (.A(_17160_),
    .Z(_11103_));
 BUF_X4 _20784_ (.A(_11103_),
    .Z(_11104_));
 BUF_X4 _20785_ (.A(_11104_),
    .Z(_11105_));
 XOR2_X1 _20786_ (.A(_17056_),
    .B(_11105_),
    .Z(_11106_));
 XNOR2_X1 _20787_ (.A(_06567_),
    .B(_08887_),
    .ZN(_11107_));
 XOR2_X1 _20788_ (.A(_11107_),
    .B(_09412_),
    .Z(_11108_));
 XNOR2_X1 _20789_ (.A(_11059_),
    .B(_01054_),
    .ZN(_11109_));
 XNOR2_X1 _20790_ (.A(_11108_),
    .B(_11109_),
    .ZN(_11110_));
 MUX2_X1 _20791_ (.A(_11106_),
    .B(_11110_),
    .S(_11091_),
    .Z(_00628_));
 BUF_X4 _20792_ (.A(_17161_),
    .Z(_11111_));
 XOR2_X1 _20793_ (.A(_17057_),
    .B(_11111_),
    .Z(_11112_));
 XNOR2_X1 _20794_ (.A(_09837_),
    .B(_01055_),
    .ZN(_11113_));
 XNOR2_X1 _20795_ (.A(_11066_),
    .B(_11113_),
    .ZN(_11114_));
 XOR2_X1 _20796_ (.A(_11059_),
    .B(_08888_),
    .Z(_11115_));
 XNOR2_X1 _20797_ (.A(_11114_),
    .B(_11115_),
    .ZN(_11116_));
 MUX2_X1 _20798_ (.A(_11112_),
    .B(_11116_),
    .S(_11091_),
    .Z(_00629_));
 XOR2_X1 _20799_ (.A(_17162_),
    .B(_17058_),
    .Z(_11117_));
 XOR2_X1 _20800_ (.A(_09616_),
    .B(_09763_),
    .Z(_11118_));
 XNOR2_X1 _20801_ (.A(_09288_),
    .B(_11118_),
    .ZN(_11119_));
 XNOR2_X1 _20802_ (.A(_11119_),
    .B(_09914_),
    .ZN(_11120_));
 XNOR2_X1 _20803_ (.A(_11120_),
    .B(_17162_),
    .ZN(_11121_));
 MUX2_X1 _20804_ (.A(_11117_),
    .B(_11121_),
    .S(_11091_),
    .Z(_00630_));
 XOR2_X1 _20805_ (.A(_17163_),
    .B(_17059_),
    .Z(_11122_));
 XNOR2_X1 _20806_ (.A(_10068_),
    .B(_10065_),
    .ZN(_11123_));
 XNOR2_X1 _20807_ (.A(_11123_),
    .B(_10401_),
    .ZN(_11124_));
 XNOR2_X1 _20808_ (.A(_11071_),
    .B(_10148_),
    .ZN(_11125_));
 XNOR2_X1 _20809_ (.A(_11124_),
    .B(_11125_),
    .ZN(_11126_));
 INV_X1 _20810_ (.A(_17163_),
    .ZN(_11127_));
 XNOR2_X1 _20811_ (.A(_11126_),
    .B(_11127_),
    .ZN(_11128_));
 MUX2_X1 _20812_ (.A(_11122_),
    .B(_11128_),
    .S(_11091_),
    .Z(_00631_));
 XOR2_X1 _20813_ (.A(_17164_),
    .B(_17060_),
    .Z(_11129_));
 XNOR2_X1 _20814_ (.A(_11081_),
    .B(_10153_),
    .ZN(_11130_));
 XNOR2_X1 _20815_ (.A(_10212_),
    .B(_10327_),
    .ZN(_11131_));
 XNOR2_X1 _20816_ (.A(_11131_),
    .B(_10616_),
    .ZN(_11132_));
 XNOR2_X1 _20817_ (.A(_11130_),
    .B(_11132_),
    .ZN(_11133_));
 XNOR2_X1 _20818_ (.A(_11133_),
    .B(_17164_),
    .ZN(_11134_));
 MUX2_X1 _20819_ (.A(_11129_),
    .B(_11134_),
    .S(_11091_),
    .Z(_00632_));
 XOR2_X1 _20820_ (.A(_17061_),
    .B(_17165_),
    .Z(_11135_));
 XNOR2_X1 _20821_ (.A(_10514_),
    .B(_01056_),
    .ZN(_11136_));
 XOR2_X1 _20822_ (.A(_11136_),
    .B(_10465_),
    .Z(_11137_));
 XNOR2_X1 _20823_ (.A(_10328_),
    .B(_10837_),
    .ZN(_11138_));
 XNOR2_X1 _20824_ (.A(_11137_),
    .B(_11138_),
    .ZN(_11139_));
 MUX2_X1 _20825_ (.A(_11135_),
    .B(_11139_),
    .S(_11091_),
    .Z(_00633_));
 XOR2_X1 _20826_ (.A(_17063_),
    .B(_17167_),
    .Z(_11140_));
 XOR2_X1 _20827_ (.A(_10717_),
    .B(_10777_),
    .Z(_11141_));
 XNOR2_X1 _20828_ (.A(_10989_),
    .B(_01057_),
    .ZN(_11142_));
 XNOR2_X1 _20829_ (.A(_11141_),
    .B(_11142_),
    .ZN(_11143_));
 XNOR2_X1 _20830_ (.A(_11143_),
    .B(_10565_),
    .ZN(_11144_));
 MUX2_X1 _20831_ (.A(_11140_),
    .B(_11144_),
    .S(_11091_),
    .Z(_00634_));
 XOR2_X1 _20832_ (.A(_17168_),
    .B(_17064_),
    .Z(_11145_));
 XNOR2_X1 _20833_ (.A(_10718_),
    .B(_10935_),
    .ZN(_11146_));
 XNOR2_X1 _20834_ (.A(_11146_),
    .B(_09093_),
    .ZN(_11147_));
 XNOR2_X1 _20835_ (.A(_11147_),
    .B(_17168_),
    .ZN(_11148_));
 BUF_X4 _20836_ (.A(_09099_),
    .Z(_11149_));
 MUX2_X1 _20837_ (.A(_11145_),
    .B(_11148_),
    .S(_11149_),
    .Z(_00635_));
 XOR2_X1 _20838_ (.A(_17240_),
    .B(_17065_),
    .Z(_11150_));
 INV_X32 _20839_ (.A(_16816_),
    .ZN(_11151_));
 AND2_X4 _20840_ (.A1(_11151_),
    .A2(_16817_),
    .ZN(_11152_));
 BUF_X16 _20841_ (.A(_11152_),
    .Z(_11153_));
 INV_X32 _20842_ (.A(_16818_),
    .ZN(_11154_));
 NOR2_X4 _20843_ (.A1(_11154_),
    .A2(_16819_),
    .ZN(_11155_));
 AND2_X4 _20844_ (.A1(_11153_),
    .A2(_11155_),
    .ZN(_11156_));
 BUF_X4 _20845_ (.A(_11156_),
    .Z(_11157_));
 NOR2_X4 _20846_ (.A1(_16814_),
    .A2(_16815_),
    .ZN(_11158_));
 BUF_X8 _20847_ (.A(_11158_),
    .Z(_11159_));
 AND2_X1 _20848_ (.A1(_11159_),
    .A2(_16812_),
    .ZN(_11160_));
 INV_X32 _20849_ (.A(_16814_),
    .ZN(_11161_));
 NOR2_X4 _20850_ (.A1(_11161_),
    .A2(_16815_),
    .ZN(_11162_));
 BUF_X4 _20851_ (.A(_11162_),
    .Z(_11163_));
 BUF_X4 _20852_ (.A(_11163_),
    .Z(_11164_));
 BUF_X4 _20853_ (.A(_11164_),
    .Z(_11165_));
 OAI21_X1 _20854_ (.A(_11157_),
    .B1(_11160_),
    .B2(_11165_),
    .ZN(_11166_));
 BUF_X2 _20855_ (.A(_11155_),
    .Z(_11167_));
 AND2_X4 _20856_ (.A1(_16817_),
    .A2(_16816_),
    .ZN(_11168_));
 BUF_X8 _20857_ (.A(_11168_),
    .Z(_11169_));
 AND2_X4 _20858_ (.A1(_11167_),
    .A2(_11169_),
    .ZN(_11170_));
 BUF_X8 _20859_ (.A(_11170_),
    .Z(_11171_));
 AND2_X4 _20860_ (.A1(_16813_),
    .A2(_16812_),
    .ZN(_11172_));
 AND2_X2 _20861_ (.A1(_11172_),
    .A2(_11158_),
    .ZN(_11173_));
 BUF_X8 _20862_ (.A(_11173_),
    .Z(_11174_));
 NAND2_X1 _20863_ (.A1(_11171_),
    .A2(_11174_),
    .ZN(_11175_));
 INV_X1 _20864_ (.A(_11171_),
    .ZN(_11176_));
 INV_X32 _20865_ (.A(_16813_),
    .ZN(_11177_));
 BUF_X16 _20866_ (.A(_11177_),
    .Z(_11178_));
 AND2_X4 _20867_ (.A1(_11159_),
    .A2(_11178_),
    .ZN(_11179_));
 INV_X1 _20868_ (.A(_11179_),
    .ZN(_11180_));
 OAI21_X1 _20869_ (.A(_11175_),
    .B1(_11176_),
    .B2(_11180_),
    .ZN(_11181_));
 INV_X32 _20870_ (.A(_16815_),
    .ZN(_11182_));
 NOR2_X4 _20871_ (.A1(_11182_),
    .A2(_16814_),
    .ZN(_11183_));
 AND2_X2 _20872_ (.A1(_11183_),
    .A2(_11172_),
    .ZN(_11184_));
 INV_X8 _20873_ (.A(_11184_),
    .ZN(_11185_));
 NOR2_X4 _20874_ (.A1(_11177_),
    .A2(_16812_),
    .ZN(_11186_));
 AND2_X4 _20875_ (.A1(_16814_),
    .A2(_16815_),
    .ZN(_11187_));
 BUF_X16 _20876_ (.A(_11187_),
    .Z(_11188_));
 AND2_X4 _20877_ (.A1(_11186_),
    .A2(_11188_),
    .ZN(_11189_));
 BUF_X16 _20878_ (.A(_11189_),
    .Z(_11190_));
 INV_X16 _20879_ (.A(_11190_),
    .ZN(_11191_));
 AOI21_X1 _20880_ (.A(_11176_),
    .B1(_11185_),
    .B2(_11191_),
    .ZN(_11192_));
 INV_X32 _20881_ (.A(_16812_),
    .ZN(_11193_));
 NOR2_X4 _20882_ (.A1(_11193_),
    .A2(_16813_),
    .ZN(_11194_));
 AND2_X4 _20883_ (.A1(_11194_),
    .A2(_11188_),
    .ZN(_11195_));
 BUF_X8 _20884_ (.A(_11195_),
    .Z(_11196_));
 AND2_X1 _20885_ (.A1(_11196_),
    .A2(_11171_),
    .ZN(_11197_));
 OR2_X1 _20886_ (.A1(_11192_),
    .A2(_11197_),
    .ZN(_11198_));
 BUF_X4 _20887_ (.A(_11171_),
    .Z(_11199_));
 NOR2_X1 _20888_ (.A1(_11193_),
    .A2(_16815_),
    .ZN(_11200_));
 AND2_X1 _20889_ (.A1(_11200_),
    .A2(_16814_),
    .ZN(_11201_));
 AOI211_X2 _20890_ (.A(_11181_),
    .B(_11198_),
    .C1(_11199_),
    .C2(_11201_),
    .ZN(_11202_));
 NOR2_X4 _20891_ (.A1(_11151_),
    .A2(_16817_),
    .ZN(_11203_));
 AND2_X2 _20892_ (.A1(_11155_),
    .A2(_11203_),
    .ZN(_11204_));
 INV_X4 _20893_ (.A(_11204_),
    .ZN(_11205_));
 AND2_X4 _20894_ (.A1(_11172_),
    .A2(_11187_),
    .ZN(_11206_));
 BUF_X8 _20895_ (.A(_11206_),
    .Z(_11207_));
 INV_X1 _20896_ (.A(_11207_),
    .ZN(_11208_));
 BUF_X4 _20897_ (.A(_16812_),
    .Z(_11209_));
 AND2_X1 _20898_ (.A1(_11183_),
    .A2(_11209_),
    .ZN(_11210_));
 INV_X1 _20899_ (.A(_11210_),
    .ZN(_11211_));
 AOI21_X1 _20900_ (.A(_11205_),
    .B1(_11208_),
    .B2(_11211_),
    .ZN(_11212_));
 BUF_X4 _20901_ (.A(_16813_),
    .Z(_11213_));
 AND2_X2 _20902_ (.A1(_11163_),
    .A2(_11213_),
    .ZN(_11214_));
 INV_X1 _20903_ (.A(_11214_),
    .ZN(_11215_));
 INV_X1 _20904_ (.A(_11158_),
    .ZN(_11216_));
 BUF_X4 _20905_ (.A(_11186_),
    .Z(_11217_));
 NOR2_X1 _20906_ (.A1(_11216_),
    .A2(_11217_),
    .ZN(_11218_));
 INV_X1 _20907_ (.A(_11218_),
    .ZN(_11219_));
 AOI21_X1 _20908_ (.A(_11205_),
    .B1(_11215_),
    .B2(_11219_),
    .ZN(_11220_));
 NOR2_X4 _20909_ (.A1(_16817_),
    .A2(_16816_),
    .ZN(_11221_));
 AND2_X2 _20910_ (.A1(_11167_),
    .A2(_11221_),
    .ZN(_11222_));
 BUF_X4 _20911_ (.A(_11222_),
    .Z(_11223_));
 INV_X1 _20912_ (.A(_11223_),
    .ZN(_11224_));
 NOR2_X4 _20913_ (.A1(_16813_),
    .A2(_16812_),
    .ZN(_11225_));
 AND2_X1 _20914_ (.A1(_11162_),
    .A2(_11225_),
    .ZN(_11226_));
 INV_X1 _20915_ (.A(_11226_),
    .ZN(_11227_));
 AOI21_X1 _20916_ (.A(_11224_),
    .B1(_11227_),
    .B2(_11180_),
    .ZN(_11228_));
 AND2_X1 _20917_ (.A1(_11187_),
    .A2(_11177_),
    .ZN(_11229_));
 BUF_X4 _20918_ (.A(_11229_),
    .Z(_11230_));
 OAI21_X1 _20919_ (.A(_11223_),
    .B1(_11190_),
    .B2(_11230_),
    .ZN(_11231_));
 BUF_X4 _20920_ (.A(_11183_),
    .Z(_11232_));
 BUF_X4 _20921_ (.A(_11209_),
    .Z(_11233_));
 BUF_X2 _20922_ (.A(_11221_),
    .Z(_11234_));
 NAND4_X1 _20923_ (.A1(_11232_),
    .A2(_11167_),
    .A3(_11233_),
    .A4(_11234_),
    .ZN(_11235_));
 NAND2_X1 _20924_ (.A1(_11231_),
    .A2(_11235_),
    .ZN(_11236_));
 NOR4_X1 _20925_ (.A1(_11212_),
    .A2(_11220_),
    .A3(_11228_),
    .A4(_11236_),
    .ZN(_11237_));
 NOR3_X2 _20926_ (.A1(_11186_),
    .A2(_16814_),
    .A3(_11182_),
    .ZN(_11238_));
 OAI21_X1 _20927_ (.A(_11157_),
    .B1(_11238_),
    .B2(_11190_),
    .ZN(_11239_));
 AND4_X1 _20928_ (.A1(_11166_),
    .A2(_11202_),
    .A3(_11237_),
    .A4(_11239_),
    .ZN(_11240_));
 NOR2_X4 _20929_ (.A1(_16819_),
    .A2(_16818_),
    .ZN(_11241_));
 AND2_X2 _20930_ (.A1(_11241_),
    .A2(_11221_),
    .ZN(_11242_));
 INV_X1 _20931_ (.A(_11242_),
    .ZN(_11243_));
 BUF_X4 _20932_ (.A(_11194_),
    .Z(_11244_));
 AND2_X2 _20933_ (.A1(_11244_),
    .A2(_11163_),
    .ZN(_11245_));
 INV_X1 _20934_ (.A(_11245_),
    .ZN(_11246_));
 AOI21_X1 _20935_ (.A(_11243_),
    .B1(_11246_),
    .B2(_11215_),
    .ZN(_11247_));
 AND2_X2 _20936_ (.A1(_11244_),
    .A2(_11183_),
    .ZN(_11248_));
 INV_X1 _20937_ (.A(_11248_),
    .ZN(_11249_));
 AND2_X1 _20938_ (.A1(_11183_),
    .A2(_16813_),
    .ZN(_11250_));
 INV_X1 _20939_ (.A(_11250_),
    .ZN(_11251_));
 AOI21_X1 _20940_ (.A(_11243_),
    .B1(_11249_),
    .B2(_11251_),
    .ZN(_11252_));
 BUF_X4 _20941_ (.A(_11242_),
    .Z(_11253_));
 AND2_X1 _20942_ (.A1(_11159_),
    .A2(_11213_),
    .ZN(_11254_));
 AND2_X1 _20943_ (.A1(_11253_),
    .A2(_11254_),
    .ZN(_11255_));
 INV_X1 _20944_ (.A(_11172_),
    .ZN(_11256_));
 BUF_X2 _20945_ (.A(_11256_),
    .Z(_11257_));
 BUF_X4 _20946_ (.A(_11188_),
    .Z(_11258_));
 INV_X1 _20947_ (.A(_11225_),
    .ZN(_11259_));
 BUF_X2 _20948_ (.A(_11259_),
    .Z(_11260_));
 AND4_X1 _20949_ (.A1(_11257_),
    .A2(_11253_),
    .A3(_11258_),
    .A4(_11260_),
    .ZN(_11261_));
 NOR4_X1 _20950_ (.A1(_11247_),
    .A2(_11252_),
    .A3(_11255_),
    .A4(_11261_),
    .ZN(_11262_));
 AND2_X2 _20951_ (.A1(_11203_),
    .A2(_11241_),
    .ZN(_11263_));
 BUF_X4 _20952_ (.A(_11263_),
    .Z(_11264_));
 BUF_X8 _20953_ (.A(_11264_),
    .Z(_11265_));
 AND4_X1 _20954_ (.A1(_11257_),
    .A2(_11265_),
    .A3(_11260_),
    .A4(_11164_),
    .ZN(_11266_));
 BUF_X2 _20955_ (.A(_11254_),
    .Z(_11267_));
 AOI21_X1 _20956_ (.A(_11266_),
    .B1(_11265_),
    .B2(_11267_),
    .ZN(_11268_));
 BUF_X4 _20957_ (.A(_11225_),
    .Z(_11269_));
 AND2_X2 _20958_ (.A1(_11232_),
    .A2(_11269_),
    .ZN(_11270_));
 NAND2_X1 _20959_ (.A1(_11265_),
    .A2(_11270_),
    .ZN(_11271_));
 NAND2_X1 _20960_ (.A1(_11265_),
    .A2(_11184_),
    .ZN(_11272_));
 AND3_X1 _20961_ (.A1(_11268_),
    .A2(_11271_),
    .A3(_11272_),
    .ZN(_11273_));
 AND2_X4 _20962_ (.A1(_11153_),
    .A2(_11241_),
    .ZN(_11274_));
 BUF_X8 _20963_ (.A(_11274_),
    .Z(_11275_));
 INV_X4 _20964_ (.A(_11275_),
    .ZN(_11276_));
 AND2_X4 _20965_ (.A1(_11188_),
    .A2(_11225_),
    .ZN(_11277_));
 INV_X2 _20966_ (.A(_11277_),
    .ZN(_11278_));
 AND2_X4 _20967_ (.A1(_11188_),
    .A2(_16813_),
    .ZN(_11279_));
 INV_X4 _20968_ (.A(_11279_),
    .ZN(_11280_));
 AOI21_X1 _20969_ (.A(_11276_),
    .B1(_11278_),
    .B2(_11280_),
    .ZN(_11281_));
 AND2_X1 _20970_ (.A1(_11256_),
    .A2(_11163_),
    .ZN(_11282_));
 AND3_X1 _20971_ (.A1(_11282_),
    .A2(_11260_),
    .A3(_11275_),
    .ZN(_11283_));
 NOR2_X1 _20972_ (.A1(_11216_),
    .A2(_11172_),
    .ZN(_11284_));
 AND2_X2 _20973_ (.A1(_11274_),
    .A2(_11284_),
    .ZN(_11285_));
 AND2_X2 _20974_ (.A1(_11259_),
    .A2(_11183_),
    .ZN(_11286_));
 AND2_X1 _20975_ (.A1(_11274_),
    .A2(_11286_),
    .ZN(_11287_));
 NOR4_X1 _20976_ (.A1(_11281_),
    .A2(_11283_),
    .A3(_11285_),
    .A4(_11287_),
    .ZN(_11288_));
 AND2_X4 _20977_ (.A1(_11169_),
    .A2(_11241_),
    .ZN(_11289_));
 INV_X1 _20978_ (.A(_11289_),
    .ZN(_11290_));
 INV_X1 _20979_ (.A(_11229_),
    .ZN(_11291_));
 AOI21_X1 _20980_ (.A(_11290_),
    .B1(_11208_),
    .B2(_11291_),
    .ZN(_11292_));
 BUF_X4 _20981_ (.A(_11289_),
    .Z(_11293_));
 AND3_X1 _20982_ (.A1(_11293_),
    .A2(_11269_),
    .A3(_11232_),
    .ZN(_11294_));
 NOR2_X1 _20983_ (.A1(_11216_),
    .A2(_11269_),
    .ZN(_11295_));
 AND2_X1 _20984_ (.A1(_11295_),
    .A2(_11289_),
    .ZN(_11296_));
 BUF_X2 _20985_ (.A(_11241_),
    .Z(_11297_));
 BUF_X4 _20986_ (.A(_11169_),
    .Z(_11298_));
 AND4_X1 _20987_ (.A1(_11297_),
    .A2(_11164_),
    .A3(_11217_),
    .A4(_11298_),
    .ZN(_11299_));
 NOR4_X1 _20988_ (.A1(_11292_),
    .A2(_11294_),
    .A3(_11296_),
    .A4(_11299_),
    .ZN(_11300_));
 AND4_X1 _20989_ (.A1(_11262_),
    .A2(_11273_),
    .A3(_11288_),
    .A4(_11300_),
    .ZN(_11301_));
 INV_X1 _20990_ (.A(_11163_),
    .ZN(_11302_));
 NOR2_X1 _20991_ (.A1(_11302_),
    .A2(_11186_),
    .ZN(_11303_));
 AND2_X4 _20992_ (.A1(_11154_),
    .A2(_16819_),
    .ZN(_11304_));
 BUF_X8 _20993_ (.A(_11304_),
    .Z(_11305_));
 AND2_X4 _20994_ (.A1(_11305_),
    .A2(_11169_),
    .ZN(_11306_));
 AND2_X1 _20995_ (.A1(_11303_),
    .A2(_11306_),
    .ZN(_11307_));
 INV_X1 _20996_ (.A(_11307_),
    .ZN(_11308_));
 BUF_X4 _20997_ (.A(_11306_),
    .Z(_11309_));
 AND2_X2 _20998_ (.A1(_11225_),
    .A2(_11158_),
    .ZN(_11310_));
 OAI21_X4 _20999_ (.A(_11309_),
    .B1(_11310_),
    .B2(_11267_),
    .ZN(_11311_));
 INV_X2 _21000_ (.A(_11306_),
    .ZN(_11312_));
 OAI211_X2 _21001_ (.A(_11308_),
    .B(_11311_),
    .C1(_11278_),
    .C2(_11312_),
    .ZN(_11313_));
 AND2_X2 _21002_ (.A1(_11305_),
    .A2(_11221_),
    .ZN(_11314_));
 BUF_X2 _21003_ (.A(_11314_),
    .Z(_11315_));
 BUF_X2 _21004_ (.A(_11279_),
    .Z(_11316_));
 OAI21_X1 _21005_ (.A(_11315_),
    .B1(_11196_),
    .B2(_11316_),
    .ZN(_11317_));
 NAND2_X1 _21006_ (.A1(_11303_),
    .A2(_11314_),
    .ZN(_11318_));
 BUF_X4 _21007_ (.A(_11305_),
    .Z(_11319_));
 BUF_X4 _21008_ (.A(_11319_),
    .Z(_11320_));
 BUF_X2 _21009_ (.A(_11193_),
    .Z(_11321_));
 BUF_X4 _21010_ (.A(_11159_),
    .Z(_11322_));
 NAND4_X1 _21011_ (.A1(_11320_),
    .A2(_11321_),
    .A3(_11234_),
    .A4(_11322_),
    .ZN(_11323_));
 NAND4_X1 _21012_ (.A1(_11320_),
    .A2(_11232_),
    .A3(_11233_),
    .A4(_11234_),
    .ZN(_11324_));
 NAND4_X1 _21013_ (.A1(_11317_),
    .A2(_11318_),
    .A3(_11323_),
    .A4(_11324_),
    .ZN(_11325_));
 BUF_X4 _21014_ (.A(_11203_),
    .Z(_11326_));
 AND2_X4 _21015_ (.A1(_11305_),
    .A2(_11326_),
    .ZN(_11327_));
 BUF_X8 _21016_ (.A(_11327_),
    .Z(_11328_));
 NAND3_X1 _21017_ (.A1(_11328_),
    .A2(_11284_),
    .A3(_11260_),
    .ZN(_11329_));
 INV_X1 _21018_ (.A(_11327_),
    .ZN(_11330_));
 OAI21_X1 _21019_ (.A(_11329_),
    .B1(_11280_),
    .B2(_11330_),
    .ZN(_11331_));
 BUF_X4 _21020_ (.A(_11153_),
    .Z(_11332_));
 OAI211_X2 _21021_ (.A(_11332_),
    .B(_11320_),
    .C1(_11207_),
    .C2(_11230_),
    .ZN(_11333_));
 NAND4_X1 _21022_ (.A1(_11332_),
    .A2(_11320_),
    .A3(_11244_),
    .A4(_11232_),
    .ZN(_11334_));
 AND2_X4 _21023_ (.A1(_11153_),
    .A2(_11305_),
    .ZN(_11335_));
 BUF_X4 _21024_ (.A(_11335_),
    .Z(_11336_));
 INV_X1 _21025_ (.A(_11336_),
    .ZN(_11337_));
 OAI211_X2 _21026_ (.A(_11333_),
    .B(_11334_),
    .C1(_11337_),
    .C2(_11227_),
    .ZN(_11338_));
 NOR4_X1 _21027_ (.A1(_11313_),
    .A2(_11325_),
    .A3(_11331_),
    .A4(_11338_),
    .ZN(_11339_));
 AND2_X4 _21028_ (.A1(_16819_),
    .A2(_16818_),
    .ZN(_11340_));
 BUF_X8 _21029_ (.A(_11340_),
    .Z(_11341_));
 AND2_X4 _21030_ (.A1(_11203_),
    .A2(_11341_),
    .ZN(_11342_));
 BUF_X8 _21031_ (.A(_11342_),
    .Z(_11343_));
 INV_X2 _21032_ (.A(_11196_),
    .ZN(_11344_));
 AND2_X2 _21033_ (.A1(_11186_),
    .A2(_11159_),
    .ZN(_11345_));
 INV_X1 _21034_ (.A(_11345_),
    .ZN(_11346_));
 NAND3_X1 _21035_ (.A1(_11246_),
    .A2(_11344_),
    .A3(_11346_),
    .ZN(_11347_));
 INV_X1 _21036_ (.A(_11186_),
    .ZN(_11348_));
 AOI21_X1 _21037_ (.A(_11182_),
    .B1(_11348_),
    .B2(_16814_),
    .ZN(_11349_));
 OAI21_X1 _21038_ (.A(_11343_),
    .B1(_11347_),
    .B2(_11349_),
    .ZN(_11350_));
 INV_X1 _21039_ (.A(_11183_),
    .ZN(_11351_));
 NOR2_X1 _21040_ (.A1(_11351_),
    .A2(_11244_),
    .ZN(_11352_));
 AND2_X4 _21041_ (.A1(_11153_),
    .A2(_11340_),
    .ZN(_11353_));
 AND2_X2 _21042_ (.A1(_11352_),
    .A2(_11353_),
    .ZN(_11354_));
 INV_X1 _21043_ (.A(_11353_),
    .ZN(_11355_));
 INV_X4 _21044_ (.A(_11174_),
    .ZN(_11356_));
 INV_X4 _21045_ (.A(_11310_),
    .ZN(_11357_));
 NAND2_X4 _21046_ (.A1(_11356_),
    .A2(_11357_),
    .ZN(_11358_));
 INV_X2 _21047_ (.A(_11358_),
    .ZN(_11359_));
 AND2_X2 _21048_ (.A1(_11162_),
    .A2(_11178_),
    .ZN(_11360_));
 INV_X1 _21049_ (.A(_11360_),
    .ZN(_11361_));
 AOI21_X1 _21050_ (.A(_11355_),
    .B1(_11359_),
    .B2(_11361_),
    .ZN(_11362_));
 BUF_X2 _21051_ (.A(_11353_),
    .Z(_11363_));
 AND2_X2 _21052_ (.A1(_11188_),
    .A2(_11209_),
    .ZN(_11364_));
 AOI211_X4 _21053_ (.A(_11354_),
    .B(_11362_),
    .C1(_11363_),
    .C2(_11364_),
    .ZN(_11365_));
 AND4_X1 _21054_ (.A1(_11234_),
    .A2(_11217_),
    .A3(_11322_),
    .A4(_11341_),
    .ZN(_11366_));
 AND2_X4 _21055_ (.A1(_11340_),
    .A2(_11221_),
    .ZN(_11367_));
 BUF_X8 _21056_ (.A(_11367_),
    .Z(_11368_));
 INV_X1 _21057_ (.A(_11368_),
    .ZN(_11369_));
 AOI21_X1 _21058_ (.A(_11369_),
    .B1(_11191_),
    .B2(_11291_),
    .ZN(_11370_));
 BUF_X4 _21059_ (.A(_11368_),
    .Z(_11371_));
 AOI211_X4 _21060_ (.A(_11366_),
    .B(_11370_),
    .C1(_11210_),
    .C2(_11371_),
    .ZN(_11372_));
 AND2_X2 _21061_ (.A1(_11168_),
    .A2(_11340_),
    .ZN(_11373_));
 NAND2_X1 _21062_ (.A1(_11226_),
    .A2(_11373_),
    .ZN(_11374_));
 BUF_X4 _21063_ (.A(_11373_),
    .Z(_11375_));
 NOR2_X1 _21064_ (.A1(_11182_),
    .A2(_16813_),
    .ZN(_11376_));
 AND2_X2 _21065_ (.A1(_11376_),
    .A2(_11161_),
    .ZN(_11377_));
 BUF_X4 _21066_ (.A(_11377_),
    .Z(_11378_));
 BUF_X2 _21067_ (.A(_11250_),
    .Z(_11379_));
 OAI21_X1 _21068_ (.A(_11375_),
    .B1(_11378_),
    .B2(_11379_),
    .ZN(_11380_));
 OAI211_X2 _21069_ (.A(_11375_),
    .B(_11322_),
    .C1(_11213_),
    .C2(_11233_),
    .ZN(_11381_));
 NAND3_X1 _21070_ (.A1(_11373_),
    .A2(_11258_),
    .A3(_11217_),
    .ZN(_11382_));
 AND4_X1 _21071_ (.A1(_11374_),
    .A2(_11380_),
    .A3(_11381_),
    .A4(_11382_),
    .ZN(_11383_));
 AND4_X1 _21072_ (.A1(_11350_),
    .A2(_11365_),
    .A3(_11372_),
    .A4(_11383_),
    .ZN(_11384_));
 NAND4_X1 _21073_ (.A1(_11240_),
    .A2(_11301_),
    .A3(_11339_),
    .A4(_11384_),
    .ZN(_11385_));
 AND2_X1 _21074_ (.A1(_11253_),
    .A2(_11310_),
    .ZN(_11386_));
 NOR2_X2 _21075_ (.A1(_11385_),
    .A2(_11386_),
    .ZN(_11387_));
 NOR2_X4 _21076_ (.A1(_16827_),
    .A2(_16826_),
    .ZN(_11388_));
 NOR2_X4 _21077_ (.A1(_16825_),
    .A2(_16824_),
    .ZN(_11389_));
 AND2_X1 _21078_ (.A1(_11388_),
    .A2(_11389_),
    .ZN(_11390_));
 BUF_X4 _21079_ (.A(_11390_),
    .Z(_11391_));
 BUF_X4 _21080_ (.A(_11391_),
    .Z(_11392_));
 NOR2_X4 _21081_ (.A1(_16822_),
    .A2(_16823_),
    .ZN(_11393_));
 BUF_X8 _21082_ (.A(_11393_),
    .Z(_11394_));
 AND2_X4 _21083_ (.A1(_11394_),
    .A2(_16821_),
    .ZN(_11395_));
 BUF_X4 _21084_ (.A(_11395_),
    .Z(_11396_));
 NAND2_X1 _21085_ (.A1(_11392_),
    .A2(_11396_),
    .ZN(_11397_));
 AND2_X4 _21086_ (.A1(_16822_),
    .A2(_16823_),
    .ZN(_11398_));
 BUF_X16 _21087_ (.A(_11398_),
    .Z(_11399_));
 INV_X8 _21088_ (.A(_11399_),
    .ZN(_11400_));
 NOR2_X4 _21089_ (.A1(_16821_),
    .A2(_16820_),
    .ZN(_11401_));
 BUF_X8 _21090_ (.A(_11401_),
    .Z(_11402_));
 NOR2_X4 _21091_ (.A1(_11400_),
    .A2(_11402_),
    .ZN(_11403_));
 AND2_X4 _21092_ (.A1(_16821_),
    .A2(_16820_),
    .ZN(_11404_));
 BUF_X8 _21093_ (.A(_11404_),
    .Z(_11405_));
 INV_X4 _21094_ (.A(_11405_),
    .ZN(_11406_));
 BUF_X8 _21095_ (.A(_11406_),
    .Z(_11407_));
 NAND3_X1 _21096_ (.A1(_11403_),
    .A2(_11407_),
    .A3(_11392_),
    .ZN(_11408_));
 INV_X32 _21097_ (.A(_16822_),
    .ZN(_11409_));
 NOR2_X2 _21098_ (.A1(_11409_),
    .A2(_16823_),
    .ZN(_11410_));
 BUF_X4 _21099_ (.A(_11410_),
    .Z(_11411_));
 BUF_X4 _21100_ (.A(_11411_),
    .Z(_11412_));
 BUF_X4 _21101_ (.A(_16821_),
    .Z(_11413_));
 BUF_X4 _21102_ (.A(_16820_),
    .Z(_11414_));
 BUF_X4 _21103_ (.A(_11414_),
    .Z(_11415_));
 OAI211_X2 _21104_ (.A(_11392_),
    .B(_11412_),
    .C1(_11413_),
    .C2(_11415_),
    .ZN(_11416_));
 INV_X32 _21105_ (.A(_16823_),
    .ZN(_11417_));
 NOR2_X4 _21106_ (.A1(_11417_),
    .A2(_16822_),
    .ZN(_11418_));
 BUF_X4 _21107_ (.A(_11418_),
    .Z(_11419_));
 BUF_X4 _21108_ (.A(_11419_),
    .Z(_11420_));
 OAI211_X2 _21109_ (.A(_11392_),
    .B(_11420_),
    .C1(_11413_),
    .C2(_11415_),
    .ZN(_11421_));
 AND4_X1 _21110_ (.A1(_11397_),
    .A2(_11408_),
    .A3(_11416_),
    .A4(_11421_),
    .ZN(_11422_));
 AND2_X4 _21111_ (.A1(_16825_),
    .A2(_16824_),
    .ZN(_11423_));
 AND2_X2 _21112_ (.A1(_11423_),
    .A2(_11388_),
    .ZN(_11424_));
 INV_X1 _21113_ (.A(_11424_),
    .ZN(_11425_));
 INV_X4 _21114_ (.A(_11402_),
    .ZN(_11426_));
 NAND2_X2 _21115_ (.A1(_11426_),
    .A2(_11394_),
    .ZN(_11427_));
 NOR2_X1 _21116_ (.A1(_11425_),
    .A2(_11427_),
    .ZN(_11428_));
 INV_X32 _21117_ (.A(_16821_),
    .ZN(_11429_));
 AND2_X4 _21118_ (.A1(_11399_),
    .A2(_11429_),
    .ZN(_11430_));
 AND2_X4 _21119_ (.A1(_11430_),
    .A2(_11424_),
    .ZN(_11431_));
 INV_X2 _21120_ (.A(_11431_),
    .ZN(_11432_));
 AND2_X4 _21121_ (.A1(_11405_),
    .A2(_11399_),
    .ZN(_11433_));
 BUF_X8 _21122_ (.A(_11433_),
    .Z(_11434_));
 NAND2_X2 _21123_ (.A1(_11434_),
    .A2(_11424_),
    .ZN(_11435_));
 AND2_X2 _21124_ (.A1(_11418_),
    .A2(_11402_),
    .ZN(_11436_));
 INV_X1 _21125_ (.A(_11436_),
    .ZN(_11437_));
 OAI211_X2 _21126_ (.A(_11432_),
    .B(_11435_),
    .C1(_11437_),
    .C2(_11425_),
    .ZN(_11438_));
 NOR2_X4 _21127_ (.A1(_11429_),
    .A2(_16820_),
    .ZN(_11439_));
 AND2_X1 _21128_ (.A1(_11410_),
    .A2(_11439_),
    .ZN(_11440_));
 BUF_X2 _21129_ (.A(_11440_),
    .Z(_11441_));
 BUF_X2 _21130_ (.A(_11424_),
    .Z(_11442_));
 AOI211_X2 _21131_ (.A(_11428_),
    .B(_11438_),
    .C1(_11441_),
    .C2(_11442_),
    .ZN(_11443_));
 INV_X32 _21132_ (.A(_16824_),
    .ZN(_11444_));
 NOR2_X4 _21133_ (.A1(_11444_),
    .A2(_16825_),
    .ZN(_11445_));
 AND2_X1 _21134_ (.A1(_11445_),
    .A2(_11388_),
    .ZN(_11446_));
 BUF_X4 _21135_ (.A(_11446_),
    .Z(_11447_));
 AND2_X1 _21136_ (.A1(_11447_),
    .A2(_11395_),
    .ZN(_11448_));
 AND2_X4 _21137_ (.A1(_11418_),
    .A2(_11404_),
    .ZN(_11449_));
 BUF_X4 _21138_ (.A(_11449_),
    .Z(_11450_));
 INV_X2 _21139_ (.A(_11450_),
    .ZN(_11451_));
 NAND2_X1 _21140_ (.A1(_11451_),
    .A2(_11437_),
    .ZN(_11452_));
 AND2_X1 _21141_ (.A1(_11452_),
    .A2(_11447_),
    .ZN(_11453_));
 BUF_X2 _21142_ (.A(_11447_),
    .Z(_11454_));
 INV_X2 _21143_ (.A(_11440_),
    .ZN(_11455_));
 INV_X32 _21144_ (.A(_16820_),
    .ZN(_11456_));
 NOR2_X4 _21145_ (.A1(_11456_),
    .A2(_16821_),
    .ZN(_11457_));
 AND2_X1 _21146_ (.A1(_11410_),
    .A2(_11457_),
    .ZN(_11458_));
 BUF_X4 _21147_ (.A(_11458_),
    .Z(_11459_));
 INV_X1 _21148_ (.A(_11459_),
    .ZN(_11460_));
 NAND2_X1 _21149_ (.A1(_11455_),
    .A2(_11460_),
    .ZN(_11461_));
 AOI211_X2 _21150_ (.A(_11448_),
    .B(_11453_),
    .C1(_11454_),
    .C2(_11461_),
    .ZN(_11462_));
 AND2_X4 _21151_ (.A1(_11444_),
    .A2(_16825_),
    .ZN(_11463_));
 BUF_X8 _21152_ (.A(_11463_),
    .Z(_11464_));
 AND2_X4 _21153_ (.A1(_11464_),
    .A2(_11388_),
    .ZN(_11465_));
 INV_X1 _21154_ (.A(_11465_),
    .ZN(_11466_));
 BUF_X16 _21155_ (.A(_11429_),
    .Z(_11467_));
 AOI211_X4 _21156_ (.A(_11400_),
    .B(_11466_),
    .C1(_11467_),
    .C2(_11414_),
    .ZN(_11468_));
 INV_X1 _21157_ (.A(_11394_),
    .ZN(_11469_));
 NOR2_X1 _21158_ (.A1(_11469_),
    .A2(_11405_),
    .ZN(_11470_));
 AND2_X1 _21159_ (.A1(_11465_),
    .A2(_11470_),
    .ZN(_11471_));
 AND2_X4 _21160_ (.A1(_11426_),
    .A2(_11418_),
    .ZN(_11472_));
 AND2_X1 _21161_ (.A1(_11465_),
    .A2(_11472_),
    .ZN(_11473_));
 AND2_X1 _21162_ (.A1(_11406_),
    .A2(_11411_),
    .ZN(_11474_));
 AND3_X1 _21163_ (.A1(_11474_),
    .A2(_11465_),
    .A3(_11426_),
    .ZN(_11475_));
 NOR4_X1 _21164_ (.A1(_11468_),
    .A2(_11471_),
    .A3(_11473_),
    .A4(_11475_),
    .ZN(_11476_));
 AND4_X2 _21165_ (.A1(_11422_),
    .A2(_11443_),
    .A3(_11462_),
    .A4(_11476_),
    .ZN(_11477_));
 AND2_X4 _21166_ (.A1(_16827_),
    .A2(_16826_),
    .ZN(_11478_));
 AND2_X2 _21167_ (.A1(_11463_),
    .A2(_11478_),
    .ZN(_11479_));
 BUF_X2 _21168_ (.A(_11479_),
    .Z(_11480_));
 AND2_X2 _21169_ (.A1(_11410_),
    .A2(_11467_),
    .ZN(_11481_));
 BUF_X4 _21170_ (.A(_11481_),
    .Z(_11482_));
 AND2_X1 _21171_ (.A1(_11480_),
    .A2(_11482_),
    .ZN(_11483_));
 INV_X1 _21172_ (.A(_11483_),
    .ZN(_11484_));
 INV_X1 _21173_ (.A(_11479_),
    .ZN(_11485_));
 AND2_X4 _21174_ (.A1(_11405_),
    .A2(_11394_),
    .ZN(_11486_));
 INV_X4 _21175_ (.A(_11486_),
    .ZN(_11487_));
 AND2_X2 _21176_ (.A1(_11393_),
    .A2(_11402_),
    .ZN(_11488_));
 INV_X2 _21177_ (.A(_11488_),
    .ZN(_11489_));
 NAND2_X1 _21178_ (.A1(_11487_),
    .A2(_11489_),
    .ZN(_11490_));
 INV_X1 _21179_ (.A(_11490_),
    .ZN(_11491_));
 OAI21_X1 _21180_ (.A(_11484_),
    .B1(_11485_),
    .B2(_11491_),
    .ZN(_11492_));
 INV_X1 _21181_ (.A(_11418_),
    .ZN(_11493_));
 NOR2_X1 _21182_ (.A1(_11493_),
    .A2(_11457_),
    .ZN(_11494_));
 AND2_X1 _21183_ (.A1(_11494_),
    .A2(_11479_),
    .ZN(_11495_));
 AND2_X2 _21184_ (.A1(_11399_),
    .A2(_11414_),
    .ZN(_11496_));
 AND2_X1 _21185_ (.A1(_11480_),
    .A2(_11496_),
    .ZN(_11497_));
 OR3_X1 _21186_ (.A1(_11492_),
    .A2(_11495_),
    .A3(_11497_),
    .ZN(_11498_));
 AND2_X1 _21187_ (.A1(_11457_),
    .A2(_11393_),
    .ZN(_11499_));
 BUF_X4 _21188_ (.A(_11499_),
    .Z(_11500_));
 AND2_X4 _21189_ (.A1(_11423_),
    .A2(_11478_),
    .ZN(_11501_));
 BUF_X4 _21190_ (.A(_11501_),
    .Z(_11502_));
 AND2_X1 _21191_ (.A1(_11500_),
    .A2(_11502_),
    .ZN(_11503_));
 INV_X1 _21192_ (.A(_11503_),
    .ZN(_11504_));
 BUF_X4 _21193_ (.A(_11502_),
    .Z(_11505_));
 NAND2_X1 _21194_ (.A1(_11505_),
    .A2(_11396_),
    .ZN(_11506_));
 AND2_X2 _21195_ (.A1(_11410_),
    .A2(_11402_),
    .ZN(_11507_));
 NAND2_X1 _21196_ (.A1(_11507_),
    .A2(_11505_),
    .ZN(_11508_));
 AND3_X2 _21197_ (.A1(_11504_),
    .A2(_11506_),
    .A3(_11508_),
    .ZN(_11509_));
 AND2_X4 _21198_ (.A1(_11439_),
    .A2(_11398_),
    .ZN(_11510_));
 BUF_X4 _21199_ (.A(_11510_),
    .Z(_11511_));
 NAND2_X1 _21200_ (.A1(_11511_),
    .A2(_11502_),
    .ZN(_11512_));
 INV_X1 _21201_ (.A(_11502_),
    .ZN(_11513_));
 OAI211_X2 _21202_ (.A(_11509_),
    .B(_11512_),
    .C1(_11493_),
    .C2(_11513_),
    .ZN(_11514_));
 AND2_X2 _21203_ (.A1(_11445_),
    .A2(_11478_),
    .ZN(_11515_));
 BUF_X4 _21204_ (.A(_11515_),
    .Z(_11516_));
 INV_X1 _21205_ (.A(_11516_),
    .ZN(_11517_));
 AOI21_X1 _21206_ (.A(_11420_),
    .B1(_11403_),
    .B2(_11407_),
    .ZN(_11518_));
 AND2_X2 _21207_ (.A1(_11439_),
    .A2(_11393_),
    .ZN(_11519_));
 NOR2_X1 _21208_ (.A1(_11459_),
    .A2(_11519_),
    .ZN(_11520_));
 AOI21_X1 _21209_ (.A(_11517_),
    .B1(_11518_),
    .B2(_11520_),
    .ZN(_11521_));
 AND2_X4 _21210_ (.A1(_11478_),
    .A2(_11389_),
    .ZN(_11522_));
 INV_X1 _21211_ (.A(_11522_),
    .ZN(_11523_));
 INV_X1 _21212_ (.A(_11510_),
    .ZN(_11524_));
 INV_X4 _21213_ (.A(_11430_),
    .ZN(_11525_));
 AOI21_X1 _21214_ (.A(_11523_),
    .B1(_11524_),
    .B2(_11525_),
    .ZN(_11526_));
 BUF_X8 _21215_ (.A(_11522_),
    .Z(_11527_));
 BUF_X4 _21216_ (.A(_11527_),
    .Z(_11528_));
 BUF_X4 _21217_ (.A(_11456_),
    .Z(_11529_));
 AND3_X1 _21218_ (.A1(_11528_),
    .A2(_11529_),
    .A3(_11396_),
    .ZN(_11530_));
 AND2_X1 _21219_ (.A1(_11419_),
    .A2(_11414_),
    .ZN(_11531_));
 AND2_X2 _21220_ (.A1(_11531_),
    .A2(_11528_),
    .ZN(_11532_));
 OR3_X4 _21221_ (.A1(_11526_),
    .A2(_11530_),
    .A3(_11532_),
    .ZN(_11533_));
 NOR4_X2 _21222_ (.A1(_11498_),
    .A2(_11514_),
    .A3(_11521_),
    .A4(_11533_),
    .ZN(_11534_));
 INV_X32 _21223_ (.A(_16826_),
    .ZN(_11535_));
 NOR2_X4 _21224_ (.A1(_11535_),
    .A2(_16827_),
    .ZN(_11536_));
 BUF_X4 _21225_ (.A(_11536_),
    .Z(_11537_));
 AND4_X1 _21226_ (.A1(_11405_),
    .A2(_11464_),
    .A3(_11537_),
    .A4(_11419_),
    .ZN(_11538_));
 AND2_X1 _21227_ (.A1(_11463_),
    .A2(_11536_),
    .ZN(_11539_));
 AND2_X2 _21228_ (.A1(_11539_),
    .A2(_11511_),
    .ZN(_11540_));
 NAND2_X4 _21229_ (.A1(_11418_),
    .A2(_11467_),
    .ZN(_11541_));
 INV_X4 _21230_ (.A(_11541_),
    .ZN(_11542_));
 BUF_X8 _21231_ (.A(_11542_),
    .Z(_11543_));
 BUF_X4 _21232_ (.A(_11539_),
    .Z(_11544_));
 AOI211_X2 _21233_ (.A(_11538_),
    .B(_11540_),
    .C1(_11543_),
    .C2(_11544_),
    .ZN(_11545_));
 BUF_X4 _21234_ (.A(_11544_),
    .Z(_11546_));
 NAND2_X1 _21235_ (.A1(_11546_),
    .A2(_11482_),
    .ZN(_11547_));
 AND2_X4 _21236_ (.A1(_11410_),
    .A2(_11405_),
    .ZN(_11548_));
 OAI21_X1 _21237_ (.A(_11546_),
    .B1(_11441_),
    .B2(_11548_),
    .ZN(_11549_));
 OAI21_X1 _21238_ (.A(_11546_),
    .B1(_11500_),
    .B2(_11486_),
    .ZN(_11550_));
 NAND4_X1 _21239_ (.A1(_11545_),
    .A2(_11547_),
    .A3(_11549_),
    .A4(_11550_),
    .ZN(_11551_));
 BUF_X2 _21240_ (.A(_11389_),
    .Z(_11552_));
 AND2_X1 _21241_ (.A1(_11536_),
    .A2(_11552_),
    .ZN(_11553_));
 BUF_X4 _21242_ (.A(_11553_),
    .Z(_11554_));
 BUF_X4 _21243_ (.A(_11554_),
    .Z(_11555_));
 BUF_X8 _21244_ (.A(_11430_),
    .Z(_11556_));
 OAI21_X1 _21245_ (.A(_11555_),
    .B1(_11511_),
    .B2(_11556_),
    .ZN(_11557_));
 NAND4_X1 _21246_ (.A1(_11537_),
    .A2(_11420_),
    .A3(_11415_),
    .A4(_11552_),
    .ZN(_11558_));
 NAND2_X1 _21247_ (.A1(_11507_),
    .A2(_11555_),
    .ZN(_11559_));
 AND2_X1 _21248_ (.A1(_11393_),
    .A2(_11429_),
    .ZN(_11560_));
 BUF_X4 _21249_ (.A(_11560_),
    .Z(_11561_));
 NAND3_X1 _21250_ (.A1(_11561_),
    .A2(_11552_),
    .A3(_11537_),
    .ZN(_11562_));
 NAND4_X1 _21251_ (.A1(_11557_),
    .A2(_11558_),
    .A3(_11559_),
    .A4(_11562_),
    .ZN(_11563_));
 AND2_X2 _21252_ (.A1(_11537_),
    .A2(_11445_),
    .ZN(_11564_));
 AND2_X4 _21253_ (.A1(_11564_),
    .A2(_11486_),
    .ZN(_11565_));
 INV_X1 _21254_ (.A(_11565_),
    .ZN(_11566_));
 BUF_X4 _21255_ (.A(_11564_),
    .Z(_11567_));
 OAI21_X1 _21256_ (.A(_11567_),
    .B1(_11531_),
    .B2(_11434_),
    .ZN(_11568_));
 NAND2_X1 _21257_ (.A1(_11567_),
    .A2(_11561_),
    .ZN(_11569_));
 AND2_X2 _21258_ (.A1(_11411_),
    .A2(_16821_),
    .ZN(_11570_));
 NAND2_X1 _21259_ (.A1(_11567_),
    .A2(_11570_),
    .ZN(_11571_));
 NAND4_X1 _21260_ (.A1(_11566_),
    .A2(_11568_),
    .A3(_11569_),
    .A4(_11571_),
    .ZN(_11572_));
 AND2_X1 _21261_ (.A1(_11536_),
    .A2(_11423_),
    .ZN(_11573_));
 BUF_X4 _21262_ (.A(_11573_),
    .Z(_11574_));
 AND2_X4 _21263_ (.A1(_11403_),
    .A2(_11407_),
    .ZN(_11575_));
 OAI21_X1 _21264_ (.A(_11574_),
    .B1(_11575_),
    .B2(_11450_),
    .ZN(_11576_));
 AND2_X1 _21265_ (.A1(_11410_),
    .A2(_11414_),
    .ZN(_11577_));
 AND2_X1 _21266_ (.A1(_11574_),
    .A2(_11577_),
    .ZN(_11578_));
 INV_X1 _21267_ (.A(_11578_),
    .ZN(_11579_));
 NAND2_X1 _21268_ (.A1(_11573_),
    .A2(_11486_),
    .ZN(_11580_));
 OAI21_X1 _21269_ (.A(_11574_),
    .B1(_11500_),
    .B2(_11488_),
    .ZN(_11581_));
 NAND4_X1 _21270_ (.A1(_11576_),
    .A2(_11579_),
    .A3(_11580_),
    .A4(_11581_),
    .ZN(_11582_));
 NOR4_X1 _21271_ (.A1(_11551_),
    .A2(_11563_),
    .A3(_11572_),
    .A4(_11582_),
    .ZN(_11583_));
 INV_X1 _21272_ (.A(_11410_),
    .ZN(_11584_));
 NOR2_X1 _21273_ (.A1(_11584_),
    .A2(_11439_),
    .ZN(_11585_));
 AND2_X4 _21274_ (.A1(_11535_),
    .A2(_16827_),
    .ZN(_11586_));
 AND2_X2 _21275_ (.A1(_11586_),
    .A2(_11423_),
    .ZN(_11587_));
 AND2_X1 _21276_ (.A1(_11585_),
    .A2(_11587_),
    .ZN(_11588_));
 AND2_X2 _21277_ (.A1(_11398_),
    .A2(_11401_),
    .ZN(_11589_));
 BUF_X4 _21278_ (.A(_11589_),
    .Z(_11590_));
 BUF_X2 _21279_ (.A(_11423_),
    .Z(_11591_));
 BUF_X4 _21280_ (.A(_11586_),
    .Z(_11592_));
 AND3_X1 _21281_ (.A1(_11590_),
    .A2(_11591_),
    .A3(_11592_),
    .ZN(_11593_));
 AND4_X1 _21282_ (.A1(_11394_),
    .A2(_11586_),
    .A3(_11402_),
    .A4(_11591_),
    .ZN(_11594_));
 AND4_X1 _21283_ (.A1(_16821_),
    .A2(_11586_),
    .A3(_11394_),
    .A4(_11591_),
    .ZN(_11595_));
 OR4_X1 _21284_ (.A1(_11588_),
    .A2(_11593_),
    .A3(_11594_),
    .A4(_11595_),
    .ZN(_11596_));
 AND2_X1 _21285_ (.A1(_11586_),
    .A2(_11445_),
    .ZN(_11597_));
 INV_X1 _21286_ (.A(_11597_),
    .ZN(_11598_));
 BUF_X4 _21287_ (.A(_11394_),
    .Z(_11599_));
 BUF_X8 _21288_ (.A(_11439_),
    .Z(_11600_));
 BUF_X4 _21289_ (.A(_11457_),
    .Z(_11601_));
 OAI21_X1 _21290_ (.A(_11599_),
    .B1(_11600_),
    .B2(_11601_),
    .ZN(_11602_));
 AND2_X4 _21291_ (.A1(_11399_),
    .A2(_16821_),
    .ZN(_11603_));
 INV_X2 _21292_ (.A(_11603_),
    .ZN(_11604_));
 AOI21_X1 _21293_ (.A(_11598_),
    .B1(_11602_),
    .B2(_11604_),
    .ZN(_11605_));
 AND2_X2 _21294_ (.A1(_11586_),
    .A2(_11552_),
    .ZN(_11606_));
 BUF_X2 _21295_ (.A(_11606_),
    .Z(_11607_));
 OAI21_X1 _21296_ (.A(_11607_),
    .B1(_11403_),
    .B2(_11531_),
    .ZN(_11608_));
 NAND2_X1 _21297_ (.A1(_11585_),
    .A2(_11606_),
    .ZN(_11609_));
 INV_X1 _21298_ (.A(_11607_),
    .ZN(_11610_));
 NAND2_X1 _21299_ (.A1(_11599_),
    .A2(_11529_),
    .ZN(_11611_));
 OAI211_X2 _21300_ (.A(_11608_),
    .B(_11609_),
    .C1(_11610_),
    .C2(_11611_),
    .ZN(_11612_));
 OAI211_X2 _21301_ (.A(_11464_),
    .B(_11592_),
    .C1(_11434_),
    .C2(_11556_),
    .ZN(_11613_));
 NAND4_X1 _21302_ (.A1(_11464_),
    .A2(_11592_),
    .A3(_11601_),
    .A4(_11420_),
    .ZN(_11614_));
 INV_X1 _21303_ (.A(_11507_),
    .ZN(_11615_));
 AND2_X2 _21304_ (.A1(_11463_),
    .A2(_11586_),
    .ZN(_11616_));
 INV_X1 _21305_ (.A(_11616_),
    .ZN(_11617_));
 OAI211_X2 _21306_ (.A(_11613_),
    .B(_11614_),
    .C1(_11615_),
    .C2(_11617_),
    .ZN(_11618_));
 NOR4_X4 _21307_ (.A1(_11596_),
    .A2(_11605_),
    .A3(_11612_),
    .A4(_11618_),
    .ZN(_11619_));
 NAND4_X1 _21308_ (.A1(_11477_),
    .A2(_11534_),
    .A3(_11583_),
    .A4(_11619_),
    .ZN(_11620_));
 OAI21_X1 _21309_ (.A(_11417_),
    .B1(_11426_),
    .B2(_16822_),
    .ZN(_11621_));
 AND3_X1 _21310_ (.A1(_11388_),
    .A2(_11552_),
    .A3(_11417_),
    .ZN(_11622_));
 AND2_X1 _21311_ (.A1(_11621_),
    .A2(_11622_),
    .ZN(_11623_));
 NOR2_X2 _21312_ (.A1(_11620_),
    .A2(_11623_),
    .ZN(_11624_));
 XNOR2_X1 _21313_ (.A(_11387_),
    .B(_11624_),
    .ZN(_11625_));
 AND2_X4 _21314_ (.A1(_16772_),
    .A2(_16773_),
    .ZN(_11626_));
 INV_X32 _21315_ (.A(_16775_),
    .ZN(_11627_));
 INV_X32 _21316_ (.A(_16774_),
    .ZN(_11628_));
 NOR3_X1 _21317_ (.A1(_11626_),
    .A2(_11627_),
    .A3(_11628_),
    .ZN(_11629_));
 INV_X32 _21318_ (.A(_16776_),
    .ZN(_11630_));
 NOR2_X4 _21319_ (.A1(_11630_),
    .A2(_16777_),
    .ZN(_11631_));
 BUF_X4 _21320_ (.A(_11631_),
    .Z(_11632_));
 AND2_X4 _21321_ (.A1(_16779_),
    .A2(_16778_),
    .ZN(_11633_));
 BUF_X8 _21322_ (.A(_11633_),
    .Z(_11634_));
 BUF_X4 _21323_ (.A(_11634_),
    .Z(_11635_));
 NOR2_X4 _21324_ (.A1(_16772_),
    .A2(_16773_),
    .ZN(_11636_));
 BUF_X8 _21325_ (.A(_11636_),
    .Z(_11637_));
 INV_X8 _21326_ (.A(_11637_),
    .ZN(_11638_));
 NAND4_X1 _21327_ (.A1(_11629_),
    .A2(_11632_),
    .A3(_11635_),
    .A4(_11638_),
    .ZN(_11639_));
 AND2_X4 _21328_ (.A1(_11631_),
    .A2(_11633_),
    .ZN(_11640_));
 BUF_X8 _21329_ (.A(_11640_),
    .Z(_11641_));
 NOR2_X4 _21330_ (.A1(_11627_),
    .A2(_16774_),
    .ZN(_11642_));
 INV_X32 _21331_ (.A(_16773_),
    .ZN(_11643_));
 AND2_X2 _21332_ (.A1(_11642_),
    .A2(_11643_),
    .ZN(_11644_));
 BUF_X4 _21333_ (.A(_11644_),
    .Z(_11645_));
 NAND2_X1 _21334_ (.A1(_11641_),
    .A2(_11645_),
    .ZN(_11646_));
 INV_X1 _21335_ (.A(_11641_),
    .ZN(_11647_));
 AND2_X2 _21336_ (.A1(_11642_),
    .A2(_16773_),
    .ZN(_11648_));
 INV_X1 _21337_ (.A(_11648_),
    .ZN(_11649_));
 OAI211_X2 _21338_ (.A(_11639_),
    .B(_11646_),
    .C1(_11647_),
    .C2(_11649_),
    .ZN(_11650_));
 INV_X32 _21339_ (.A(_16772_),
    .ZN(_11651_));
 NOR2_X4 _21340_ (.A1(_11651_),
    .A2(_16773_),
    .ZN(_11652_));
 NOR2_X4 _21341_ (.A1(_11628_),
    .A2(_16775_),
    .ZN(_11653_));
 AND2_X4 _21342_ (.A1(_11652_),
    .A2(_11653_),
    .ZN(_11654_));
 BUF_X8 _21343_ (.A(_11654_),
    .Z(_11655_));
 NAND2_X1 _21344_ (.A1(_11655_),
    .A2(_11641_),
    .ZN(_11656_));
 NOR2_X4 _21345_ (.A1(_11643_),
    .A2(_16772_),
    .ZN(_11657_));
 NOR2_X4 _21346_ (.A1(_16775_),
    .A2(_16774_),
    .ZN(_11658_));
 AND2_X2 _21347_ (.A1(_11657_),
    .A2(_11658_),
    .ZN(_11659_));
 NAND2_X2 _21348_ (.A1(_11659_),
    .A2(_11641_),
    .ZN(_11660_));
 NAND2_X1 _21349_ (.A1(_11656_),
    .A2(_11660_),
    .ZN(_11661_));
 NOR2_X4 _21350_ (.A1(_16777_),
    .A2(_16776_),
    .ZN(_11662_));
 BUF_X8 _21351_ (.A(_11662_),
    .Z(_11663_));
 AND2_X4 _21352_ (.A1(_11634_),
    .A2(_11663_),
    .ZN(_11664_));
 BUF_X32 _21353_ (.A(_16772_),
    .Z(_11665_));
 BUF_X4 _21354_ (.A(_11642_),
    .Z(_11666_));
 NAND3_X1 _21355_ (.A1(_11664_),
    .A2(_11665_),
    .A3(_11666_),
    .ZN(_11667_));
 AND2_X4 _21356_ (.A1(_16775_),
    .A2(_16774_),
    .ZN(_11668_));
 BUF_X16 _21357_ (.A(_11668_),
    .Z(_11669_));
 AND2_X4 _21358_ (.A1(_11669_),
    .A2(_11643_),
    .ZN(_11670_));
 NAND2_X2 _21359_ (.A1(_11664_),
    .A2(_11670_),
    .ZN(_11671_));
 BUF_X4 _21360_ (.A(_11657_),
    .Z(_11672_));
 BUF_X16 _21361_ (.A(_11669_),
    .Z(_11673_));
 NAND4_X1 _21362_ (.A1(_11672_),
    .A2(_11634_),
    .A3(_11673_),
    .A4(_11663_),
    .ZN(_11674_));
 NAND3_X1 _21363_ (.A1(_11667_),
    .A2(_11671_),
    .A3(_11674_),
    .ZN(_11675_));
 BUF_X8 _21364_ (.A(_11658_),
    .Z(_11676_));
 AND4_X1 _21365_ (.A1(_11634_),
    .A2(_11672_),
    .A3(_11676_),
    .A4(_11663_),
    .ZN(_11677_));
 NOR4_X1 _21366_ (.A1(_11650_),
    .A2(_11661_),
    .A3(_11675_),
    .A4(_11677_),
    .ZN(_11678_));
 INV_X1 _21367_ (.A(_11642_),
    .ZN(_11679_));
 NOR2_X1 _21368_ (.A1(_11679_),
    .A2(_11652_),
    .ZN(_11680_));
 AND2_X4 _21369_ (.A1(_11630_),
    .A2(_16777_),
    .ZN(_11681_));
 AND2_X4 _21370_ (.A1(_11681_),
    .A2(_11634_),
    .ZN(_11682_));
 AND2_X1 _21371_ (.A1(_11680_),
    .A2(_11682_),
    .ZN(_11683_));
 INV_X4 _21372_ (.A(_11682_),
    .ZN(_11684_));
 AND2_X4 _21373_ (.A1(_11626_),
    .A2(_11658_),
    .ZN(_11685_));
 INV_X4 _21374_ (.A(_11685_),
    .ZN(_11686_));
 AND2_X4 _21375_ (.A1(_11658_),
    .A2(_11636_),
    .ZN(_11687_));
 INV_X4 _21376_ (.A(_11687_),
    .ZN(_11688_));
 NAND2_X4 _21377_ (.A1(_11686_),
    .A2(_11688_),
    .ZN(_11689_));
 INV_X2 _21378_ (.A(_11689_),
    .ZN(_11690_));
 AND2_X4 _21379_ (.A1(_11653_),
    .A2(_11643_),
    .ZN(_11691_));
 INV_X1 _21380_ (.A(_11691_),
    .ZN(_11692_));
 AOI21_X2 _21381_ (.A(_11684_),
    .B1(_11690_),
    .B2(_11692_),
    .ZN(_11693_));
 BUF_X4 _21382_ (.A(_11682_),
    .Z(_11694_));
 AND2_X4 _21383_ (.A1(_11669_),
    .A2(_11665_),
    .ZN(_11695_));
 AOI211_X2 _21384_ (.A(_11683_),
    .B(_11693_),
    .C1(_11694_),
    .C2(_11695_),
    .ZN(_11696_));
 AND2_X4 _21385_ (.A1(_16777_),
    .A2(_16776_),
    .ZN(_11697_));
 AND2_X4 _21386_ (.A1(_11634_),
    .A2(_11697_),
    .ZN(_11698_));
 BUF_X4 _21387_ (.A(_11652_),
    .Z(_11699_));
 AND3_X1 _21388_ (.A1(_11698_),
    .A2(_11699_),
    .A3(_11676_),
    .ZN(_11700_));
 BUF_X8 _21389_ (.A(_11653_),
    .Z(_11701_));
 AND2_X4 _21390_ (.A1(_11701_),
    .A2(_11636_),
    .ZN(_11702_));
 AND2_X4 _21391_ (.A1(_11702_),
    .A2(_11698_),
    .ZN(_11703_));
 AND2_X4 _21392_ (.A1(_11658_),
    .A2(_16773_),
    .ZN(_11704_));
 BUF_X4 _21393_ (.A(_11698_),
    .Z(_11705_));
 AOI211_X2 _21394_ (.A(_11700_),
    .B(_11703_),
    .C1(_11704_),
    .C2(_11705_),
    .ZN(_11706_));
 AND3_X1 _21395_ (.A1(_11698_),
    .A2(_11672_),
    .A3(_11669_),
    .ZN(_11707_));
 AND2_X1 _21396_ (.A1(_11648_),
    .A2(_11698_),
    .ZN(_11708_));
 AOI211_X2 _21397_ (.A(_11707_),
    .B(_11708_),
    .C1(_11645_),
    .C2(_11698_),
    .ZN(_11709_));
 AND4_X2 _21398_ (.A1(_11678_),
    .A2(_11696_),
    .A3(_11706_),
    .A4(_11709_),
    .ZN(_11710_));
 NOR2_X4 _21399_ (.A1(_16779_),
    .A2(_16778_),
    .ZN(_11711_));
 BUF_X4 _21400_ (.A(_11711_),
    .Z(_11712_));
 AND2_X2 _21401_ (.A1(_11632_),
    .A2(_11712_),
    .ZN(_11713_));
 INV_X1 _21402_ (.A(_11713_),
    .ZN(_11714_));
 INV_X1 _21403_ (.A(_11654_),
    .ZN(_11715_));
 AND2_X2 _21404_ (.A1(_11657_),
    .A2(_11653_),
    .ZN(_11716_));
 INV_X1 _21405_ (.A(_11716_),
    .ZN(_11717_));
 NAND2_X1 _21406_ (.A1(_11715_),
    .A2(_11717_),
    .ZN(_11718_));
 INV_X1 _21407_ (.A(_11718_),
    .ZN(_11719_));
 INV_X1 _21408_ (.A(_11704_),
    .ZN(_11720_));
 AOI21_X1 _21409_ (.A(_11714_),
    .B1(_11719_),
    .B2(_11720_),
    .ZN(_11721_));
 AND2_X4 _21410_ (.A1(_11666_),
    .A2(_11637_),
    .ZN(_11722_));
 INV_X1 _21411_ (.A(_11722_),
    .ZN(_11723_));
 AND2_X2 _21412_ (.A1(_11642_),
    .A2(_11626_),
    .ZN(_11724_));
 INV_X1 _21413_ (.A(_11724_),
    .ZN(_11725_));
 NAND2_X1 _21414_ (.A1(_11723_),
    .A2(_11725_),
    .ZN(_11726_));
 BUF_X4 _21415_ (.A(_11713_),
    .Z(_11727_));
 AND2_X1 _21416_ (.A1(_11726_),
    .A2(_11727_),
    .ZN(_11728_));
 OR2_X1 _21417_ (.A1(_11721_),
    .A2(_11728_),
    .ZN(_11729_));
 AND2_X4 _21418_ (.A1(_11711_),
    .A2(_11662_),
    .ZN(_11730_));
 BUF_X8 _21419_ (.A(_11730_),
    .Z(_11731_));
 BUF_X4 _21420_ (.A(_11731_),
    .Z(_11732_));
 BUF_X4 _21421_ (.A(_11665_),
    .Z(_11733_));
 BUF_X4 _21422_ (.A(_16773_),
    .Z(_11734_));
 BUF_X4 _21423_ (.A(_11666_),
    .Z(_11735_));
 OAI221_X1 _21424_ (.A(_11732_),
    .B1(_11733_),
    .B2(_11734_),
    .C1(_11629_),
    .C2(_11735_),
    .ZN(_11736_));
 BUF_X4 _21425_ (.A(_11701_),
    .Z(_11737_));
 OAI211_X2 _21426_ (.A(_11732_),
    .B(_11737_),
    .C1(_11733_),
    .C2(_11734_),
    .ZN(_11738_));
 INV_X1 _21427_ (.A(_11731_),
    .ZN(_11739_));
 OAI211_X2 _21428_ (.A(_11736_),
    .B(_11738_),
    .C1(_11739_),
    .C2(_11720_),
    .ZN(_11740_));
 INV_X1 _21429_ (.A(_11653_),
    .ZN(_11741_));
 NOR2_X1 _21430_ (.A1(_11741_),
    .A2(_11626_),
    .ZN(_11742_));
 AND2_X2 _21431_ (.A1(_11681_),
    .A2(_11711_),
    .ZN(_11743_));
 BUF_X4 _21432_ (.A(_11743_),
    .Z(_11744_));
 NAND3_X1 _21433_ (.A1(_11742_),
    .A2(_11744_),
    .A3(_11638_),
    .ZN(_11745_));
 AND2_X4 _21434_ (.A1(_11668_),
    .A2(_11636_),
    .ZN(_11746_));
 BUF_X4 _21435_ (.A(_11746_),
    .Z(_11747_));
 AND2_X4 _21436_ (.A1(_11669_),
    .A2(_11734_),
    .ZN(_11748_));
 BUF_X8 _21437_ (.A(_11748_),
    .Z(_11749_));
 OAI21_X4 _21438_ (.A(_11744_),
    .B1(_11747_),
    .B2(_11749_),
    .ZN(_11750_));
 AND2_X4 _21439_ (.A1(_11638_),
    .A2(_11666_),
    .ZN(_11751_));
 NAND2_X1 _21440_ (.A1(_11743_),
    .A2(_11751_),
    .ZN(_11752_));
 NOR3_X1 _21441_ (.A1(_11626_),
    .A2(_16775_),
    .A3(_16774_),
    .ZN(_11753_));
 NAND2_X1 _21442_ (.A1(_11743_),
    .A2(_11753_),
    .ZN(_11754_));
 NAND4_X1 _21443_ (.A1(_11745_),
    .A2(_11750_),
    .A3(_11752_),
    .A4(_11754_),
    .ZN(_11755_));
 AND2_X4 _21444_ (.A1(_11697_),
    .A2(_11711_),
    .ZN(_11756_));
 AND2_X2 _21445_ (.A1(_11659_),
    .A2(_11756_),
    .ZN(_11757_));
 AND2_X4 _21446_ (.A1(_11658_),
    .A2(_11665_),
    .ZN(_11758_));
 AND2_X2 _21447_ (.A1(_11756_),
    .A2(_11758_),
    .ZN(_11759_));
 NOR2_X1 _21448_ (.A1(_11757_),
    .A2(_11759_),
    .ZN(_11760_));
 BUF_X4 _21449_ (.A(_11672_),
    .Z(_11761_));
 BUF_X4 _21450_ (.A(_11697_),
    .Z(_11762_));
 NAND4_X1 _21451_ (.A1(_11761_),
    .A2(_11737_),
    .A3(_11712_),
    .A4(_11762_),
    .ZN(_11763_));
 BUF_X4 _21452_ (.A(_11756_),
    .Z(_11764_));
 BUF_X8 _21453_ (.A(_11643_),
    .Z(_11765_));
 OAI211_X2 _21454_ (.A(_11764_),
    .B(_11673_),
    .C1(_11733_),
    .C2(_11765_),
    .ZN(_11766_));
 NAND3_X1 _21455_ (.A1(_11764_),
    .A2(_11735_),
    .A3(_11637_),
    .ZN(_11767_));
 NAND4_X1 _21456_ (.A1(_11760_),
    .A2(_11763_),
    .A3(_11766_),
    .A4(_11767_),
    .ZN(_11768_));
 NOR4_X2 _21457_ (.A1(_11729_),
    .A2(_11740_),
    .A3(_11755_),
    .A4(_11768_),
    .ZN(_11769_));
 INV_X32 _21458_ (.A(_16779_),
    .ZN(_11770_));
 AND2_X4 _21459_ (.A1(_11770_),
    .A2(_16778_),
    .ZN(_11771_));
 AND2_X4 _21460_ (.A1(_11771_),
    .A2(_11663_),
    .ZN(_11772_));
 AND2_X1 _21461_ (.A1(_11772_),
    .A2(_11702_),
    .ZN(_11773_));
 AND2_X4 _21462_ (.A1(_11657_),
    .A2(_11668_),
    .ZN(_11774_));
 BUF_X8 _21463_ (.A(_11774_),
    .Z(_11775_));
 OAI21_X2 _21464_ (.A(_11772_),
    .B1(_11775_),
    .B2(_11670_),
    .ZN(_11776_));
 BUF_X4 _21465_ (.A(_11771_),
    .Z(_11777_));
 NAND4_X1 _21466_ (.A1(_11777_),
    .A2(_11665_),
    .A3(_11666_),
    .A4(_11663_),
    .ZN(_11778_));
 NAND2_X1 _21467_ (.A1(_11776_),
    .A2(_11778_),
    .ZN(_11779_));
 BUF_X4 _21468_ (.A(_11772_),
    .Z(_11780_));
 AND2_X2 _21469_ (.A1(_11658_),
    .A2(_11643_),
    .ZN(_11781_));
 BUF_X4 _21470_ (.A(_11781_),
    .Z(_11782_));
 AOI211_X2 _21471_ (.A(_11773_),
    .B(_11779_),
    .C1(_11780_),
    .C2(_11782_),
    .ZN(_11783_));
 AND2_X4 _21472_ (.A1(_11771_),
    .A2(_11681_),
    .ZN(_11784_));
 AND2_X4 _21473_ (.A1(_11784_),
    .A2(_11775_),
    .ZN(_11785_));
 INV_X2 _21474_ (.A(_11785_),
    .ZN(_11786_));
 NOR2_X2 _21475_ (.A1(_11679_),
    .A2(_11672_),
    .ZN(_11787_));
 INV_X1 _21476_ (.A(_11787_),
    .ZN(_11788_));
 INV_X2 _21477_ (.A(_11784_),
    .ZN(_11789_));
 OAI21_X1 _21478_ (.A(_11786_),
    .B1(_11788_),
    .B2(_11789_),
    .ZN(_11790_));
 BUF_X8 _21479_ (.A(_11784_),
    .Z(_11791_));
 BUF_X8 _21480_ (.A(_11685_),
    .Z(_11792_));
 AND2_X1 _21481_ (.A1(_11791_),
    .A2(_11792_),
    .ZN(_11793_));
 AND2_X2 _21482_ (.A1(_11653_),
    .A2(_16773_),
    .ZN(_11794_));
 INV_X1 _21483_ (.A(_11794_),
    .ZN(_11795_));
 AOI21_X1 _21484_ (.A(_11789_),
    .B1(_11795_),
    .B2(_11692_),
    .ZN(_11796_));
 AND2_X4 _21485_ (.A1(_11652_),
    .A2(_11676_),
    .ZN(_11797_));
 AND2_X2 _21486_ (.A1(_11791_),
    .A2(_11797_),
    .ZN(_11798_));
 NOR4_X1 _21487_ (.A1(_11790_),
    .A2(_11793_),
    .A3(_11796_),
    .A4(_11798_),
    .ZN(_11799_));
 AND2_X4 _21488_ (.A1(_11771_),
    .A2(_11632_),
    .ZN(_11800_));
 AND2_X1 _21489_ (.A1(_11800_),
    .A2(_11794_),
    .ZN(_11801_));
 INV_X1 _21490_ (.A(_11801_),
    .ZN(_11802_));
 BUF_X8 _21491_ (.A(_11800_),
    .Z(_11803_));
 AND2_X1 _21492_ (.A1(_11666_),
    .A2(_11665_),
    .ZN(_11804_));
 AND2_X4 _21493_ (.A1(_11668_),
    .A2(_11626_),
    .ZN(_11805_));
 OAI21_X1 _21494_ (.A(_11803_),
    .B1(_11804_),
    .B2(_11805_),
    .ZN(_11806_));
 NAND2_X2 _21495_ (.A1(_11803_),
    .A2(_11781_),
    .ZN(_11807_));
 NAND2_X1 _21496_ (.A1(_11800_),
    .A2(_11792_),
    .ZN(_11808_));
 AND4_X1 _21497_ (.A1(_11802_),
    .A2(_11806_),
    .A3(_11807_),
    .A4(_11808_),
    .ZN(_11809_));
 AND2_X4 _21498_ (.A1(_11771_),
    .A2(_11697_),
    .ZN(_11810_));
 NAND3_X1 _21499_ (.A1(_11810_),
    .A2(_11638_),
    .A3(_11629_),
    .ZN(_11811_));
 NAND3_X1 _21500_ (.A1(_11724_),
    .A2(_11762_),
    .A3(_11777_),
    .ZN(_11812_));
 NAND2_X1 _21501_ (.A1(_11811_),
    .A2(_11812_),
    .ZN(_11813_));
 INV_X4 _21502_ (.A(_11810_),
    .ZN(_11814_));
 INV_X1 _21503_ (.A(_11781_),
    .ZN(_11815_));
 AOI21_X1 _21504_ (.A(_11814_),
    .B1(_11686_),
    .B2(_11815_),
    .ZN(_11816_));
 BUF_X8 _21505_ (.A(_11810_),
    .Z(_11817_));
 AND2_X4 _21506_ (.A1(_11701_),
    .A2(_11665_),
    .ZN(_11818_));
 AOI211_X2 _21507_ (.A(_11813_),
    .B(_11816_),
    .C1(_11817_),
    .C2(_11818_),
    .ZN(_11819_));
 AND4_X2 _21508_ (.A1(_11783_),
    .A2(_11799_),
    .A3(_11809_),
    .A4(_11819_),
    .ZN(_11820_));
 NOR2_X4 _21509_ (.A1(_11770_),
    .A2(_16778_),
    .ZN(_11821_));
 AND2_X2 _21510_ (.A1(_11631_),
    .A2(_11821_),
    .ZN(_11822_));
 BUF_X4 _21511_ (.A(_11822_),
    .Z(_11823_));
 AND3_X1 _21512_ (.A1(_11823_),
    .A2(_11638_),
    .A3(_11753_),
    .ZN(_11824_));
 AOI21_X1 _21513_ (.A(_11824_),
    .B1(_11823_),
    .B2(_11749_),
    .ZN(_11825_));
 CLKBUF_X3 _21514_ (.A(_11821_),
    .Z(_11826_));
 AND4_X1 _21515_ (.A1(_11665_),
    .A2(_11666_),
    .A3(_11826_),
    .A4(_11663_),
    .ZN(_11827_));
 NOR2_X2 _21516_ (.A1(_11741_),
    .A2(_11657_),
    .ZN(_11828_));
 AND2_X4 _21517_ (.A1(_11821_),
    .A2(_11663_),
    .ZN(_11829_));
 NAND2_X2 _21518_ (.A1(_11828_),
    .A2(_11829_),
    .ZN(_11830_));
 INV_X1 _21519_ (.A(_11829_),
    .ZN(_11831_));
 AND2_X4 _21520_ (.A1(_11676_),
    .A2(_11651_),
    .ZN(_11832_));
 INV_X4 _21521_ (.A(_11832_),
    .ZN(_11833_));
 OAI21_X2 _21522_ (.A(_11830_),
    .B1(_11831_),
    .B2(_11833_),
    .ZN(_11834_));
 NOR3_X1 _21523_ (.A1(_11636_),
    .A2(_11627_),
    .A3(_11628_),
    .ZN(_11835_));
 AOI211_X4 _21524_ (.A(_11827_),
    .B(_11834_),
    .C1(_11829_),
    .C2(_11835_),
    .ZN(_11836_));
 AND2_X2 _21525_ (.A1(_11681_),
    .A2(_11821_),
    .ZN(_11837_));
 BUF_X4 _21526_ (.A(_11837_),
    .Z(_11838_));
 BUF_X8 _21527_ (.A(_11670_),
    .Z(_11839_));
 OAI21_X2 _21528_ (.A(_11838_),
    .B1(_11839_),
    .B2(_11805_),
    .ZN(_11840_));
 BUF_X4 _21529_ (.A(_11681_),
    .Z(_11841_));
 NAND4_X1 _21530_ (.A1(_11841_),
    .A2(_11735_),
    .A3(_11699_),
    .A4(_11826_),
    .ZN(_11842_));
 NAND2_X1 _21531_ (.A1(_11840_),
    .A2(_11842_),
    .ZN(_11843_));
 AND2_X1 _21532_ (.A1(_11837_),
    .A2(_11702_),
    .ZN(_11844_));
 NOR2_X1 _21533_ (.A1(_11843_),
    .A2(_11844_),
    .ZN(_11845_));
 AND2_X2 _21534_ (.A1(_11821_),
    .A2(_11697_),
    .ZN(_11846_));
 INV_X2 _21535_ (.A(_11658_),
    .ZN(_11847_));
 NOR2_X2 _21536_ (.A1(_11847_),
    .A2(_11652_),
    .ZN(_11848_));
 AND2_X1 _21537_ (.A1(_11846_),
    .A2(_11848_),
    .ZN(_11849_));
 INV_X1 _21538_ (.A(_11657_),
    .ZN(_11850_));
 AND3_X1 _21539_ (.A1(_11846_),
    .A2(_11850_),
    .A3(_11701_),
    .ZN(_11851_));
 BUF_X4 _21540_ (.A(_11846_),
    .Z(_11852_));
 AOI211_X2 _21541_ (.A(_11849_),
    .B(_11851_),
    .C1(_11747_),
    .C2(_11852_),
    .ZN(_11853_));
 AND4_X4 _21542_ (.A1(_11825_),
    .A2(_11836_),
    .A3(_11845_),
    .A4(_11853_),
    .ZN(_11854_));
 NAND4_X1 _21543_ (.A1(_11710_),
    .A2(_11769_),
    .A3(_11820_),
    .A4(_11854_),
    .ZN(_11855_));
 AND2_X1 _21544_ (.A1(_11732_),
    .A2(_11687_),
    .ZN(_11856_));
 NOR2_X2 _21545_ (.A1(_11855_),
    .A2(_11856_),
    .ZN(_11857_));
 AND2_X2 _21546_ (.A1(_11642_),
    .A2(_11652_),
    .ZN(_11858_));
 AND2_X1 _21547_ (.A1(_11858_),
    .A2(_11698_),
    .ZN(_11859_));
 INV_X1 _21548_ (.A(_11859_),
    .ZN(_11860_));
 AOI211_X2 _21549_ (.A(_11847_),
    .B(_11684_),
    .C1(_11665_),
    .C2(_11734_),
    .ZN(_11861_));
 INV_X4 _21550_ (.A(_11805_),
    .ZN(_11862_));
 INV_X2 _21551_ (.A(_11746_),
    .ZN(_11863_));
 NAND2_X4 _21552_ (.A1(_11862_),
    .A2(_11863_),
    .ZN(_11864_));
 AND2_X4 _21553_ (.A1(_11864_),
    .A2(_11682_),
    .ZN(_11865_));
 NAND2_X2 _21554_ (.A1(_11682_),
    .A2(_11794_),
    .ZN(_11866_));
 OAI21_X2 _21555_ (.A(_11866_),
    .B1(_11684_),
    .B2(_11715_),
    .ZN(_11867_));
 NOR4_X2 _21556_ (.A1(_11861_),
    .A2(_11683_),
    .A3(_11865_),
    .A4(_11867_),
    .ZN(_11868_));
 AND2_X4 _21557_ (.A1(_11669_),
    .A2(_11651_),
    .ZN(_11869_));
 NAND2_X1 _21558_ (.A1(_11705_),
    .A2(_11869_),
    .ZN(_11870_));
 OAI21_X1 _21559_ (.A(_11705_),
    .B1(_11691_),
    .B2(_11753_),
    .ZN(_11871_));
 AND4_X2 _21560_ (.A1(_11860_),
    .A2(_11868_),
    .A3(_11870_),
    .A4(_11871_),
    .ZN(_11872_));
 AND2_X1 _21561_ (.A1(_11644_),
    .A2(_11664_),
    .ZN(_11873_));
 INV_X1 _21562_ (.A(_11873_),
    .ZN(_11874_));
 AND2_X2 _21563_ (.A1(_11641_),
    .A2(_11724_),
    .ZN(_11875_));
 NAND2_X2 _21564_ (.A1(_11716_),
    .A2(_11641_),
    .ZN(_11876_));
 NAND2_X1 _21565_ (.A1(_11660_),
    .A2(_11876_),
    .ZN(_11877_));
 AND2_X4 _21566_ (.A1(_11850_),
    .A2(_11669_),
    .ZN(_11878_));
 AOI211_X2 _21567_ (.A(_11875_),
    .B(_11877_),
    .C1(_11641_),
    .C2(_11878_),
    .ZN(_11879_));
 BUF_X4 _21568_ (.A(_11664_),
    .Z(_11880_));
 NOR3_X1 _21569_ (.A1(_11637_),
    .A2(_16775_),
    .A3(_11628_),
    .ZN(_11881_));
 OAI21_X1 _21570_ (.A(_11880_),
    .B1(_11881_),
    .B2(_11687_),
    .ZN(_11882_));
 OAI211_X2 _21571_ (.A(_11880_),
    .B(_11673_),
    .C1(_11733_),
    .C2(_11734_),
    .ZN(_11883_));
 AND4_X4 _21572_ (.A1(_11874_),
    .A2(_11879_),
    .A3(_11882_),
    .A4(_11883_),
    .ZN(_11884_));
 OAI21_X1 _21573_ (.A(_11823_),
    .B1(_11794_),
    .B2(_11758_),
    .ZN(_11885_));
 INV_X4 _21574_ (.A(_11858_),
    .ZN(_11886_));
 AND2_X2 _21575_ (.A1(_11642_),
    .A2(_11657_),
    .ZN(_11887_));
 INV_X1 _21576_ (.A(_11887_),
    .ZN(_11888_));
 NAND2_X2 _21577_ (.A1(_11886_),
    .A2(_11888_),
    .ZN(_11889_));
 OAI21_X1 _21578_ (.A(_11823_),
    .B1(_11889_),
    .B2(_11864_),
    .ZN(_11890_));
 AND2_X1 _21579_ (.A1(_11644_),
    .A2(_11829_),
    .ZN(_11891_));
 INV_X1 _21580_ (.A(_11891_),
    .ZN(_11892_));
 AND4_X1 _21581_ (.A1(_11699_),
    .A2(_11701_),
    .A3(_11826_),
    .A4(_11663_),
    .ZN(_11893_));
 AOI21_X1 _21582_ (.A(_11893_),
    .B1(_11689_),
    .B2(_11829_),
    .ZN(_11894_));
 AND4_X1 _21583_ (.A1(_11885_),
    .A2(_11890_),
    .A3(_11892_),
    .A4(_11894_),
    .ZN(_11895_));
 NOR2_X1 _21584_ (.A1(_11775_),
    .A2(_11648_),
    .ZN(_11896_));
 INV_X1 _21585_ (.A(_11852_),
    .ZN(_11897_));
 NOR2_X1 _21586_ (.A1(_11896_),
    .A2(_11897_),
    .ZN(_11898_));
 INV_X1 _21587_ (.A(_11898_),
    .ZN(_11899_));
 AND2_X1 _21588_ (.A1(_11838_),
    .A2(_11687_),
    .ZN(_11900_));
 INV_X1 _21589_ (.A(_11900_),
    .ZN(_11901_));
 BUF_X4 _21590_ (.A(_11651_),
    .Z(_11902_));
 OAI221_X1 _21591_ (.A(_11838_),
    .B1(_11902_),
    .B2(_11765_),
    .C1(_11735_),
    .C2(_11673_),
    .ZN(_11903_));
 OAI21_X1 _21592_ (.A(_11852_),
    .B1(_11828_),
    .B2(_11781_),
    .ZN(_11904_));
 AND4_X1 _21593_ (.A1(_11899_),
    .A2(_11901_),
    .A3(_11903_),
    .A4(_11904_),
    .ZN(_11905_));
 NAND4_X4 _21594_ (.A1(_11872_),
    .A2(_11884_),
    .A3(_11895_),
    .A4(_11905_),
    .ZN(_11906_));
 AND2_X2 _21595_ (.A1(_11817_),
    .A2(_11644_),
    .ZN(_11907_));
 AND2_X1 _21596_ (.A1(_11810_),
    .A2(_11887_),
    .ZN(_11908_));
 AND2_X1 _21597_ (.A1(_11810_),
    .A2(_11835_),
    .ZN(_11909_));
 OR3_X4 _21598_ (.A1(_11907_),
    .A2(_11908_),
    .A3(_11909_),
    .ZN(_11910_));
 AND2_X2 _21599_ (.A1(_11653_),
    .A2(_11626_),
    .ZN(_11911_));
 NAND2_X1 _21600_ (.A1(_11817_),
    .A2(_11911_),
    .ZN(_11912_));
 NAND2_X1 _21601_ (.A1(_11817_),
    .A2(_11691_),
    .ZN(_11913_));
 INV_X4 _21602_ (.A(_11758_),
    .ZN(_11914_));
 OAI211_X2 _21603_ (.A(_11912_),
    .B(_11913_),
    .C1(_11814_),
    .C2(_11914_),
    .ZN(_11915_));
 NAND2_X1 _21604_ (.A1(_11791_),
    .A2(_11704_),
    .ZN(_11916_));
 NAND2_X2 _21605_ (.A1(_11791_),
    .A2(_11911_),
    .ZN(_11917_));
 OAI211_X2 _21606_ (.A(_11916_),
    .B(_11917_),
    .C1(_11789_),
    .C2(_11815_),
    .ZN(_11918_));
 INV_X2 _21607_ (.A(_11748_),
    .ZN(_11919_));
 AOI21_X1 _21608_ (.A(_11789_),
    .B1(_11886_),
    .B2(_11919_),
    .ZN(_11920_));
 NOR4_X4 _21609_ (.A1(_11910_),
    .A2(_11915_),
    .A3(_11918_),
    .A4(_11920_),
    .ZN(_11921_));
 INV_X2 _21610_ (.A(_11800_),
    .ZN(_11922_));
 INV_X1 _21611_ (.A(_11889_),
    .ZN(_11923_));
 AOI21_X1 _21612_ (.A(_11922_),
    .B1(_11923_),
    .B2(_11862_),
    .ZN(_11924_));
 INV_X1 _21613_ (.A(_11772_),
    .ZN(_11925_));
 INV_X1 _21614_ (.A(_11797_),
    .ZN(_11926_));
 INV_X1 _21615_ (.A(_11911_),
    .ZN(_11927_));
 AOI21_X1 _21616_ (.A(_11925_),
    .B1(_11926_),
    .B2(_11927_),
    .ZN(_11928_));
 INV_X1 _21617_ (.A(_11695_),
    .ZN(_11929_));
 AOI21_X1 _21618_ (.A(_11925_),
    .B1(_11649_),
    .B2(_11929_),
    .ZN(_11930_));
 OAI21_X2 _21619_ (.A(_11800_),
    .B1(_11655_),
    .B2(_11716_),
    .ZN(_11931_));
 OAI21_X1 _21620_ (.A(_11931_),
    .B1(_11914_),
    .B2(_11922_),
    .ZN(_11932_));
 NOR4_X1 _21621_ (.A1(_11924_),
    .A2(_11928_),
    .A3(_11930_),
    .A4(_11932_),
    .ZN(_11933_));
 AND2_X1 _21622_ (.A1(_11743_),
    .A2(_11794_),
    .ZN(_11934_));
 INV_X1 _21623_ (.A(_11934_),
    .ZN(_11935_));
 AND2_X4 _21624_ (.A1(_11652_),
    .A2(_11669_),
    .ZN(_11936_));
 AND3_X4 _21625_ (.A1(_11936_),
    .A2(_11712_),
    .A3(_11681_),
    .ZN(_11937_));
 INV_X1 _21626_ (.A(_11937_),
    .ZN(_11938_));
 NAND4_X1 _21627_ (.A1(_11935_),
    .A2(_11938_),
    .A3(_11752_),
    .A4(_11754_),
    .ZN(_11939_));
 AND2_X1 _21628_ (.A1(_11818_),
    .A2(_11756_),
    .ZN(_11940_));
 INV_X1 _21629_ (.A(_11756_),
    .ZN(_11941_));
 INV_X4 _21630_ (.A(_11869_),
    .ZN(_11942_));
 AOI21_X1 _21631_ (.A(_11941_),
    .B1(_11649_),
    .B2(_11942_),
    .ZN(_11943_));
 NOR4_X1 _21632_ (.A1(_11939_),
    .A2(_11759_),
    .A3(_11940_),
    .A4(_11943_),
    .ZN(_11944_));
 INV_X1 _21633_ (.A(_11652_),
    .ZN(_11945_));
 NAND4_X1 _21634_ (.A1(_11731_),
    .A2(_11850_),
    .A3(_11945_),
    .A4(_11737_),
    .ZN(_11946_));
 NAND2_X1 _21635_ (.A1(_11670_),
    .A2(_11731_),
    .ZN(_11947_));
 NAND3_X1 _21636_ (.A1(_11731_),
    .A2(_11672_),
    .A3(_11669_),
    .ZN(_11948_));
 AND3_X1 _21637_ (.A1(_11946_),
    .A2(_11947_),
    .A3(_11948_),
    .ZN(_11949_));
 NAND3_X1 _21638_ (.A1(_11828_),
    .A2(_11945_),
    .A3(_11713_),
    .ZN(_11950_));
 NAND3_X1 _21639_ (.A1(_11781_),
    .A2(_11632_),
    .A3(_11712_),
    .ZN(_11951_));
 NAND4_X1 _21640_ (.A1(_11632_),
    .A2(_11672_),
    .A3(_11676_),
    .A4(_11712_),
    .ZN(_11952_));
 AND3_X1 _21641_ (.A1(_11950_),
    .A2(_11951_),
    .A3(_11952_),
    .ZN(_11953_));
 OAI21_X1 _21642_ (.A(_11727_),
    .B1(_11645_),
    .B2(_11648_),
    .ZN(_11954_));
 OAI21_X1 _21643_ (.A(_11713_),
    .B1(_11805_),
    .B2(_11670_),
    .ZN(_11955_));
 AND4_X1 _21644_ (.A1(_11949_),
    .A2(_11953_),
    .A3(_11954_),
    .A4(_11955_),
    .ZN(_11956_));
 NAND4_X2 _21645_ (.A1(_11921_),
    .A2(_11933_),
    .A3(_11944_),
    .A4(_11956_),
    .ZN(_11957_));
 NOR2_X4 _21646_ (.A1(_11906_),
    .A2(_11957_),
    .ZN(_11958_));
 XOR2_X2 _21647_ (.A(_11857_),
    .B(_11958_),
    .Z(_11959_));
 XNOR2_X1 _21648_ (.A(_11625_),
    .B(_11959_),
    .ZN(_11960_));
 AND2_X4 _21649_ (.A1(_16867_),
    .A2(_16866_),
    .ZN(_11961_));
 NOR2_X4 _21650_ (.A1(_16865_),
    .A2(_16864_),
    .ZN(_11962_));
 AND2_X2 _21651_ (.A1(_11961_),
    .A2(_11962_),
    .ZN(_11963_));
 BUF_X4 _21652_ (.A(_11963_),
    .Z(_11964_));
 INV_X32 _21653_ (.A(_16862_),
    .ZN(_11965_));
 NOR2_X4 _21654_ (.A1(_11965_),
    .A2(_16863_),
    .ZN(_11966_));
 BUF_X4 _21655_ (.A(_11966_),
    .Z(_11967_));
 BUF_X32 _21656_ (.A(_16860_),
    .Z(_11968_));
 BUF_X4 _21657_ (.A(_11968_),
    .Z(_11969_));
 BUF_X4 _21658_ (.A(_16861_),
    .Z(_11970_));
 OAI211_X2 _21659_ (.A(_11964_),
    .B(_11967_),
    .C1(_11969_),
    .C2(_11970_),
    .ZN(_11971_));
 AND2_X4 _21660_ (.A1(_16863_),
    .A2(_16862_),
    .ZN(_11972_));
 AND2_X1 _21661_ (.A1(_11972_),
    .A2(_16861_),
    .ZN(_11973_));
 AND2_X4 _21662_ (.A1(_11963_),
    .A2(_11973_),
    .ZN(_11974_));
 INV_X32 _21663_ (.A(_16863_),
    .ZN(_11975_));
 NOR2_X4 _21664_ (.A1(_11975_),
    .A2(_16862_),
    .ZN(_11976_));
 INV_X32 _21665_ (.A(_16861_),
    .ZN(_11977_));
 AND2_X4 _21666_ (.A1(_11976_),
    .A2(_11977_),
    .ZN(_11978_));
 AND2_X1 _21667_ (.A1(_11978_),
    .A2(_11963_),
    .ZN(_11979_));
 INV_X32 _21668_ (.A(_16860_),
    .ZN(_11980_));
 NOR2_X2 _21669_ (.A1(_11980_),
    .A2(_16861_),
    .ZN(_11981_));
 BUF_X8 _21670_ (.A(_11972_),
    .Z(_11982_));
 AND2_X1 _21671_ (.A1(_11981_),
    .A2(_11982_),
    .ZN(_11983_));
 AOI211_X4 _21672_ (.A(_11974_),
    .B(_11979_),
    .C1(_11983_),
    .C2(_11963_),
    .ZN(_11984_));
 BUF_X4 _21673_ (.A(_11961_),
    .Z(_11985_));
 NOR2_X4 _21674_ (.A1(_11968_),
    .A2(_16861_),
    .ZN(_11986_));
 BUF_X8 _21675_ (.A(_11986_),
    .Z(_11987_));
 NOR2_X1 _21676_ (.A1(_16863_),
    .A2(_16862_),
    .ZN(_11988_));
 BUF_X4 _21677_ (.A(_11988_),
    .Z(_11989_));
 BUF_X4 _21678_ (.A(_11989_),
    .Z(_11990_));
 NAND4_X1 _21679_ (.A1(_11985_),
    .A2(_11987_),
    .A3(_11990_),
    .A4(_11962_),
    .ZN(_11991_));
 INV_X32 _21680_ (.A(_16865_),
    .ZN(_11992_));
 AND2_X4 _21681_ (.A1(_11992_),
    .A2(_16864_),
    .ZN(_11993_));
 AND2_X1 _21682_ (.A1(_11993_),
    .A2(_11961_),
    .ZN(_11994_));
 BUF_X4 _21683_ (.A(_11994_),
    .Z(_11995_));
 NOR2_X4 _21684_ (.A1(_11977_),
    .A2(_11968_),
    .ZN(_11996_));
 AND2_X2 _21685_ (.A1(_11996_),
    .A2(_11989_),
    .ZN(_11997_));
 NAND2_X1 _21686_ (.A1(_11995_),
    .A2(_11997_),
    .ZN(_11998_));
 BUF_X4 _21687_ (.A(_11982_),
    .Z(_11999_));
 BUF_X4 _21688_ (.A(_11977_),
    .Z(_12000_));
 OAI211_X2 _21689_ (.A(_11994_),
    .B(_11999_),
    .C1(_11968_),
    .C2(_12000_),
    .ZN(_12001_));
 AND2_X1 _21690_ (.A1(_11996_),
    .A2(_11966_),
    .ZN(_12002_));
 NAND2_X1 _21691_ (.A1(_11995_),
    .A2(_12002_),
    .ZN(_12003_));
 AND2_X4 _21692_ (.A1(_11968_),
    .A2(_16861_),
    .ZN(_12004_));
 AND2_X4 _21693_ (.A1(_11976_),
    .A2(_12004_),
    .ZN(_12005_));
 NAND2_X1 _21694_ (.A1(_11995_),
    .A2(_12005_),
    .ZN(_12006_));
 AND4_X1 _21695_ (.A1(_11998_),
    .A2(_12001_),
    .A3(_12003_),
    .A4(_12006_),
    .ZN(_12007_));
 AND4_X1 _21696_ (.A1(_11971_),
    .A2(_11984_),
    .A3(_11991_),
    .A4(_12007_),
    .ZN(_12008_));
 AND2_X1 _21697_ (.A1(_11966_),
    .A2(_16861_),
    .ZN(_12009_));
 NOR2_X4 _21698_ (.A1(_11992_),
    .A2(_16864_),
    .ZN(_12010_));
 AND2_X4 _21699_ (.A1(_12010_),
    .A2(_11985_),
    .ZN(_12011_));
 BUF_X4 _21700_ (.A(_12011_),
    .Z(_12012_));
 AND2_X1 _21701_ (.A1(_12009_),
    .A2(_12012_),
    .ZN(_12013_));
 INV_X1 _21702_ (.A(_12013_),
    .ZN(_12014_));
 AND2_X2 _21703_ (.A1(_11989_),
    .A2(_12000_),
    .ZN(_12015_));
 AND2_X1 _21704_ (.A1(_12012_),
    .A2(_12015_),
    .ZN(_12016_));
 INV_X1 _21705_ (.A(_12016_),
    .ZN(_12017_));
 NAND2_X1 _21706_ (.A1(_11997_),
    .A2(_12012_),
    .ZN(_12018_));
 AND2_X2 _21707_ (.A1(_11981_),
    .A2(_11966_),
    .ZN(_12019_));
 NAND2_X1 _21708_ (.A1(_12019_),
    .A2(_12012_),
    .ZN(_12020_));
 NAND4_X1 _21709_ (.A1(_12014_),
    .A2(_12017_),
    .A3(_12018_),
    .A4(_12020_),
    .ZN(_12021_));
 AND2_X4 _21710_ (.A1(_11972_),
    .A2(_11987_),
    .ZN(_12022_));
 AND2_X1 _21711_ (.A1(_12011_),
    .A2(_12022_),
    .ZN(_12023_));
 BUF_X8 _21712_ (.A(_12004_),
    .Z(_12024_));
 AND2_X4 _21713_ (.A1(_12024_),
    .A2(_11982_),
    .ZN(_12025_));
 BUF_X2 _21714_ (.A(_12010_),
    .Z(_12026_));
 AND3_X1 _21715_ (.A1(_12025_),
    .A2(_12026_),
    .A3(_11985_),
    .ZN(_12027_));
 NOR2_X1 _21716_ (.A1(_12023_),
    .A2(_12027_),
    .ZN(_12028_));
 INV_X1 _21717_ (.A(_12028_),
    .ZN(_12029_));
 BUF_X8 _21718_ (.A(_11976_),
    .Z(_12030_));
 BUF_X4 _21719_ (.A(_11996_),
    .Z(_12031_));
 OAI211_X2 _21720_ (.A(_12012_),
    .B(_12030_),
    .C1(_12024_),
    .C2(_12031_),
    .ZN(_12032_));
 NAND4_X1 _21721_ (.A1(_12026_),
    .A2(_12030_),
    .A3(_11987_),
    .A4(_11985_),
    .ZN(_12033_));
 NAND2_X1 _21722_ (.A1(_12032_),
    .A2(_12033_),
    .ZN(_12034_));
 AND2_X4 _21723_ (.A1(_16865_),
    .A2(_16864_),
    .ZN(_12035_));
 AND2_X1 _21724_ (.A1(_11985_),
    .A2(_12035_),
    .ZN(_12036_));
 BUF_X4 _21725_ (.A(_12036_),
    .Z(_12037_));
 AND2_X4 _21726_ (.A1(_11976_),
    .A2(_11981_),
    .ZN(_12038_));
 BUF_X4 _21727_ (.A(_12038_),
    .Z(_12039_));
 AND2_X1 _21728_ (.A1(_11982_),
    .A2(_11980_),
    .ZN(_12040_));
 OAI21_X1 _21729_ (.A(_12037_),
    .B1(_12039_),
    .B2(_12040_),
    .ZN(_12041_));
 OAI211_X2 _21730_ (.A(_12037_),
    .B(_11989_),
    .C1(_11980_),
    .C2(_12000_),
    .ZN(_12042_));
 INV_X1 _21731_ (.A(_12036_),
    .ZN(_12043_));
 AND2_X2 _21732_ (.A1(_11966_),
    .A2(_11977_),
    .ZN(_12044_));
 INV_X2 _21733_ (.A(_12044_),
    .ZN(_12045_));
 OAI211_X2 _21734_ (.A(_12041_),
    .B(_12042_),
    .C1(_12043_),
    .C2(_12045_),
    .ZN(_12046_));
 NOR4_X2 _21735_ (.A1(_12021_),
    .A2(_12029_),
    .A3(_12034_),
    .A4(_12046_),
    .ZN(_12047_));
 AND2_X4 _21736_ (.A1(_12004_),
    .A2(_11989_),
    .ZN(_12048_));
 INV_X1 _21737_ (.A(_12048_),
    .ZN(_12049_));
 AND2_X2 _21738_ (.A1(_11987_),
    .A2(_11989_),
    .ZN(_12050_));
 INV_X1 _21739_ (.A(_12050_),
    .ZN(_12051_));
 NAND2_X1 _21740_ (.A1(_12049_),
    .A2(_12051_),
    .ZN(_12052_));
 INV_X32 _21741_ (.A(_16866_),
    .ZN(_12053_));
 AND2_X2 _21742_ (.A1(_12053_),
    .A2(_16867_),
    .ZN(_12054_));
 AND2_X1 _21743_ (.A1(_12054_),
    .A2(_11962_),
    .ZN(_12055_));
 BUF_X2 _21744_ (.A(_12055_),
    .Z(_12056_));
 NAND2_X1 _21745_ (.A1(_12052_),
    .A2(_12056_),
    .ZN(_12057_));
 INV_X1 _21746_ (.A(_12055_),
    .ZN(_12058_));
 INV_X1 _21747_ (.A(_12019_),
    .ZN(_12059_));
 OAI21_X1 _21748_ (.A(_12057_),
    .B1(_12058_),
    .B2(_12059_),
    .ZN(_12060_));
 AND2_X4 _21749_ (.A1(_12054_),
    .A2(_11993_),
    .ZN(_12061_));
 BUF_X8 _21750_ (.A(_12061_),
    .Z(_12062_));
 INV_X1 _21751_ (.A(_12062_),
    .ZN(_12063_));
 INV_X4 _21752_ (.A(_11986_),
    .ZN(_12064_));
 NAND2_X1 _21753_ (.A1(_12064_),
    .A2(_11976_),
    .ZN(_12065_));
 NOR2_X1 _21754_ (.A1(_12065_),
    .A2(_12024_),
    .ZN(_12066_));
 INV_X1 _21755_ (.A(_12066_),
    .ZN(_12067_));
 BUF_X4 _21756_ (.A(_12022_),
    .Z(_12068_));
 NOR2_X4 _21757_ (.A1(_12025_),
    .A2(_12068_),
    .ZN(_12069_));
 AOI21_X1 _21758_ (.A(_12063_),
    .B1(_12067_),
    .B2(_12069_),
    .ZN(_12070_));
 AND2_X1 _21759_ (.A1(_11988_),
    .A2(_11968_),
    .ZN(_12071_));
 INV_X1 _21760_ (.A(_12071_),
    .ZN(_12072_));
 INV_X1 _21761_ (.A(_12009_),
    .ZN(_12073_));
 AOI21_X1 _21762_ (.A(_12063_),
    .B1(_12072_),
    .B2(_12073_),
    .ZN(_12074_));
 BUF_X2 _21763_ (.A(_11978_),
    .Z(_12075_));
 AND2_X1 _21764_ (.A1(_12056_),
    .A2(_12075_),
    .ZN(_12076_));
 NOR4_X1 _21765_ (.A1(_12060_),
    .A2(_12070_),
    .A3(_12074_),
    .A4(_12076_),
    .ZN(_12077_));
 AND2_X1 _21766_ (.A1(_12054_),
    .A2(_12035_),
    .ZN(_12078_));
 BUF_X4 _21767_ (.A(_12078_),
    .Z(_12079_));
 AND2_X2 _21768_ (.A1(_12030_),
    .A2(_11970_),
    .ZN(_12080_));
 AND2_X1 _21769_ (.A1(_12079_),
    .A2(_12080_),
    .ZN(_12081_));
 AND2_X2 _21770_ (.A1(_11996_),
    .A2(_11982_),
    .ZN(_12082_));
 AND2_X1 _21771_ (.A1(_12079_),
    .A2(_12082_),
    .ZN(_12083_));
 NOR2_X1 _21772_ (.A1(_12081_),
    .A2(_12083_),
    .ZN(_12084_));
 AND2_X2 _21773_ (.A1(_12054_),
    .A2(_12026_),
    .ZN(_12085_));
 AND2_X1 _21774_ (.A1(_12085_),
    .A2(_12050_),
    .ZN(_12086_));
 INV_X1 _21775_ (.A(_12086_),
    .ZN(_12087_));
 BUF_X4 _21776_ (.A(_12085_),
    .Z(_12088_));
 BUF_X4 _21777_ (.A(_11980_),
    .Z(_12089_));
 BUF_X4 _21778_ (.A(_12030_),
    .Z(_12090_));
 OAI221_X1 _21779_ (.A(_12088_),
    .B1(_12089_),
    .B2(_12000_),
    .C1(_12090_),
    .C2(_11999_),
    .ZN(_12091_));
 INV_X1 _21780_ (.A(_11966_),
    .ZN(_12092_));
 NOR2_X1 _21781_ (.A1(_12092_),
    .A2(_11996_),
    .ZN(_12093_));
 OAI21_X1 _21782_ (.A(_12079_),
    .B1(_12093_),
    .B2(_12015_),
    .ZN(_12094_));
 AND4_X1 _21783_ (.A1(_12084_),
    .A2(_12087_),
    .A3(_12091_),
    .A4(_12094_),
    .ZN(_12095_));
 NAND4_X1 _21784_ (.A1(_12008_),
    .A2(_12047_),
    .A3(_12077_),
    .A4(_12095_),
    .ZN(_12096_));
 NOR2_X1 _21785_ (.A1(_12053_),
    .A2(_16867_),
    .ZN(_12097_));
 AND2_X4 _21786_ (.A1(_12097_),
    .A2(_12035_),
    .ZN(_12098_));
 AND2_X1 _21787_ (.A1(_11978_),
    .A2(_12098_),
    .ZN(_12099_));
 AND2_X1 _21788_ (.A1(_11976_),
    .A2(_11996_),
    .ZN(_12100_));
 AND2_X1 _21789_ (.A1(_12098_),
    .A2(_11982_),
    .ZN(_12101_));
 AOI221_X1 _21790_ (.A(_12099_),
    .B1(_12100_),
    .B2(_12098_),
    .C1(_12064_),
    .C2(_12101_),
    .ZN(_12102_));
 AND2_X1 _21791_ (.A1(_12098_),
    .A2(_12071_),
    .ZN(_12103_));
 INV_X1 _21792_ (.A(_12103_),
    .ZN(_12104_));
 OAI211_X2 _21793_ (.A(_12098_),
    .B(_11967_),
    .C1(_11968_),
    .C2(_12000_),
    .ZN(_12105_));
 AND2_X1 _21794_ (.A1(_12104_),
    .A2(_12105_),
    .ZN(_12106_));
 AND2_X1 _21795_ (.A1(_12026_),
    .A2(_12097_),
    .ZN(_12107_));
 BUF_X4 _21796_ (.A(_12107_),
    .Z(_12108_));
 AND2_X2 _21797_ (.A1(_11966_),
    .A2(_12004_),
    .ZN(_12109_));
 OAI21_X1 _21798_ (.A(_12108_),
    .B1(_12109_),
    .B2(_11990_),
    .ZN(_12110_));
 OAI21_X1 _21799_ (.A(_12108_),
    .B1(_12039_),
    .B2(_11973_),
    .ZN(_12111_));
 AND4_X1 _21800_ (.A1(_12102_),
    .A2(_12106_),
    .A3(_12110_),
    .A4(_12111_),
    .ZN(_12112_));
 NOR2_X4 _21801_ (.A1(_16867_),
    .A2(_16866_),
    .ZN(_12113_));
 AND2_X2 _21802_ (.A1(_11993_),
    .A2(_12113_),
    .ZN(_12114_));
 AND2_X1 _21803_ (.A1(_12114_),
    .A2(_12080_),
    .ZN(_12115_));
 INV_X1 _21804_ (.A(_12115_),
    .ZN(_12116_));
 BUF_X4 _21805_ (.A(_12114_),
    .Z(_12117_));
 AND2_X4 _21806_ (.A1(_11982_),
    .A2(_11977_),
    .ZN(_12118_));
 BUF_X4 _21807_ (.A(_12118_),
    .Z(_12119_));
 NAND2_X1 _21808_ (.A1(_12117_),
    .A2(_12119_),
    .ZN(_12120_));
 NAND2_X1 _21809_ (.A1(_12117_),
    .A2(_12025_),
    .ZN(_12121_));
 AND2_X2 _21810_ (.A1(_11976_),
    .A2(_11987_),
    .ZN(_12122_));
 OAI21_X1 _21811_ (.A(_12114_),
    .B1(_12039_),
    .B2(_12122_),
    .ZN(_12123_));
 NAND4_X1 _21812_ (.A1(_12116_),
    .A2(_12120_),
    .A3(_12121_),
    .A4(_12123_),
    .ZN(_12124_));
 AND2_X2 _21813_ (.A1(_12113_),
    .A2(_11962_),
    .ZN(_12125_));
 AND2_X1 _21814_ (.A1(_12082_),
    .A2(_12125_),
    .ZN(_12126_));
 INV_X1 _21815_ (.A(_12126_),
    .ZN(_12127_));
 AND2_X4 _21816_ (.A1(_11966_),
    .A2(_11987_),
    .ZN(_12128_));
 OAI21_X1 _21817_ (.A(_12125_),
    .B1(_12109_),
    .B2(_12128_),
    .ZN(_12129_));
 INV_X1 _21818_ (.A(_12118_),
    .ZN(_12130_));
 INV_X1 _21819_ (.A(_12125_),
    .ZN(_12131_));
 OAI211_X2 _21820_ (.A(_12127_),
    .B(_12129_),
    .C1(_12130_),
    .C2(_12131_),
    .ZN(_12132_));
 INV_X1 _21821_ (.A(_12109_),
    .ZN(_12133_));
 INV_X1 _21822_ (.A(_12128_),
    .ZN(_12134_));
 NAND2_X1 _21823_ (.A1(_12133_),
    .A2(_12134_),
    .ZN(_12135_));
 AND2_X1 _21824_ (.A1(_12135_),
    .A2(_12114_),
    .ZN(_12136_));
 NAND2_X1 _21825_ (.A1(_12114_),
    .A2(_12015_),
    .ZN(_12137_));
 INV_X1 _21826_ (.A(_12114_),
    .ZN(_12138_));
 INV_X1 _21827_ (.A(_11997_),
    .ZN(_12139_));
 OAI21_X1 _21828_ (.A(_12137_),
    .B1(_12138_),
    .B2(_12139_),
    .ZN(_12140_));
 NOR4_X1 _21829_ (.A1(_12124_),
    .A2(_12132_),
    .A3(_12136_),
    .A4(_12140_),
    .ZN(_12141_));
 AND2_X2 _21830_ (.A1(_11993_),
    .A2(_12097_),
    .ZN(_12142_));
 INV_X2 _21831_ (.A(_12142_),
    .ZN(_12143_));
 INV_X2 _21832_ (.A(_12025_),
    .ZN(_12144_));
 AOI21_X1 _21833_ (.A(_12143_),
    .B1(_12067_),
    .B2(_12144_),
    .ZN(_12145_));
 NAND2_X1 _21834_ (.A1(_12142_),
    .A2(_12019_),
    .ZN(_12146_));
 NAND3_X1 _21835_ (.A1(_12002_),
    .A2(_11993_),
    .A3(_12097_),
    .ZN(_12147_));
 OAI211_X2 _21836_ (.A(_12146_),
    .B(_12147_),
    .C1(_12143_),
    .C2(_12072_),
    .ZN(_12148_));
 AND2_X2 _21837_ (.A1(_12097_),
    .A2(_11962_),
    .ZN(_12149_));
 BUF_X4 _21838_ (.A(_12149_),
    .Z(_12150_));
 INV_X2 _21839_ (.A(_12150_),
    .ZN(_12151_));
 AND2_X2 _21840_ (.A1(_11981_),
    .A2(_11989_),
    .ZN(_12152_));
 INV_X1 _21841_ (.A(_12152_),
    .ZN(_12153_));
 AOI21_X1 _21842_ (.A(_12151_),
    .B1(_12153_),
    .B2(_12133_),
    .ZN(_12154_));
 INV_X1 _21843_ (.A(_12080_),
    .ZN(_12155_));
 AND2_X2 _21844_ (.A1(_11982_),
    .A2(_11968_),
    .ZN(_12156_));
 INV_X1 _21845_ (.A(_12156_),
    .ZN(_12157_));
 AOI21_X1 _21846_ (.A(_12151_),
    .B1(_12155_),
    .B2(_12157_),
    .ZN(_12158_));
 NOR4_X1 _21847_ (.A1(_12145_),
    .A2(_12148_),
    .A3(_12154_),
    .A4(_12158_),
    .ZN(_12159_));
 AND2_X4 _21848_ (.A1(_12035_),
    .A2(_12113_),
    .ZN(_12160_));
 BUF_X4 _21849_ (.A(_12160_),
    .Z(_12161_));
 BUF_X4 _21850_ (.A(_12161_),
    .Z(_12162_));
 BUF_X4 _21851_ (.A(_12080_),
    .Z(_12163_));
 OAI21_X1 _21852_ (.A(_12162_),
    .B1(_12163_),
    .B2(_12040_),
    .ZN(_12164_));
 AND2_X4 _21853_ (.A1(_12026_),
    .A2(_12113_),
    .ZN(_12165_));
 AND3_X1 _21854_ (.A1(_12165_),
    .A2(_12030_),
    .A3(_12064_),
    .ZN(_12166_));
 BUF_X4 _21855_ (.A(_12165_),
    .Z(_12167_));
 BUF_X4 _21856_ (.A(_11983_),
    .Z(_12168_));
 AOI21_X1 _21857_ (.A(_12166_),
    .B1(_12167_),
    .B2(_12168_),
    .ZN(_12169_));
 NOR3_X1 _21858_ (.A1(_12024_),
    .A2(_16863_),
    .A3(_16862_),
    .ZN(_12170_));
 OAI21_X1 _21859_ (.A(_12167_),
    .B1(_12009_),
    .B2(_12170_),
    .ZN(_12171_));
 OAI211_X2 _21860_ (.A(_12161_),
    .B(_11969_),
    .C1(_11990_),
    .C2(_11967_),
    .ZN(_12172_));
 AND4_X1 _21861_ (.A1(_12164_),
    .A2(_12169_),
    .A3(_12171_),
    .A4(_12172_),
    .ZN(_12173_));
 NAND4_X1 _21862_ (.A1(_12112_),
    .A2(_12141_),
    .A3(_12159_),
    .A4(_12173_),
    .ZN(_12174_));
 NOR2_X4 _21863_ (.A1(_12096_),
    .A2(_12174_),
    .ZN(_12175_));
 INV_X1 _21864_ (.A(_12175_),
    .ZN(_12176_));
 XNOR2_X1 _21865_ (.A(_11960_),
    .B(_12176_),
    .ZN(_12177_));
 XNOR2_X1 _21866_ (.A(_12177_),
    .B(_17240_),
    .ZN(_12178_));
 MUX2_X1 _21867_ (.A(_11150_),
    .B(_12178_),
    .S(_11149_),
    .Z(_00716_));
 XOR2_X1 _21868_ (.A(_17251_),
    .B(_17066_),
    .Z(_12179_));
 NAND2_X1 _21869_ (.A1(_11641_),
    .A2(_11794_),
    .ZN(_12180_));
 OAI211_X2 _21870_ (.A(_11656_),
    .B(_12180_),
    .C1(_11647_),
    .C2(_11914_),
    .ZN(_12181_));
 AOI21_X1 _21871_ (.A(_11647_),
    .B1(_11863_),
    .B2(_11862_),
    .ZN(_12182_));
 AND4_X1 _21872_ (.A1(_11632_),
    .A2(_11735_),
    .A3(_11672_),
    .A4(_11635_),
    .ZN(_12183_));
 NOR3_X1 _21873_ (.A1(_12181_),
    .A2(_12182_),
    .A3(_12183_),
    .ZN(_12184_));
 INV_X2 _21874_ (.A(_11865_),
    .ZN(_12185_));
 NAND3_X1 _21875_ (.A1(_11887_),
    .A2(_11635_),
    .A3(_11841_),
    .ZN(_12186_));
 INV_X1 _21876_ (.A(_11644_),
    .ZN(_12187_));
 OAI211_X2 _21877_ (.A(_12185_),
    .B(_12186_),
    .C1(_12187_),
    .C2(_11684_),
    .ZN(_12188_));
 AND2_X2 _21878_ (.A1(_11682_),
    .A2(_11716_),
    .ZN(_12189_));
 INV_X4 _21879_ (.A(_11698_),
    .ZN(_12190_));
 AOI21_X1 _21880_ (.A(_12190_),
    .B1(_11717_),
    .B2(_11692_),
    .ZN(_12191_));
 AOI21_X1 _21881_ (.A(_12190_),
    .B1(_11725_),
    .B2(_11919_),
    .ZN(_12192_));
 NOR4_X1 _21882_ (.A1(_12188_),
    .A2(_12189_),
    .A3(_12191_),
    .A4(_12192_),
    .ZN(_12193_));
 OAI21_X1 _21883_ (.A(_11880_),
    .B1(_11689_),
    .B2(_11818_),
    .ZN(_12194_));
 AND2_X1 _21884_ (.A1(_11746_),
    .A2(_11664_),
    .ZN(_12195_));
 AND2_X1 _21885_ (.A1(_11724_),
    .A2(_11664_),
    .ZN(_12196_));
 AOI211_X2 _21886_ (.A(_12195_),
    .B(_12196_),
    .C1(_11748_),
    .C2(_11664_),
    .ZN(_12197_));
 AND4_X2 _21887_ (.A1(_12184_),
    .A2(_12193_),
    .A3(_12194_),
    .A4(_12197_),
    .ZN(_12198_));
 OAI21_X1 _21888_ (.A(_11780_),
    .B1(_11742_),
    .B2(_11758_),
    .ZN(_12199_));
 BUF_X4 _21889_ (.A(_11648_),
    .Z(_12200_));
 OAI21_X1 _21890_ (.A(_11780_),
    .B1(_11645_),
    .B2(_12200_),
    .ZN(_12201_));
 BUF_X4 _21891_ (.A(_11936_),
    .Z(_12202_));
 OAI21_X1 _21892_ (.A(_11780_),
    .B1(_11775_),
    .B2(_12202_),
    .ZN(_12203_));
 AND3_X1 _21893_ (.A1(_12199_),
    .A2(_12201_),
    .A3(_12203_),
    .ZN(_12204_));
 NOR2_X1 _21894_ (.A1(_11847_),
    .A2(_11636_),
    .ZN(_12205_));
 AND2_X1 _21895_ (.A1(_11784_),
    .A2(_12205_),
    .ZN(_12206_));
 OAI21_X1 _21896_ (.A(_11786_),
    .B1(_11649_),
    .B2(_11789_),
    .ZN(_12207_));
 AND2_X1 _21897_ (.A1(_11737_),
    .A2(_11651_),
    .ZN(_12208_));
 AOI211_X2 _21898_ (.A(_12206_),
    .B(_12207_),
    .C1(_11791_),
    .C2(_12208_),
    .ZN(_12209_));
 AOI21_X1 _21899_ (.A(_11922_),
    .B1(_11927_),
    .B2(_11688_),
    .ZN(_12210_));
 AND4_X1 _21900_ (.A1(_11850_),
    .A2(_11800_),
    .A3(_11673_),
    .A4(_11945_),
    .ZN(_12211_));
 AND2_X1 _21901_ (.A1(_11800_),
    .A2(_11887_),
    .ZN(_12212_));
 AND2_X1 _21902_ (.A1(_11800_),
    .A2(_11644_),
    .ZN(_12213_));
 NOR4_X1 _21903_ (.A1(_12210_),
    .A2(_12211_),
    .A3(_12212_),
    .A4(_12213_),
    .ZN(_12214_));
 NAND4_X1 _21904_ (.A1(_11771_),
    .A2(_11701_),
    .A3(_11637_),
    .A4(_11762_),
    .ZN(_12215_));
 OAI21_X1 _21905_ (.A(_12215_),
    .B1(_11814_),
    .B2(_11914_),
    .ZN(_12216_));
 AOI211_X2 _21906_ (.A(_11909_),
    .B(_12216_),
    .C1(_11817_),
    .C2(_11889_),
    .ZN(_12217_));
 AND4_X2 _21907_ (.A1(_12204_),
    .A2(_12209_),
    .A3(_12214_),
    .A4(_12217_),
    .ZN(_12218_));
 AOI211_X2 _21908_ (.A(_11627_),
    .B(_11739_),
    .C1(_11643_),
    .C2(_11628_),
    .ZN(_12219_));
 AND2_X1 _21909_ (.A1(_11731_),
    .A2(_11704_),
    .ZN(_12220_));
 AND2_X1 _21910_ (.A1(_11691_),
    .A2(_11731_),
    .ZN(_12221_));
 AND3_X1 _21911_ (.A1(_11730_),
    .A2(_11657_),
    .A3(_11701_),
    .ZN(_12222_));
 NOR4_X1 _21912_ (.A1(_12219_),
    .A2(_12220_),
    .A3(_12221_),
    .A4(_12222_),
    .ZN(_12223_));
 NAND2_X1 _21913_ (.A1(_11727_),
    .A2(_12200_),
    .ZN(_12224_));
 NAND2_X1 _21914_ (.A1(_11727_),
    .A2(_11775_),
    .ZN(_12225_));
 NAND4_X1 _21915_ (.A1(_11632_),
    .A2(_11737_),
    .A3(_11902_),
    .A4(_11712_),
    .ZN(_12226_));
 AND4_X1 _21916_ (.A1(_11951_),
    .A2(_12224_),
    .A3(_12225_),
    .A4(_12226_),
    .ZN(_12227_));
 OAI21_X1 _21917_ (.A(_11744_),
    .B1(_11742_),
    .B2(_11848_),
    .ZN(_12228_));
 NAND2_X1 _21918_ (.A1(_11818_),
    .A2(_11764_),
    .ZN(_12229_));
 OAI211_X2 _21919_ (.A(_11764_),
    .B(_11666_),
    .C1(_11665_),
    .C2(_11765_),
    .ZN(_12230_));
 OAI211_X2 _21920_ (.A(_11756_),
    .B(_11673_),
    .C1(_11902_),
    .C2(_11765_),
    .ZN(_12231_));
 AND4_X1 _21921_ (.A1(_11760_),
    .A2(_12229_),
    .A3(_12230_),
    .A4(_12231_),
    .ZN(_12232_));
 AND4_X4 _21922_ (.A1(_12223_),
    .A2(_12227_),
    .A3(_12228_),
    .A4(_12232_),
    .ZN(_12233_));
 AND2_X1 _21923_ (.A1(_11838_),
    .A2(_11655_),
    .ZN(_12234_));
 AND2_X2 _21924_ (.A1(_11837_),
    .A2(_11704_),
    .ZN(_12235_));
 AND2_X2 _21925_ (.A1(_11787_),
    .A2(_11837_),
    .ZN(_12236_));
 AND2_X1 _21926_ (.A1(_11837_),
    .A2(_11797_),
    .ZN(_12237_));
 OR4_X4 _21927_ (.A1(_12234_),
    .A2(_12235_),
    .A3(_12236_),
    .A4(_12237_),
    .ZN(_12238_));
 AND2_X1 _21928_ (.A1(_11823_),
    .A2(_11691_),
    .ZN(_12239_));
 AND2_X1 _21929_ (.A1(_11822_),
    .A2(_11659_),
    .ZN(_12240_));
 AND2_X2 _21930_ (.A1(_11822_),
    .A2(_11669_),
    .ZN(_12241_));
 AND2_X1 _21931_ (.A1(_11822_),
    .A2(_11644_),
    .ZN(_12242_));
 OR4_X4 _21932_ (.A1(_12239_),
    .A2(_12240_),
    .A3(_12241_),
    .A4(_12242_),
    .ZN(_12243_));
 BUF_X4 _21933_ (.A(_11829_),
    .Z(_12244_));
 OAI211_X2 _21934_ (.A(_12244_),
    .B(_11735_),
    .C1(_11761_),
    .C2(_11699_),
    .ZN(_12245_));
 BUF_X2 _21935_ (.A(_11663_),
    .Z(_12246_));
 NAND4_X1 _21936_ (.A1(_11672_),
    .A2(_11826_),
    .A3(_11676_),
    .A4(_12246_),
    .ZN(_12247_));
 NAND2_X1 _21937_ (.A1(_12244_),
    .A2(_11805_),
    .ZN(_12248_));
 NAND4_X1 _21938_ (.A1(_12245_),
    .A2(_11830_),
    .A3(_12247_),
    .A4(_12248_),
    .ZN(_12249_));
 AND2_X2 _21939_ (.A1(_11629_),
    .A2(_11638_),
    .ZN(_12250_));
 OAI21_X2 _21940_ (.A(_11852_),
    .B1(_12250_),
    .B2(_11804_),
    .ZN(_12251_));
 NAND2_X1 _21941_ (.A1(_11716_),
    .A2(_11852_),
    .ZN(_12252_));
 OAI211_X2 _21942_ (.A(_12251_),
    .B(_12252_),
    .C1(_11897_),
    .C2(_11833_),
    .ZN(_12253_));
 NOR4_X4 _21943_ (.A1(_12238_),
    .A2(_12243_),
    .A3(_12249_),
    .A4(_12253_),
    .ZN(_12254_));
 NAND4_X4 _21944_ (.A1(_12198_),
    .A2(_12218_),
    .A3(_12233_),
    .A4(_12254_),
    .ZN(_12255_));
 NOR2_X2 _21945_ (.A1(_12255_),
    .A2(_11856_),
    .ZN(_12256_));
 AND3_X4 _21946_ (.A1(_11277_),
    .A2(_11203_),
    .A3(_11340_),
    .ZN(_12257_));
 AND3_X1 _21947_ (.A1(_11207_),
    .A2(_11203_),
    .A3(_11340_),
    .ZN(_12258_));
 AND2_X4 _21948_ (.A1(_16813_),
    .A2(_16815_),
    .ZN(_12259_));
 NOR2_X1 _21949_ (.A1(_16812_),
    .A2(_16814_),
    .ZN(_12260_));
 AND2_X2 _21950_ (.A1(_12259_),
    .A2(_12260_),
    .ZN(_12261_));
 BUF_X8 _21951_ (.A(_12261_),
    .Z(_12262_));
 AOI211_X2 _21952_ (.A(_12257_),
    .B(_12258_),
    .C1(_12262_),
    .C2(_11342_),
    .ZN(_12263_));
 NAND4_X1 _21953_ (.A1(_11326_),
    .A2(_11209_),
    .A3(_11341_),
    .A4(_11322_),
    .ZN(_12264_));
 BUF_X4 _21954_ (.A(_11163_),
    .Z(_12265_));
 OAI211_X2 _21955_ (.A(_11342_),
    .B(_12265_),
    .C1(_11213_),
    .C2(_11209_),
    .ZN(_12266_));
 AND3_X1 _21956_ (.A1(_12263_),
    .A2(_12264_),
    .A3(_12266_),
    .ZN(_12267_));
 INV_X1 _21957_ (.A(_11201_),
    .ZN(_12268_));
 AOI21_X1 _21958_ (.A(_11369_),
    .B1(_11359_),
    .B2(_12268_),
    .ZN(_12269_));
 AND2_X1 _21959_ (.A1(_11184_),
    .A2(_11368_),
    .ZN(_12270_));
 AND2_X1 _21960_ (.A1(_11277_),
    .A2(_11368_),
    .ZN(_12271_));
 AND2_X1 _21961_ (.A1(_11279_),
    .A2(_11368_),
    .ZN(_12272_));
 NOR4_X1 _21962_ (.A1(_12269_),
    .A2(_12270_),
    .A3(_12271_),
    .A4(_12272_),
    .ZN(_12273_));
 INV_X1 _21963_ (.A(_11244_),
    .ZN(_12274_));
 INV_X8 _21964_ (.A(_11188_),
    .ZN(_12275_));
 NOR2_X2 _21965_ (.A1(_12275_),
    .A2(_11186_),
    .ZN(_12276_));
 AND3_X1 _21966_ (.A1(_11353_),
    .A2(_12274_),
    .A3(_12276_),
    .ZN(_12277_));
 NAND2_X1 _21967_ (.A1(_11353_),
    .A2(_11377_),
    .ZN(_12278_));
 INV_X4 _21968_ (.A(_12262_),
    .ZN(_12279_));
 OAI21_X2 _21969_ (.A(_12278_),
    .B1(_11355_),
    .B2(_12279_),
    .ZN(_12280_));
 AND2_X1 _21970_ (.A1(_11162_),
    .A2(_11186_),
    .ZN(_12281_));
 BUF_X2 _21971_ (.A(_12281_),
    .Z(_12282_));
 AOI211_X2 _21972_ (.A(_12277_),
    .B(_12280_),
    .C1(_12282_),
    .C2(_11353_),
    .ZN(_12283_));
 AND2_X1 _21973_ (.A1(_11360_),
    .A2(_11373_),
    .ZN(_12284_));
 INV_X4 _21974_ (.A(_11373_),
    .ZN(_12285_));
 AOI21_X1 _21975_ (.A(_12285_),
    .B1(_11185_),
    .B2(_11280_),
    .ZN(_12286_));
 AOI211_X2 _21976_ (.A(_12284_),
    .B(_12286_),
    .C1(_12281_),
    .C2(_11373_),
    .ZN(_12287_));
 AND4_X2 _21977_ (.A1(_12267_),
    .A2(_12273_),
    .A3(_12283_),
    .A4(_12287_),
    .ZN(_12288_));
 OAI21_X1 _21978_ (.A(_11222_),
    .B1(_11282_),
    .B2(_11160_),
    .ZN(_12289_));
 OAI21_X1 _21979_ (.A(_11222_),
    .B1(_11377_),
    .B2(_11379_),
    .ZN(_12290_));
 OAI211_X2 _21980_ (.A(_11222_),
    .B(_11258_),
    .C1(_11244_),
    .C2(_11217_),
    .ZN(_12291_));
 AND3_X1 _21981_ (.A1(_12289_),
    .A2(_12290_),
    .A3(_12291_),
    .ZN(_12292_));
 AND2_X1 _21982_ (.A1(_11156_),
    .A2(_11295_),
    .ZN(_12293_));
 NAND2_X4 _21983_ (.A1(_11156_),
    .A2(_11190_),
    .ZN(_12294_));
 INV_X4 _21984_ (.A(_11156_),
    .ZN(_12295_));
 OAI21_X2 _21985_ (.A(_12294_),
    .B1(_12295_),
    .B2(_11251_),
    .ZN(_12296_));
 AND2_X1 _21986_ (.A1(_11163_),
    .A2(_11321_),
    .ZN(_12297_));
 AOI211_X2 _21987_ (.A(_12293_),
    .B(_12296_),
    .C1(_11156_),
    .C2(_12297_),
    .ZN(_12298_));
 NAND2_X1 _21988_ (.A1(_11204_),
    .A2(_11377_),
    .ZN(_12299_));
 OAI21_X1 _21989_ (.A(_12299_),
    .B1(_11205_),
    .B2(_12279_),
    .ZN(_12300_));
 AND2_X2 _21990_ (.A1(_11162_),
    .A2(_11172_),
    .ZN(_12301_));
 INV_X1 _21991_ (.A(_12301_),
    .ZN(_12302_));
 AOI21_X1 _21992_ (.A(_11205_),
    .B1(_11357_),
    .B2(_12302_),
    .ZN(_12303_));
 NAND2_X1 _21993_ (.A1(_11208_),
    .A2(_11278_),
    .ZN(_12304_));
 AOI211_X2 _21994_ (.A(_12300_),
    .B(_12303_),
    .C1(_11204_),
    .C2(_12304_),
    .ZN(_12305_));
 AND2_X1 _21995_ (.A1(_11170_),
    .A2(_11160_),
    .ZN(_12306_));
 INV_X1 _21996_ (.A(_12306_),
    .ZN(_12307_));
 NOR2_X1 _21997_ (.A1(_12275_),
    .A2(_11269_),
    .ZN(_12308_));
 NAND2_X1 _21998_ (.A1(_12308_),
    .A2(_11171_),
    .ZN(_12309_));
 NAND4_X1 _21999_ (.A1(_12265_),
    .A2(_11167_),
    .A3(_11269_),
    .A4(_11169_),
    .ZN(_12310_));
 NAND3_X1 _22000_ (.A1(_11286_),
    .A2(_11171_),
    .A3(_11256_),
    .ZN(_12311_));
 AND4_X2 _22001_ (.A1(_12307_),
    .A2(_12309_),
    .A3(_12310_),
    .A4(_12311_),
    .ZN(_12312_));
 AND4_X2 _22002_ (.A1(_12292_),
    .A2(_12298_),
    .A3(_12305_),
    .A4(_12312_),
    .ZN(_12313_));
 NOR2_X1 _22003_ (.A1(_11216_),
    .A2(_11244_),
    .ZN(_12314_));
 OAI21_X1 _22004_ (.A(_11275_),
    .B1(_11282_),
    .B2(_12314_),
    .ZN(_12315_));
 INV_X1 _22005_ (.A(_11377_),
    .ZN(_12316_));
 AOI21_X1 _22006_ (.A(_11290_),
    .B1(_12316_),
    .B2(_11185_),
    .ZN(_12317_));
 AOI21_X1 _22007_ (.A(_11290_),
    .B1(_11191_),
    .B2(_11291_),
    .ZN(_12318_));
 AND2_X1 _22008_ (.A1(_11201_),
    .A2(_11289_),
    .ZN(_12319_));
 NOR4_X1 _22009_ (.A1(_12317_),
    .A2(_12318_),
    .A3(_11296_),
    .A4(_12319_),
    .ZN(_12320_));
 AND2_X1 _22010_ (.A1(_11282_),
    .A2(_11253_),
    .ZN(_12321_));
 AND2_X1 _22011_ (.A1(_11229_),
    .A2(_11242_),
    .ZN(_12322_));
 AND2_X1 _22012_ (.A1(_11242_),
    .A2(_12259_),
    .ZN(_12323_));
 NOR4_X1 _22013_ (.A1(_12321_),
    .A2(_11255_),
    .A3(_12322_),
    .A4(_12323_),
    .ZN(_12324_));
 AND2_X1 _22014_ (.A1(_11264_),
    .A2(_11379_),
    .ZN(_12325_));
 AND2_X1 _22015_ (.A1(_11264_),
    .A2(_11190_),
    .ZN(_12326_));
 BUF_X8 _22016_ (.A(_11179_),
    .Z(_12327_));
 AND2_X1 _22017_ (.A1(_11264_),
    .A2(_12327_),
    .ZN(_12328_));
 AND4_X1 _22018_ (.A1(_11321_),
    .A2(_11163_),
    .A3(_11326_),
    .A4(_11297_),
    .ZN(_12329_));
 NOR4_X2 _22019_ (.A1(_12325_),
    .A2(_12326_),
    .A3(_12328_),
    .A4(_12329_),
    .ZN(_12330_));
 AND4_X2 _22020_ (.A1(_12315_),
    .A2(_12320_),
    .A3(_12324_),
    .A4(_12330_),
    .ZN(_12331_));
 AOI21_X1 _22021_ (.A(_11312_),
    .B1(_11344_),
    .B2(_11191_),
    .ZN(_12332_));
 NAND4_X1 _22022_ (.A1(_11305_),
    .A2(_11321_),
    .A3(_11169_),
    .A4(_11159_),
    .ZN(_12333_));
 INV_X1 _22023_ (.A(_12281_),
    .ZN(_12334_));
 OAI21_X1 _22024_ (.A(_12333_),
    .B1(_12334_),
    .B2(_11312_),
    .ZN(_12335_));
 AND4_X1 _22025_ (.A1(_11209_),
    .A2(_11305_),
    .A3(_11232_),
    .A4(_11169_),
    .ZN(_12336_));
 OR3_X1 _22026_ (.A1(_12332_),
    .A2(_12335_),
    .A3(_12336_),
    .ZN(_12337_));
 NAND4_X1 _22027_ (.A1(_11305_),
    .A2(_11186_),
    .A3(_11221_),
    .A4(_11159_),
    .ZN(_12338_));
 AND2_X2 _22028_ (.A1(_11318_),
    .A2(_12338_),
    .ZN(_12339_));
 NAND3_X1 _22029_ (.A1(_11314_),
    .A2(_11286_),
    .A3(_11257_),
    .ZN(_12340_));
 INV_X1 _22030_ (.A(_11314_),
    .ZN(_12341_));
 OAI211_X2 _22031_ (.A(_12339_),
    .B(_12340_),
    .C1(_11208_),
    .C2(_12341_),
    .ZN(_12342_));
 BUF_X4 _22032_ (.A(_11360_),
    .Z(_12343_));
 OAI21_X1 _22033_ (.A(_11328_),
    .B1(_11345_),
    .B2(_12343_),
    .ZN(_12344_));
 NAND2_X1 _22034_ (.A1(_11328_),
    .A2(_11378_),
    .ZN(_12345_));
 OAI211_X2 _22035_ (.A(_12344_),
    .B(_12345_),
    .C1(_12275_),
    .C2(_11330_),
    .ZN(_12346_));
 AND2_X1 _22036_ (.A1(_11335_),
    .A2(_11238_),
    .ZN(_12347_));
 INV_X1 _22037_ (.A(_12347_),
    .ZN(_12348_));
 AND2_X4 _22038_ (.A1(_11244_),
    .A2(_11159_),
    .ZN(_12349_));
 BUF_X4 _22039_ (.A(_12349_),
    .Z(_12350_));
 NAND2_X1 _22040_ (.A1(_11336_),
    .A2(_12350_),
    .ZN(_12351_));
 NAND2_X1 _22041_ (.A1(_11335_),
    .A2(_11254_),
    .ZN(_12352_));
 NAND2_X2 _22042_ (.A1(_11336_),
    .A2(_11245_),
    .ZN(_12353_));
 NAND4_X1 _22043_ (.A1(_12348_),
    .A2(_12351_),
    .A3(_12352_),
    .A4(_12353_),
    .ZN(_12354_));
 NOR4_X4 _22044_ (.A1(_12337_),
    .A2(_12342_),
    .A3(_12346_),
    .A4(_12354_),
    .ZN(_12355_));
 NAND4_X2 _22045_ (.A1(_12288_),
    .A2(_12313_),
    .A3(_12331_),
    .A4(_12355_),
    .ZN(_12356_));
 NOR2_X2 _22046_ (.A1(_12356_),
    .A2(_11386_),
    .ZN(_12357_));
 XOR2_X2 _22047_ (.A(_12256_),
    .B(_12357_),
    .Z(_12358_));
 XOR2_X1 _22048_ (.A(_12358_),
    .B(_11959_),
    .Z(_12359_));
 AND2_X1 _22049_ (.A1(_11603_),
    .A2(_11527_),
    .ZN(_12360_));
 INV_X1 _22050_ (.A(_11577_),
    .ZN(_12361_));
 AOI21_X1 _22051_ (.A(_11523_),
    .B1(_11491_),
    .B2(_12361_),
    .ZN(_12362_));
 AND2_X1 _22052_ (.A1(_11590_),
    .A2(_11527_),
    .ZN(_12363_));
 AND2_X1 _22053_ (.A1(_11450_),
    .A2(_11527_),
    .ZN(_12364_));
 OR4_X1 _22054_ (.A1(_12360_),
    .A2(_12362_),
    .A3(_12363_),
    .A4(_12364_),
    .ZN(_12365_));
 AND2_X1 _22055_ (.A1(_11480_),
    .A2(_11441_),
    .ZN(_12366_));
 BUF_X8 _22056_ (.A(_11603_),
    .Z(_12367_));
 OAI21_X4 _22057_ (.A(_11502_),
    .B1(_11450_),
    .B2(_12367_),
    .ZN(_12368_));
 NAND2_X1 _22058_ (.A1(_11482_),
    .A2(_11501_),
    .ZN(_12369_));
 OAI211_X2 _22059_ (.A(_12368_),
    .B(_12369_),
    .C1(_11455_),
    .C2(_11513_),
    .ZN(_12370_));
 AND2_X4 _22060_ (.A1(_11600_),
    .A2(_11418_),
    .ZN(_12371_));
 INV_X1 _22061_ (.A(_12371_),
    .ZN(_12372_));
 AOI21_X1 _22062_ (.A(_11485_),
    .B1(_12372_),
    .B2(_11541_),
    .ZN(_12373_));
 NAND3_X1 _22063_ (.A1(_11434_),
    .A2(_11464_),
    .A3(_11478_),
    .ZN(_12374_));
 NAND3_X1 _22064_ (.A1(_11590_),
    .A2(_11464_),
    .A3(_11478_),
    .ZN(_12375_));
 NAND2_X2 _22065_ (.A1(_12374_),
    .A2(_12375_),
    .ZN(_12376_));
 OR4_X2 _22066_ (.A1(_12366_),
    .A2(_12370_),
    .A3(_12373_),
    .A4(_12376_),
    .ZN(_12377_));
 OAI211_X2 _22067_ (.A(_11516_),
    .B(_11412_),
    .C1(_11413_),
    .C2(_11415_),
    .ZN(_12378_));
 AND2_X2 _22068_ (.A1(_11393_),
    .A2(_11414_),
    .ZN(_12379_));
 INV_X1 _22069_ (.A(_12379_),
    .ZN(_12380_));
 OAI21_X1 _22070_ (.A(_12378_),
    .B1(_12380_),
    .B2(_11517_),
    .ZN(_12381_));
 NAND3_X1 _22071_ (.A1(_11590_),
    .A2(_11445_),
    .A3(_11478_),
    .ZN(_12382_));
 NAND2_X1 _22072_ (.A1(_11515_),
    .A2(_12367_),
    .ZN(_12383_));
 OAI221_X1 _22073_ (.A(_12382_),
    .B1(_12372_),
    .B2(_11517_),
    .C1(_11529_),
    .C2(_12383_),
    .ZN(_12384_));
 NOR4_X2 _22074_ (.A1(_12365_),
    .A2(_12377_),
    .A3(_12381_),
    .A4(_12384_),
    .ZN(_12385_));
 AND2_X1 _22075_ (.A1(_11457_),
    .A2(_11418_),
    .ZN(_12386_));
 INV_X1 _22076_ (.A(_12386_),
    .ZN(_12387_));
 AOI21_X1 _22077_ (.A(_11425_),
    .B1(_12387_),
    .B2(_11437_),
    .ZN(_12388_));
 AND2_X1 _22078_ (.A1(_11450_),
    .A2(_11424_),
    .ZN(_12389_));
 AND2_X1 _22079_ (.A1(_11511_),
    .A2(_11424_),
    .ZN(_12390_));
 NOR4_X1 _22080_ (.A1(_12388_),
    .A2(_12389_),
    .A3(_12390_),
    .A4(_11431_),
    .ZN(_12391_));
 BUF_X4 _22081_ (.A(_11465_),
    .Z(_12392_));
 INV_X1 _22082_ (.A(_11457_),
    .ZN(_12393_));
 NAND3_X1 _22083_ (.A1(_12392_),
    .A2(_11599_),
    .A3(_12393_),
    .ZN(_12394_));
 OAI21_X1 _22084_ (.A(_12392_),
    .B1(_11441_),
    .B2(_11482_),
    .ZN(_12395_));
 INV_X1 _22085_ (.A(_11427_),
    .ZN(_12396_));
 OAI21_X1 _22086_ (.A(_11442_),
    .B1(_12396_),
    .B2(_11577_),
    .ZN(_12397_));
 NAND4_X1 _22087_ (.A1(_12391_),
    .A2(_12394_),
    .A3(_12395_),
    .A4(_12397_),
    .ZN(_12398_));
 OAI21_X1 _22088_ (.A(_11392_),
    .B1(_11459_),
    .B2(_11507_),
    .ZN(_12399_));
 INV_X4 _22089_ (.A(_11391_),
    .ZN(_12400_));
 OAI211_X2 _22090_ (.A(_12399_),
    .B(_11397_),
    .C1(_12400_),
    .C2(_11455_),
    .ZN(_12401_));
 NAND2_X1 _22091_ (.A1(_11449_),
    .A2(_11391_),
    .ZN(_12402_));
 NAND3_X1 _22092_ (.A1(_11391_),
    .A2(_11600_),
    .A3(_11419_),
    .ZN(_12403_));
 AND2_X1 _22093_ (.A1(_12402_),
    .A2(_12403_),
    .ZN(_12404_));
 NAND2_X1 _22094_ (.A1(_12367_),
    .A2(_11392_),
    .ZN(_12405_));
 OAI211_X2 _22095_ (.A(_12404_),
    .B(_12405_),
    .C1(_12400_),
    .C2(_11525_),
    .ZN(_12406_));
 AND2_X1 _22096_ (.A1(_11454_),
    .A2(_11511_),
    .ZN(_12407_));
 INV_X1 _22097_ (.A(_12407_),
    .ZN(_12408_));
 AND2_X2 _22098_ (.A1(_11419_),
    .A2(_16821_),
    .ZN(_12409_));
 AND2_X1 _22099_ (.A1(_11447_),
    .A2(_12409_),
    .ZN(_12410_));
 INV_X1 _22100_ (.A(_12410_),
    .ZN(_12411_));
 AND2_X2 _22101_ (.A1(_11411_),
    .A2(_11456_),
    .ZN(_12412_));
 OAI21_X1 _22102_ (.A(_11454_),
    .B1(_12412_),
    .B2(_11561_),
    .ZN(_12413_));
 NAND3_X1 _22103_ (.A1(_12408_),
    .A2(_12411_),
    .A3(_12413_),
    .ZN(_12414_));
 NOR4_X1 _22104_ (.A1(_12398_),
    .A2(_12401_),
    .A3(_12406_),
    .A4(_12414_),
    .ZN(_12415_));
 NAND2_X1 _22105_ (.A1(_11474_),
    .A2(_11555_),
    .ZN(_12416_));
 BUF_X2 _22106_ (.A(_12409_),
    .Z(_12417_));
 OAI21_X1 _22107_ (.A(_11554_),
    .B1(_11543_),
    .B2(_12417_),
    .ZN(_12418_));
 OAI211_X2 _22108_ (.A(_11554_),
    .B(_11399_),
    .C1(_11600_),
    .C2(_11601_),
    .ZN(_12419_));
 NAND4_X1 _22109_ (.A1(_11537_),
    .A2(_11414_),
    .A3(_11599_),
    .A4(_11552_),
    .ZN(_12420_));
 AND4_X1 _22110_ (.A1(_12416_),
    .A2(_12418_),
    .A3(_12419_),
    .A4(_12420_),
    .ZN(_12421_));
 AND2_X1 _22111_ (.A1(_12396_),
    .A2(_11539_),
    .ZN(_12422_));
 INV_X1 _22112_ (.A(_11539_),
    .ZN(_12423_));
 INV_X1 _22113_ (.A(_12409_),
    .ZN(_12424_));
 AOI21_X1 _22114_ (.A(_12423_),
    .B1(_11524_),
    .B2(_12424_),
    .ZN(_12425_));
 AOI211_X4 _22115_ (.A(_12422_),
    .B(_12425_),
    .C1(_11544_),
    .C2(_12412_),
    .ZN(_12426_));
 INV_X1 _22116_ (.A(_11564_),
    .ZN(_12427_));
 INV_X1 _22117_ (.A(_11548_),
    .ZN(_12428_));
 AOI21_X1 _22118_ (.A(_12427_),
    .B1(_12428_),
    .B2(_11489_),
    .ZN(_12429_));
 NOR2_X2 _22119_ (.A1(_11400_),
    .A2(_11600_),
    .ZN(_12430_));
 AND3_X1 _22120_ (.A1(_11564_),
    .A2(_12430_),
    .A3(_12393_),
    .ZN(_12431_));
 AND2_X1 _22121_ (.A1(_11542_),
    .A2(_11564_),
    .ZN(_12432_));
 AND2_X1 _22122_ (.A1(_12371_),
    .A2(_11564_),
    .ZN(_12433_));
 NOR4_X1 _22123_ (.A1(_12429_),
    .A2(_12431_),
    .A3(_12432_),
    .A4(_12433_),
    .ZN(_12434_));
 AND3_X1 _22124_ (.A1(_11472_),
    .A2(_11407_),
    .A3(_11574_),
    .ZN(_12435_));
 AND2_X1 _22125_ (.A1(_11403_),
    .A2(_11573_),
    .ZN(_12436_));
 AND2_X1 _22126_ (.A1(_11573_),
    .A2(_12379_),
    .ZN(_12437_));
 AND4_X1 _22127_ (.A1(_11411_),
    .A2(_11537_),
    .A3(_11402_),
    .A4(_11591_),
    .ZN(_12438_));
 NOR4_X1 _22128_ (.A1(_12435_),
    .A2(_12436_),
    .A3(_12437_),
    .A4(_12438_),
    .ZN(_12439_));
 AND4_X1 _22129_ (.A1(_12421_),
    .A2(_12426_),
    .A3(_12434_),
    .A4(_12439_),
    .ZN(_12440_));
 AND2_X4 _22130_ (.A1(_11457_),
    .A2(_11398_),
    .ZN(_12441_));
 AND2_X1 _22131_ (.A1(_11587_),
    .A2(_12441_),
    .ZN(_12442_));
 INV_X1 _22132_ (.A(_12442_),
    .ZN(_12443_));
 BUF_X4 _22133_ (.A(_11587_),
    .Z(_12444_));
 INV_X1 _22134_ (.A(_12444_),
    .ZN(_12445_));
 OAI21_X1 _22135_ (.A(_12443_),
    .B1(_11524_),
    .B2(_12445_),
    .ZN(_12446_));
 AOI21_X1 _22136_ (.A(_12445_),
    .B1(_11455_),
    .B2(_11611_),
    .ZN(_12447_));
 AND4_X1 _22137_ (.A1(_11414_),
    .A2(_11592_),
    .A3(_11420_),
    .A4(_11591_),
    .ZN(_12448_));
 NOR3_X1 _22138_ (.A1(_12446_),
    .A2(_12447_),
    .A3(_12448_),
    .ZN(_12449_));
 NAND4_X1 _22139_ (.A1(_11586_),
    .A2(_11394_),
    .A3(_11600_),
    .A4(_11552_),
    .ZN(_12450_));
 AND2_X1 _22140_ (.A1(_11609_),
    .A2(_12450_),
    .ZN(_12451_));
 INV_X1 _22141_ (.A(_12451_),
    .ZN(_12452_));
 AND2_X1 _22142_ (.A1(_11607_),
    .A2(_11434_),
    .ZN(_12453_));
 AND3_X1 _22143_ (.A1(_11606_),
    .A2(_11472_),
    .A3(_11407_),
    .ZN(_12454_));
 NOR3_X1 _22144_ (.A1(_12452_),
    .A2(_12453_),
    .A3(_12454_),
    .ZN(_12455_));
 BUF_X2 _22145_ (.A(_11597_),
    .Z(_12456_));
 AND2_X1 _22146_ (.A1(_12456_),
    .A2(_11519_),
    .ZN(_12457_));
 AND2_X1 _22147_ (.A1(_12456_),
    .A2(_11399_),
    .ZN(_12458_));
 AND2_X1 _22148_ (.A1(_11597_),
    .A2(_11482_),
    .ZN(_12459_));
 AND2_X1 _22149_ (.A1(_12456_),
    .A2(_11543_),
    .ZN(_12460_));
 NOR4_X1 _22150_ (.A1(_12457_),
    .A2(_12458_),
    .A3(_12459_),
    .A4(_12460_),
    .ZN(_12461_));
 NAND3_X1 _22151_ (.A1(_11459_),
    .A2(_11464_),
    .A3(_11592_),
    .ZN(_12462_));
 BUF_X4 _22152_ (.A(_11616_),
    .Z(_12463_));
 AND2_X1 _22153_ (.A1(_12463_),
    .A2(_11543_),
    .ZN(_12464_));
 INV_X1 _22154_ (.A(_12464_),
    .ZN(_12465_));
 AND2_X1 _22155_ (.A1(_11616_),
    .A2(_11450_),
    .ZN(_12466_));
 INV_X1 _22156_ (.A(_12466_),
    .ZN(_12467_));
 OAI211_X2 _22157_ (.A(_11464_),
    .B(_11592_),
    .C1(_11500_),
    .C2(_11396_),
    .ZN(_12468_));
 AND4_X1 _22158_ (.A1(_12462_),
    .A2(_12465_),
    .A3(_12467_),
    .A4(_12468_),
    .ZN(_12469_));
 AND4_X1 _22159_ (.A1(_12449_),
    .A2(_12455_),
    .A3(_12461_),
    .A4(_12469_),
    .ZN(_12470_));
 NAND4_X1 _22160_ (.A1(_12385_),
    .A2(_12415_),
    .A3(_12440_),
    .A4(_12470_),
    .ZN(_12471_));
 NOR2_X2 _22161_ (.A1(_12471_),
    .A2(_11623_),
    .ZN(_12472_));
 XNOR2_X1 _22162_ (.A(_12359_),
    .B(_12472_),
    .ZN(_12473_));
 AND2_X1 _22163_ (.A1(_12093_),
    .A2(_12055_),
    .ZN(_12474_));
 NAND2_X2 _22164_ (.A1(_12064_),
    .A2(_11982_),
    .ZN(_12475_));
 AND2_X1 _22165_ (.A1(_12030_),
    .A2(_11968_),
    .ZN(_12476_));
 INV_X1 _22166_ (.A(_12476_),
    .ZN(_12477_));
 AOI21_X1 _22167_ (.A(_12058_),
    .B1(_12475_),
    .B2(_12477_),
    .ZN(_12478_));
 AND2_X2 _22168_ (.A1(_11988_),
    .A2(_11980_),
    .ZN(_12479_));
 AOI211_X4 _22169_ (.A(_12474_),
    .B(_12478_),
    .C1(_12056_),
    .C2(_12479_),
    .ZN(_12480_));
 AND2_X1 _22170_ (.A1(_12079_),
    .A2(_12022_),
    .ZN(_12481_));
 INV_X1 _22171_ (.A(_12078_),
    .ZN(_12482_));
 AND2_X1 _22172_ (.A1(_11988_),
    .A2(_16861_),
    .ZN(_12483_));
 BUF_X4 _22173_ (.A(_12483_),
    .Z(_12484_));
 NOR2_X1 _22174_ (.A1(_12484_),
    .A2(_12479_),
    .ZN(_12485_));
 NOR2_X1 _22175_ (.A1(_12482_),
    .A2(_12485_),
    .ZN(_12486_));
 BUF_X4 _22176_ (.A(_12079_),
    .Z(_12487_));
 AOI211_X4 _22177_ (.A(_12481_),
    .B(_12486_),
    .C1(_12487_),
    .C2(_12093_),
    .ZN(_12488_));
 NAND2_X1 _22178_ (.A1(_12064_),
    .A2(_11989_),
    .ZN(_12489_));
 INV_X1 _22179_ (.A(_12489_),
    .ZN(_12490_));
 INV_X1 _22180_ (.A(_12004_),
    .ZN(_12491_));
 AND3_X1 _22181_ (.A1(_12062_),
    .A2(_12490_),
    .A3(_12491_),
    .ZN(_12492_));
 BUF_X4 _22182_ (.A(_11973_),
    .Z(_12493_));
 AOI21_X1 _22183_ (.A(_12492_),
    .B1(_12493_),
    .B2(_12062_),
    .ZN(_12494_));
 OAI21_X1 _22184_ (.A(_12088_),
    .B1(_12025_),
    .B2(_12119_),
    .ZN(_12495_));
 BUF_X4 _22185_ (.A(_12054_),
    .Z(_12496_));
 NAND3_X1 _22186_ (.A1(_12039_),
    .A2(_12026_),
    .A3(_12496_),
    .ZN(_12497_));
 NAND2_X1 _22187_ (.A1(_12085_),
    .A2(_12128_),
    .ZN(_12498_));
 AND3_X1 _22188_ (.A1(_12495_),
    .A2(_12497_),
    .A3(_12498_),
    .ZN(_12499_));
 AND4_X1 _22189_ (.A1(_12480_),
    .A2(_12488_),
    .A3(_12494_),
    .A4(_12499_),
    .ZN(_12500_));
 NAND3_X1 _22190_ (.A1(_12125_),
    .A2(_12090_),
    .A3(_11981_),
    .ZN(_12501_));
 NAND2_X1 _22191_ (.A1(_12163_),
    .A2(_12125_),
    .ZN(_12502_));
 NOR2_X2 _22192_ (.A1(_12475_),
    .A2(_12024_),
    .ZN(_12503_));
 INV_X1 _22193_ (.A(_12503_),
    .ZN(_12504_));
 OAI211_X2 _22194_ (.A(_12501_),
    .B(_12502_),
    .C1(_12504_),
    .C2(_12131_),
    .ZN(_12505_));
 NAND2_X1 _22195_ (.A1(_12491_),
    .A2(_11966_),
    .ZN(_12506_));
 NOR2_X1 _22196_ (.A1(_12506_),
    .A2(_11987_),
    .ZN(_12507_));
 INV_X1 _22197_ (.A(_12507_),
    .ZN(_12508_));
 INV_X1 _22198_ (.A(_12484_),
    .ZN(_12509_));
 AOI21_X1 _22199_ (.A(_12138_),
    .B1(_12508_),
    .B2(_12509_),
    .ZN(_12510_));
 NAND2_X1 _22200_ (.A1(_12114_),
    .A2(_12122_),
    .ZN(_12511_));
 NAND2_X1 _22201_ (.A1(_12117_),
    .A2(_12005_),
    .ZN(_12512_));
 NAND2_X1 _22202_ (.A1(_12511_),
    .A2(_12512_),
    .ZN(_12513_));
 NAND2_X1 _22203_ (.A1(_12125_),
    .A2(_12484_),
    .ZN(_12514_));
 NAND3_X1 _22204_ (.A1(_12125_),
    .A2(_11981_),
    .A3(_11967_),
    .ZN(_12515_));
 OAI211_X2 _22205_ (.A(_12514_),
    .B(_12515_),
    .C1(_12073_),
    .C2(_12131_),
    .ZN(_12516_));
 NOR4_X1 _22206_ (.A1(_12505_),
    .A2(_12510_),
    .A3(_12513_),
    .A4(_12516_),
    .ZN(_12517_));
 OAI21_X1 _22207_ (.A(_12167_),
    .B1(_12507_),
    .B2(_12170_),
    .ZN(_12518_));
 AND2_X1 _22208_ (.A1(_12165_),
    .A2(_12022_),
    .ZN(_12519_));
 AOI211_X4 _22209_ (.A(_12166_),
    .B(_12519_),
    .C1(_12167_),
    .C2(_12493_),
    .ZN(_12520_));
 NAND3_X1 _22210_ (.A1(_12162_),
    .A2(_12031_),
    .A3(_11967_),
    .ZN(_12521_));
 NAND2_X1 _22211_ (.A1(_12490_),
    .A2(_12162_),
    .ZN(_12522_));
 OAI211_X2 _22212_ (.A(_12162_),
    .B(_11999_),
    .C1(_11969_),
    .C2(_12000_),
    .ZN(_12523_));
 NAND2_X1 _22213_ (.A1(_12122_),
    .A2(_12161_),
    .ZN(_12524_));
 AND4_X1 _22214_ (.A1(_12521_),
    .A2(_12522_),
    .A3(_12523_),
    .A4(_12524_),
    .ZN(_12525_));
 AND4_X1 _22215_ (.A1(_12517_),
    .A2(_12518_),
    .A3(_12520_),
    .A4(_12525_),
    .ZN(_12526_));
 BUF_X4 _22216_ (.A(_12108_),
    .Z(_12527_));
 BUF_X4 _22217_ (.A(_11967_),
    .Z(_12528_));
 OAI21_X1 _22218_ (.A(_12527_),
    .B1(_12071_),
    .B2(_12528_),
    .ZN(_12529_));
 AOI21_X1 _22219_ (.A(_12143_),
    .B1(_12144_),
    .B2(_12477_),
    .ZN(_12530_));
 NAND2_X1 _22220_ (.A1(_12142_),
    .A2(_12009_),
    .ZN(_12531_));
 INV_X1 _22221_ (.A(_11996_),
    .ZN(_12532_));
 NAND2_X1 _22222_ (.A1(_12532_),
    .A2(_11989_),
    .ZN(_12533_));
 OAI21_X1 _22223_ (.A(_12531_),
    .B1(_12143_),
    .B2(_12533_),
    .ZN(_12534_));
 INV_X1 _22224_ (.A(_12015_),
    .ZN(_12535_));
 AOI21_X1 _22225_ (.A(_12151_),
    .B1(_12535_),
    .B2(_12134_),
    .ZN(_12536_));
 OAI21_X4 _22226_ (.A(_12150_),
    .B1(_12082_),
    .B2(_12119_),
    .ZN(_12537_));
 NAND4_X1 _22227_ (.A1(_12030_),
    .A2(_12097_),
    .A3(_11969_),
    .A4(_11962_),
    .ZN(_12538_));
 NAND2_X1 _22228_ (.A1(_12537_),
    .A2(_12538_),
    .ZN(_12539_));
 NOR4_X1 _22229_ (.A1(_12530_),
    .A2(_12534_),
    .A3(_12536_),
    .A4(_12539_),
    .ZN(_12540_));
 NOR3_X1 _22230_ (.A1(_12031_),
    .A2(_11975_),
    .A3(_16862_),
    .ZN(_12541_));
 OAI21_X1 _22231_ (.A(_12527_),
    .B1(_12541_),
    .B2(_12082_),
    .ZN(_12542_));
 INV_X1 _22232_ (.A(_12475_),
    .ZN(_12543_));
 BUF_X8 _22233_ (.A(_12098_),
    .Z(_12544_));
 NAND3_X1 _22234_ (.A1(_12543_),
    .A2(_12491_),
    .A3(_12544_),
    .ZN(_12545_));
 NAND2_X1 _22235_ (.A1(_12005_),
    .A2(_12544_),
    .ZN(_12546_));
 NAND2_X1 _22236_ (.A1(_12545_),
    .A2(_12546_),
    .ZN(_12547_));
 NAND2_X1 _22237_ (.A1(_12152_),
    .A2(_12098_),
    .ZN(_12548_));
 INV_X1 _22238_ (.A(_12098_),
    .ZN(_12549_));
 OAI21_X1 _22239_ (.A(_12548_),
    .B1(_12549_),
    .B2(_12051_),
    .ZN(_12550_));
 AND2_X2 _22240_ (.A1(_12544_),
    .A2(_12048_),
    .ZN(_12551_));
 AND2_X2 _22241_ (.A1(_11966_),
    .A2(_11968_),
    .ZN(_12552_));
 AND2_X1 _22242_ (.A1(_12552_),
    .A2(_12098_),
    .ZN(_12553_));
 NOR4_X1 _22243_ (.A1(_12547_),
    .A2(_12550_),
    .A3(_12551_),
    .A4(_12553_),
    .ZN(_12554_));
 AND4_X2 _22244_ (.A1(_12529_),
    .A2(_12540_),
    .A3(_12542_),
    .A4(_12554_),
    .ZN(_12555_));
 AND2_X1 _22245_ (.A1(_11997_),
    .A2(_11964_),
    .ZN(_12556_));
 AND2_X1 _22246_ (.A1(_12476_),
    .A2(_11963_),
    .ZN(_12557_));
 AND3_X1 _22247_ (.A1(_11963_),
    .A2(_12031_),
    .A3(_11999_),
    .ZN(_12558_));
 AND2_X1 _22248_ (.A1(_12119_),
    .A2(_11963_),
    .ZN(_12559_));
 NOR4_X1 _22249_ (.A1(_12556_),
    .A2(_12557_),
    .A3(_12558_),
    .A4(_12559_),
    .ZN(_12560_));
 INV_X1 _22250_ (.A(_12012_),
    .ZN(_12561_));
 NOR3_X1 _22251_ (.A1(_12561_),
    .A2(_11981_),
    .A3(_12533_),
    .ZN(_12562_));
 AND2_X1 _22252_ (.A1(_12011_),
    .A2(_12156_),
    .ZN(_12563_));
 AND2_X1 _22253_ (.A1(_12012_),
    .A2(_12044_),
    .ZN(_12564_));
 NOR4_X1 _22254_ (.A1(_12034_),
    .A2(_12562_),
    .A3(_12563_),
    .A4(_12564_),
    .ZN(_12565_));
 INV_X1 _22255_ (.A(_11995_),
    .ZN(_12566_));
 OAI21_X1 _22256_ (.A(_11998_),
    .B1(_12566_),
    .B2(_12059_),
    .ZN(_12567_));
 AND3_X1 _22257_ (.A1(_12543_),
    .A2(_11995_),
    .A3(_12491_),
    .ZN(_12568_));
 AND2_X1 _22258_ (.A1(_11995_),
    .A2(_12080_),
    .ZN(_12569_));
 AND2_X1 _22259_ (.A1(_11995_),
    .A2(_12075_),
    .ZN(_12570_));
 NOR4_X1 _22260_ (.A1(_12567_),
    .A2(_12568_),
    .A3(_12569_),
    .A4(_12570_),
    .ZN(_12571_));
 AND2_X1 _22261_ (.A1(_12128_),
    .A2(_12037_),
    .ZN(_12572_));
 INV_X1 _22262_ (.A(_12572_),
    .ZN(_12573_));
 NAND2_X1 _22263_ (.A1(_12082_),
    .A2(_12037_),
    .ZN(_12574_));
 OAI211_X2 _22264_ (.A(_12037_),
    .B(_11990_),
    .C1(_11969_),
    .C2(_11970_),
    .ZN(_12575_));
 OAI21_X1 _22265_ (.A(_12037_),
    .B1(_12163_),
    .B2(_12075_),
    .ZN(_12576_));
 AND4_X1 _22266_ (.A1(_12573_),
    .A2(_12574_),
    .A3(_12575_),
    .A4(_12576_),
    .ZN(_12577_));
 AND4_X1 _22267_ (.A1(_12560_),
    .A2(_12565_),
    .A3(_12571_),
    .A4(_12577_),
    .ZN(_12578_));
 NAND4_X2 _22268_ (.A1(_12500_),
    .A2(_12526_),
    .A3(_12555_),
    .A4(_12578_),
    .ZN(_12579_));
 OAI21_X1 _22269_ (.A(_11975_),
    .B1(_12064_),
    .B2(_16862_),
    .ZN(_12580_));
 AND3_X1 _22270_ (.A1(_12113_),
    .A2(_11962_),
    .A3(_11975_),
    .ZN(_12581_));
 AND2_X1 _22271_ (.A1(_12580_),
    .A2(_12581_),
    .ZN(_12582_));
 NOR2_X4 _22272_ (.A1(_12579_),
    .A2(_12582_),
    .ZN(_12583_));
 XNOR2_X2 _22273_ (.A(_12583_),
    .B(_12176_),
    .ZN(_12584_));
 XNOR2_X1 _22274_ (.A(_12473_),
    .B(_12584_),
    .ZN(_12585_));
 XNOR2_X1 _22275_ (.A(_12585_),
    .B(_17251_),
    .ZN(_12586_));
 MUX2_X1 _22276_ (.A(_12179_),
    .B(_12586_),
    .S(_11149_),
    .Z(_00717_));
 XOR2_X1 _22277_ (.A(_17262_),
    .B(_17067_),
    .Z(_12587_));
 OAI21_X1 _22278_ (.A(_12244_),
    .B1(_11794_),
    .B2(_11691_),
    .ZN(_12588_));
 AND2_X1 _22279_ (.A1(_11823_),
    .A2(_11704_),
    .ZN(_12589_));
 INV_X1 _22280_ (.A(_11822_),
    .ZN(_12590_));
 AOI21_X1 _22281_ (.A(_12590_),
    .B1(_12187_),
    .B2(_11725_),
    .ZN(_12591_));
 AOI211_X4 _22282_ (.A(_12589_),
    .B(_12591_),
    .C1(_11839_),
    .C2(_11823_),
    .ZN(_12592_));
 OAI21_X1 _22283_ (.A(_11829_),
    .B1(_11792_),
    .B2(_11782_),
    .ZN(_12593_));
 OAI211_X2 _22284_ (.A(_12244_),
    .B(_16775_),
    .C1(_11765_),
    .C2(_11628_),
    .ZN(_12594_));
 AND4_X2 _22285_ (.A1(_12588_),
    .A2(_12592_),
    .A3(_12593_),
    .A4(_12594_),
    .ZN(_12595_));
 OAI21_X1 _22286_ (.A(_11694_),
    .B1(_11889_),
    .B2(_11878_),
    .ZN(_12596_));
 OAI21_X1 _22287_ (.A(_11705_),
    .B1(_12200_),
    .B2(_11695_),
    .ZN(_12597_));
 OAI21_X1 _22288_ (.A(_11705_),
    .B1(_11689_),
    .B2(_11691_),
    .ZN(_12598_));
 AND4_X1 _22289_ (.A1(_11866_),
    .A2(_12596_),
    .A3(_12597_),
    .A4(_12598_),
    .ZN(_12599_));
 OAI211_X2 _22290_ (.A(_11880_),
    .B(_11735_),
    .C1(_11733_),
    .C2(_11734_),
    .ZN(_12600_));
 NAND2_X1 _22291_ (.A1(_12202_),
    .A2(_11880_),
    .ZN(_12601_));
 NAND2_X2 _22292_ (.A1(_12600_),
    .A2(_12601_),
    .ZN(_12602_));
 INV_X1 _22293_ (.A(_12602_),
    .ZN(_12603_));
 BUF_X8 _22294_ (.A(_11641_),
    .Z(_12604_));
 BUF_X4 _22295_ (.A(_11735_),
    .Z(_12605_));
 OAI211_X2 _22296_ (.A(_12604_),
    .B(_12605_),
    .C1(_11761_),
    .C2(_11699_),
    .ZN(_12606_));
 NAND3_X1 _22297_ (.A1(_11747_),
    .A2(_11632_),
    .A3(_11635_),
    .ZN(_12607_));
 NAND2_X1 _22298_ (.A1(_12604_),
    .A2(_11748_),
    .ZN(_12608_));
 AND3_X1 _22299_ (.A1(_12606_),
    .A2(_12607_),
    .A3(_12608_),
    .ZN(_12609_));
 BUF_X4 _22300_ (.A(_11737_),
    .Z(_12610_));
 OAI21_X1 _22301_ (.A(_11880_),
    .B1(_11704_),
    .B2(_12610_),
    .ZN(_12611_));
 NAND2_X1 _22302_ (.A1(_11797_),
    .A2(_12604_),
    .ZN(_12612_));
 NAND2_X1 _22303_ (.A1(_12604_),
    .A2(_11704_),
    .ZN(_12613_));
 AND3_X1 _22304_ (.A1(_12180_),
    .A2(_12612_),
    .A3(_12613_),
    .ZN(_12614_));
 AND4_X1 _22305_ (.A1(_12603_),
    .A2(_12609_),
    .A3(_12611_),
    .A4(_12614_),
    .ZN(_12615_));
 OAI21_X1 _22306_ (.A(_11838_),
    .B1(_12250_),
    .B2(_11887_),
    .ZN(_12616_));
 NAND2_X1 _22307_ (.A1(_11838_),
    .A2(_11655_),
    .ZN(_12617_));
 INV_X1 _22308_ (.A(_11837_),
    .ZN(_12618_));
 OAI211_X2 _22309_ (.A(_12616_),
    .B(_12617_),
    .C1(_11795_),
    .C2(_12618_),
    .ZN(_12619_));
 BUF_X4 _22310_ (.A(_11852_),
    .Z(_12620_));
 NAND2_X1 _22311_ (.A1(_11645_),
    .A2(_12620_),
    .ZN(_12621_));
 NAND4_X1 _22312_ (.A1(_12605_),
    .A2(_11761_),
    .A3(_11826_),
    .A4(_11762_),
    .ZN(_12622_));
 OAI211_X2 _22313_ (.A(_12621_),
    .B(_12622_),
    .C1(_11942_),
    .C2(_11897_),
    .ZN(_12623_));
 OAI21_X1 _22314_ (.A(_12252_),
    .B1(_11692_),
    .B2(_11897_),
    .ZN(_12624_));
 NOR4_X1 _22315_ (.A1(_12619_),
    .A2(_12623_),
    .A3(_12624_),
    .A4(_11849_),
    .ZN(_12625_));
 NAND4_X1 _22316_ (.A1(_12595_),
    .A2(_12599_),
    .A3(_12615_),
    .A4(_12625_),
    .ZN(_12626_));
 NOR2_X1 _22317_ (.A1(_11847_),
    .A2(_11761_),
    .ZN(_12627_));
 NAND2_X1 _22318_ (.A1(_11744_),
    .A2(_12627_),
    .ZN(_12628_));
 INV_X1 _22319_ (.A(_11743_),
    .ZN(_12629_));
 OAI211_X2 _22320_ (.A(_11935_),
    .B(_12628_),
    .C1(_11692_),
    .C2(_12629_),
    .ZN(_12630_));
 AOI21_X1 _22321_ (.A(_11941_),
    .B1(_11719_),
    .B2(_11815_),
    .ZN(_12631_));
 AOI21_X1 _22322_ (.A(_11941_),
    .B1(_11723_),
    .B2(_11929_),
    .ZN(_12632_));
 NAND2_X1 _22323_ (.A1(_11744_),
    .A2(_11645_),
    .ZN(_12633_));
 NAND3_X1 _22324_ (.A1(_11887_),
    .A2(_11712_),
    .A3(_11841_),
    .ZN(_12634_));
 OAI211_X2 _22325_ (.A(_12633_),
    .B(_12634_),
    .C1(_12629_),
    .C2(_11862_),
    .ZN(_12635_));
 NOR4_X1 _22326_ (.A1(_12630_),
    .A2(_12631_),
    .A3(_12632_),
    .A4(_12635_),
    .ZN(_12636_));
 NOR2_X1 _22327_ (.A1(_11775_),
    .A2(_11724_),
    .ZN(_12637_));
 NOR2_X4 _22328_ (.A1(_11722_),
    .A2(_11936_),
    .ZN(_12638_));
 AOI21_X1 _22329_ (.A(_11789_),
    .B1(_12637_),
    .B2(_12638_),
    .ZN(_12639_));
 NAND2_X1 _22330_ (.A1(_11791_),
    .A2(_11655_),
    .ZN(_12640_));
 OAI211_X2 _22331_ (.A(_11917_),
    .B(_12640_),
    .C1(_11789_),
    .C2(_11926_),
    .ZN(_12641_));
 INV_X1 _22332_ (.A(_12202_),
    .ZN(_12642_));
 AOI21_X1 _22333_ (.A(_11814_),
    .B1(_12642_),
    .B2(_12187_),
    .ZN(_12643_));
 INV_X1 _22334_ (.A(_11818_),
    .ZN(_12644_));
 AOI21_X1 _22335_ (.A(_11814_),
    .B1(_11686_),
    .B2(_12644_),
    .ZN(_12645_));
 NOR4_X1 _22336_ (.A1(_12639_),
    .A2(_12641_),
    .A3(_12643_),
    .A4(_12645_),
    .ZN(_12646_));
 OAI21_X1 _22337_ (.A(_11780_),
    .B1(_11655_),
    .B2(_11659_),
    .ZN(_12647_));
 OAI21_X1 _22338_ (.A(_11780_),
    .B1(_11887_),
    .B2(_11749_),
    .ZN(_12648_));
 OAI21_X1 _22339_ (.A(_11803_),
    .B1(_11655_),
    .B2(_11792_),
    .ZN(_12649_));
 OAI21_X1 _22340_ (.A(_11803_),
    .B1(_11887_),
    .B2(_11695_),
    .ZN(_12650_));
 AND4_X1 _22341_ (.A1(_12647_),
    .A2(_12648_),
    .A3(_12649_),
    .A4(_12650_),
    .ZN(_12651_));
 AOI21_X1 _22342_ (.A(_11839_),
    .B1(_12605_),
    .B2(_11850_),
    .ZN(_12652_));
 NOR2_X1 _22343_ (.A1(_11716_),
    .A2(_11685_),
    .ZN(_12653_));
 AOI21_X1 _22344_ (.A(_11714_),
    .B1(_12652_),
    .B2(_12653_),
    .ZN(_12654_));
 OAI21_X1 _22345_ (.A(_11732_),
    .B1(_11805_),
    .B2(_11839_),
    .ZN(_12655_));
 OAI21_X1 _22346_ (.A(_12655_),
    .B1(_11888_),
    .B2(_11739_),
    .ZN(_12656_));
 AND2_X1 _22347_ (.A1(_11794_),
    .A2(_11732_),
    .ZN(_12657_));
 AND3_X1 _22348_ (.A1(_11753_),
    .A2(_11638_),
    .A3(_11732_),
    .ZN(_12658_));
 NOR4_X1 _22349_ (.A1(_12654_),
    .A2(_12656_),
    .A3(_12657_),
    .A4(_12658_),
    .ZN(_12659_));
 NAND4_X1 _22350_ (.A1(_12636_),
    .A2(_12646_),
    .A3(_12651_),
    .A4(_12659_),
    .ZN(_12660_));
 NOR2_X2 _22351_ (.A1(_12626_),
    .A2(_12660_),
    .ZN(_12661_));
 AND2_X1 _22352_ (.A1(_11238_),
    .A2(_12274_),
    .ZN(_12662_));
 AND2_X1 _22353_ (.A1(_12308_),
    .A2(_11257_),
    .ZN(_12663_));
 OAI21_X1 _22354_ (.A(_11157_),
    .B1(_12662_),
    .B2(_12663_),
    .ZN(_12664_));
 AND2_X1 _22355_ (.A1(_11157_),
    .A2(_12350_),
    .ZN(_12665_));
 INV_X1 _22356_ (.A(_12665_),
    .ZN(_12666_));
 OAI211_X2 _22357_ (.A(_12664_),
    .B(_12666_),
    .C1(_12295_),
    .C2(_12268_),
    .ZN(_12667_));
 NAND2_X1 _22358_ (.A1(_11199_),
    .A2(_11201_),
    .ZN(_12668_));
 NAND2_X1 _22359_ (.A1(_12668_),
    .A2(_11175_),
    .ZN(_12669_));
 AND2_X1 _22360_ (.A1(_11377_),
    .A2(_11171_),
    .ZN(_12670_));
 NOR4_X1 _22361_ (.A1(_12667_),
    .A2(_12669_),
    .A3(_11197_),
    .A4(_12670_),
    .ZN(_12671_));
 AOI21_X1 _22362_ (.A(_11276_),
    .B1(_11215_),
    .B2(_11361_),
    .ZN(_12672_));
 NAND4_X1 _22363_ (.A1(_11332_),
    .A2(_11297_),
    .A3(_12259_),
    .A4(_12260_),
    .ZN(_12673_));
 NAND4_X1 _22364_ (.A1(_11332_),
    .A2(_11172_),
    .A3(_11258_),
    .A4(_11297_),
    .ZN(_12674_));
 OAI211_X2 _22365_ (.A(_12673_),
    .B(_12674_),
    .C1(_11276_),
    .C2(_12316_),
    .ZN(_12675_));
 OAI21_X1 _22366_ (.A(_11293_),
    .B1(_11270_),
    .B2(_11364_),
    .ZN(_12676_));
 NAND4_X1 _22367_ (.A1(_11298_),
    .A2(_11297_),
    .A3(_11322_),
    .A4(_11178_),
    .ZN(_12677_));
 NAND4_X1 _22368_ (.A1(_11293_),
    .A2(_11257_),
    .A3(_11260_),
    .A4(_11165_),
    .ZN(_12678_));
 NAND3_X1 _22369_ (.A1(_12676_),
    .A2(_12677_),
    .A3(_12678_),
    .ZN(_12679_));
 AND2_X2 _22370_ (.A1(_11275_),
    .A2(_11218_),
    .ZN(_12680_));
 NOR4_X1 _22371_ (.A1(_12672_),
    .A2(_12675_),
    .A3(_12679_),
    .A4(_12680_),
    .ZN(_12681_));
 OAI21_X1 _22372_ (.A(_11223_),
    .B1(_11245_),
    .B2(_11345_),
    .ZN(_12682_));
 BUF_X2 _22373_ (.A(_11204_),
    .Z(_12683_));
 OAI21_X1 _22374_ (.A(_12683_),
    .B1(_11245_),
    .B2(_11174_),
    .ZN(_12684_));
 OAI21_X1 _22375_ (.A(_11223_),
    .B1(_12262_),
    .B2(_11316_),
    .ZN(_12685_));
 OAI21_X1 _22376_ (.A(_12683_),
    .B1(_12262_),
    .B2(_11364_),
    .ZN(_12686_));
 AND4_X1 _22377_ (.A1(_12682_),
    .A2(_12684_),
    .A3(_12685_),
    .A4(_12686_),
    .ZN(_12687_));
 AOI22_X1 _22378_ (.A1(_11348_),
    .A2(_11258_),
    .B1(_12260_),
    .B2(_12259_),
    .ZN(_12688_));
 NOR2_X1 _22379_ (.A1(_12688_),
    .A2(_11243_),
    .ZN(_12689_));
 INV_X1 _22380_ (.A(_12689_),
    .ZN(_12690_));
 NAND2_X1 _22381_ (.A1(_11295_),
    .A2(_11253_),
    .ZN(_12691_));
 INV_X1 _22382_ (.A(_12691_),
    .ZN(_12692_));
 AOI22_X1 _22383_ (.A1(_12692_),
    .A2(_11257_),
    .B1(_11253_),
    .B2(_11214_),
    .ZN(_12693_));
 OAI21_X1 _22384_ (.A(_11265_),
    .B1(_12282_),
    .B2(_11174_),
    .ZN(_12694_));
 NAND2_X1 _22385_ (.A1(_11265_),
    .A2(_11378_),
    .ZN(_12695_));
 NAND3_X1 _22386_ (.A1(_11230_),
    .A2(_11297_),
    .A3(_11326_),
    .ZN(_12696_));
 AND3_X1 _22387_ (.A1(_11272_),
    .A2(_12695_),
    .A3(_12696_),
    .ZN(_12697_));
 AND4_X1 _22388_ (.A1(_12690_),
    .A2(_12693_),
    .A3(_12694_),
    .A4(_12697_),
    .ZN(_12698_));
 NAND4_X1 _22389_ (.A1(_12671_),
    .A2(_12681_),
    .A3(_12687_),
    .A4(_12698_),
    .ZN(_12699_));
 AND2_X1 _22390_ (.A1(_11214_),
    .A2(_11342_),
    .ZN(_12700_));
 AND2_X1 _22391_ (.A1(_12349_),
    .A2(_11342_),
    .ZN(_12701_));
 AOI211_X4 _22392_ (.A(_12700_),
    .B(_12701_),
    .C1(_11267_),
    .C2(_11343_),
    .ZN(_12702_));
 AND2_X1 _22393_ (.A1(_11343_),
    .A2(_11316_),
    .ZN(_12703_));
 AND2_X2 _22394_ (.A1(_11286_),
    .A2(_11256_),
    .ZN(_12704_));
 AOI211_X2 _22395_ (.A(_12257_),
    .B(_12703_),
    .C1(_11343_),
    .C2(_12704_),
    .ZN(_12705_));
 OAI21_X1 _22396_ (.A(_11371_),
    .B1(_11267_),
    .B2(_11165_),
    .ZN(_12706_));
 OAI211_X2 _22397_ (.A(_11371_),
    .B(_11232_),
    .C1(_11213_),
    .C2(_11233_),
    .ZN(_12707_));
 NAND2_X4 _22398_ (.A1(_11196_),
    .A2(_11368_),
    .ZN(_12708_));
 NAND2_X1 _22399_ (.A1(_12707_),
    .A2(_12708_),
    .ZN(_12709_));
 INV_X1 _22400_ (.A(_12709_),
    .ZN(_12710_));
 AND4_X4 _22401_ (.A1(_12702_),
    .A2(_12705_),
    .A3(_12706_),
    .A4(_12710_),
    .ZN(_12711_));
 OAI21_X1 _22402_ (.A(_11375_),
    .B1(_11379_),
    .B2(_11364_),
    .ZN(_12712_));
 OAI21_X1 _22403_ (.A(_11363_),
    .B1(_12704_),
    .B2(_12276_),
    .ZN(_12713_));
 OAI21_X1 _22404_ (.A(_11375_),
    .B1(_11358_),
    .B2(_12343_),
    .ZN(_12714_));
 NAND3_X1 _22405_ (.A1(_11214_),
    .A2(_11332_),
    .A3(_11341_),
    .ZN(_12715_));
 AND4_X1 _22406_ (.A1(_12712_),
    .A2(_12713_),
    .A3(_12714_),
    .A4(_12715_),
    .ZN(_12716_));
 NAND2_X1 _22407_ (.A1(_11327_),
    .A2(_11267_),
    .ZN(_12717_));
 NAND2_X1 _22408_ (.A1(_11328_),
    .A2(_11230_),
    .ZN(_12718_));
 NAND3_X1 _22409_ (.A1(_11184_),
    .A2(_11320_),
    .A3(_11326_),
    .ZN(_12719_));
 NAND4_X1 _22410_ (.A1(_12717_),
    .A2(_12345_),
    .A3(_12718_),
    .A4(_12719_),
    .ZN(_12720_));
 AOI21_X1 _22411_ (.A(_12341_),
    .B1(_11356_),
    .B2(_11180_),
    .ZN(_12721_));
 NAND2_X1 _22412_ (.A1(_11315_),
    .A2(_11378_),
    .ZN(_12722_));
 NAND2_X1 _22413_ (.A1(_11315_),
    .A2(_11379_),
    .ZN(_12723_));
 NAND3_X1 _22414_ (.A1(_11230_),
    .A2(_11320_),
    .A3(_11234_),
    .ZN(_12724_));
 NAND3_X1 _22415_ (.A1(_12722_),
    .A2(_12723_),
    .A3(_12724_),
    .ZN(_12725_));
 AND3_X1 _22416_ (.A1(_11320_),
    .A2(_11165_),
    .A3(_11234_),
    .ZN(_12726_));
 NOR4_X1 _22417_ (.A1(_12720_),
    .A2(_12721_),
    .A3(_12725_),
    .A4(_12726_),
    .ZN(_12727_));
 OAI21_X1 _22418_ (.A(_11309_),
    .B1(_12282_),
    .B2(_12343_),
    .ZN(_12728_));
 OAI21_X1 _22419_ (.A(_11309_),
    .B1(_11378_),
    .B2(_12262_),
    .ZN(_12729_));
 NAND4_X1 _22420_ (.A1(_11319_),
    .A2(_11258_),
    .A3(_11298_),
    .A4(_11321_),
    .ZN(_12730_));
 AND4_X1 _22421_ (.A1(_11311_),
    .A2(_12728_),
    .A3(_12729_),
    .A4(_12730_),
    .ZN(_12731_));
 NAND4_X1 _22422_ (.A1(_11332_),
    .A2(_11320_),
    .A3(_11165_),
    .A4(_11213_),
    .ZN(_12732_));
 OAI21_X1 _22423_ (.A(_11336_),
    .B1(_12663_),
    .B2(_12262_),
    .ZN(_12733_));
 AND4_X1 _22424_ (.A1(_12353_),
    .A2(_12731_),
    .A3(_12732_),
    .A4(_12733_),
    .ZN(_12734_));
 NAND4_X1 _22425_ (.A1(_12711_),
    .A2(_12716_),
    .A3(_12727_),
    .A4(_12734_),
    .ZN(_12735_));
 NOR2_X2 _22426_ (.A1(_12699_),
    .A2(_12735_),
    .ZN(_12736_));
 XNOR2_X1 _22427_ (.A(_12661_),
    .B(_12736_),
    .ZN(_12737_));
 AND2_X1 _22428_ (.A1(_11452_),
    .A2(_11544_),
    .ZN(_12738_));
 OAI22_X1 _22429_ (.A1(_11400_),
    .A2(_11426_),
    .B1(_11469_),
    .B2(_11601_),
    .ZN(_12739_));
 AND2_X1 _22430_ (.A1(_12739_),
    .A2(_12444_),
    .ZN(_12740_));
 BUF_X8 _22431_ (.A(_12441_),
    .Z(_12741_));
 NAND2_X1 _22432_ (.A1(_12741_),
    .A2(_11574_),
    .ZN(_12742_));
 NAND4_X1 _22433_ (.A1(_11566_),
    .A2(_12742_),
    .A3(_12462_),
    .A4(_12382_),
    .ZN(_12743_));
 OR3_X1 _22434_ (.A1(_12738_),
    .A2(_12740_),
    .A3(_12743_),
    .ZN(_12744_));
 AND3_X1 _22435_ (.A1(_12463_),
    .A2(_11407_),
    .A3(_11403_),
    .ZN(_12745_));
 INV_X2 _22436_ (.A(_11574_),
    .ZN(_12746_));
 OAI21_X1 _22437_ (.A(_12369_),
    .B1(_12746_),
    .B2(_11541_),
    .ZN(_12747_));
 AOI22_X1 _22438_ (.A1(_11485_),
    .A2(_12445_),
    .B1(_12372_),
    .B2(_12387_),
    .ZN(_12748_));
 NOR4_X2 _22439_ (.A1(_12744_),
    .A2(_12745_),
    .A3(_12747_),
    .A4(_12748_),
    .ZN(_12749_));
 NAND2_X1 _22440_ (.A1(_11597_),
    .A2(_11396_),
    .ZN(_12750_));
 OAI21_X1 _22441_ (.A(_12750_),
    .B1(_11598_),
    .B2(_11541_),
    .ZN(_12751_));
 AND2_X1 _22442_ (.A1(_11587_),
    .A2(_11511_),
    .ZN(_12752_));
 NOR3_X1 _22443_ (.A1(_12751_),
    .A2(_12433_),
    .A3(_12752_),
    .ZN(_12753_));
 AND2_X1 _22444_ (.A1(_11480_),
    .A2(_12430_),
    .ZN(_12754_));
 INV_X1 _22445_ (.A(_12754_),
    .ZN(_12755_));
 AND2_X1 _22446_ (.A1(_11616_),
    .A2(_12371_),
    .ZN(_12756_));
 INV_X1 _22447_ (.A(_12756_),
    .ZN(_12757_));
 AND2_X1 _22448_ (.A1(_11606_),
    .A2(_12409_),
    .ZN(_12758_));
 INV_X1 _22449_ (.A(_12758_),
    .ZN(_12759_));
 NAND2_X1 _22450_ (.A1(_11459_),
    .A2(_11567_),
    .ZN(_12760_));
 AND4_X1 _22451_ (.A1(_12755_),
    .A2(_12757_),
    .A3(_12759_),
    .A4(_12760_),
    .ZN(_12761_));
 NAND2_X1 _22452_ (.A1(_11546_),
    .A2(_11500_),
    .ZN(_12762_));
 NAND2_X1 _22453_ (.A1(_11528_),
    .A2(_11396_),
    .ZN(_12763_));
 NAND2_X1 _22454_ (.A1(_11539_),
    .A2(_11548_),
    .ZN(_12764_));
 AND4_X1 _22455_ (.A1(_12762_),
    .A2(_11579_),
    .A3(_12763_),
    .A4(_12764_),
    .ZN(_12765_));
 AND2_X1 _22456_ (.A1(_11570_),
    .A2(_11392_),
    .ZN(_12766_));
 AND3_X1 _22457_ (.A1(_11454_),
    .A2(_11409_),
    .A3(_11405_),
    .ZN(_12767_));
 AND2_X1 _22458_ (.A1(_12417_),
    .A2(_11505_),
    .ZN(_12768_));
 AND2_X2 _22459_ (.A1(_11446_),
    .A2(_11556_),
    .ZN(_12769_));
 NOR4_X1 _22460_ (.A1(_12766_),
    .A2(_12767_),
    .A3(_12768_),
    .A4(_12769_),
    .ZN(_12770_));
 AND4_X1 _22461_ (.A1(_12753_),
    .A2(_12761_),
    .A3(_12765_),
    .A4(_12770_),
    .ZN(_12771_));
 AND2_X1 _22462_ (.A1(_11546_),
    .A2(_12741_),
    .ZN(_12772_));
 NOR2_X1 _22463_ (.A1(_11540_),
    .A2(_12772_),
    .ZN(_12773_));
 OAI21_X1 _22464_ (.A(_11555_),
    .B1(_11459_),
    .B2(_11519_),
    .ZN(_12774_));
 OAI21_X1 _22465_ (.A(_11555_),
    .B1(_12371_),
    .B2(_12367_),
    .ZN(_12775_));
 AND2_X1 _22466_ (.A1(_12774_),
    .A2(_12775_),
    .ZN(_12776_));
 AND2_X1 _22467_ (.A1(_12741_),
    .A2(_11527_),
    .ZN(_12777_));
 AND4_X1 _22468_ (.A1(_11426_),
    .A2(_11420_),
    .A3(_11552_),
    .A4(_11478_),
    .ZN(_12778_));
 NOR2_X1 _22469_ (.A1(_12777_),
    .A2(_12778_),
    .ZN(_12779_));
 OAI21_X1 _22470_ (.A(_11505_),
    .B1(_11490_),
    .B2(_11496_),
    .ZN(_12780_));
 AND4_X1 _22471_ (.A1(_12773_),
    .A2(_12776_),
    .A3(_12779_),
    .A4(_12780_),
    .ZN(_12781_));
 AND2_X1 _22472_ (.A1(_11606_),
    .A2(_11543_),
    .ZN(_12782_));
 AND3_X1 _22473_ (.A1(_11516_),
    .A2(_11413_),
    .A3(_11493_),
    .ZN(_12783_));
 AND2_X1 _22474_ (.A1(_11441_),
    .A2(_11447_),
    .ZN(_12784_));
 AND2_X1 _22475_ (.A1(_11499_),
    .A2(_11515_),
    .ZN(_12785_));
 OR4_X1 _22476_ (.A1(_12782_),
    .A2(_12783_),
    .A3(_12784_),
    .A4(_12785_),
    .ZN(_12786_));
 NOR2_X1 _22477_ (.A1(_11469_),
    .A2(_11600_),
    .ZN(_12787_));
 AND2_X1 _22478_ (.A1(_11606_),
    .A2(_12787_),
    .ZN(_12788_));
 INV_X1 _22479_ (.A(_12788_),
    .ZN(_12789_));
 AOI22_X1 _22480_ (.A1(_11570_),
    .A2(_12463_),
    .B1(_11465_),
    .B2(_11482_),
    .ZN(_12790_));
 OAI211_X2 _22481_ (.A(_12789_),
    .B(_12790_),
    .C1(_11525_),
    .C2(_11610_),
    .ZN(_12791_));
 NAND3_X1 _22482_ (.A1(_11527_),
    .A2(_11411_),
    .A3(_11601_),
    .ZN(_12792_));
 NAND3_X1 _22483_ (.A1(_11527_),
    .A2(_11413_),
    .A3(_11411_),
    .ZN(_12793_));
 AND2_X1 _22484_ (.A1(_12792_),
    .A2(_12793_),
    .ZN(_12794_));
 AND2_X1 _22485_ (.A1(_11542_),
    .A2(_11446_),
    .ZN(_12795_));
 INV_X1 _22486_ (.A(_12795_),
    .ZN(_12796_));
 NAND2_X1 _22487_ (.A1(_12444_),
    .A2(_11436_),
    .ZN(_12797_));
 NAND2_X1 _22488_ (.A1(_12392_),
    .A2(_12787_),
    .ZN(_12798_));
 NAND4_X1 _22489_ (.A1(_12794_),
    .A2(_12796_),
    .A3(_12797_),
    .A4(_12798_),
    .ZN(_12799_));
 NAND2_X1 _22490_ (.A1(_11546_),
    .A2(_11459_),
    .ZN(_12800_));
 NAND2_X1 _22491_ (.A1(_11507_),
    .A2(_11527_),
    .ZN(_12801_));
 NAND3_X1 _22492_ (.A1(_11496_),
    .A2(_11537_),
    .A3(_11445_),
    .ZN(_12802_));
 NAND4_X1 _22493_ (.A1(_12800_),
    .A2(_11580_),
    .A3(_12801_),
    .A4(_12802_),
    .ZN(_12803_));
 NOR4_X1 _22494_ (.A1(_12786_),
    .A2(_12791_),
    .A3(_12799_),
    .A4(_12803_),
    .ZN(_12804_));
 NAND4_X1 _22495_ (.A1(_12749_),
    .A2(_12771_),
    .A3(_12781_),
    .A4(_12804_),
    .ZN(_12805_));
 AOI21_X1 _22496_ (.A(_11466_),
    .B1(_12372_),
    .B2(_11541_),
    .ZN(_12806_));
 AOI221_X4 _22497_ (.A(_12806_),
    .B1(_11412_),
    .B2(_11607_),
    .C1(_11434_),
    .C2(_12392_),
    .ZN(_12807_));
 OAI21_X1 _22498_ (.A(_11442_),
    .B1(_11436_),
    .B2(_11496_),
    .ZN(_12808_));
 NAND4_X1 _22499_ (.A1(_11591_),
    .A2(_11599_),
    .A3(_11388_),
    .A4(_11467_),
    .ZN(_12809_));
 NAND4_X1 _22500_ (.A1(_11442_),
    .A2(_11412_),
    .A3(_11407_),
    .A4(_11426_),
    .ZN(_12810_));
 AND3_X1 _22501_ (.A1(_12808_),
    .A2(_12809_),
    .A3(_12810_),
    .ZN(_12811_));
 AND2_X2 _22502_ (.A1(_11472_),
    .A2(_11406_),
    .ZN(_12812_));
 AOI22_X1 _22503_ (.A1(_12812_),
    .A2(_11516_),
    .B1(_11474_),
    .B2(_12444_),
    .ZN(_12813_));
 NAND2_X1 _22504_ (.A1(_12430_),
    .A2(_11391_),
    .ZN(_12814_));
 AND2_X1 _22505_ (.A1(_12814_),
    .A2(_12403_),
    .ZN(_12815_));
 OAI21_X1 _22506_ (.A(_12456_),
    .B1(_11450_),
    .B2(_11556_),
    .ZN(_12816_));
 AND3_X1 _22507_ (.A1(_12813_),
    .A2(_12815_),
    .A3(_12816_),
    .ZN(_12817_));
 AND2_X1 _22508_ (.A1(_11479_),
    .A2(_11570_),
    .ZN(_12818_));
 AND2_X1 _22509_ (.A1(_11465_),
    .A2(_11570_),
    .ZN(_12819_));
 NOR2_X1 _22510_ (.A1(_12400_),
    .A2(_11602_),
    .ZN(_12820_));
 NOR3_X1 _22511_ (.A1(_12818_),
    .A2(_12819_),
    .A3(_12820_),
    .ZN(_12821_));
 NAND4_X1 _22512_ (.A1(_12807_),
    .A2(_12811_),
    .A3(_12817_),
    .A4(_12821_),
    .ZN(_12822_));
 NOR2_X4 _22513_ (.A1(_12805_),
    .A2(_12822_),
    .ZN(_12823_));
 XNOR2_X1 _22514_ (.A(_12737_),
    .B(_12823_),
    .ZN(_12824_));
 AND2_X1 _22515_ (.A1(_12114_),
    .A2(_12082_),
    .ZN(_12825_));
 INV_X1 _22516_ (.A(_12825_),
    .ZN(_12826_));
 NAND2_X1 _22517_ (.A1(_12005_),
    .A2(_12037_),
    .ZN(_12827_));
 AOI22_X1 _22518_ (.A1(_11995_),
    .A2(_12100_),
    .B1(_12165_),
    .B2(_12048_),
    .ZN(_12828_));
 AND4_X1 _22519_ (.A1(_12524_),
    .A2(_12826_),
    .A3(_12827_),
    .A4(_12828_),
    .ZN(_12829_));
 CLKBUF_X2 _22520_ (.A(_12125_),
    .Z(_12830_));
 AOI22_X1 _22521_ (.A1(_12163_),
    .A2(_12830_),
    .B1(_12119_),
    .B2(_12162_),
    .ZN(_12831_));
 AOI221_X4 _22522_ (.A(_11974_),
    .B1(_12036_),
    .B2(_12044_),
    .C1(_12552_),
    .C2(_12161_),
    .ZN(_12832_));
 AND4_X1 _22523_ (.A1(_12514_),
    .A2(_12829_),
    .A3(_12831_),
    .A4(_12832_),
    .ZN(_12833_));
 BUF_X4 _22524_ (.A(_12002_),
    .Z(_12834_));
 NAND2_X1 _22525_ (.A1(_12079_),
    .A2(_12834_),
    .ZN(_12835_));
 NAND2_X1 _22526_ (.A1(_12085_),
    .A2(_12152_),
    .ZN(_12836_));
 INV_X1 _22527_ (.A(_12085_),
    .ZN(_12837_));
 OAI211_X2 _22528_ (.A(_12835_),
    .B(_12836_),
    .C1(_12837_),
    .C2(_12059_),
    .ZN(_12838_));
 INV_X2 _22529_ (.A(_12161_),
    .ZN(_12839_));
 INV_X1 _22530_ (.A(_12082_),
    .ZN(_12840_));
 AOI21_X1 _22531_ (.A(_12839_),
    .B1(_12477_),
    .B2(_12840_),
    .ZN(_12841_));
 AND2_X1 _22532_ (.A1(_12142_),
    .A2(_12100_),
    .ZN(_12842_));
 OR3_X2 _22533_ (.A1(_12838_),
    .A2(_12841_),
    .A3(_12842_),
    .ZN(_12843_));
 OAI21_X1 _22534_ (.A(_12028_),
    .B1(_12566_),
    .B2(_12069_),
    .ZN(_12844_));
 NAND3_X1 _22535_ (.A1(_12479_),
    .A2(_12026_),
    .A3(_12113_),
    .ZN(_12845_));
 NAND4_X1 _22536_ (.A1(_12116_),
    .A2(_12104_),
    .A3(_12137_),
    .A4(_12845_),
    .ZN(_12846_));
 NAND3_X1 _22537_ (.A1(_12108_),
    .A2(_12089_),
    .A3(_11973_),
    .ZN(_12847_));
 NAND2_X1 _22538_ (.A1(_12068_),
    .A2(_11963_),
    .ZN(_12848_));
 INV_X1 _22539_ (.A(_12005_),
    .ZN(_12849_));
 INV_X2 _22540_ (.A(_11963_),
    .ZN(_12850_));
 OAI211_X2 _22541_ (.A(_12847_),
    .B(_12848_),
    .C1(_12849_),
    .C2(_12850_),
    .ZN(_12851_));
 NOR4_X1 _22542_ (.A1(_12843_),
    .A2(_12844_),
    .A3(_12846_),
    .A4(_12851_),
    .ZN(_12852_));
 INV_X4 _22543_ (.A(_12165_),
    .ZN(_12853_));
 NOR2_X1 _22544_ (.A1(_12853_),
    .A2(_12506_),
    .ZN(_12854_));
 NOR2_X1 _22545_ (.A1(_12839_),
    .A2(_12489_),
    .ZN(_12855_));
 AND3_X1 _22546_ (.A1(_12125_),
    .A2(_12491_),
    .A3(_11967_),
    .ZN(_12856_));
 AND2_X2 _22547_ (.A1(_12125_),
    .A2(_11999_),
    .ZN(_12857_));
 NOR4_X1 _22548_ (.A1(_12854_),
    .A2(_12855_),
    .A3(_12856_),
    .A4(_12857_),
    .ZN(_12858_));
 NAND2_X1 _22549_ (.A1(_12543_),
    .A2(_12544_),
    .ZN(_12859_));
 BUF_X4 _22550_ (.A(_12012_),
    .Z(_12860_));
 BUF_X4 _22551_ (.A(_12100_),
    .Z(_12861_));
 AOI22_X1 _22552_ (.A1(_12860_),
    .A2(_12861_),
    .B1(_12834_),
    .B2(_12037_),
    .ZN(_12862_));
 BUF_X4 _22553_ (.A(_11993_),
    .Z(_12863_));
 NAND3_X1 _22554_ (.A1(_11997_),
    .A2(_12863_),
    .A3(_12496_),
    .ZN(_12864_));
 NAND2_X1 _22555_ (.A1(_12834_),
    .A2(_12860_),
    .ZN(_12865_));
 AND4_X1 _22556_ (.A1(_12859_),
    .A2(_12862_),
    .A3(_12864_),
    .A4(_12865_),
    .ZN(_12866_));
 AND4_X1 _22557_ (.A1(_12833_),
    .A2(_12852_),
    .A3(_12858_),
    .A4(_12866_),
    .ZN(_12867_));
 NAND3_X1 _22558_ (.A1(_12019_),
    .A2(_12863_),
    .A3(_11985_),
    .ZN(_12868_));
 AND4_X1 _22559_ (.A1(_11989_),
    .A2(_12054_),
    .A3(_12031_),
    .A4(_11962_),
    .ZN(_12869_));
 NOR2_X1 _22560_ (.A1(_12474_),
    .A2(_12869_),
    .ZN(_12870_));
 NAND4_X1 _22561_ (.A1(_12863_),
    .A2(_11969_),
    .A3(_11985_),
    .A4(_11990_),
    .ZN(_12871_));
 NAND3_X1 _22562_ (.A1(_12009_),
    .A2(_12863_),
    .A3(_11985_),
    .ZN(_12872_));
 AND4_X1 _22563_ (.A1(_12868_),
    .A2(_12870_),
    .A3(_12871_),
    .A4(_12872_),
    .ZN(_12873_));
 AND2_X1 _22564_ (.A1(_12062_),
    .A2(_12075_),
    .ZN(_12874_));
 AOI221_X4 _22565_ (.A(_12874_),
    .B1(_12484_),
    .B2(_12085_),
    .C1(_12037_),
    .C2(_12493_),
    .ZN(_12875_));
 AND2_X1 _22566_ (.A1(_11967_),
    .A2(_11980_),
    .ZN(_12876_));
 INV_X1 _22567_ (.A(_12876_),
    .ZN(_12877_));
 OAI22_X1 _22568_ (.A1(_12063_),
    .A2(_12045_),
    .B1(_12138_),
    .B2(_12877_),
    .ZN(_12878_));
 AND2_X1 _22569_ (.A1(_12142_),
    .A2(_12075_),
    .ZN(_12879_));
 AND3_X1 _22570_ (.A1(_12012_),
    .A2(_12000_),
    .A3(_12030_),
    .ZN(_12880_));
 AND3_X1 _22571_ (.A1(_12479_),
    .A2(_12035_),
    .A3(_12496_),
    .ZN(_12881_));
 NOR4_X1 _22572_ (.A1(_12878_),
    .A2(_12879_),
    .A3(_12880_),
    .A4(_12881_),
    .ZN(_12882_));
 INV_X1 _22573_ (.A(_12582_),
    .ZN(_12883_));
 NAND4_X1 _22574_ (.A1(_12873_),
    .A2(_12875_),
    .A3(_12882_),
    .A4(_12883_),
    .ZN(_12884_));
 AND2_X1 _22575_ (.A1(_12150_),
    .A2(_12090_),
    .ZN(_12885_));
 AOI21_X1 _22576_ (.A(_12151_),
    .B1(_12504_),
    .B2(_12072_),
    .ZN(_12886_));
 NOR2_X1 _22577_ (.A1(_12109_),
    .A2(_12050_),
    .ZN(_12887_));
 AOI21_X1 _22578_ (.A(_12143_),
    .B1(_12887_),
    .B2(_12069_),
    .ZN(_12888_));
 NOR2_X1 _22579_ (.A1(_12151_),
    .A2(_12506_),
    .ZN(_12889_));
 OR4_X4 _22580_ (.A1(_12885_),
    .A2(_12886_),
    .A3(_12888_),
    .A4(_12889_),
    .ZN(_12890_));
 AND2_X1 _22581_ (.A1(_12490_),
    .A2(_12108_),
    .ZN(_12891_));
 INV_X1 _22582_ (.A(_12891_),
    .ZN(_12892_));
 OAI21_X1 _22583_ (.A(_12056_),
    .B1(_12066_),
    .B2(_12025_),
    .ZN(_12893_));
 OAI21_X1 _22584_ (.A(_12544_),
    .B1(_12066_),
    .B2(_12128_),
    .ZN(_12894_));
 OAI21_X1 _22585_ (.A(_12527_),
    .B1(_12163_),
    .B2(_12876_),
    .ZN(_12895_));
 NAND4_X1 _22586_ (.A1(_12892_),
    .A2(_12893_),
    .A3(_12894_),
    .A4(_12895_),
    .ZN(_12896_));
 OAI21_X1 _22587_ (.A(_11964_),
    .B1(_12052_),
    .B2(_12552_),
    .ZN(_12897_));
 AND2_X1 _22588_ (.A1(_12062_),
    .A2(_11999_),
    .ZN(_12898_));
 INV_X1 _22589_ (.A(_12898_),
    .ZN(_12899_));
 NAND2_X1 _22590_ (.A1(_12088_),
    .A2(_12541_),
    .ZN(_12900_));
 OAI21_X1 _22591_ (.A(_12487_),
    .B1(_12503_),
    .B2(_12476_),
    .ZN(_12901_));
 NAND4_X1 _22592_ (.A1(_12897_),
    .A2(_12899_),
    .A3(_12900_),
    .A4(_12901_),
    .ZN(_12902_));
 NOR4_X4 _22593_ (.A1(_12884_),
    .A2(_12890_),
    .A3(_12896_),
    .A4(_12902_),
    .ZN(_12903_));
 NAND2_X2 _22594_ (.A1(_12867_),
    .A2(_12903_),
    .ZN(_12904_));
 XOR2_X1 _22595_ (.A(_12256_),
    .B(_12904_),
    .Z(_12905_));
 XNOR2_X1 _22596_ (.A(_12824_),
    .B(_12905_),
    .ZN(_12906_));
 XNOR2_X1 _22597_ (.A(_12906_),
    .B(_17262_),
    .ZN(_12907_));
 MUX2_X1 _22598_ (.A(_12587_),
    .B(_12907_),
    .S(_11149_),
    .Z(_00718_));
 XOR2_X1 _22599_ (.A(_17265_),
    .B(_17068_),
    .Z(_12908_));
 XOR2_X1 _22600_ (.A(_11958_),
    .B(_12661_),
    .Z(_12909_));
 OAI211_X2 _22601_ (.A(_11502_),
    .B(_11411_),
    .C1(_11405_),
    .C2(_11402_),
    .ZN(_12910_));
 OAI211_X2 _22602_ (.A(_11502_),
    .B(_11419_),
    .C1(_11413_),
    .C2(_11414_),
    .ZN(_12911_));
 OAI21_X1 _22603_ (.A(_11502_),
    .B1(_11488_),
    .B2(_11396_),
    .ZN(_12912_));
 AND4_X1 _22604_ (.A1(_11512_),
    .A2(_12910_),
    .A3(_12911_),
    .A4(_12912_),
    .ZN(_12913_));
 AND3_X1 _22605_ (.A1(_11590_),
    .A2(_11464_),
    .A3(_11478_),
    .ZN(_12914_));
 AOI21_X1 _22606_ (.A(_11485_),
    .B1(_11451_),
    .B2(_11541_),
    .ZN(_12915_));
 AOI211_X4 _22607_ (.A(_12914_),
    .B(_12915_),
    .C1(_12367_),
    .C2(_11479_),
    .ZN(_12916_));
 OAI21_X1 _22608_ (.A(_11480_),
    .B1(_11519_),
    .B2(_11500_),
    .ZN(_12917_));
 OAI21_X1 _22609_ (.A(_11480_),
    .B1(_11441_),
    .B2(_11482_),
    .ZN(_12918_));
 AND4_X4 _22610_ (.A1(_12913_),
    .A2(_12916_),
    .A3(_12917_),
    .A4(_12918_),
    .ZN(_12919_));
 AND2_X1 _22611_ (.A1(_11527_),
    .A2(_11560_),
    .ZN(_12920_));
 INV_X1 _22612_ (.A(_12920_),
    .ZN(_12921_));
 NAND2_X1 _22613_ (.A1(_11486_),
    .A2(_11527_),
    .ZN(_12922_));
 AND3_X1 _22614_ (.A1(_12921_),
    .A2(_12922_),
    .A3(_12801_),
    .ZN(_12923_));
 AND3_X1 _22615_ (.A1(_11585_),
    .A2(_12393_),
    .A3(_11515_),
    .ZN(_12924_));
 NAND2_X1 _22616_ (.A1(_11449_),
    .A2(_11515_),
    .ZN(_12925_));
 NAND2_X1 _22617_ (.A1(_12925_),
    .A2(_12383_),
    .ZN(_12926_));
 NOR3_X1 _22618_ (.A1(_12924_),
    .A2(_12926_),
    .A3(_12785_),
    .ZN(_12927_));
 OAI21_X1 _22619_ (.A(_11528_),
    .B1(_11556_),
    .B2(_12367_),
    .ZN(_12928_));
 OAI211_X2 _22620_ (.A(_11528_),
    .B(_11420_),
    .C1(_11467_),
    .C2(_11415_),
    .ZN(_12929_));
 AND4_X1 _22621_ (.A1(_12923_),
    .A2(_12927_),
    .A3(_12928_),
    .A4(_12929_),
    .ZN(_12930_));
 NAND2_X1 _22622_ (.A1(_11575_),
    .A2(_11607_),
    .ZN(_12931_));
 NAND2_X1 _22623_ (.A1(_11607_),
    .A2(_11507_),
    .ZN(_12932_));
 NAND4_X1 _22624_ (.A1(_12759_),
    .A2(_12789_),
    .A3(_12931_),
    .A4(_12932_),
    .ZN(_12933_));
 AND2_X1 _22625_ (.A1(_12812_),
    .A2(_12456_),
    .ZN(_12934_));
 OAI21_X1 _22626_ (.A(_12750_),
    .B1(_11598_),
    .B2(_12361_),
    .ZN(_12935_));
 NOR4_X1 _22627_ (.A1(_12933_),
    .A2(_12458_),
    .A3(_12934_),
    .A4(_12935_),
    .ZN(_12936_));
 NAND4_X1 _22628_ (.A1(_11592_),
    .A2(_11415_),
    .A3(_11599_),
    .A4(_11591_),
    .ZN(_12937_));
 NAND2_X1 _22629_ (.A1(_12463_),
    .A2(_11434_),
    .ZN(_12938_));
 AND2_X1 _22630_ (.A1(_11616_),
    .A2(_11507_),
    .ZN(_12939_));
 AND2_X1 _22631_ (.A1(_11616_),
    .A2(_11548_),
    .ZN(_12940_));
 NOR2_X1 _22632_ (.A1(_12939_),
    .A2(_12940_),
    .ZN(_12941_));
 NAND2_X1 _22633_ (.A1(_11616_),
    .A2(_11396_),
    .ZN(_12942_));
 AND4_X1 _22634_ (.A1(_12938_),
    .A2(_12941_),
    .A3(_12942_),
    .A4(_12757_),
    .ZN(_12943_));
 OAI211_X2 _22635_ (.A(_12444_),
    .B(_11412_),
    .C1(_11413_),
    .C2(_11529_),
    .ZN(_12944_));
 INV_X1 _22636_ (.A(_11600_),
    .ZN(_12945_));
 AND3_X1 _22637_ (.A1(_11494_),
    .A2(_11587_),
    .A3(_12945_),
    .ZN(_12946_));
 AOI211_X4 _22638_ (.A(_12442_),
    .B(_12946_),
    .C1(_12367_),
    .C2(_11587_),
    .ZN(_12947_));
 AND4_X1 _22639_ (.A1(_12937_),
    .A2(_12943_),
    .A3(_12944_),
    .A4(_12947_),
    .ZN(_12948_));
 NAND4_X1 _22640_ (.A1(_12919_),
    .A2(_12930_),
    .A3(_12936_),
    .A4(_12948_),
    .ZN(_12949_));
 NAND2_X1 _22641_ (.A1(_11454_),
    .A2(_11482_),
    .ZN(_12950_));
 AOI21_X1 _22642_ (.A(_12400_),
    .B1(_11455_),
    .B2(_11460_),
    .ZN(_12951_));
 NAND2_X1 _22643_ (.A1(_11589_),
    .A2(_11391_),
    .ZN(_12952_));
 OAI211_X2 _22644_ (.A(_12402_),
    .B(_12952_),
    .C1(_11524_),
    .C2(_12400_),
    .ZN(_12953_));
 AOI211_X2 _22645_ (.A(_12951_),
    .B(_12953_),
    .C1(_12379_),
    .C2(_11391_),
    .ZN(_12954_));
 AND4_X1 _22646_ (.A1(_11394_),
    .A2(_11445_),
    .A3(_11402_),
    .A4(_11388_),
    .ZN(_12955_));
 NOR2_X1 _22647_ (.A1(_11448_),
    .A2(_12955_),
    .ZN(_12956_));
 OAI21_X1 _22648_ (.A(_11454_),
    .B1(_11452_),
    .B2(_11590_),
    .ZN(_12957_));
 AND4_X1 _22649_ (.A1(_12950_),
    .A2(_12954_),
    .A3(_12956_),
    .A4(_12957_),
    .ZN(_12958_));
 NAND2_X1 _22650_ (.A1(_11544_),
    .A2(_11531_),
    .ZN(_12959_));
 NAND4_X1 _22651_ (.A1(_11573_),
    .A2(_11411_),
    .A3(_11406_),
    .A4(_11426_),
    .ZN(_12960_));
 NAND4_X1 _22652_ (.A1(_11537_),
    .A2(_11419_),
    .A3(_11529_),
    .A4(_11591_),
    .ZN(_12961_));
 AND4_X1 _22653_ (.A1(_12742_),
    .A2(_12960_),
    .A3(_11580_),
    .A4(_12961_),
    .ZN(_12962_));
 OAI21_X1 _22654_ (.A(_11544_),
    .B1(_12396_),
    .B2(_11459_),
    .ZN(_12963_));
 OAI21_X1 _22655_ (.A(_11544_),
    .B1(_12741_),
    .B2(_12367_),
    .ZN(_12964_));
 AND4_X1 _22656_ (.A1(_12959_),
    .A2(_12962_),
    .A3(_12963_),
    .A4(_12964_),
    .ZN(_12965_));
 OAI21_X1 _22657_ (.A(_11564_),
    .B1(_11510_),
    .B2(_11433_),
    .ZN(_12966_));
 OAI21_X1 _22658_ (.A(_12966_),
    .B1(_11525_),
    .B2(_12427_),
    .ZN(_12967_));
 AOI21_X1 _22659_ (.A(_12427_),
    .B1(_11487_),
    .B2(_12361_),
    .ZN(_12968_));
 AND2_X1 _22660_ (.A1(_11564_),
    .A2(_12409_),
    .ZN(_12969_));
 NOR4_X1 _22661_ (.A1(_12967_),
    .A2(_12968_),
    .A3(_12432_),
    .A4(_12969_),
    .ZN(_12970_));
 OAI211_X2 _22662_ (.A(_11554_),
    .B(_11599_),
    .C1(_11413_),
    .C2(_11529_),
    .ZN(_12971_));
 AND2_X1 _22663_ (.A1(_11399_),
    .A2(_11456_),
    .ZN(_12972_));
 OAI21_X1 _22664_ (.A(_11554_),
    .B1(_12386_),
    .B2(_12972_),
    .ZN(_12973_));
 AND4_X1 _22665_ (.A1(_12416_),
    .A2(_12970_),
    .A3(_12971_),
    .A4(_12973_),
    .ZN(_12974_));
 INV_X1 _22666_ (.A(_11500_),
    .ZN(_12975_));
 AOI21_X1 _22667_ (.A(_11466_),
    .B1(_12975_),
    .B2(_12361_),
    .ZN(_12976_));
 AND3_X1 _22668_ (.A1(_11585_),
    .A2(_12393_),
    .A3(_11424_),
    .ZN(_12977_));
 AND2_X1 _22669_ (.A1(_11465_),
    .A2(_12741_),
    .ZN(_12978_));
 AND2_X1 _22670_ (.A1(_11590_),
    .A2(_11424_),
    .ZN(_12979_));
 NOR4_X1 _22671_ (.A1(_12976_),
    .A2(_12977_),
    .A3(_12978_),
    .A4(_12979_),
    .ZN(_12980_));
 NAND4_X1 _22672_ (.A1(_12958_),
    .A2(_12965_),
    .A3(_12974_),
    .A4(_12980_),
    .ZN(_12981_));
 NOR2_X2 _22673_ (.A1(_12949_),
    .A2(_12981_),
    .ZN(_12982_));
 INV_X2 _22674_ (.A(_12982_),
    .ZN(_12983_));
 XNOR2_X1 _22675_ (.A(_12909_),
    .B(_12983_),
    .ZN(_12984_));
 AOI21_X1 _22676_ (.A(_12721_),
    .B1(_11226_),
    .B2(_11315_),
    .ZN(_12985_));
 NAND4_X1 _22677_ (.A1(_12308_),
    .A2(_11257_),
    .A3(_11319_),
    .A4(_11234_),
    .ZN(_12986_));
 NAND3_X1 _22678_ (.A1(_12985_),
    .A2(_12723_),
    .A3(_12986_),
    .ZN(_12987_));
 AND2_X1 _22679_ (.A1(_12704_),
    .A2(_11328_),
    .ZN(_12988_));
 AND2_X1 _22680_ (.A1(_11327_),
    .A2(_11188_),
    .ZN(_12989_));
 OAI21_X1 _22681_ (.A(_12717_),
    .B1(_11330_),
    .B2(_12268_),
    .ZN(_12990_));
 NOR4_X1 _22682_ (.A1(_12987_),
    .A2(_12988_),
    .A3(_12989_),
    .A4(_12990_),
    .ZN(_12991_));
 OAI21_X1 _22683_ (.A(_11363_),
    .B1(_11345_),
    .B2(_12350_),
    .ZN(_12992_));
 OAI21_X1 _22684_ (.A(_11363_),
    .B1(_12282_),
    .B2(_12343_),
    .ZN(_12993_));
 OAI21_X1 _22685_ (.A(_11363_),
    .B1(_11378_),
    .B2(_11184_),
    .ZN(_12994_));
 OAI21_X1 _22686_ (.A(_11353_),
    .B1(_11277_),
    .B2(_11316_),
    .ZN(_12995_));
 NAND4_X1 _22687_ (.A1(_12992_),
    .A2(_12993_),
    .A3(_12994_),
    .A4(_12995_),
    .ZN(_12996_));
 NAND2_X1 _22688_ (.A1(_11248_),
    .A2(_11375_),
    .ZN(_12997_));
 OAI211_X2 _22689_ (.A(_12997_),
    .B(_11382_),
    .C1(_11251_),
    .C2(_12285_),
    .ZN(_12998_));
 INV_X1 _22690_ (.A(_11254_),
    .ZN(_12999_));
 AOI21_X1 _22691_ (.A(_12285_),
    .B1(_11357_),
    .B2(_12999_),
    .ZN(_13000_));
 OAI21_X1 _22692_ (.A(_11374_),
    .B1(_12302_),
    .B2(_12285_),
    .ZN(_13001_));
 NOR4_X1 _22693_ (.A1(_12996_),
    .A2(_12998_),
    .A3(_13000_),
    .A4(_13001_),
    .ZN(_13002_));
 OAI21_X1 _22694_ (.A(_11371_),
    .B1(_11230_),
    .B2(_11316_),
    .ZN(_13003_));
 OAI211_X2 _22695_ (.A(_11368_),
    .B(_11232_),
    .C1(_11178_),
    .C2(_11233_),
    .ZN(_13004_));
 OAI21_X1 _22696_ (.A(_11368_),
    .B1(_11174_),
    .B2(_12327_),
    .ZN(_13005_));
 NAND4_X1 _22697_ (.A1(_12265_),
    .A2(_11269_),
    .A3(_11341_),
    .A4(_11234_),
    .ZN(_13006_));
 NAND4_X1 _22698_ (.A1(_13003_),
    .A2(_13004_),
    .A3(_13005_),
    .A4(_13006_),
    .ZN(_13007_));
 INV_X1 _22699_ (.A(_11342_),
    .ZN(_13008_));
 AOI21_X1 _22700_ (.A(_13008_),
    .B1(_11185_),
    .B2(_11280_),
    .ZN(_13009_));
 AND4_X1 _22701_ (.A1(_12274_),
    .A2(_11342_),
    .A3(_12265_),
    .A4(_11348_),
    .ZN(_13010_));
 NOR4_X1 _22702_ (.A1(_13007_),
    .A2(_13009_),
    .A3(_13010_),
    .A4(_12701_),
    .ZN(_13011_));
 NAND4_X1 _22703_ (.A1(_11238_),
    .A2(_11319_),
    .A3(_12274_),
    .A4(_11298_),
    .ZN(_13012_));
 NAND3_X1 _22704_ (.A1(_11196_),
    .A2(_11319_),
    .A3(_11298_),
    .ZN(_13013_));
 OAI211_X2 _22705_ (.A(_13012_),
    .B(_13013_),
    .C1(_11280_),
    .C2(_11312_),
    .ZN(_13014_));
 OAI211_X2 _22706_ (.A(_11153_),
    .B(_11305_),
    .C1(_11207_),
    .C2(_12262_),
    .ZN(_13015_));
 NAND2_X1 _22707_ (.A1(_11336_),
    .A2(_11226_),
    .ZN(_13016_));
 NAND2_X1 _22708_ (.A1(_11336_),
    .A2(_12301_),
    .ZN(_13017_));
 NAND4_X1 _22709_ (.A1(_13015_),
    .A2(_13016_),
    .A3(_13017_),
    .A4(_12352_),
    .ZN(_13018_));
 AOI21_X1 _22710_ (.A(_11312_),
    .B1(_11215_),
    .B2(_11227_),
    .ZN(_13019_));
 AND4_X1 _22711_ (.A1(_11209_),
    .A2(_11305_),
    .A3(_11159_),
    .A4(_11169_),
    .ZN(_13020_));
 NOR4_X1 _22712_ (.A1(_13014_),
    .A2(_13018_),
    .A3(_13019_),
    .A4(_13020_),
    .ZN(_13021_));
 NAND4_X1 _22713_ (.A1(_12991_),
    .A2(_13002_),
    .A3(_13011_),
    .A4(_13021_),
    .ZN(_13022_));
 AND4_X1 _22714_ (.A1(_11172_),
    .A2(_11183_),
    .A3(_11241_),
    .A4(_11221_),
    .ZN(_13023_));
 AOI221_X1 _22715_ (.A(_13023_),
    .B1(_11242_),
    .B2(_11189_),
    .C1(_12322_),
    .C2(_11321_),
    .ZN(_13024_));
 NAND4_X1 _22716_ (.A1(_11297_),
    .A2(_11221_),
    .A3(_11159_),
    .A4(_11209_),
    .ZN(_13025_));
 OAI211_X2 _22717_ (.A(_11242_),
    .B(_12265_),
    .C1(_11244_),
    .C2(_11217_),
    .ZN(_13026_));
 AND3_X1 _22718_ (.A1(_13024_),
    .A2(_13025_),
    .A3(_13026_),
    .ZN(_13027_));
 NAND2_X1 _22719_ (.A1(_11265_),
    .A2(_12343_),
    .ZN(_13028_));
 OAI21_X1 _22720_ (.A(_11264_),
    .B1(_11310_),
    .B2(_11267_),
    .ZN(_13029_));
 OAI21_X1 _22721_ (.A(_11264_),
    .B1(_12662_),
    .B2(_11277_),
    .ZN(_13030_));
 AND4_X2 _22722_ (.A1(_13027_),
    .A2(_13028_),
    .A3(_13029_),
    .A4(_13030_),
    .ZN(_13031_));
 AND2_X1 _22723_ (.A1(_12260_),
    .A2(_16815_),
    .ZN(_13032_));
 OAI21_X1 _22724_ (.A(_11199_),
    .B1(_11196_),
    .B2(_13032_),
    .ZN(_13033_));
 NAND4_X1 _22725_ (.A1(_11171_),
    .A2(_11256_),
    .A3(_11260_),
    .A4(_12265_),
    .ZN(_13034_));
 AND2_X1 _22726_ (.A1(_13034_),
    .A2(_11175_),
    .ZN(_13035_));
 OAI21_X1 _22727_ (.A(_11157_),
    .B1(_11245_),
    .B2(_11295_),
    .ZN(_13036_));
 OAI21_X1 _22728_ (.A(_11157_),
    .B1(_12308_),
    .B2(_11210_),
    .ZN(_13037_));
 AND4_X1 _22729_ (.A1(_13033_),
    .A2(_13035_),
    .A3(_13036_),
    .A4(_13037_),
    .ZN(_13038_));
 AND2_X4 _22730_ (.A1(_11188_),
    .A2(_11321_),
    .ZN(_13039_));
 OAI21_X1 _22731_ (.A(_11223_),
    .B1(_11248_),
    .B2(_13039_),
    .ZN(_13040_));
 OAI21_X1 _22732_ (.A(_11223_),
    .B1(_11310_),
    .B2(_11267_),
    .ZN(_13041_));
 NAND4_X1 _22733_ (.A1(_11164_),
    .A2(_11167_),
    .A3(_11178_),
    .A4(_11234_),
    .ZN(_13042_));
 NAND2_X1 _22734_ (.A1(_12282_),
    .A2(_11223_),
    .ZN(_13043_));
 NAND4_X1 _22735_ (.A1(_13040_),
    .A2(_13041_),
    .A3(_13042_),
    .A4(_13043_),
    .ZN(_13044_));
 NAND2_X1 _22736_ (.A1(_11204_),
    .A2(_11379_),
    .ZN(_13045_));
 OAI211_X2 _22737_ (.A(_12299_),
    .B(_13045_),
    .C1(_11205_),
    .C2(_12275_),
    .ZN(_13046_));
 NAND2_X1 _22738_ (.A1(_12683_),
    .A2(_11201_),
    .ZN(_13047_));
 NAND2_X1 _22739_ (.A1(_12683_),
    .A2(_11174_),
    .ZN(_13048_));
 NAND2_X1 _22740_ (.A1(_13047_),
    .A2(_13048_),
    .ZN(_13049_));
 NOR3_X1 _22741_ (.A1(_13044_),
    .A2(_13046_),
    .A3(_13049_),
    .ZN(_13050_));
 NAND3_X1 _22742_ (.A1(_12350_),
    .A2(_11153_),
    .A3(_11297_),
    .ZN(_13051_));
 OAI21_X1 _22743_ (.A(_13051_),
    .B1(_11276_),
    .B2(_12268_),
    .ZN(_13052_));
 AND3_X1 _22744_ (.A1(_11303_),
    .A2(_12274_),
    .A3(_11293_),
    .ZN(_13053_));
 AND2_X1 _22745_ (.A1(_11274_),
    .A2(_11195_),
    .ZN(_13054_));
 AND2_X1 _22746_ (.A1(_11277_),
    .A2(_11293_),
    .ZN(_13055_));
 NOR4_X1 _22747_ (.A1(_13052_),
    .A2(_13053_),
    .A3(_13054_),
    .A4(_13055_),
    .ZN(_13056_));
 NAND4_X2 _22748_ (.A1(_13031_),
    .A2(_13038_),
    .A3(_13050_),
    .A4(_13056_),
    .ZN(_13057_));
 NOR2_X4 _22749_ (.A1(_13022_),
    .A2(_13057_),
    .ZN(_13058_));
 INV_X2 _22750_ (.A(_11703_),
    .ZN(_13059_));
 OAI21_X1 _22751_ (.A(_13059_),
    .B1(_11927_),
    .B2(_12190_),
    .ZN(_13060_));
 AOI21_X1 _22752_ (.A(_12190_),
    .B1(_11886_),
    .B2(_11649_),
    .ZN(_13061_));
 AOI21_X1 _22753_ (.A(_12190_),
    .B1(_11720_),
    .B2(_11688_),
    .ZN(_13062_));
 NOR4_X1 _22754_ (.A1(_13060_),
    .A2(_11707_),
    .A3(_13061_),
    .A4(_13062_),
    .ZN(_13063_));
 AND2_X2 _22755_ (.A1(_11694_),
    .A2(_11691_),
    .ZN(_13064_));
 AND3_X1 _22756_ (.A1(_11659_),
    .A2(_11634_),
    .A3(_11681_),
    .ZN(_13065_));
 AND3_X1 _22757_ (.A1(_11797_),
    .A2(_11634_),
    .A3(_11681_),
    .ZN(_13066_));
 NOR4_X1 _22758_ (.A1(_13064_),
    .A2(_13065_),
    .A3(_12189_),
    .A4(_13066_),
    .ZN(_13067_));
 OAI21_X1 _22759_ (.A(_11694_),
    .B1(_11645_),
    .B2(_11724_),
    .ZN(_13068_));
 OAI21_X1 _22760_ (.A(_11694_),
    .B1(_11747_),
    .B2(_11748_),
    .ZN(_13069_));
 AND4_X1 _22761_ (.A1(_13063_),
    .A2(_13067_),
    .A3(_13068_),
    .A4(_13069_),
    .ZN(_13070_));
 INV_X1 _22762_ (.A(_11875_),
    .ZN(_13071_));
 NAND3_X1 _22763_ (.A1(_11828_),
    .A2(_12604_),
    .A3(_11945_),
    .ZN(_13072_));
 NAND4_X1 _22764_ (.A1(_13071_),
    .A2(_12612_),
    .A3(_12608_),
    .A4(_13072_),
    .ZN(_13073_));
 NAND4_X1 _22765_ (.A1(_11635_),
    .A2(_11626_),
    .A3(_11676_),
    .A4(_12246_),
    .ZN(_13074_));
 NAND4_X1 _22766_ (.A1(_11737_),
    .A2(_11634_),
    .A3(_11637_),
    .A4(_12246_),
    .ZN(_13075_));
 INV_X1 _22767_ (.A(_11664_),
    .ZN(_13076_));
 OAI211_X2 _22768_ (.A(_13074_),
    .B(_13075_),
    .C1(_13076_),
    .C2(_11815_),
    .ZN(_13077_));
 OAI21_X1 _22769_ (.A(_11671_),
    .B1(_11919_),
    .B2(_13076_),
    .ZN(_13078_));
 AOI21_X1 _22770_ (.A(_13076_),
    .B1(_12187_),
    .B2(_11725_),
    .ZN(_13079_));
 NOR4_X2 _22771_ (.A1(_13073_),
    .A2(_13077_),
    .A3(_13078_),
    .A4(_13079_),
    .ZN(_13080_));
 OAI21_X1 _22772_ (.A(_12244_),
    .B1(_12250_),
    .B2(_12200_),
    .ZN(_13081_));
 NAND4_X1 _22773_ (.A1(_11737_),
    .A2(_11826_),
    .A3(_11637_),
    .A4(_12246_),
    .ZN(_13082_));
 NAND3_X1 _22774_ (.A1(_13081_),
    .A2(_12593_),
    .A3(_13082_),
    .ZN(_13083_));
 AND2_X1 _22775_ (.A1(_11889_),
    .A2(_11823_),
    .ZN(_13084_));
 AOI21_X1 _22776_ (.A(_12590_),
    .B1(_11720_),
    .B2(_12644_),
    .ZN(_13085_));
 NOR4_X2 _22777_ (.A1(_13083_),
    .A2(_13084_),
    .A3(_12241_),
    .A4(_13085_),
    .ZN(_13086_));
 AND4_X1 _22778_ (.A1(_11701_),
    .A2(_11821_),
    .A3(_11637_),
    .A4(_11762_),
    .ZN(_13087_));
 AND4_X1 _22779_ (.A1(_16773_),
    .A2(_11701_),
    .A3(_11821_),
    .A4(_11762_),
    .ZN(_13088_));
 AOI211_X2 _22780_ (.A(_13087_),
    .B(_13088_),
    .C1(_11758_),
    .C2(_11852_),
    .ZN(_13089_));
 AOI21_X1 _22781_ (.A(_12618_),
    .B1(_11888_),
    .B2(_11862_),
    .ZN(_13090_));
 AND2_X2 _22782_ (.A1(_11837_),
    .A2(_11911_),
    .ZN(_13091_));
 NOR4_X1 _22783_ (.A1(_13090_),
    .A2(_11844_),
    .A3(_12235_),
    .A4(_13091_),
    .ZN(_13092_));
 NAND4_X1 _22784_ (.A1(_11852_),
    .A2(_11735_),
    .A3(_11850_),
    .A4(_11945_),
    .ZN(_13093_));
 OAI21_X1 _22785_ (.A(_11852_),
    .B1(_12202_),
    .B2(_11748_),
    .ZN(_13094_));
 AND4_X2 _22786_ (.A1(_13089_),
    .A2(_13092_),
    .A3(_13093_),
    .A4(_13094_),
    .ZN(_13095_));
 NAND4_X2 _22787_ (.A1(_13070_),
    .A2(_13080_),
    .A3(_13086_),
    .A4(_13095_),
    .ZN(_13096_));
 AOI21_X1 _22788_ (.A(_11925_),
    .B1(_11720_),
    .B2(_11688_),
    .ZN(_13097_));
 AOI21_X1 _22789_ (.A(_11925_),
    .B1(_11886_),
    .B2(_11942_),
    .ZN(_13098_));
 AND2_X2 _22790_ (.A1(_11742_),
    .A2(_11780_),
    .ZN(_13099_));
 OR3_X4 _22791_ (.A1(_13097_),
    .A2(_13098_),
    .A3(_13099_),
    .ZN(_13100_));
 AND2_X1 _22792_ (.A1(_11803_),
    .A2(_11673_),
    .ZN(_13101_));
 AOI21_X1 _22793_ (.A(_11922_),
    .B1(_12187_),
    .B2(_11649_),
    .ZN(_13102_));
 OAI21_X1 _22794_ (.A(_11808_),
    .B1(_11922_),
    .B2(_12644_),
    .ZN(_13103_));
 NOR4_X4 _22795_ (.A1(_13100_),
    .A2(_13101_),
    .A3(_13102_),
    .A4(_13103_),
    .ZN(_13104_));
 AND2_X1 _22796_ (.A1(_11666_),
    .A2(_11902_),
    .ZN(_13105_));
 OAI21_X1 _22797_ (.A(_11817_),
    .B1(_12202_),
    .B2(_13105_),
    .ZN(_13106_));
 OAI21_X1 _22798_ (.A(_11817_),
    .B1(_11718_),
    .B2(_11792_),
    .ZN(_13107_));
 OAI211_X2 _22799_ (.A(_11777_),
    .B(_11681_),
    .C1(_11936_),
    .C2(_11748_),
    .ZN(_13108_));
 NAND2_X1 _22800_ (.A1(_11791_),
    .A2(_11804_),
    .ZN(_13109_));
 AND2_X1 _22801_ (.A1(_13108_),
    .A2(_13109_),
    .ZN(_13110_));
 OAI21_X1 _22802_ (.A(_11791_),
    .B1(_11655_),
    .B2(_12205_),
    .ZN(_13111_));
 AND4_X1 _22803_ (.A1(_13106_),
    .A2(_13107_),
    .A3(_13110_),
    .A4(_13111_),
    .ZN(_13112_));
 AND3_X1 _22804_ (.A1(_11731_),
    .A2(_11652_),
    .A3(_11701_),
    .ZN(_13113_));
 AOI211_X2 _22805_ (.A(_13113_),
    .B(_12222_),
    .C1(_11731_),
    .C2(_11758_),
    .ZN(_13114_));
 NAND2_X1 _22806_ (.A1(_11747_),
    .A2(_11731_),
    .ZN(_13115_));
 NAND4_X1 _22807_ (.A1(_11666_),
    .A2(_11626_),
    .A3(_11712_),
    .A4(_11663_),
    .ZN(_13116_));
 AND3_X1 _22808_ (.A1(_11948_),
    .A2(_13115_),
    .A3(_13116_),
    .ZN(_13117_));
 AND2_X1 _22809_ (.A1(_11713_),
    .A2(_11691_),
    .ZN(_13118_));
 AND2_X1 _22810_ (.A1(_11713_),
    .A2(_11848_),
    .ZN(_13119_));
 NOR2_X1 _22811_ (.A1(_13118_),
    .A2(_13119_),
    .ZN(_13120_));
 OAI21_X1 _22812_ (.A(_11727_),
    .B1(_11726_),
    .B2(_11747_),
    .ZN(_13121_));
 AND4_X2 _22813_ (.A1(_13114_),
    .A2(_13117_),
    .A3(_13120_),
    .A4(_13121_),
    .ZN(_13122_));
 NAND3_X1 _22814_ (.A1(_11797_),
    .A2(_11712_),
    .A3(_11841_),
    .ZN(_13123_));
 OAI21_X1 _22815_ (.A(_13123_),
    .B1(_12629_),
    .B2(_12644_),
    .ZN(_13124_));
 AND3_X1 _22816_ (.A1(_11828_),
    .A2(_11945_),
    .A3(_11764_),
    .ZN(_13125_));
 AND2_X2 _22817_ (.A1(_11747_),
    .A2(_11764_),
    .ZN(_13126_));
 NOR4_X1 _22818_ (.A1(_13124_),
    .A2(_13125_),
    .A3(_11937_),
    .A4(_13126_),
    .ZN(_13127_));
 NAND4_X4 _22819_ (.A1(_13104_),
    .A2(_13112_),
    .A3(_13122_),
    .A4(_13127_),
    .ZN(_13128_));
 NOR2_X4 _22820_ (.A1(_13096_),
    .A2(_13128_),
    .ZN(_13129_));
 XOR2_X1 _22821_ (.A(_13058_),
    .B(_13129_),
    .Z(_13130_));
 AOI211_X4 _22822_ (.A(_12023_),
    .B(_12563_),
    .C1(_12860_),
    .C2(_12066_),
    .ZN(_13131_));
 BUF_X4 _22823_ (.A(_12037_),
    .Z(_13132_));
 OAI21_X1 _22824_ (.A(_13132_),
    .B1(_12163_),
    .B2(_12156_),
    .ZN(_13133_));
 OAI21_X1 _22825_ (.A(_13132_),
    .B1(_12052_),
    .B2(_12044_),
    .ZN(_13134_));
 AND4_X1 _22826_ (.A1(_12014_),
    .A2(_13131_),
    .A3(_13133_),
    .A4(_13134_),
    .ZN(_13135_));
 AND2_X1 _22827_ (.A1(_12062_),
    .A2(_12119_),
    .ZN(_13136_));
 AND2_X1 _22828_ (.A1(_12061_),
    .A2(_12484_),
    .ZN(_13137_));
 AND3_X1 _22829_ (.A1(_12005_),
    .A2(_11993_),
    .A3(_12496_),
    .ZN(_13138_));
 OR4_X2 _22830_ (.A1(_13136_),
    .A2(_12874_),
    .A3(_13137_),
    .A4(_13138_),
    .ZN(_13139_));
 NOR2_X1 _22831_ (.A1(_12058_),
    .A2(_12533_),
    .ZN(_13140_));
 AND2_X1 _22832_ (.A1(_12056_),
    .A2(_12528_),
    .ZN(_13141_));
 AOI211_X4 _22833_ (.A(_11975_),
    .B(_12058_),
    .C1(_11970_),
    .C2(_16862_),
    .ZN(_13142_));
 NOR4_X1 _22834_ (.A1(_13139_),
    .A2(_13140_),
    .A3(_13141_),
    .A4(_13142_),
    .ZN(_13143_));
 BUF_X4 _22835_ (.A(_11995_),
    .Z(_13144_));
 OAI21_X1 _22836_ (.A(_13144_),
    .B1(_12861_),
    .B2(_12039_),
    .ZN(_13145_));
 OAI21_X1 _22837_ (.A(_13144_),
    .B1(_12152_),
    .B2(_12484_),
    .ZN(_13146_));
 OAI21_X1 _22838_ (.A(_13144_),
    .B1(_12068_),
    .B2(_12493_),
    .ZN(_13147_));
 NAND4_X1 _22839_ (.A1(_13145_),
    .A2(_13146_),
    .A3(_13147_),
    .A4(_12872_),
    .ZN(_13148_));
 OAI21_X1 _22840_ (.A(_11964_),
    .B1(_12476_),
    .B2(_12168_),
    .ZN(_13149_));
 NAND2_X1 _22841_ (.A1(_12861_),
    .A2(_11964_),
    .ZN(_13150_));
 NAND2_X1 _22842_ (.A1(_13149_),
    .A2(_13150_),
    .ZN(_13151_));
 AOI21_X1 _22843_ (.A(_12850_),
    .B1(_12509_),
    .B2(_12092_),
    .ZN(_13152_));
 NOR3_X1 _22844_ (.A1(_13148_),
    .A2(_13151_),
    .A3(_13152_),
    .ZN(_13153_));
 INV_X1 _22845_ (.A(_12486_),
    .ZN(_13154_));
 OAI21_X1 _22846_ (.A(_12487_),
    .B1(_12082_),
    .B2(_12068_),
    .ZN(_13155_));
 OAI21_X1 _22847_ (.A(_12079_),
    .B1(_12834_),
    .B2(_12044_),
    .ZN(_13156_));
 OAI21_X1 _22848_ (.A(_12079_),
    .B1(_12861_),
    .B2(_12075_),
    .ZN(_13157_));
 AND4_X1 _22849_ (.A1(_13154_),
    .A2(_13155_),
    .A3(_13156_),
    .A4(_13157_),
    .ZN(_13158_));
 OAI211_X2 _22850_ (.A(_12088_),
    .B(_12528_),
    .C1(_11969_),
    .C2(_11970_),
    .ZN(_13159_));
 OAI21_X1 _22851_ (.A(_12088_),
    .B1(_12503_),
    .B2(_12861_),
    .ZN(_13160_));
 AND3_X1 _22852_ (.A1(_13158_),
    .A2(_13159_),
    .A3(_13160_),
    .ZN(_13161_));
 AND4_X1 _22853_ (.A1(_13135_),
    .A2(_13143_),
    .A3(_13153_),
    .A4(_13161_),
    .ZN(_13162_));
 AND2_X1 _22854_ (.A1(_12009_),
    .A2(_12830_),
    .ZN(_13163_));
 BUF_X8 _22855_ (.A(_12048_),
    .Z(_13164_));
 OAI21_X2 _22856_ (.A(_12117_),
    .B1(_12834_),
    .B2(_13164_),
    .ZN(_13165_));
 NAND4_X1 _22857_ (.A1(_12123_),
    .A2(_13165_),
    .A3(_12120_),
    .A4(_12512_),
    .ZN(_13166_));
 NAND2_X1 _22858_ (.A1(_12857_),
    .A2(_12532_),
    .ZN(_13167_));
 NAND3_X1 _22859_ (.A1(_12830_),
    .A2(_12090_),
    .A3(_12031_),
    .ZN(_13168_));
 NAND2_X1 _22860_ (.A1(_13167_),
    .A2(_13168_),
    .ZN(_13169_));
 NOR3_X1 _22861_ (.A1(_12131_),
    .A2(_12024_),
    .A3(_12489_),
    .ZN(_13170_));
 OR4_X1 _22862_ (.A1(_13163_),
    .A2(_13166_),
    .A3(_13169_),
    .A4(_13170_),
    .ZN(_13171_));
 AND2_X1 _22863_ (.A1(_12108_),
    .A2(_12109_),
    .ZN(_13172_));
 AND2_X1 _22864_ (.A1(_12107_),
    .A2(_12019_),
    .ZN(_13173_));
 AOI211_X2 _22865_ (.A(_13172_),
    .B(_13173_),
    .C1(_12152_),
    .C2(_12527_),
    .ZN(_13174_));
 AND2_X1 _22866_ (.A1(_11983_),
    .A2(_12544_),
    .ZN(_13175_));
 NOR4_X1 _22867_ (.A1(_12553_),
    .A2(_12099_),
    .A3(_13175_),
    .A4(_12551_),
    .ZN(_13176_));
 INV_X1 _22868_ (.A(_12108_),
    .ZN(_13177_));
 INV_X1 _22869_ (.A(_12168_),
    .ZN(_13178_));
 AOI21_X1 _22870_ (.A(_13177_),
    .B1(_13178_),
    .B2(_12840_),
    .ZN(_13179_));
 INV_X1 _22871_ (.A(_12122_),
    .ZN(_13180_));
 NAND2_X1 _22872_ (.A1(_12849_),
    .A2(_13180_),
    .ZN(_13181_));
 AOI21_X1 _22873_ (.A(_13179_),
    .B1(_12527_),
    .B2(_13181_),
    .ZN(_13182_));
 OAI21_X1 _22874_ (.A(_12150_),
    .B1(_12019_),
    .B2(_11997_),
    .ZN(_13183_));
 OAI21_X1 _22875_ (.A(_12142_),
    .B1(_12019_),
    .B2(_13164_),
    .ZN(_13184_));
 OAI21_X1 _22876_ (.A(_12142_),
    .B1(_12861_),
    .B2(_12156_),
    .ZN(_13185_));
 OAI21_X1 _22877_ (.A(_12150_),
    .B1(_12861_),
    .B2(_12493_),
    .ZN(_13186_));
 AND4_X1 _22878_ (.A1(_13183_),
    .A2(_13184_),
    .A3(_13185_),
    .A4(_13186_),
    .ZN(_13187_));
 NAND4_X1 _22879_ (.A1(_13174_),
    .A2(_13176_),
    .A3(_13182_),
    .A4(_13187_),
    .ZN(_13188_));
 NOR2_X1 _22880_ (.A1(_12853_),
    .A2(_12533_),
    .ZN(_13189_));
 NAND4_X1 _22881_ (.A1(_12026_),
    .A2(_12090_),
    .A3(_12031_),
    .A4(_12113_),
    .ZN(_13190_));
 INV_X4 _22882_ (.A(_12075_),
    .ZN(_13191_));
 OAI21_X1 _22883_ (.A(_13190_),
    .B1(_12853_),
    .B2(_13191_),
    .ZN(_13192_));
 AOI21_X1 _22884_ (.A(_12853_),
    .B1(_12073_),
    .B2(_12045_),
    .ZN(_13193_));
 AND4_X1 _22885_ (.A1(_12026_),
    .A2(_12113_),
    .A3(_12024_),
    .A4(_11999_),
    .ZN(_13194_));
 OR4_X1 _22886_ (.A1(_13189_),
    .A2(_13192_),
    .A3(_13193_),
    .A4(_13194_),
    .ZN(_13195_));
 OAI21_X1 _22887_ (.A(_12162_),
    .B1(_12507_),
    .B2(_12015_),
    .ZN(_13196_));
 OAI211_X2 _22888_ (.A(_13196_),
    .B(_12524_),
    .C1(_12157_),
    .C2(_12839_),
    .ZN(_13197_));
 NOR4_X4 _22889_ (.A1(_13171_),
    .A2(_13188_),
    .A3(_13195_),
    .A4(_13197_),
    .ZN(_13198_));
 NAND2_X2 _22890_ (.A1(_13162_),
    .A2(_13198_),
    .ZN(_13199_));
 XNOR2_X2 _22891_ (.A(_13199_),
    .B(_12175_),
    .ZN(_13200_));
 XNOR2_X2 _22892_ (.A(_13130_),
    .B(_13200_),
    .ZN(_13201_));
 XNOR2_X1 _22893_ (.A(_12984_),
    .B(_13201_),
    .ZN(_13202_));
 XNOR2_X1 _22894_ (.A(_13202_),
    .B(_17265_),
    .ZN(_13203_));
 MUX2_X1 _22895_ (.A(_12908_),
    .B(_13203_),
    .S(_11149_),
    .Z(_00719_));
 XOR2_X1 _22896_ (.A(_17266_),
    .B(_17069_),
    .Z(_13204_));
 AND4_X1 _22897_ (.A1(_11970_),
    .A2(_12054_),
    .A3(_12035_),
    .A4(_11982_),
    .ZN(_13205_));
 AND2_X1 _22898_ (.A1(_12079_),
    .A2(_11983_),
    .ZN(_13206_));
 AOI211_X4 _22899_ (.A(_13205_),
    .B(_13206_),
    .C1(_12079_),
    .C2(_13181_),
    .ZN(_13207_));
 NAND4_X1 _22900_ (.A1(_12496_),
    .A2(_11969_),
    .A3(_11990_),
    .A4(_12035_),
    .ZN(_13208_));
 OAI211_X2 _22901_ (.A(_12487_),
    .B(_12528_),
    .C1(_12089_),
    .C2(_11970_),
    .ZN(_13209_));
 NAND3_X1 _22902_ (.A1(_13207_),
    .A2(_13208_),
    .A3(_13209_),
    .ZN(_13210_));
 AND2_X1 _22903_ (.A1(_12085_),
    .A2(_12109_),
    .ZN(_13211_));
 INV_X1 _22904_ (.A(_13211_),
    .ZN(_13212_));
 AND2_X1 _22905_ (.A1(_13212_),
    .A2(_12498_),
    .ZN(_13213_));
 OAI21_X1 _22906_ (.A(_12088_),
    .B1(_12861_),
    .B2(_12025_),
    .ZN(_13214_));
 OAI211_X2 _22907_ (.A(_13213_),
    .B(_13214_),
    .C1(_12509_),
    .C2(_12837_),
    .ZN(_13215_));
 AND2_X4 _22908_ (.A1(_12503_),
    .A2(_12055_),
    .ZN(_13216_));
 AND2_X1 _22909_ (.A1(_12055_),
    .A2(_12128_),
    .ZN(_13217_));
 AND2_X1 _22910_ (.A1(_12055_),
    .A2(_12080_),
    .ZN(_13218_));
 OR4_X4 _22911_ (.A1(_13140_),
    .A2(_13216_),
    .A3(_13217_),
    .A4(_13218_),
    .ZN(_13219_));
 AND2_X1 _22912_ (.A1(_12066_),
    .A2(_12062_),
    .ZN(_13220_));
 AND3_X1 _22913_ (.A1(_12552_),
    .A2(_11993_),
    .A3(_12054_),
    .ZN(_13221_));
 OR4_X4 _22914_ (.A1(_13220_),
    .A2(_12898_),
    .A3(_13137_),
    .A4(_13221_),
    .ZN(_13222_));
 OR4_X4 _22915_ (.A1(_13210_),
    .A2(_13215_),
    .A3(_13219_),
    .A4(_13222_),
    .ZN(_13223_));
 OAI211_X2 _22916_ (.A(_13132_),
    .B(_12090_),
    .C1(_11969_),
    .C2(_11970_),
    .ZN(_13224_));
 OAI211_X2 _22917_ (.A(_13132_),
    .B(_12528_),
    .C1(_12024_),
    .C2(_11987_),
    .ZN(_13225_));
 OAI21_X1 _22918_ (.A(_13132_),
    .B1(_12050_),
    .B2(_12484_),
    .ZN(_13226_));
 NAND4_X1 _22919_ (.A1(_13224_),
    .A2(_13225_),
    .A3(_12574_),
    .A4(_13226_),
    .ZN(_13227_));
 OAI211_X2 _22920_ (.A(_12860_),
    .B(_12528_),
    .C1(_12089_),
    .C2(_12000_),
    .ZN(_13228_));
 OAI211_X2 _22921_ (.A(_12860_),
    .B(_11990_),
    .C1(_11981_),
    .C2(_12031_),
    .ZN(_13229_));
 OAI211_X2 _22922_ (.A(_12860_),
    .B(_12090_),
    .C1(_11969_),
    .C2(_12000_),
    .ZN(_13230_));
 OAI21_X1 _22923_ (.A(_12860_),
    .B1(_12068_),
    .B2(_12493_),
    .ZN(_13231_));
 NAND4_X1 _22924_ (.A1(_13228_),
    .A2(_13229_),
    .A3(_13230_),
    .A4(_13231_),
    .ZN(_13232_));
 OAI21_X1 _22925_ (.A(_13144_),
    .B1(_12135_),
    .B2(_12152_),
    .ZN(_13233_));
 NAND2_X1 _22926_ (.A1(_13144_),
    .A2(_12493_),
    .ZN(_13234_));
 AND3_X1 _22927_ (.A1(_13233_),
    .A2(_12006_),
    .A3(_13234_),
    .ZN(_13235_));
 NAND3_X1 _22928_ (.A1(_11964_),
    .A2(_11987_),
    .A3(_11967_),
    .ZN(_13236_));
 NAND2_X1 _22929_ (.A1(_13164_),
    .A2(_11964_),
    .ZN(_13237_));
 OAI211_X2 _22930_ (.A(_13236_),
    .B(_13237_),
    .C1(_12535_),
    .C2(_12850_),
    .ZN(_13238_));
 AOI21_X1 _22931_ (.A(_12850_),
    .B1(_12849_),
    .B2(_13191_),
    .ZN(_13239_));
 NOR4_X1 _22932_ (.A1(_13238_),
    .A2(_13239_),
    .A3(_12559_),
    .A4(_11974_),
    .ZN(_13240_));
 NAND2_X1 _22933_ (.A1(_13235_),
    .A2(_13240_),
    .ZN(_13241_));
 NOR4_X4 _22934_ (.A1(_13223_),
    .A2(_13227_),
    .A3(_13232_),
    .A4(_13241_),
    .ZN(_13242_));
 AND4_X1 _22935_ (.A1(_12491_),
    .A2(_12544_),
    .A3(_12064_),
    .A4(_11967_),
    .ZN(_13243_));
 AND4_X1 _22936_ (.A1(_11980_),
    .A2(_12030_),
    .A3(_12097_),
    .A4(_12035_),
    .ZN(_13244_));
 OR4_X2 _22937_ (.A1(_12551_),
    .A2(_13243_),
    .A3(_13175_),
    .A4(_13244_),
    .ZN(_13245_));
 INV_X1 _22938_ (.A(_13173_),
    .ZN(_13246_));
 NAND2_X1 _22939_ (.A1(_12527_),
    .A2(_12476_),
    .ZN(_13247_));
 OAI21_X1 _22940_ (.A(_12527_),
    .B1(_12168_),
    .B2(_12493_),
    .ZN(_13248_));
 NAND4_X1 _22941_ (.A1(_12892_),
    .A2(_13246_),
    .A3(_13247_),
    .A4(_13248_),
    .ZN(_13249_));
 OR2_X1 _22942_ (.A1(_13245_),
    .A2(_13249_),
    .ZN(_13250_));
 AOI21_X1 _22943_ (.A(_12131_),
    .B1(_12508_),
    .B2(_12072_),
    .ZN(_13251_));
 AND3_X1 _22944_ (.A1(_12830_),
    .A2(_12090_),
    .A3(_12024_),
    .ZN(_13252_));
 AND2_X1 _22945_ (.A1(_12068_),
    .A2(_12830_),
    .ZN(_13253_));
 NOR4_X1 _22946_ (.A1(_13251_),
    .A2(_12126_),
    .A3(_13252_),
    .A4(_13253_),
    .ZN(_13254_));
 OAI21_X1 _22947_ (.A(_12117_),
    .B1(_12484_),
    .B2(_12479_),
    .ZN(_13255_));
 NAND3_X1 _22948_ (.A1(_12044_),
    .A2(_12113_),
    .A3(_12863_),
    .ZN(_13256_));
 AND2_X1 _22949_ (.A1(_13255_),
    .A2(_13256_),
    .ZN(_13257_));
 AND3_X1 _22950_ (.A1(_12068_),
    .A2(_12113_),
    .A3(_12863_),
    .ZN(_13258_));
 AOI21_X1 _22951_ (.A(_13258_),
    .B1(_13181_),
    .B2(_12117_),
    .ZN(_13259_));
 NAND2_X1 _22952_ (.A1(_12168_),
    .A2(_12167_),
    .ZN(_13260_));
 OAI21_X1 _22953_ (.A(_12162_),
    .B1(_12109_),
    .B2(_12128_),
    .ZN(_13261_));
 OAI21_X1 _22954_ (.A(_12167_),
    .B1(_12152_),
    .B2(_12552_),
    .ZN(_13262_));
 NAND2_X1 _22955_ (.A1(_12022_),
    .A2(_12161_),
    .ZN(_13263_));
 AND4_X1 _22956_ (.A1(_13260_),
    .A2(_13261_),
    .A3(_13262_),
    .A4(_13263_),
    .ZN(_13264_));
 NAND4_X1 _22957_ (.A1(_13254_),
    .A2(_13257_),
    .A3(_13259_),
    .A4(_13264_),
    .ZN(_13265_));
 OAI211_X2 _22958_ (.A(_12150_),
    .B(_11990_),
    .C1(_12089_),
    .C2(_11970_),
    .ZN(_13266_));
 OAI21_X1 _22959_ (.A(_12150_),
    .B1(_12039_),
    .B2(_12040_),
    .ZN(_13267_));
 OAI211_X2 _22960_ (.A(_13266_),
    .B(_13267_),
    .C1(_12151_),
    .C2(_12506_),
    .ZN(_13268_));
 AND2_X1 _22961_ (.A1(_12142_),
    .A2(_12552_),
    .ZN(_13269_));
 AOI21_X1 _22962_ (.A(_12143_),
    .B1(_12155_),
    .B2(_13191_),
    .ZN(_13270_));
 AND2_X1 _22963_ (.A1(_12142_),
    .A2(_13164_),
    .ZN(_13271_));
 AND3_X1 _22964_ (.A1(_12863_),
    .A2(_12097_),
    .A3(_11999_),
    .ZN(_13272_));
 OR4_X1 _22965_ (.A1(_13269_),
    .A2(_13270_),
    .A3(_13271_),
    .A4(_13272_),
    .ZN(_13273_));
 NOR4_X1 _22966_ (.A1(_13250_),
    .A2(_13265_),
    .A3(_13268_),
    .A4(_13273_),
    .ZN(_13274_));
 AND2_X4 _22967_ (.A1(_13242_),
    .A2(_13274_),
    .ZN(_13275_));
 XNOR2_X2 _22968_ (.A(_13275_),
    .B(_12176_),
    .ZN(_13276_));
 AND4_X1 _22969_ (.A1(_11643_),
    .A2(_11634_),
    .A3(_11673_),
    .A4(_11762_),
    .ZN(_13277_));
 AOI211_X2 _22970_ (.A(_13277_),
    .B(_11859_),
    .C1(_11749_),
    .C2(_11705_),
    .ZN(_13278_));
 OAI21_X1 _22971_ (.A(_11694_),
    .B1(_11818_),
    .B2(_12205_),
    .ZN(_13279_));
 OAI21_X1 _22972_ (.A(_11694_),
    .B1(_11645_),
    .B2(_11695_),
    .ZN(_13280_));
 AND4_X1 _22973_ (.A1(_13059_),
    .A2(_13278_),
    .A3(_13279_),
    .A4(_13280_),
    .ZN(_13281_));
 OAI21_X1 _22974_ (.A(_12620_),
    .B1(_11655_),
    .B2(_11659_),
    .ZN(_13282_));
 OAI211_X2 _22975_ (.A(_11852_),
    .B(_12605_),
    .C1(_11761_),
    .C2(_11699_),
    .ZN(_13283_));
 NAND2_X1 _22976_ (.A1(_12202_),
    .A2(_12620_),
    .ZN(_13284_));
 AND3_X1 _22977_ (.A1(_13282_),
    .A2(_13283_),
    .A3(_13284_),
    .ZN(_13285_));
 AND2_X1 _22978_ (.A1(_11878_),
    .A2(_11822_),
    .ZN(_13286_));
 NOR2_X1 _22979_ (.A1(_12653_),
    .A2(_12590_),
    .ZN(_13287_));
 AOI211_X2 _22980_ (.A(_13286_),
    .B(_13287_),
    .C1(_12200_),
    .C2(_11823_),
    .ZN(_13288_));
 OAI21_X1 _22981_ (.A(_12244_),
    .B1(_12200_),
    .B2(_11835_),
    .ZN(_13289_));
 AND3_X1 _22982_ (.A1(_13289_),
    .A2(_11830_),
    .A3(_12247_),
    .ZN(_13290_));
 AND2_X1 _22983_ (.A1(_11838_),
    .A2(_11659_),
    .ZN(_13291_));
 NOR4_X1 _22984_ (.A1(_11843_),
    .A2(_12237_),
    .A3(_13091_),
    .A4(_13291_),
    .ZN(_13292_));
 AND4_X1 _22985_ (.A1(_13285_),
    .A2(_13288_),
    .A3(_13290_),
    .A4(_13292_),
    .ZN(_13293_));
 AND4_X1 _22986_ (.A1(_11902_),
    .A2(_11737_),
    .A3(_11635_),
    .A4(_12246_),
    .ZN(_13294_));
 AOI211_X4 _22987_ (.A(_13294_),
    .B(_12602_),
    .C1(_11782_),
    .C2(_11880_),
    .ZN(_13295_));
 OAI21_X1 _22988_ (.A(_12604_),
    .B1(_11751_),
    .B2(_11749_),
    .ZN(_13296_));
 NAND2_X1 _22989_ (.A1(_12604_),
    .A2(_11782_),
    .ZN(_13297_));
 AND4_X1 _22990_ (.A1(_11660_),
    .A2(_13296_),
    .A3(_11876_),
    .A4(_13297_),
    .ZN(_13298_));
 AND4_X4 _22991_ (.A1(_13281_),
    .A2(_13293_),
    .A3(_13295_),
    .A4(_13298_),
    .ZN(_13299_));
 AND2_X1 _22992_ (.A1(_11803_),
    .A2(_11782_),
    .ZN(_13300_));
 AOI211_X4 _22993_ (.A(_11801_),
    .B(_13300_),
    .C1(_11655_),
    .C2(_11803_),
    .ZN(_13301_));
 AND4_X1 _22994_ (.A1(_11676_),
    .A2(_11777_),
    .A3(_11626_),
    .A4(_12246_),
    .ZN(_13302_));
 AOI211_X4 _22995_ (.A(_13302_),
    .B(_11773_),
    .C1(_11716_),
    .C2(_11780_),
    .ZN(_13303_));
 OAI21_X1 _22996_ (.A(_11803_),
    .B1(_11775_),
    .B2(_12200_),
    .ZN(_13304_));
 NAND4_X1 _22997_ (.A1(_13301_),
    .A2(_13303_),
    .A3(_12201_),
    .A4(_13304_),
    .ZN(_13305_));
 OAI211_X2 _22998_ (.A(_11777_),
    .B(_11841_),
    .C1(_11775_),
    .C2(_11839_),
    .ZN(_13306_));
 NAND2_X1 _22999_ (.A1(_11791_),
    .A2(_11716_),
    .ZN(_13307_));
 NAND4_X1 _23000_ (.A1(_11848_),
    .A2(_11850_),
    .A3(_11777_),
    .A4(_11841_),
    .ZN(_13308_));
 AND4_X1 _23001_ (.A1(_13109_),
    .A2(_13306_),
    .A3(_13307_),
    .A4(_13308_),
    .ZN(_13309_));
 NOR2_X1 _23002_ (.A1(_11907_),
    .A2(_11908_),
    .ZN(_13310_));
 OAI21_X1 _23003_ (.A(_11817_),
    .B1(_11839_),
    .B2(_11749_),
    .ZN(_13311_));
 NAND2_X1 _23004_ (.A1(_11817_),
    .A2(_11794_),
    .ZN(_13312_));
 NAND4_X1 _23005_ (.A1(_11777_),
    .A2(_11676_),
    .A3(_11637_),
    .A4(_11762_),
    .ZN(_13313_));
 AND3_X1 _23006_ (.A1(_11913_),
    .A2(_13312_),
    .A3(_13313_),
    .ZN(_13314_));
 NAND4_X1 _23007_ (.A1(_13309_),
    .A2(_13310_),
    .A3(_13311_),
    .A4(_13314_),
    .ZN(_13315_));
 NAND2_X1 _23008_ (.A1(_11727_),
    .A2(_11792_),
    .ZN(_13316_));
 OAI211_X2 _23009_ (.A(_11727_),
    .B(_12610_),
    .C1(_11733_),
    .C2(_11765_),
    .ZN(_13317_));
 OAI21_X1 _23010_ (.A(_11727_),
    .B1(_11775_),
    .B2(_11747_),
    .ZN(_13318_));
 NAND2_X1 _23011_ (.A1(_11858_),
    .A2(_11727_),
    .ZN(_13319_));
 AND4_X1 _23012_ (.A1(_13316_),
    .A2(_13317_),
    .A3(_13318_),
    .A4(_13319_),
    .ZN(_13320_));
 NAND2_X1 _23013_ (.A1(_11722_),
    .A2(_11732_),
    .ZN(_13321_));
 OAI21_X1 _23014_ (.A(_11732_),
    .B1(_11702_),
    .B2(_12205_),
    .ZN(_13322_));
 NAND4_X1 _23015_ (.A1(_13320_),
    .A2(_12655_),
    .A3(_13321_),
    .A4(_13322_),
    .ZN(_13323_));
 OAI21_X1 _23016_ (.A(_11764_),
    .B1(_11858_),
    .B2(_11749_),
    .ZN(_13324_));
 OAI211_X2 _23017_ (.A(_11764_),
    .B(_12610_),
    .C1(_11733_),
    .C2(_11765_),
    .ZN(_13325_));
 AND2_X1 _23018_ (.A1(_13324_),
    .A2(_13325_),
    .ZN(_13326_));
 OAI21_X1 _23019_ (.A(_11744_),
    .B1(_11722_),
    .B2(_11724_),
    .ZN(_13327_));
 OAI21_X1 _23020_ (.A(_11744_),
    .B1(_11742_),
    .B2(_11753_),
    .ZN(_13328_));
 OAI21_X1 _23021_ (.A(_11744_),
    .B1(_11839_),
    .B2(_11749_),
    .ZN(_13329_));
 NAND4_X1 _23022_ (.A1(_13326_),
    .A2(_13327_),
    .A3(_13328_),
    .A4(_13329_),
    .ZN(_13330_));
 NOR4_X1 _23023_ (.A1(_13305_),
    .A2(_13315_),
    .A3(_13323_),
    .A4(_13330_),
    .ZN(_13331_));
 AND2_X2 _23024_ (.A1(_13299_),
    .A2(_13331_),
    .ZN(_13332_));
 AND2_X1 _23025_ (.A1(_11171_),
    .A2(_12262_),
    .ZN(_13333_));
 NOR2_X1 _23026_ (.A1(_12670_),
    .A2(_13333_),
    .ZN(_13334_));
 OAI21_X1 _23027_ (.A(_12294_),
    .B1(_12295_),
    .B2(_11291_),
    .ZN(_13335_));
 AND3_X1 _23028_ (.A1(_11156_),
    .A2(_11348_),
    .A3(_12314_),
    .ZN(_13336_));
 AND2_X2 _23029_ (.A1(_11157_),
    .A2(_12282_),
    .ZN(_13337_));
 AND2_X1 _23030_ (.A1(_11156_),
    .A2(_11210_),
    .ZN(_13338_));
 NOR4_X2 _23031_ (.A1(_13335_),
    .A2(_13336_),
    .A3(_13337_),
    .A4(_13338_),
    .ZN(_13339_));
 OAI21_X1 _23032_ (.A(_11199_),
    .B1(_11230_),
    .B2(_11316_),
    .ZN(_13340_));
 NAND2_X1 _23033_ (.A1(_12343_),
    .A2(_11199_),
    .ZN(_13341_));
 NAND2_X1 _23034_ (.A1(_11214_),
    .A2(_11199_),
    .ZN(_13342_));
 NAND4_X1 _23035_ (.A1(_11167_),
    .A2(_11269_),
    .A3(_11298_),
    .A4(_11322_),
    .ZN(_13343_));
 AND3_X1 _23036_ (.A1(_13341_),
    .A2(_13342_),
    .A3(_13343_),
    .ZN(_13344_));
 AND4_X2 _23037_ (.A1(_13334_),
    .A2(_13339_),
    .A3(_13340_),
    .A4(_13344_),
    .ZN(_13345_));
 OAI21_X1 _23038_ (.A(_11275_),
    .B1(_12662_),
    .B2(_11258_),
    .ZN(_13346_));
 OAI211_X2 _23039_ (.A(_11293_),
    .B(_11165_),
    .C1(_11178_),
    .C2(_11233_),
    .ZN(_13347_));
 OAI21_X1 _23040_ (.A(_11293_),
    .B1(_11248_),
    .B2(_11316_),
    .ZN(_13348_));
 OAI21_X1 _23041_ (.A(_11275_),
    .B1(_11282_),
    .B2(_11284_),
    .ZN(_13349_));
 AND4_X1 _23042_ (.A1(_13346_),
    .A2(_13347_),
    .A3(_13348_),
    .A4(_13349_),
    .ZN(_13350_));
 OAI211_X2 _23043_ (.A(_11223_),
    .B(_11165_),
    .C1(_11269_),
    .C2(_11217_),
    .ZN(_13351_));
 NAND4_X1 _23044_ (.A1(_11167_),
    .A2(_11172_),
    .A3(_11234_),
    .A4(_11322_),
    .ZN(_13352_));
 NAND3_X1 _23045_ (.A1(_12290_),
    .A2(_13351_),
    .A3(_13352_),
    .ZN(_13353_));
 AOI21_X1 _23046_ (.A(_11205_),
    .B1(_11215_),
    .B2(_11246_),
    .ZN(_13354_));
 OAI21_X1 _23047_ (.A(_13045_),
    .B1(_11205_),
    .B2(_11191_),
    .ZN(_13355_));
 AND2_X1 _23048_ (.A1(_12683_),
    .A2(_12327_),
    .ZN(_13356_));
 NOR4_X1 _23049_ (.A1(_13353_),
    .A2(_13354_),
    .A3(_13355_),
    .A4(_13356_),
    .ZN(_13357_));
 NAND2_X1 _23050_ (.A1(_11264_),
    .A2(_11174_),
    .ZN(_13358_));
 OAI211_X2 _23051_ (.A(_11264_),
    .B(_12265_),
    .C1(_11178_),
    .C2(_11209_),
    .ZN(_13359_));
 OAI21_X1 _23052_ (.A(_11264_),
    .B1(_11190_),
    .B2(_11277_),
    .ZN(_13360_));
 NAND2_X1 _23053_ (.A1(_11248_),
    .A2(_11264_),
    .ZN(_13361_));
 AND4_X1 _23054_ (.A1(_13358_),
    .A2(_13359_),
    .A3(_13360_),
    .A4(_13361_),
    .ZN(_13362_));
 NAND3_X1 _23055_ (.A1(_11253_),
    .A2(_11269_),
    .A3(_11165_),
    .ZN(_13363_));
 OAI21_X1 _23056_ (.A(_11253_),
    .B1(_12276_),
    .B2(_11270_),
    .ZN(_13364_));
 AND4_X1 _23057_ (.A1(_12691_),
    .A2(_13362_),
    .A3(_13363_),
    .A4(_13364_),
    .ZN(_13365_));
 AND4_X2 _23058_ (.A1(_13345_),
    .A2(_13350_),
    .A3(_13357_),
    .A4(_13365_),
    .ZN(_13366_));
 AND2_X1 _23059_ (.A1(_12989_),
    .A2(_11348_),
    .ZN(_13367_));
 AOI21_X1 _23060_ (.A(_11330_),
    .B1(_11356_),
    .B2(_12334_),
    .ZN(_13368_));
 AND4_X1 _23061_ (.A1(_11213_),
    .A2(_11319_),
    .A3(_11232_),
    .A4(_11326_),
    .ZN(_13369_));
 NOR3_X1 _23062_ (.A1(_13367_),
    .A2(_13368_),
    .A3(_13369_),
    .ZN(_13370_));
 NAND4_X1 _23063_ (.A1(_13370_),
    .A2(_11317_),
    .A3(_12339_),
    .A4(_12723_),
    .ZN(_13371_));
 OAI21_X1 _23064_ (.A(_11363_),
    .B1(_11267_),
    .B2(_11200_),
    .ZN(_13372_));
 OAI21_X1 _23065_ (.A(_11363_),
    .B1(_11378_),
    .B2(_11364_),
    .ZN(_13373_));
 OAI21_X1 _23066_ (.A(_11375_),
    .B1(_11248_),
    .B2(_11258_),
    .ZN(_13374_));
 NAND4_X1 _23067_ (.A1(_13372_),
    .A2(_13373_),
    .A3(_13374_),
    .A4(_11374_),
    .ZN(_13375_));
 OAI21_X1 _23068_ (.A(_11309_),
    .B1(_11347_),
    .B2(_12704_),
    .ZN(_13376_));
 OAI21_X1 _23069_ (.A(_11336_),
    .B1(_11345_),
    .B2(_12350_),
    .ZN(_13377_));
 AND2_X1 _23070_ (.A1(_13377_),
    .A2(_13017_),
    .ZN(_13378_));
 NAND4_X1 _23071_ (.A1(_13376_),
    .A2(_11334_),
    .A3(_11333_),
    .A4(_13378_),
    .ZN(_13379_));
 NAND2_X1 _23072_ (.A1(_11345_),
    .A2(_11343_),
    .ZN(_13380_));
 NAND2_X1 _23073_ (.A1(_12282_),
    .A2(_11343_),
    .ZN(_13381_));
 NAND2_X1 _23074_ (.A1(_13380_),
    .A2(_13381_),
    .ZN(_13382_));
 AND2_X1 _23075_ (.A1(_11342_),
    .A2(_12327_),
    .ZN(_13383_));
 NOR2_X1 _23076_ (.A1(_13382_),
    .A2(_13383_),
    .ZN(_13384_));
 OAI21_X1 _23077_ (.A(_11371_),
    .B1(_12297_),
    .B2(_12327_),
    .ZN(_13385_));
 OAI21_X1 _23078_ (.A(_11343_),
    .B1(_11286_),
    .B2(_11316_),
    .ZN(_13386_));
 NAND4_X1 _23079_ (.A1(_13384_),
    .A2(_12710_),
    .A3(_13385_),
    .A4(_13386_),
    .ZN(_13387_));
 NOR4_X1 _23080_ (.A1(_13371_),
    .A2(_13375_),
    .A3(_13379_),
    .A4(_13387_),
    .ZN(_13388_));
 AND2_X4 _23081_ (.A1(_13366_),
    .A2(_13388_),
    .ZN(_13389_));
 XOR2_X2 _23082_ (.A(_13332_),
    .B(_13389_),
    .Z(_13390_));
 XNOR2_X1 _23083_ (.A(_13276_),
    .B(_13390_),
    .ZN(_13391_));
 XOR2_X2 _23084_ (.A(_11958_),
    .B(_13129_),
    .Z(_13392_));
 OAI211_X2 _23085_ (.A(_11546_),
    .B(_11399_),
    .C1(_11467_),
    .C2(_11529_),
    .ZN(_13393_));
 NAND2_X1 _23086_ (.A1(_11546_),
    .A2(_11441_),
    .ZN(_13394_));
 NAND3_X1 _23087_ (.A1(_11546_),
    .A2(_12393_),
    .A3(_12787_),
    .ZN(_13395_));
 NAND4_X1 _23088_ (.A1(_13393_),
    .A2(_12959_),
    .A3(_13394_),
    .A4(_13395_),
    .ZN(_13396_));
 AOI21_X1 _23089_ (.A(_12746_),
    .B1(_11525_),
    .B2(_11604_),
    .ZN(_13397_));
 AND3_X1 _23090_ (.A1(_11573_),
    .A2(_11406_),
    .A3(_11419_),
    .ZN(_13398_));
 AOI21_X1 _23091_ (.A(_12746_),
    .B1(_11584_),
    .B2(_11489_),
    .ZN(_13399_));
 NOR4_X1 _23092_ (.A1(_13396_),
    .A2(_13397_),
    .A3(_13398_),
    .A4(_13399_),
    .ZN(_13400_));
 OAI21_X1 _23093_ (.A(_12392_),
    .B1(_11450_),
    .B2(_11436_),
    .ZN(_13401_));
 AND3_X1 _23094_ (.A1(_11424_),
    .A2(_11457_),
    .A3(_11419_),
    .ZN(_13402_));
 OAI21_X1 _23095_ (.A(_11435_),
    .B1(_11524_),
    .B2(_11425_),
    .ZN(_13403_));
 AOI211_X2 _23096_ (.A(_13402_),
    .B(_13403_),
    .C1(_11442_),
    .C2(_11585_),
    .ZN(_13404_));
 OAI221_X1 _23097_ (.A(_12392_),
    .B1(_11467_),
    .B2(_11600_),
    .C1(_11412_),
    .C2(_11599_),
    .ZN(_13405_));
 OAI21_X1 _23098_ (.A(_12392_),
    .B1(_11556_),
    .B2(_12367_),
    .ZN(_13406_));
 AND4_X1 _23099_ (.A1(_13401_),
    .A2(_13404_),
    .A3(_13405_),
    .A4(_13406_),
    .ZN(_13407_));
 INV_X1 _23100_ (.A(_11555_),
    .ZN(_13408_));
 OAI21_X1 _23101_ (.A(_11559_),
    .B1(_11455_),
    .B2(_13408_),
    .ZN(_13409_));
 AOI21_X1 _23102_ (.A(_13409_),
    .B1(_11486_),
    .B2(_11555_),
    .ZN(_13410_));
 AND3_X1 _23103_ (.A1(_12760_),
    .A2(_11571_),
    .A3(_11569_),
    .ZN(_13411_));
 OAI21_X1 _23104_ (.A(_11567_),
    .B1(_11511_),
    .B2(_12417_),
    .ZN(_13412_));
 AND4_X1 _23105_ (.A1(_12418_),
    .A2(_13410_),
    .A3(_13411_),
    .A4(_13412_),
    .ZN(_13413_));
 NAND2_X1 _23106_ (.A1(_12396_),
    .A2(_11392_),
    .ZN(_13414_));
 NAND2_X1 _23107_ (.A1(_11454_),
    .A2(_11486_),
    .ZN(_13415_));
 OAI21_X1 _23108_ (.A(_11454_),
    .B1(_11511_),
    .B2(_11590_),
    .ZN(_13416_));
 NAND2_X1 _23109_ (.A1(_11585_),
    .A2(_11447_),
    .ZN(_13417_));
 NAND2_X1 _23110_ (.A1(_12386_),
    .A2(_11447_),
    .ZN(_13418_));
 AND4_X1 _23111_ (.A1(_13415_),
    .A2(_13416_),
    .A3(_13417_),
    .A4(_13418_),
    .ZN(_13419_));
 NAND3_X1 _23112_ (.A1(_11392_),
    .A2(_11412_),
    .A3(_11402_),
    .ZN(_13420_));
 OAI21_X1 _23113_ (.A(_11392_),
    .B1(_12430_),
    .B2(_11436_),
    .ZN(_13421_));
 AND4_X1 _23114_ (.A1(_13414_),
    .A2(_13419_),
    .A3(_13420_),
    .A4(_13421_),
    .ZN(_13422_));
 AND4_X1 _23115_ (.A1(_13400_),
    .A2(_13407_),
    .A3(_13413_),
    .A4(_13422_),
    .ZN(_13423_));
 OAI21_X1 _23116_ (.A(_11480_),
    .B1(_12396_),
    .B2(_11577_),
    .ZN(_13424_));
 OAI211_X2 _23117_ (.A(_11505_),
    .B(_16823_),
    .C1(_16822_),
    .C2(_11601_),
    .ZN(_13425_));
 OAI21_X1 _23118_ (.A(_11480_),
    .B1(_11543_),
    .B2(_11496_),
    .ZN(_13426_));
 AND4_X1 _23119_ (.A1(_11508_),
    .A2(_13424_),
    .A3(_13425_),
    .A4(_13426_),
    .ZN(_13427_));
 AND2_X1 _23120_ (.A1(_11519_),
    .A2(_11515_),
    .ZN(_13428_));
 AND2_X1 _23121_ (.A1(_11440_),
    .A2(_11515_),
    .ZN(_13429_));
 AOI211_X4 _23122_ (.A(_13428_),
    .B(_13429_),
    .C1(_11516_),
    .C2(_11561_),
    .ZN(_13430_));
 AOI21_X1 _23123_ (.A(_12926_),
    .B1(_11516_),
    .B2(_12812_),
    .ZN(_13431_));
 OAI21_X1 _23124_ (.A(_11528_),
    .B1(_12412_),
    .B2(_11561_),
    .ZN(_13432_));
 AND4_X1 _23125_ (.A1(_12779_),
    .A2(_13430_),
    .A3(_13431_),
    .A4(_13432_),
    .ZN(_13433_));
 NAND2_X1 _23126_ (.A1(_12812_),
    .A2(_12444_),
    .ZN(_13434_));
 OAI211_X2 _23127_ (.A(_13434_),
    .B(_12443_),
    .C1(_11520_),
    .C2(_12445_),
    .ZN(_13435_));
 NAND2_X1 _23128_ (.A1(_11613_),
    .A2(_11614_),
    .ZN(_13436_));
 NOR2_X1 _23129_ (.A1(_11617_),
    .A2(_11602_),
    .ZN(_13437_));
 NOR4_X1 _23130_ (.A1(_13435_),
    .A2(_13436_),
    .A3(_13437_),
    .A4(_12940_),
    .ZN(_13438_));
 AOI22_X1 _23131_ (.A1(_12458_),
    .A2(_12945_),
    .B1(_12417_),
    .B2(_12456_),
    .ZN(_13439_));
 OAI21_X1 _23132_ (.A(_12456_),
    .B1(_11441_),
    .B2(_11486_),
    .ZN(_13440_));
 OAI21_X1 _23133_ (.A(_11607_),
    .B1(_11403_),
    .B2(_12417_),
    .ZN(_13441_));
 AND4_X1 _23134_ (.A1(_12451_),
    .A2(_13439_),
    .A3(_13440_),
    .A4(_13441_),
    .ZN(_13442_));
 AND4_X1 _23135_ (.A1(_13427_),
    .A2(_13433_),
    .A3(_13438_),
    .A4(_13442_),
    .ZN(_13443_));
 NAND2_X1 _23136_ (.A1(_13423_),
    .A2(_13443_),
    .ZN(_13444_));
 XNOR2_X1 _23137_ (.A(_13392_),
    .B(_13444_),
    .ZN(_13445_));
 XNOR2_X1 _23138_ (.A(_13391_),
    .B(_13445_),
    .ZN(_13446_));
 XNOR2_X1 _23139_ (.A(_13446_),
    .B(_17266_),
    .ZN(_13447_));
 MUX2_X1 _23140_ (.A(_13204_),
    .B(_13447_),
    .S(_11149_),
    .Z(_00720_));
 XOR2_X1 _23141_ (.A(_17267_),
    .B(_17070_),
    .Z(_13448_));
 NAND2_X1 _23142_ (.A1(_12205_),
    .A2(_11732_),
    .ZN(_13449_));
 INV_X1 _23143_ (.A(_13449_),
    .ZN(_13450_));
 NOR3_X1 _23144_ (.A1(_13450_),
    .A2(_12221_),
    .A3(_12222_),
    .ZN(_13451_));
 NAND2_X1 _23145_ (.A1(_11742_),
    .A2(_11744_),
    .ZN(_13452_));
 AND2_X4 _23146_ (.A1(_11743_),
    .A2(_11869_),
    .ZN(_13453_));
 AND2_X1 _23147_ (.A1(_11743_),
    .A2(_11648_),
    .ZN(_13454_));
 AOI211_X2 _23148_ (.A(_13453_),
    .B(_13454_),
    .C1(_11645_),
    .C2(_11743_),
    .ZN(_13455_));
 AND2_X1 _23149_ (.A1(_11724_),
    .A2(_11756_),
    .ZN(_13456_));
 AOI211_X2 _23150_ (.A(_11757_),
    .B(_13456_),
    .C1(_11673_),
    .C2(_11764_),
    .ZN(_13457_));
 AND4_X2 _23151_ (.A1(_13452_),
    .A2(_13455_),
    .A3(_12628_),
    .A4(_13457_),
    .ZN(_13458_));
 OAI221_X1 _23152_ (.A(_11732_),
    .B1(_11902_),
    .B2(_11734_),
    .C1(_12605_),
    .C2(_11673_),
    .ZN(_13459_));
 AND3_X1 _23153_ (.A1(_11828_),
    .A2(_11945_),
    .A3(_11713_),
    .ZN(_13460_));
 AOI21_X1 _23154_ (.A(_11714_),
    .B1(_11896_),
    .B2(_12638_),
    .ZN(_13461_));
 AOI211_X2 _23155_ (.A(_13460_),
    .B(_13461_),
    .C1(_11727_),
    .C2(_11792_),
    .ZN(_13462_));
 AND4_X2 _23156_ (.A1(_13451_),
    .A2(_13458_),
    .A3(_13459_),
    .A4(_13462_),
    .ZN(_13463_));
 INV_X1 _23157_ (.A(_12206_),
    .ZN(_13464_));
 NAND3_X1 _23158_ (.A1(_11695_),
    .A2(_11777_),
    .A3(_11841_),
    .ZN(_13465_));
 NAND4_X1 _23159_ (.A1(_13464_),
    .A2(_13465_),
    .A3(_13109_),
    .A4(_13307_),
    .ZN(_13466_));
 OAI21_X1 _23160_ (.A(_11803_),
    .B1(_11716_),
    .B2(_11691_),
    .ZN(_13467_));
 OAI21_X1 _23161_ (.A(_11803_),
    .B1(_11722_),
    .B2(_12200_),
    .ZN(_13468_));
 NAND3_X1 _23162_ (.A1(_13467_),
    .A2(_13468_),
    .A3(_11808_),
    .ZN(_13469_));
 OAI21_X1 _23163_ (.A(_11817_),
    .B1(_11645_),
    .B2(_11724_),
    .ZN(_13470_));
 NAND3_X1 _23164_ (.A1(_11797_),
    .A2(_11762_),
    .A3(_11777_),
    .ZN(_13471_));
 NAND4_X1 _23165_ (.A1(_13470_),
    .A2(_11811_),
    .A3(_13471_),
    .A4(_13312_),
    .ZN(_13472_));
 OAI21_X1 _23166_ (.A(_11780_),
    .B1(_11659_),
    .B2(_11818_),
    .ZN(_13473_));
 NAND3_X1 _23167_ (.A1(_13473_),
    .A2(_11776_),
    .A3(_11778_),
    .ZN(_13474_));
 NOR4_X1 _23168_ (.A1(_13466_),
    .A2(_13469_),
    .A3(_13472_),
    .A4(_13474_),
    .ZN(_13475_));
 AND4_X1 _23169_ (.A1(_11672_),
    .A2(_11841_),
    .A3(_11737_),
    .A4(_11826_),
    .ZN(_13476_));
 AOI221_X4 _23170_ (.A(_13476_),
    .B1(_11838_),
    .B2(_11782_),
    .C1(_12235_),
    .C2(_11902_),
    .ZN(_13477_));
 OAI21_X1 _23171_ (.A(_12244_),
    .B1(_11805_),
    .B2(_11747_),
    .ZN(_13478_));
 NAND2_X1 _23172_ (.A1(_12244_),
    .A2(_12200_),
    .ZN(_13479_));
 NAND4_X1 _23173_ (.A1(_11735_),
    .A2(_11699_),
    .A3(_11826_),
    .A4(_12246_),
    .ZN(_13480_));
 NAND3_X1 _23174_ (.A1(_13478_),
    .A2(_13479_),
    .A3(_13480_),
    .ZN(_13481_));
 AOI21_X1 _23175_ (.A(_12590_),
    .B1(_11692_),
    .B2(_11688_),
    .ZN(_13482_));
 AND3_X1 _23176_ (.A1(_11792_),
    .A2(_12246_),
    .A3(_11826_),
    .ZN(_13483_));
 NOR4_X1 _23177_ (.A1(_13084_),
    .A2(_13481_),
    .A3(_13482_),
    .A4(_13483_),
    .ZN(_13484_));
 OAI21_X1 _23178_ (.A(_11838_),
    .B1(_12200_),
    .B2(_11749_),
    .ZN(_13485_));
 NAND2_X1 _23179_ (.A1(_11775_),
    .A2(_12620_),
    .ZN(_13486_));
 OAI211_X2 _23180_ (.A(_12620_),
    .B(_12605_),
    .C1(_11902_),
    .C2(_11734_),
    .ZN(_13487_));
 OAI21_X1 _23181_ (.A(_12620_),
    .B1(_11911_),
    .B2(_11848_),
    .ZN(_13488_));
 NAND2_X1 _23182_ (.A1(_12620_),
    .A2(_11839_),
    .ZN(_13489_));
 AND4_X1 _23183_ (.A1(_13486_),
    .A2(_13487_),
    .A3(_13488_),
    .A4(_13489_),
    .ZN(_13490_));
 AND4_X1 _23184_ (.A1(_13477_),
    .A2(_13484_),
    .A3(_13485_),
    .A4(_13490_),
    .ZN(_13491_));
 OAI21_X1 _23185_ (.A(_11880_),
    .B1(_12202_),
    .B2(_13105_),
    .ZN(_13492_));
 OAI21_X1 _23186_ (.A(_11880_),
    .B1(_11704_),
    .B2(_11782_),
    .ZN(_13493_));
 OAI211_X2 _23187_ (.A(_11880_),
    .B(_12610_),
    .C1(_11761_),
    .C2(_11699_),
    .ZN(_13494_));
 AND3_X1 _23188_ (.A1(_13492_),
    .A2(_13493_),
    .A3(_13494_),
    .ZN(_13495_));
 NOR2_X1 _23189_ (.A1(_12637_),
    .A2(_11684_),
    .ZN(_13496_));
 AND2_X1 _23190_ (.A1(_11694_),
    .A2(_11782_),
    .ZN(_13497_));
 AND4_X1 _23191_ (.A1(_11635_),
    .A2(_11841_),
    .A3(_12610_),
    .A4(_11637_),
    .ZN(_13498_));
 NOR3_X1 _23192_ (.A1(_13496_),
    .A2(_13497_),
    .A3(_13498_),
    .ZN(_13499_));
 OAI211_X2 _23193_ (.A(_12604_),
    .B(_12605_),
    .C1(_11733_),
    .C2(_11765_),
    .ZN(_13500_));
 AND4_X1 _23194_ (.A1(_11876_),
    .A2(_13500_),
    .A3(_13297_),
    .A4(_12613_),
    .ZN(_13501_));
 NAND3_X1 _23195_ (.A1(_11705_),
    .A2(_11699_),
    .A3(_11676_),
    .ZN(_13502_));
 OAI211_X2 _23196_ (.A(_11705_),
    .B(_12610_),
    .C1(_11733_),
    .C2(_11765_),
    .ZN(_13503_));
 NAND4_X1 _23197_ (.A1(_12605_),
    .A2(_11761_),
    .A3(_11635_),
    .A4(_11762_),
    .ZN(_13504_));
 AND4_X1 _23198_ (.A1(_13502_),
    .A2(_13503_),
    .A3(_11870_),
    .A4(_13504_),
    .ZN(_13505_));
 AND4_X1 _23199_ (.A1(_13495_),
    .A2(_13499_),
    .A3(_13501_),
    .A4(_13505_),
    .ZN(_13506_));
 NAND4_X1 _23200_ (.A1(_13463_),
    .A2(_13475_),
    .A3(_13491_),
    .A4(_13506_),
    .ZN(_13507_));
 NOR2_X2 _23201_ (.A1(_13507_),
    .A2(_11856_),
    .ZN(_13508_));
 AND2_X1 _23202_ (.A1(_11282_),
    .A2(_11275_),
    .ZN(_13509_));
 AOI21_X1 _23203_ (.A(_11276_),
    .B1(_12316_),
    .B2(_11251_),
    .ZN(_13510_));
 AND4_X1 _23204_ (.A1(_11321_),
    .A2(_11153_),
    .A3(_11258_),
    .A4(_11297_),
    .ZN(_13511_));
 OR4_X4 _23205_ (.A1(_13509_),
    .A2(_13510_),
    .A3(_12680_),
    .A4(_13511_),
    .ZN(_13512_));
 AOI221_X1 _23206_ (.A(_11243_),
    .B1(_11178_),
    .B2(_11260_),
    .C1(_12275_),
    .C2(_11351_),
    .ZN(_13513_));
 OR3_X1 _23207_ (.A1(_13513_),
    .A2(_12692_),
    .A3(_12321_),
    .ZN(_13514_));
 AOI21_X1 _23208_ (.A(_11290_),
    .B1(_11291_),
    .B2(_11280_),
    .ZN(_13515_));
 AND2_X4 _23209_ (.A1(_11184_),
    .A2(_11293_),
    .ZN(_13516_));
 AND4_X1 _23210_ (.A1(_11297_),
    .A2(_11217_),
    .A3(_11322_),
    .A4(_11169_),
    .ZN(_13517_));
 OR3_X1 _23211_ (.A1(_13515_),
    .A2(_13516_),
    .A3(_13517_),
    .ZN(_13518_));
 OAI21_X1 _23212_ (.A(_11265_),
    .B1(_12663_),
    .B2(_11352_),
    .ZN(_13519_));
 NAND2_X1 _23213_ (.A1(_12302_),
    .A2(_11227_),
    .ZN(_13520_));
 NAND2_X1 _23214_ (.A1(_13520_),
    .A2(_11263_),
    .ZN(_13521_));
 NAND3_X1 _23215_ (.A1(_13519_),
    .A2(_13358_),
    .A3(_13521_),
    .ZN(_13522_));
 NOR4_X4 _23216_ (.A1(_13512_),
    .A2(_13514_),
    .A3(_13518_),
    .A4(_13522_),
    .ZN(_13523_));
 OAI21_X1 _23217_ (.A(_12683_),
    .B1(_12282_),
    .B2(_12343_),
    .ZN(_13524_));
 OAI21_X1 _23218_ (.A(_12683_),
    .B1(_11270_),
    .B2(_11379_),
    .ZN(_13525_));
 AND3_X1 _23219_ (.A1(_13524_),
    .A2(_13525_),
    .A3(_13048_),
    .ZN(_13526_));
 AND3_X1 _23220_ (.A1(_11364_),
    .A2(_11332_),
    .A3(_11167_),
    .ZN(_13527_));
 NOR4_X1 _23221_ (.A1(_12293_),
    .A2(_13337_),
    .A3(_13338_),
    .A4(_13527_),
    .ZN(_13528_));
 AOI21_X1 _23222_ (.A(_11224_),
    .B1(_11346_),
    .B2(_12268_),
    .ZN(_13529_));
 NOR2_X1 _23223_ (.A1(_13529_),
    .A2(_11236_),
    .ZN(_13530_));
 NAND3_X1 _23224_ (.A1(_12308_),
    .A2(_11199_),
    .A3(_11257_),
    .ZN(_13531_));
 OAI211_X2 _23225_ (.A(_11199_),
    .B(_11232_),
    .C1(_11178_),
    .C2(_11233_),
    .ZN(_13532_));
 NAND2_X1 _23226_ (.A1(_12350_),
    .A2(_11199_),
    .ZN(_13533_));
 AND4_X1 _23227_ (.A1(_13531_),
    .A2(_13532_),
    .A3(_13533_),
    .A4(_13342_),
    .ZN(_13534_));
 AND4_X1 _23228_ (.A1(_13526_),
    .A2(_13528_),
    .A3(_13530_),
    .A4(_13534_),
    .ZN(_13535_));
 OAI21_X1 _23229_ (.A(_11315_),
    .B1(_12304_),
    .B2(_11286_),
    .ZN(_13536_));
 NAND2_X1 _23230_ (.A1(_12704_),
    .A2(_11328_),
    .ZN(_13537_));
 NAND2_X1 _23231_ (.A1(_11315_),
    .A2(_11174_),
    .ZN(_13538_));
 OAI21_X1 _23232_ (.A(_11328_),
    .B1(_12343_),
    .B2(_11310_),
    .ZN(_13539_));
 NAND4_X1 _23233_ (.A1(_13536_),
    .A2(_13537_),
    .A3(_13538_),
    .A4(_13539_),
    .ZN(_13540_));
 NAND4_X1 _23234_ (.A1(_11332_),
    .A2(_11320_),
    .A3(_11164_),
    .A4(_11217_),
    .ZN(_13541_));
 OAI221_X1 _23235_ (.A(_13541_),
    .B1(_11337_),
    .B2(_11180_),
    .C1(_11233_),
    .C2(_12352_),
    .ZN(_13542_));
 AOI21_X1 _23236_ (.A(_11337_),
    .B1(_11251_),
    .B2(_11280_),
    .ZN(_13543_));
 OAI21_X1 _23237_ (.A(_11309_),
    .B1(_11270_),
    .B2(_11379_),
    .ZN(_13544_));
 OAI21_X1 _23238_ (.A(_11309_),
    .B1(_11190_),
    .B2(_11230_),
    .ZN(_13545_));
 NAND2_X1 _23239_ (.A1(_11309_),
    .A2(_12301_),
    .ZN(_13546_));
 NAND4_X1 _23240_ (.A1(_13544_),
    .A2(_13545_),
    .A3(_11311_),
    .A4(_13546_),
    .ZN(_13547_));
 NOR4_X1 _23241_ (.A1(_13540_),
    .A2(_13542_),
    .A3(_13543_),
    .A4(_13547_),
    .ZN(_13548_));
 AND3_X1 _23242_ (.A1(_11267_),
    .A2(_11326_),
    .A3(_11341_),
    .ZN(_13549_));
 AOI21_X1 _23243_ (.A(_13008_),
    .B1(_12316_),
    .B2(_11185_),
    .ZN(_13550_));
 AND2_X2 _23244_ (.A1(_12282_),
    .A2(_11343_),
    .ZN(_13551_));
 OR4_X4 _23245_ (.A1(_13549_),
    .A2(_13550_),
    .A3(_13383_),
    .A4(_13551_),
    .ZN(_13552_));
 AND2_X1 _23246_ (.A1(_12350_),
    .A2(_11375_),
    .ZN(_13553_));
 NAND2_X1 _23247_ (.A1(_11373_),
    .A2(_13039_),
    .ZN(_13554_));
 OAI21_X1 _23248_ (.A(_13554_),
    .B1(_12285_),
    .B2(_12279_),
    .ZN(_13555_));
 AND3_X1 _23249_ (.A1(_11373_),
    .A2(_11172_),
    .A3(_12265_),
    .ZN(_13556_));
 OR4_X2 _23250_ (.A1(_13553_),
    .A2(_13555_),
    .A3(_12284_),
    .A4(_13556_),
    .ZN(_13557_));
 OAI21_X1 _23251_ (.A(_11363_),
    .B1(_11184_),
    .B2(_11190_),
    .ZN(_13558_));
 NAND2_X1 _23252_ (.A1(_11353_),
    .A2(_12327_),
    .ZN(_13559_));
 NAND4_X1 _23253_ (.A1(_11332_),
    .A2(_11164_),
    .A3(_11269_),
    .A4(_11341_),
    .ZN(_13560_));
 NAND3_X1 _23254_ (.A1(_13558_),
    .A2(_13559_),
    .A3(_13560_),
    .ZN(_13561_));
 OAI21_X1 _23255_ (.A(_11371_),
    .B1(_11196_),
    .B2(_13032_),
    .ZN(_13562_));
 OAI21_X1 _23256_ (.A(_11371_),
    .B1(_11267_),
    .B2(_12327_),
    .ZN(_13563_));
 NAND4_X1 _23257_ (.A1(_11371_),
    .A2(_11257_),
    .A3(_11260_),
    .A4(_11164_),
    .ZN(_13564_));
 NAND3_X1 _23258_ (.A1(_13562_),
    .A2(_13563_),
    .A3(_13564_),
    .ZN(_13565_));
 NOR4_X2 _23259_ (.A1(_13552_),
    .A2(_13557_),
    .A3(_13561_),
    .A4(_13565_),
    .ZN(_13566_));
 NAND4_X1 _23260_ (.A1(_13523_),
    .A2(_13535_),
    .A3(_13548_),
    .A4(_13566_),
    .ZN(_13567_));
 NOR2_X2 _23261_ (.A1(_13567_),
    .A2(_11386_),
    .ZN(_13568_));
 XNOR2_X2 _23262_ (.A(_13508_),
    .B(_13568_),
    .ZN(_13569_));
 OAI21_X1 _23263_ (.A(_12167_),
    .B1(_12005_),
    .B2(_12122_),
    .ZN(_13570_));
 AND2_X1 _23264_ (.A1(_11973_),
    .A2(_12161_),
    .ZN(_13571_));
 AND2_X1 _23265_ (.A1(_12039_),
    .A2(_12161_),
    .ZN(_13572_));
 AOI211_X2 _23266_ (.A(_13571_),
    .B(_13572_),
    .C1(_12162_),
    .C2(_12093_),
    .ZN(_13573_));
 OAI211_X2 _23267_ (.A(_12167_),
    .B(_12491_),
    .C1(_11990_),
    .C2(_12528_),
    .ZN(_13574_));
 OAI21_X1 _23268_ (.A(_12167_),
    .B1(_12119_),
    .B2(_12493_),
    .ZN(_13575_));
 AND4_X1 _23269_ (.A1(_13570_),
    .A2(_13573_),
    .A3(_13574_),
    .A4(_13575_),
    .ZN(_13576_));
 NAND2_X1 _23270_ (.A1(_12052_),
    .A2(_12527_),
    .ZN(_13577_));
 NAND2_X1 _23271_ (.A1(_12834_),
    .A2(_12108_),
    .ZN(_13578_));
 OAI211_X2 _23272_ (.A(_12527_),
    .B(_11999_),
    .C1(_12089_),
    .C2(_12000_),
    .ZN(_13579_));
 NAND4_X1 _23273_ (.A1(_13577_),
    .A2(_13247_),
    .A3(_13578_),
    .A4(_13579_),
    .ZN(_13580_));
 AND2_X1 _23274_ (.A1(_12100_),
    .A2(_12544_),
    .ZN(_13581_));
 OR2_X1 _23275_ (.A1(_12099_),
    .A2(_13581_),
    .ZN(_13582_));
 NAND2_X1 _23276_ (.A1(_12544_),
    .A2(_12479_),
    .ZN(_13583_));
 OAI22_X1 _23277_ (.A1(_13583_),
    .A2(_11970_),
    .B1(_12549_),
    .B2(_12092_),
    .ZN(_13584_));
 NOR4_X1 _23278_ (.A1(_13580_),
    .A2(_13582_),
    .A3(_12101_),
    .A4(_13584_),
    .ZN(_13585_));
 OAI211_X2 _23279_ (.A(_12146_),
    .B(_12531_),
    .C1(_12143_),
    .C2(_12535_),
    .ZN(_13586_));
 AOI21_X1 _23280_ (.A(_12143_),
    .B1(_12155_),
    .B2(_12840_),
    .ZN(_13587_));
 AOI21_X1 _23281_ (.A(_12151_),
    .B1(_12049_),
    .B2(_12877_),
    .ZN(_13588_));
 NOR4_X1 _23282_ (.A1(_13586_),
    .A2(_13587_),
    .A3(_13588_),
    .A4(_12885_),
    .ZN(_13589_));
 AND2_X1 _23283_ (.A1(_12122_),
    .A2(_12830_),
    .ZN(_13590_));
 INV_X1 _23284_ (.A(_13590_),
    .ZN(_13591_));
 NAND2_X1 _23285_ (.A1(_12117_),
    .A2(_12039_),
    .ZN(_13592_));
 OAI21_X1 _23286_ (.A(_12117_),
    .B1(_12109_),
    .B2(_12044_),
    .ZN(_13593_));
 OAI21_X1 _23287_ (.A(_12117_),
    .B1(_12082_),
    .B2(_12068_),
    .ZN(_13594_));
 NAND2_X1 _23288_ (.A1(_12117_),
    .A2(_13164_),
    .ZN(_13595_));
 AND4_X1 _23289_ (.A1(_13592_),
    .A2(_13593_),
    .A3(_13594_),
    .A4(_13595_),
    .ZN(_13596_));
 OAI21_X1 _23290_ (.A(_12830_),
    .B1(_12490_),
    .B2(_12128_),
    .ZN(_13597_));
 AND4_X1 _23291_ (.A1(_13591_),
    .A2(_13596_),
    .A3(_13167_),
    .A4(_13597_),
    .ZN(_13598_));
 NAND4_X1 _23292_ (.A1(_13576_),
    .A2(_13585_),
    .A3(_13589_),
    .A4(_13598_),
    .ZN(_13599_));
 AND2_X1 _23293_ (.A1(_12495_),
    .A2(_12497_),
    .ZN(_13600_));
 NAND3_X1 _23294_ (.A1(_11997_),
    .A2(_12026_),
    .A3(_12496_),
    .ZN(_13601_));
 AND3_X1 _23295_ (.A1(_13212_),
    .A2(_12836_),
    .A3(_13601_),
    .ZN(_13602_));
 OAI21_X1 _23296_ (.A(_12487_),
    .B1(_12019_),
    .B2(_11997_),
    .ZN(_13603_));
 OAI21_X1 _23297_ (.A(_12487_),
    .B1(_12066_),
    .B2(_12168_),
    .ZN(_13604_));
 AND4_X1 _23298_ (.A1(_13600_),
    .A2(_13602_),
    .A3(_13603_),
    .A4(_13604_),
    .ZN(_13605_));
 OAI21_X1 _23299_ (.A(_12860_),
    .B1(_12490_),
    .B2(_12552_),
    .ZN(_13606_));
 OAI211_X2 _23300_ (.A(_13132_),
    .B(_16863_),
    .C1(_16862_),
    .C2(_11981_),
    .ZN(_13607_));
 OAI21_X1 _23301_ (.A(_12860_),
    .B1(_12075_),
    .B2(_12156_),
    .ZN(_13608_));
 AND4_X1 _23302_ (.A1(_12573_),
    .A2(_13606_),
    .A3(_13607_),
    .A4(_13608_),
    .ZN(_13609_));
 NAND2_X1 _23303_ (.A1(_13144_),
    .A2(_12015_),
    .ZN(_13610_));
 NAND3_X1 _23304_ (.A1(_11998_),
    .A2(_12003_),
    .A3(_13610_),
    .ZN(_13611_));
 NAND2_X1 _23305_ (.A1(_13144_),
    .A2(_12039_),
    .ZN(_13612_));
 OAI211_X2 _23306_ (.A(_13612_),
    .B(_13234_),
    .C1(_12566_),
    .C2(_12155_),
    .ZN(_13613_));
 AOI21_X1 _23307_ (.A(_12850_),
    .B1(_12877_),
    .B2(_12535_),
    .ZN(_13614_));
 NOR4_X1 _23308_ (.A1(_13611_),
    .A2(_13613_),
    .A3(_13151_),
    .A4(_13614_),
    .ZN(_13615_));
 AOI22_X1 _23309_ (.A1(_12898_),
    .A2(_12532_),
    .B1(_12163_),
    .B2(_12062_),
    .ZN(_13616_));
 OAI21_X1 _23310_ (.A(_12056_),
    .B1(_12543_),
    .B2(_12163_),
    .ZN(_13617_));
 OAI21_X1 _23311_ (.A(_12062_),
    .B1(_12834_),
    .B2(_13164_),
    .ZN(_13618_));
 AND4_X1 _23312_ (.A1(_12870_),
    .A2(_13616_),
    .A3(_13617_),
    .A4(_13618_),
    .ZN(_13619_));
 NAND4_X1 _23313_ (.A1(_13605_),
    .A2(_13609_),
    .A3(_13615_),
    .A4(_13619_),
    .ZN(_13620_));
 NOR2_X4 _23314_ (.A1(_13599_),
    .A2(_13620_),
    .ZN(_13621_));
 XOR2_X1 _23315_ (.A(_13569_),
    .B(_13621_),
    .Z(_13622_));
 AND2_X1 _23316_ (.A1(_11454_),
    .A2(_11436_),
    .ZN(_13623_));
 OAI21_X1 _23317_ (.A(_13415_),
    .B1(_13417_),
    .B2(_11601_),
    .ZN(_13624_));
 AND3_X1 _23318_ (.A1(_11403_),
    .A2(_11447_),
    .A3(_11407_),
    .ZN(_13625_));
 OR4_X2 _23319_ (.A1(_13623_),
    .A2(_13624_),
    .A3(_12410_),
    .A4(_13625_),
    .ZN(_13626_));
 AND2_X1 _23320_ (.A1(_11519_),
    .A2(_11442_),
    .ZN(_13627_));
 NOR4_X1 _23321_ (.A1(_13403_),
    .A2(_13627_),
    .A3(_12389_),
    .A4(_11431_),
    .ZN(_13628_));
 OAI21_X1 _23322_ (.A(_12392_),
    .B1(_11420_),
    .B2(_12972_),
    .ZN(_13629_));
 NAND4_X1 _23323_ (.A1(_13628_),
    .A2(_12395_),
    .A3(_12798_),
    .A4(_13629_),
    .ZN(_13630_));
 OAI211_X2 _23324_ (.A(_12399_),
    .B(_13414_),
    .C1(_12400_),
    .C2(_11455_),
    .ZN(_13631_));
 AOI221_X4 _23325_ (.A(_12400_),
    .B1(_11467_),
    .B2(_11415_),
    .C1(_11493_),
    .C2(_11400_),
    .ZN(_13632_));
 NOR4_X1 _23326_ (.A1(_13626_),
    .A2(_13630_),
    .A3(_13631_),
    .A4(_13632_),
    .ZN(_13633_));
 AND2_X1 _23327_ (.A1(_11441_),
    .A2(_11564_),
    .ZN(_13634_));
 AOI211_X4 _23328_ (.A(_11565_),
    .B(_13634_),
    .C1(_11567_),
    .C2(_11482_),
    .ZN(_13635_));
 OAI21_X1 _23329_ (.A(_11567_),
    .B1(_11436_),
    .B2(_12417_),
    .ZN(_13636_));
 NAND2_X1 _23330_ (.A1(_13635_),
    .A2(_13636_),
    .ZN(_13637_));
 NAND2_X1 _23331_ (.A1(_11519_),
    .A2(_11555_),
    .ZN(_13638_));
 NAND4_X1 _23332_ (.A1(_11412_),
    .A2(_11537_),
    .A3(_11415_),
    .A4(_11552_),
    .ZN(_13639_));
 NAND4_X1 _23333_ (.A1(_11557_),
    .A2(_11558_),
    .A3(_13638_),
    .A4(_13639_),
    .ZN(_13640_));
 INV_X1 _23334_ (.A(_12422_),
    .ZN(_13641_));
 NAND2_X1 _23335_ (.A1(_11546_),
    .A2(_11496_),
    .ZN(_13642_));
 NAND4_X1 _23336_ (.A1(_13641_),
    .A2(_12959_),
    .A3(_13394_),
    .A4(_13642_),
    .ZN(_13643_));
 OAI211_X2 _23337_ (.A(_11574_),
    .B(_11420_),
    .C1(_11467_),
    .C2(_11415_),
    .ZN(_13644_));
 NAND3_X1 _23338_ (.A1(_11403_),
    .A2(_11574_),
    .A3(_11407_),
    .ZN(_13645_));
 NAND2_X1 _23339_ (.A1(_11500_),
    .A2(_11574_),
    .ZN(_13646_));
 NAND2_X1 _23340_ (.A1(_11570_),
    .A2(_11574_),
    .ZN(_13647_));
 NAND4_X1 _23341_ (.A1(_13644_),
    .A2(_13645_),
    .A3(_13646_),
    .A4(_13647_),
    .ZN(_13648_));
 NOR4_X1 _23342_ (.A1(_13637_),
    .A2(_13640_),
    .A3(_13643_),
    .A4(_13648_),
    .ZN(_13649_));
 AND2_X1 _23343_ (.A1(_11548_),
    .A2(_11505_),
    .ZN(_13650_));
 INV_X1 _23344_ (.A(_13650_),
    .ZN(_13651_));
 OAI21_X1 _23345_ (.A(_11505_),
    .B1(_12371_),
    .B2(_12972_),
    .ZN(_13652_));
 NAND4_X1 _23346_ (.A1(_11504_),
    .A2(_13651_),
    .A3(_12369_),
    .A4(_13652_),
    .ZN(_13653_));
 INV_X1 _23347_ (.A(_13429_),
    .ZN(_13654_));
 NAND2_X1 _23348_ (.A1(_11543_),
    .A2(_11516_),
    .ZN(_13655_));
 OAI21_X1 _23349_ (.A(_11516_),
    .B1(_11396_),
    .B2(_11561_),
    .ZN(_13656_));
 NAND4_X1 _23350_ (.A1(_13654_),
    .A2(_13655_),
    .A3(_12925_),
    .A4(_13656_),
    .ZN(_13657_));
 AND2_X1 _23351_ (.A1(_11419_),
    .A2(_11456_),
    .ZN(_13658_));
 OAI21_X1 _23352_ (.A(_11528_),
    .B1(_12741_),
    .B2(_13658_),
    .ZN(_13659_));
 NAND4_X1 _23353_ (.A1(_11528_),
    .A2(_11412_),
    .A3(_11407_),
    .A4(_11426_),
    .ZN(_13660_));
 NAND4_X1 _23354_ (.A1(_12921_),
    .A2(_13659_),
    .A3(_12763_),
    .A4(_13660_),
    .ZN(_13661_));
 OAI21_X1 _23355_ (.A(_11480_),
    .B1(_11450_),
    .B2(_11511_),
    .ZN(_13662_));
 NAND2_X1 _23356_ (.A1(_11480_),
    .A2(_11507_),
    .ZN(_13663_));
 INV_X1 _23357_ (.A(_11561_),
    .ZN(_13664_));
 OAI211_X2 _23358_ (.A(_13662_),
    .B(_13663_),
    .C1(_11485_),
    .C2(_13664_),
    .ZN(_13665_));
 NOR4_X1 _23359_ (.A1(_13653_),
    .A2(_13657_),
    .A3(_13661_),
    .A4(_13665_),
    .ZN(_13666_));
 AOI211_X2 _23360_ (.A(_11594_),
    .B(_11595_),
    .C1(_11548_),
    .C2(_12444_),
    .ZN(_13667_));
 INV_X1 _23361_ (.A(_12752_),
    .ZN(_13668_));
 OAI21_X1 _23362_ (.A(_12444_),
    .B1(_11436_),
    .B2(_12417_),
    .ZN(_13669_));
 OAI21_X1 _23363_ (.A(_12444_),
    .B1(_12741_),
    .B2(_11590_),
    .ZN(_13670_));
 NAND4_X1 _23364_ (.A1(_13667_),
    .A2(_13668_),
    .A3(_13669_),
    .A4(_13670_),
    .ZN(_13671_));
 AND3_X1 _23365_ (.A1(_11488_),
    .A2(_11445_),
    .A3(_11592_),
    .ZN(_13672_));
 OR3_X1 _23366_ (.A1(_12934_),
    .A2(_12459_),
    .A3(_13672_),
    .ZN(_13673_));
 AND3_X1 _23367_ (.A1(_11606_),
    .A2(_12393_),
    .A3(_12430_),
    .ZN(_13674_));
 AND4_X1 _23368_ (.A1(_11601_),
    .A2(_11592_),
    .A3(_11552_),
    .A4(_11420_),
    .ZN(_13675_));
 NOR3_X1 _23369_ (.A1(_13674_),
    .A2(_12758_),
    .A3(_13675_),
    .ZN(_13676_));
 OAI21_X1 _23370_ (.A(_13676_),
    .B1(_11487_),
    .B2(_11610_),
    .ZN(_13677_));
 OAI211_X2 _23371_ (.A(_12463_),
    .B(_11599_),
    .C1(_11467_),
    .C2(_11529_),
    .ZN(_13678_));
 NAND2_X1 _23372_ (.A1(_12463_),
    .A2(_11441_),
    .ZN(_13679_));
 OAI21_X1 _23373_ (.A(_12463_),
    .B1(_12371_),
    .B2(_11450_),
    .ZN(_13680_));
 NAND2_X1 _23374_ (.A1(_12463_),
    .A2(_12367_),
    .ZN(_13681_));
 NAND4_X1 _23375_ (.A1(_13678_),
    .A2(_13679_),
    .A3(_13680_),
    .A4(_13681_),
    .ZN(_13682_));
 NOR4_X1 _23376_ (.A1(_13671_),
    .A2(_13673_),
    .A3(_13677_),
    .A4(_13682_),
    .ZN(_13683_));
 NAND4_X1 _23377_ (.A1(_13633_),
    .A2(_13649_),
    .A3(_13666_),
    .A4(_13683_),
    .ZN(_13684_));
 NOR2_X2 _23378_ (.A1(_13684_),
    .A2(_11623_),
    .ZN(_13685_));
 XOR2_X1 _23379_ (.A(_13332_),
    .B(_13685_),
    .Z(_13686_));
 XNOR2_X1 _23380_ (.A(_13622_),
    .B(_13686_),
    .ZN(_13687_));
 XNOR2_X1 _23381_ (.A(_13687_),
    .B(_17267_),
    .ZN(_13688_));
 MUX2_X1 _23382_ (.A(_13448_),
    .B(_13688_),
    .S(_11149_),
    .Z(_00721_));
 XOR2_X1 _23383_ (.A(_17268_),
    .B(_17071_),
    .Z(_13689_));
 AND4_X1 _23384_ (.A1(_11394_),
    .A2(_11586_),
    .A3(_11405_),
    .A4(_11591_),
    .ZN(_13690_));
 AND2_X2 _23385_ (.A1(_11587_),
    .A2(_11560_),
    .ZN(_13691_));
 AOI211_X2 _23386_ (.A(_13690_),
    .B(_13691_),
    .C1(_11461_),
    .C2(_11587_),
    .ZN(_13692_));
 OAI21_X1 _23387_ (.A(_12444_),
    .B1(_11543_),
    .B2(_12417_),
    .ZN(_13693_));
 AND3_X1 _23388_ (.A1(_13692_),
    .A2(_13670_),
    .A3(_13693_),
    .ZN(_13694_));
 OAI21_X1 _23389_ (.A(_11516_),
    .B1(_11490_),
    .B2(_12412_),
    .ZN(_13695_));
 OAI21_X1 _23390_ (.A(_11516_),
    .B1(_12741_),
    .B2(_13658_),
    .ZN(_13696_));
 INV_X1 _23391_ (.A(_12815_),
    .ZN(_13697_));
 NOR4_X1 _23392_ (.A1(_13697_),
    .A2(_12967_),
    .A3(_11623_),
    .A4(_12432_),
    .ZN(_13698_));
 AND4_X1 _23393_ (.A1(_13694_),
    .A2(_13695_),
    .A3(_13696_),
    .A4(_13698_),
    .ZN(_13699_));
 NAND4_X1 _23394_ (.A1(_12465_),
    .A2(_12956_),
    .A3(_12467_),
    .A4(_12755_),
    .ZN(_13700_));
 AND2_X1 _23395_ (.A1(_12463_),
    .A2(_11488_),
    .ZN(_13701_));
 AND2_X2 _23396_ (.A1(_11446_),
    .A2(_11433_),
    .ZN(_13702_));
 OR3_X1 _23397_ (.A1(_13701_),
    .A2(_13702_),
    .A3(_13672_),
    .ZN(_13703_));
 NOR3_X1 _23398_ (.A1(_13700_),
    .A2(_13703_),
    .A3(_12436_),
    .ZN(_13704_));
 OAI22_X1 _23399_ (.A1(_11485_),
    .A2(_11451_),
    .B1(_12372_),
    .B2(_12746_),
    .ZN(_13705_));
 AND2_X1 _23400_ (.A1(_11544_),
    .A2(_11590_),
    .ZN(_13706_));
 AND2_X1 _23401_ (.A1(_11548_),
    .A2(_11573_),
    .ZN(_13707_));
 OR4_X2 _23402_ (.A1(_13650_),
    .A2(_13705_),
    .A3(_13706_),
    .A4(_13707_),
    .ZN(_13708_));
 OAI221_X1 _23403_ (.A(_11566_),
    .B1(_12427_),
    .B2(_13664_),
    .C1(_12959_),
    .C2(_11413_),
    .ZN(_13709_));
 OAI21_X1 _23404_ (.A(_11607_),
    .B1(_12412_),
    .B2(_13658_),
    .ZN(_13710_));
 NAND2_X1 _23405_ (.A1(_12456_),
    .A2(_11556_),
    .ZN(_13711_));
 NAND4_X1 _23406_ (.A1(_11592_),
    .A2(_11405_),
    .A3(_11445_),
    .A4(_11399_),
    .ZN(_13712_));
 NAND4_X1 _23407_ (.A1(_13710_),
    .A2(_13711_),
    .A3(_13417_),
    .A4(_13712_),
    .ZN(_13713_));
 NOR4_X2 _23408_ (.A1(_13708_),
    .A2(_12738_),
    .A3(_13709_),
    .A4(_13713_),
    .ZN(_13714_));
 NAND2_X1 _23409_ (.A1(_11461_),
    .A2(_11555_),
    .ZN(_13715_));
 NAND2_X1 _23410_ (.A1(_11442_),
    .A2(_12379_),
    .ZN(_13716_));
 NAND4_X1 _23411_ (.A1(_13715_),
    .A2(_11484_),
    .A3(_13716_),
    .A4(_11547_),
    .ZN(_13717_));
 AND2_X1 _23412_ (.A1(_11607_),
    .A2(_11556_),
    .ZN(_13718_));
 NOR4_X1 _23413_ (.A1(_13717_),
    .A2(_12819_),
    .A3(_12751_),
    .A4(_13718_),
    .ZN(_13719_));
 NAND4_X2 _23414_ (.A1(_13699_),
    .A2(_13704_),
    .A3(_13714_),
    .A4(_13719_),
    .ZN(_13720_));
 AND3_X1 _23415_ (.A1(_11447_),
    .A2(_12412_),
    .A3(_11413_),
    .ZN(_13721_));
 OAI21_X1 _23416_ (.A(_13418_),
    .B1(_12372_),
    .B2(_11523_),
    .ZN(_13722_));
 AOI211_X2 _23417_ (.A(_13721_),
    .B(_13722_),
    .C1(_11529_),
    .C2(_11431_),
    .ZN(_13723_));
 AOI221_X1 _23418_ (.A(_12363_),
    .B1(_11486_),
    .B2(_11544_),
    .C1(_11434_),
    .C2(_11606_),
    .ZN(_13724_));
 AOI22_X1 _23419_ (.A1(_12392_),
    .A2(_12417_),
    .B1(_11434_),
    .B2(_11442_),
    .ZN(_13725_));
 AOI22_X1 _23420_ (.A1(_11500_),
    .A2(_12392_),
    .B1(_12741_),
    .B2(_11555_),
    .ZN(_13726_));
 AND4_X1 _23421_ (.A1(_13723_),
    .A2(_13724_),
    .A3(_13725_),
    .A4(_13726_),
    .ZN(_13727_));
 AOI221_X4 _23422_ (.A(_12389_),
    .B1(_11454_),
    .B2(_11511_),
    .C1(_11461_),
    .C2(_11505_),
    .ZN(_13728_));
 OR2_X1 _23423_ (.A1(_12400_),
    .A2(_11621_),
    .ZN(_13729_));
 OAI21_X1 _23424_ (.A(_13681_),
    .B1(_12423_),
    .B2(_13664_),
    .ZN(_13730_));
 AND2_X1 _23425_ (.A1(_11465_),
    .A2(_11556_),
    .ZN(_13731_));
 AND2_X1 _23426_ (.A1(_11479_),
    .A2(_11561_),
    .ZN(_13732_));
 AND2_X1 _23427_ (.A1(_11554_),
    .A2(_13658_),
    .ZN(_13733_));
 NOR4_X1 _23428_ (.A1(_13730_),
    .A2(_13731_),
    .A3(_13732_),
    .A4(_13733_),
    .ZN(_13734_));
 OAI21_X1 _23429_ (.A(_11528_),
    .B1(_11500_),
    .B2(_11548_),
    .ZN(_13735_));
 NAND3_X1 _23430_ (.A1(_11607_),
    .A2(_12393_),
    .A3(_12787_),
    .ZN(_13736_));
 AND4_X1 _23431_ (.A1(_13729_),
    .A2(_13734_),
    .A3(_13735_),
    .A4(_13736_),
    .ZN(_13737_));
 OR2_X1 _23432_ (.A1(_12746_),
    .A2(_11611_),
    .ZN(_13738_));
 OAI21_X1 _23433_ (.A(_11505_),
    .B1(_11436_),
    .B2(_12741_),
    .ZN(_13739_));
 AOI22_X1 _23434_ (.A1(_11543_),
    .A2(_11528_),
    .B1(_11567_),
    .B2(_11577_),
    .ZN(_13740_));
 AND4_X1 _23435_ (.A1(_13738_),
    .A2(_12941_),
    .A3(_13739_),
    .A4(_13740_),
    .ZN(_13741_));
 NAND4_X2 _23436_ (.A1(_13727_),
    .A2(_13728_),
    .A3(_13737_),
    .A4(_13741_),
    .ZN(_13742_));
 NOR2_X4 _23437_ (.A1(_13720_),
    .A2(_13742_),
    .ZN(_13743_));
 XNOR2_X1 _23438_ (.A(_13508_),
    .B(_13743_),
    .ZN(_13744_));
 AND4_X1 _23439_ (.A1(_11321_),
    .A2(_11167_),
    .A3(_11322_),
    .A4(_11298_),
    .ZN(_13745_));
 AOI21_X1 _23440_ (.A(_13745_),
    .B1(_12301_),
    .B2(_11199_),
    .ZN(_13746_));
 AND2_X1 _23441_ (.A1(_13520_),
    .A2(_11336_),
    .ZN(_13747_));
 AOI21_X1 _23442_ (.A(_12295_),
    .B1(_11278_),
    .B2(_11361_),
    .ZN(_13748_));
 NAND2_X1 _23443_ (.A1(_12717_),
    .A2(_13047_),
    .ZN(_13749_));
 NOR4_X1 _23444_ (.A1(_13747_),
    .A2(_13748_),
    .A3(_13749_),
    .A4(_13336_),
    .ZN(_13750_));
 OAI21_X1 _23445_ (.A(_11315_),
    .B1(_12297_),
    .B2(_13032_),
    .ZN(_13751_));
 AOI221_X1 _23446_ (.A(_13367_),
    .B1(_11336_),
    .B2(_11310_),
    .C1(_11363_),
    .C2(_12327_),
    .ZN(_13752_));
 AND4_X1 _23447_ (.A1(_13746_),
    .A2(_13750_),
    .A3(_13751_),
    .A4(_13752_),
    .ZN(_13753_));
 AOI21_X1 _23448_ (.A(_12271_),
    .B1(_11207_),
    .B2(_11315_),
    .ZN(_13754_));
 AND3_X1 _23449_ (.A1(_13754_),
    .A2(_12309_),
    .A3(_12348_),
    .ZN(_13755_));
 OAI21_X1 _23450_ (.A(_12299_),
    .B1(_11185_),
    .B2(_11290_),
    .ZN(_13756_));
 AOI221_X4 _23451_ (.A(_13756_),
    .B1(_11378_),
    .B2(_11328_),
    .C1(_12683_),
    .C2(_11218_),
    .ZN(_13757_));
 OAI22_X1 _23452_ (.A1(_11355_),
    .A2(_11361_),
    .B1(_11243_),
    .B2(_11357_),
    .ZN(_13758_));
 AOI221_X4 _23453_ (.A(_13758_),
    .B1(_11207_),
    .B2(_11293_),
    .C1(_11238_),
    .C2(_11157_),
    .ZN(_13759_));
 AND2_X1 _23454_ (.A1(_11274_),
    .A2(_11214_),
    .ZN(_13760_));
 AND2_X1 _23455_ (.A1(_11363_),
    .A2(_12276_),
    .ZN(_13761_));
 NOR3_X1 _23456_ (.A1(_12689_),
    .A2(_13760_),
    .A3(_13761_),
    .ZN(_13762_));
 AND4_X1 _23457_ (.A1(_13755_),
    .A2(_13757_),
    .A3(_13759_),
    .A4(_13762_),
    .ZN(_13763_));
 AND3_X1 _23458_ (.A1(_11315_),
    .A2(_12314_),
    .A3(_11348_),
    .ZN(_13764_));
 AND2_X1 _23459_ (.A1(_11289_),
    .A2(_11160_),
    .ZN(_13765_));
 NOR2_X1 _23460_ (.A1(_13764_),
    .A2(_13765_),
    .ZN(_13766_));
 OAI21_X1 _23461_ (.A(_11265_),
    .B1(_11214_),
    .B2(_12343_),
    .ZN(_13767_));
 OAI21_X1 _23462_ (.A(_11265_),
    .B1(_11248_),
    .B2(_11316_),
    .ZN(_13768_));
 AND3_X1 _23463_ (.A1(_13767_),
    .A2(_13768_),
    .A3(_13029_),
    .ZN(_13769_));
 AND2_X1 _23464_ (.A1(_11275_),
    .A2(_11379_),
    .ZN(_13770_));
 OAI22_X1 _23465_ (.A1(_13770_),
    .A2(_11230_),
    .B1(_11275_),
    .B2(_11315_),
    .ZN(_13771_));
 OR2_X1 _23466_ (.A1(_12350_),
    .A2(_12301_),
    .ZN(_13772_));
 OAI21_X1 _23467_ (.A(_11371_),
    .B1(_13772_),
    .B2(_12262_),
    .ZN(_13773_));
 AND4_X1 _23468_ (.A1(_13766_),
    .A2(_13769_),
    .A3(_13771_),
    .A4(_13773_),
    .ZN(_13774_));
 OAI22_X1 _23469_ (.A1(_11330_),
    .A2(_11357_),
    .B1(_11176_),
    .B2(_12279_),
    .ZN(_13775_));
 AOI221_X4 _23470_ (.A(_13775_),
    .B1(_11336_),
    .B2(_11316_),
    .C1(_11253_),
    .C2(_11164_),
    .ZN(_13776_));
 AOI22_X1 _23471_ (.A1(_11157_),
    .A2(_12350_),
    .B1(_11295_),
    .B2(_11253_),
    .ZN(_13777_));
 AOI22_X1 _23472_ (.A1(_11258_),
    .A2(_12683_),
    .B1(_11378_),
    .B2(_11371_),
    .ZN(_13778_));
 NAND3_X1 _23473_ (.A1(_11184_),
    .A2(_11332_),
    .A3(_11341_),
    .ZN(_13779_));
 AOI22_X1 _23474_ (.A1(_11275_),
    .A2(_12350_),
    .B1(_11277_),
    .B2(_11293_),
    .ZN(_13780_));
 OAI21_X1 _23475_ (.A(_11375_),
    .B1(_11270_),
    .B2(_11196_),
    .ZN(_13781_));
 OAI211_X2 _23476_ (.A(_11375_),
    .B(_11164_),
    .C1(_11213_),
    .C2(_11233_),
    .ZN(_13782_));
 AND4_X1 _23477_ (.A1(_13779_),
    .A2(_13780_),
    .A3(_13781_),
    .A4(_13782_),
    .ZN(_13783_));
 AND4_X1 _23478_ (.A1(_13776_),
    .A2(_13777_),
    .A3(_13778_),
    .A4(_13783_),
    .ZN(_13784_));
 NAND4_X1 _23479_ (.A1(_13753_),
    .A2(_13763_),
    .A3(_13774_),
    .A4(_13784_),
    .ZN(_13785_));
 OAI211_X2 _23480_ (.A(_11309_),
    .B(_16815_),
    .C1(_11178_),
    .C2(_11161_),
    .ZN(_13786_));
 OAI211_X2 _23481_ (.A(_11320_),
    .B(_11298_),
    .C1(_11174_),
    .C2(_12327_),
    .ZN(_13787_));
 OAI21_X1 _23482_ (.A(_11309_),
    .B1(_12282_),
    .B2(_11245_),
    .ZN(_13788_));
 AND3_X1 _23483_ (.A1(_13786_),
    .A2(_13787_),
    .A3(_13788_),
    .ZN(_13789_));
 OAI21_X1 _23484_ (.A(_11343_),
    .B1(_11196_),
    .B2(_13032_),
    .ZN(_13790_));
 NAND3_X1 _23485_ (.A1(_11343_),
    .A2(_12314_),
    .A3(_11348_),
    .ZN(_13791_));
 NAND4_X1 _23486_ (.A1(_11165_),
    .A2(_11326_),
    .A3(_11321_),
    .A4(_11341_),
    .ZN(_13792_));
 AND3_X1 _23487_ (.A1(_13790_),
    .A2(_13791_),
    .A3(_13792_),
    .ZN(_13793_));
 NAND4_X1 _23488_ (.A1(_11223_),
    .A2(_11257_),
    .A3(_11260_),
    .A4(_11165_),
    .ZN(_13794_));
 OAI21_X1 _23489_ (.A(_11223_),
    .B1(_11196_),
    .B2(_13032_),
    .ZN(_13795_));
 NAND4_X1 _23490_ (.A1(_13789_),
    .A2(_13793_),
    .A3(_13794_),
    .A4(_13795_),
    .ZN(_13796_));
 NOR2_X4 _23491_ (.A1(_13785_),
    .A2(_13796_),
    .ZN(_13797_));
 NOR3_X1 _23492_ (.A1(_11844_),
    .A2(_11900_),
    .A3(_13091_),
    .ZN(_13798_));
 NAND2_X1 _23493_ (.A1(_11838_),
    .A2(_11749_),
    .ZN(_13799_));
 OAI211_X2 _23494_ (.A(_13798_),
    .B(_13799_),
    .C1(_11788_),
    .C2(_12618_),
    .ZN(_13800_));
 AND2_X1 _23495_ (.A1(_11823_),
    .A2(_11687_),
    .ZN(_13801_));
 OR4_X2 _23496_ (.A1(_12589_),
    .A2(_13286_),
    .A3(_12242_),
    .A4(_13801_),
    .ZN(_13802_));
 OAI211_X2 _23497_ (.A(_12620_),
    .B(_12610_),
    .C1(_11761_),
    .C2(_11699_),
    .ZN(_13803_));
 OAI211_X2 _23498_ (.A(_12620_),
    .B(_16775_),
    .C1(_11765_),
    .C2(_11628_),
    .ZN(_13804_));
 OAI21_X1 _23499_ (.A(_12620_),
    .B1(_11792_),
    .B2(_11782_),
    .ZN(_13805_));
 NAND3_X1 _23500_ (.A1(_13803_),
    .A2(_13804_),
    .A3(_13805_),
    .ZN(_13806_));
 OAI21_X1 _23501_ (.A(_12244_),
    .B1(_11689_),
    .B2(_12208_),
    .ZN(_13807_));
 NAND4_X1 _23502_ (.A1(_12605_),
    .A2(_11826_),
    .A3(_11902_),
    .A4(_12246_),
    .ZN(_13808_));
 OAI21_X1 _23503_ (.A(_12244_),
    .B1(_11805_),
    .B2(_11839_),
    .ZN(_13809_));
 NAND3_X1 _23504_ (.A1(_13807_),
    .A2(_13808_),
    .A3(_13809_),
    .ZN(_13810_));
 NOR4_X2 _23505_ (.A1(_13800_),
    .A2(_13802_),
    .A3(_13806_),
    .A4(_13810_),
    .ZN(_13811_));
 NOR4_X1 _23506_ (.A1(_12656_),
    .A2(_12657_),
    .A3(_13450_),
    .A4(_12221_),
    .ZN(_13812_));
 OAI21_X1 _23507_ (.A(_13123_),
    .B1(_12629_),
    .B2(_11795_),
    .ZN(_13813_));
 AOI211_X4 _23508_ (.A(_13454_),
    .B(_13813_),
    .C1(_11839_),
    .C2(_11744_),
    .ZN(_13814_));
 OAI21_X1 _23509_ (.A(_13319_),
    .B1(_11714_),
    .B2(_11919_),
    .ZN(_13815_));
 AND4_X1 _23510_ (.A1(_11734_),
    .A2(_11632_),
    .A3(_12610_),
    .A4(_11712_),
    .ZN(_13816_));
 NOR4_X1 _23511_ (.A1(_13815_),
    .A2(_13118_),
    .A3(_13119_),
    .A4(_13816_),
    .ZN(_13817_));
 AND2_X1 _23512_ (.A1(_11805_),
    .A2(_11764_),
    .ZN(_13818_));
 NOR4_X1 _23513_ (.A1(_13818_),
    .A2(_13456_),
    .A3(_13126_),
    .A4(_11759_),
    .ZN(_13819_));
 AND4_X1 _23514_ (.A1(_13812_),
    .A2(_13814_),
    .A3(_13817_),
    .A4(_13819_),
    .ZN(_13820_));
 OAI211_X2 _23515_ (.A(_11807_),
    .B(_11808_),
    .C1(_11922_),
    .C2(_12644_),
    .ZN(_13821_));
 OR3_X1 _23516_ (.A1(_13821_),
    .A2(_12213_),
    .A3(_13101_),
    .ZN(_13822_));
 OAI21_X1 _23517_ (.A(_11912_),
    .B1(_11814_),
    .B2(_11833_),
    .ZN(_13823_));
 OR3_X1 _23518_ (.A1(_13823_),
    .A2(_11908_),
    .A3(_11909_),
    .ZN(_13824_));
 OAI21_X1 _23519_ (.A(_11780_),
    .B1(_12202_),
    .B2(_13105_),
    .ZN(_13825_));
 OAI21_X1 _23520_ (.A(_13825_),
    .B1(_11719_),
    .B2(_11925_),
    .ZN(_13826_));
 OAI21_X1 _23521_ (.A(_11791_),
    .B1(_11787_),
    .B2(_11747_),
    .ZN(_13827_));
 OAI211_X2 _23522_ (.A(_11777_),
    .B(_11841_),
    .C1(_11792_),
    .C2(_11782_),
    .ZN(_13828_));
 OAI211_X2 _23523_ (.A(_13827_),
    .B(_13828_),
    .C1(_11692_),
    .C2(_11789_),
    .ZN(_13829_));
 NOR4_X1 _23524_ (.A1(_13822_),
    .A2(_13824_),
    .A3(_13826_),
    .A4(_13829_),
    .ZN(_13830_));
 OAI21_X1 _23525_ (.A(_12604_),
    .B1(_12202_),
    .B2(_13105_),
    .ZN(_13831_));
 NAND3_X1 _23526_ (.A1(_12604_),
    .A2(_11848_),
    .A3(_11850_),
    .ZN(_13832_));
 NAND4_X1 _23527_ (.A1(_11632_),
    .A2(_12610_),
    .A3(_11902_),
    .A4(_11635_),
    .ZN(_13833_));
 AND3_X1 _23528_ (.A1(_13831_),
    .A2(_13832_),
    .A3(_13833_),
    .ZN(_13834_));
 AND2_X1 _23529_ (.A1(_11878_),
    .A2(_11694_),
    .ZN(_13835_));
 AND2_X1 _23530_ (.A1(_11694_),
    .A2(_11724_),
    .ZN(_13836_));
 NOR4_X1 _23531_ (.A1(_13064_),
    .A2(_13835_),
    .A3(_13836_),
    .A4(_13497_),
    .ZN(_13837_));
 OAI21_X1 _23532_ (.A(_11705_),
    .B1(_12202_),
    .B2(_11722_),
    .ZN(_13838_));
 OAI211_X2 _23533_ (.A(_11705_),
    .B(_12610_),
    .C1(_11733_),
    .C2(_11734_),
    .ZN(_13839_));
 AND2_X1 _23534_ (.A1(_13838_),
    .A2(_13839_),
    .ZN(_13840_));
 AOI21_X1 _23535_ (.A(_13076_),
    .B1(_11926_),
    .B2(_11927_),
    .ZN(_13841_));
 AND4_X1 _23536_ (.A1(_11635_),
    .A2(_12605_),
    .A3(_11761_),
    .A4(_12246_),
    .ZN(_13842_));
 NOR4_X1 _23537_ (.A1(_13841_),
    .A2(_11873_),
    .A3(_12195_),
    .A4(_13842_),
    .ZN(_13843_));
 AND4_X1 _23538_ (.A1(_13834_),
    .A2(_13837_),
    .A3(_13840_),
    .A4(_13843_),
    .ZN(_13844_));
 NAND4_X1 _23539_ (.A1(_13811_),
    .A2(_13820_),
    .A3(_13830_),
    .A4(_13844_),
    .ZN(_13845_));
 OR2_X2 _23540_ (.A1(_13845_),
    .A2(_11856_),
    .ZN(_13846_));
 XNOR2_X2 _23541_ (.A(_13797_),
    .B(_13846_),
    .ZN(_13847_));
 XNOR2_X1 _23542_ (.A(_13744_),
    .B(_13847_),
    .ZN(_13848_));
 OAI21_X1 _23543_ (.A(_13132_),
    .B1(_12044_),
    .B2(_12040_),
    .ZN(_13849_));
 OAI21_X1 _23544_ (.A(_12006_),
    .B1(_12153_),
    .B2(_12043_),
    .ZN(_13850_));
 AOI221_X1 _23545_ (.A(_13850_),
    .B1(_13144_),
    .B2(_12834_),
    .C1(_12168_),
    .C2(_11964_),
    .ZN(_13851_));
 AOI221_X2 _23546_ (.A(_12016_),
    .B1(_11995_),
    .B2(_12075_),
    .C1(_12119_),
    .C2(_12162_),
    .ZN(_13852_));
 AND4_X1 _23547_ (.A1(_13849_),
    .A2(_13851_),
    .A3(_12116_),
    .A4(_13852_),
    .ZN(_13853_));
 AOI21_X1 _23548_ (.A(_12561_),
    .B1(_12840_),
    .B2(_12849_),
    .ZN(_13854_));
 NAND2_X1 _23549_ (.A1(_12088_),
    .A2(_12493_),
    .ZN(_13855_));
 NAND2_X1 _23550_ (.A1(_12487_),
    .A2(_12119_),
    .ZN(_13856_));
 NAND2_X1 _23551_ (.A1(_13855_),
    .A2(_13856_),
    .ZN(_13857_));
 NOR3_X1 _23552_ (.A1(_12539_),
    .A2(_13854_),
    .A3(_13857_),
    .ZN(_13858_));
 AOI22_X1 _23553_ (.A1(_12062_),
    .A2(_12044_),
    .B1(_13144_),
    .B2(_12484_),
    .ZN(_13859_));
 OAI211_X2 _23554_ (.A(_13859_),
    .B(_13247_),
    .C1(_12509_),
    .C2(_12850_),
    .ZN(_13860_));
 AND2_X1 _23555_ (.A1(_12025_),
    .A2(_12830_),
    .ZN(_13861_));
 OR2_X1 _23556_ (.A1(_12126_),
    .A2(_13861_),
    .ZN(_13862_));
 OAI211_X2 _23557_ (.A(_12511_),
    .B(_12548_),
    .C1(_13191_),
    .C2(_12549_),
    .ZN(_13863_));
 NOR4_X1 _23558_ (.A1(_13860_),
    .A2(_12136_),
    .A3(_13862_),
    .A4(_13863_),
    .ZN(_13864_));
 INV_X1 _23559_ (.A(_13220_),
    .ZN(_13865_));
 OAI221_X1 _23560_ (.A(_13865_),
    .B1(_12535_),
    .B2(_12850_),
    .C1(_12073_),
    .C2(_12549_),
    .ZN(_13866_));
 INV_X1 _23561_ (.A(_13571_),
    .ZN(_13867_));
 OAI21_X1 _23562_ (.A(_13867_),
    .B1(_12138_),
    .B2(_12504_),
    .ZN(_13868_));
 AND2_X1 _23563_ (.A1(_12527_),
    .A2(_12156_),
    .ZN(_13869_));
 NAND3_X1 _23564_ (.A1(_12836_),
    .A2(_13610_),
    .A3(_13601_),
    .ZN(_13870_));
 NOR4_X1 _23565_ (.A1(_13866_),
    .A2(_13868_),
    .A3(_13869_),
    .A4(_13870_),
    .ZN(_13871_));
 NAND4_X1 _23566_ (.A1(_13853_),
    .A2(_13858_),
    .A3(_13864_),
    .A4(_13871_),
    .ZN(_13872_));
 OAI21_X1 _23567_ (.A(_12167_),
    .B1(_12040_),
    .B2(_12090_),
    .ZN(_13873_));
 AOI21_X1 _23568_ (.A(_12143_),
    .B1(_12155_),
    .B2(_13180_),
    .ZN(_13874_));
 OAI21_X1 _23569_ (.A(_12147_),
    .B1(_12143_),
    .B2(_12045_),
    .ZN(_13875_));
 NOR4_X1 _23570_ (.A1(_13874_),
    .A2(_13875_),
    .A3(_13271_),
    .A4(_12582_),
    .ZN(_13876_));
 OAI21_X1 _23571_ (.A(_12056_),
    .B1(_12039_),
    .B2(_12163_),
    .ZN(_13877_));
 OAI21_X1 _23572_ (.A(_12056_),
    .B1(_12068_),
    .B2(_12025_),
    .ZN(_13878_));
 AND4_X1 _23573_ (.A1(_13873_),
    .A2(_13876_),
    .A3(_13877_),
    .A4(_13878_),
    .ZN(_13879_));
 OR2_X1 _23574_ (.A1(_12853_),
    .A2(_12533_),
    .ZN(_13880_));
 OAI21_X1 _23575_ (.A(_12150_),
    .B1(_11997_),
    .B2(_12552_),
    .ZN(_13881_));
 OAI21_X1 _23576_ (.A(_13881_),
    .B1(_13177_),
    .B2(_12489_),
    .ZN(_13882_));
 NOR4_X1 _23577_ (.A1(_13882_),
    .A2(_12486_),
    .A3(_12856_),
    .A4(_12854_),
    .ZN(_13883_));
 AND2_X1 _23578_ (.A1(_12030_),
    .A2(_12089_),
    .ZN(_13884_));
 OAI21_X1 _23579_ (.A(_11964_),
    .B1(_12507_),
    .B2(_13884_),
    .ZN(_13885_));
 AOI22_X1 _23580_ (.A1(_12834_),
    .A2(_12088_),
    .B1(_12056_),
    .B2(_13164_),
    .ZN(_13886_));
 NAND2_X1 _23581_ (.A1(_12088_),
    .A2(_12005_),
    .ZN(_13887_));
 NAND2_X1 _23582_ (.A1(_12487_),
    .A2(_12122_),
    .ZN(_13888_));
 AND3_X1 _23583_ (.A1(_13886_),
    .A2(_13887_),
    .A3(_13888_),
    .ZN(_13889_));
 AND4_X1 _23584_ (.A1(_13880_),
    .A2(_13883_),
    .A3(_13885_),
    .A4(_13889_),
    .ZN(_13890_));
 NOR2_X1 _23585_ (.A1(_12547_),
    .A2(_13590_),
    .ZN(_13891_));
 NAND2_X1 _23586_ (.A1(_12490_),
    .A2(_12830_),
    .ZN(_13892_));
 AND4_X1 _23587_ (.A1(_12084_),
    .A2(_13891_),
    .A3(_13892_),
    .A4(_12502_),
    .ZN(_13893_));
 AOI22_X1 _23588_ (.A1(_12860_),
    .A2(_12128_),
    .B1(_12861_),
    .B2(_13132_),
    .ZN(_13894_));
 NAND2_X1 _23589_ (.A1(_12005_),
    .A2(_12161_),
    .ZN(_13895_));
 OAI211_X2 _23590_ (.A(_13894_),
    .B(_13895_),
    .C1(_12139_),
    .C2(_12839_),
    .ZN(_13896_));
 OAI221_X1 _23591_ (.A(_13578_),
    .B1(_12133_),
    .B2(_12043_),
    .C1(_12063_),
    .C2(_12051_),
    .ZN(_13897_));
 OAI21_X1 _23592_ (.A(_12088_),
    .B1(_12861_),
    .B2(_12050_),
    .ZN(_13898_));
 OAI211_X2 _23593_ (.A(_13898_),
    .B(_13595_),
    .C1(_12133_),
    .C2(_12482_),
    .ZN(_13899_));
 AND3_X1 _23594_ (.A1(_12830_),
    .A2(_11987_),
    .A3(_11999_),
    .ZN(_13900_));
 NOR4_X1 _23595_ (.A1(_13896_),
    .A2(_13897_),
    .A3(_13899_),
    .A4(_13900_),
    .ZN(_13901_));
 NAND4_X1 _23596_ (.A1(_13879_),
    .A2(_13890_),
    .A3(_13893_),
    .A4(_13901_),
    .ZN(_13902_));
 NOR2_X4 _23597_ (.A1(_13872_),
    .A2(_13902_),
    .ZN(_13903_));
 XNOR2_X1 _23598_ (.A(_13848_),
    .B(_13903_),
    .ZN(_13904_));
 INV_X1 _23599_ (.A(_17268_),
    .ZN(_13905_));
 XNOR2_X1 _23600_ (.A(_13904_),
    .B(_13905_),
    .ZN(_13906_));
 MUX2_X1 _23601_ (.A(_13689_),
    .B(_13906_),
    .S(_11149_),
    .Z(_00722_));
 XOR2_X1 _23602_ (.A(_17269_),
    .B(_17072_),
    .Z(_13907_));
 OAI21_X1 _23603_ (.A(_13559_),
    .B1(_11355_),
    .B2(_11346_),
    .ZN(_13908_));
 AND3_X1 _23604_ (.A1(_11353_),
    .A2(_11260_),
    .A3(_11163_),
    .ZN(_13909_));
 NOR4_X1 _23605_ (.A1(_13908_),
    .A2(_12277_),
    .A3(_13909_),
    .A4(_11354_),
    .ZN(_13910_));
 OAI21_X1 _23606_ (.A(_11375_),
    .B1(_12343_),
    .B2(_11284_),
    .ZN(_13911_));
 AND4_X1 _23607_ (.A1(_12997_),
    .A2(_13910_),
    .A3(_13554_),
    .A4(_13911_),
    .ZN(_13912_));
 AND2_X1 _23608_ (.A1(_11184_),
    .A2(_11342_),
    .ZN(_13913_));
 INV_X1 _23609_ (.A(_13913_),
    .ZN(_13914_));
 NAND3_X1 _23610_ (.A1(_11207_),
    .A2(_11326_),
    .A3(_11341_),
    .ZN(_13915_));
 OAI211_X2 _23611_ (.A(_13914_),
    .B(_13915_),
    .C1(_11291_),
    .C2(_13008_),
    .ZN(_13916_));
 OAI211_X2 _23612_ (.A(_11368_),
    .B(_12265_),
    .C1(_11213_),
    .C2(_11209_),
    .ZN(_13917_));
 OAI21_X1 _23613_ (.A(_13917_),
    .B1(_11357_),
    .B2(_11369_),
    .ZN(_13918_));
 NAND2_X1 _23614_ (.A1(_11368_),
    .A2(_11279_),
    .ZN(_13919_));
 OAI211_X2 _23615_ (.A(_12708_),
    .B(_13919_),
    .C1(_12316_),
    .C2(_11369_),
    .ZN(_13920_));
 NOR4_X2 _23616_ (.A1(_13916_),
    .A2(_13382_),
    .A3(_13918_),
    .A4(_13920_),
    .ZN(_13921_));
 OAI21_X1 _23617_ (.A(_11328_),
    .B1(_12704_),
    .B2(_12304_),
    .ZN(_13922_));
 OAI21_X1 _23618_ (.A(_11328_),
    .B1(_11214_),
    .B2(_11160_),
    .ZN(_13923_));
 OAI21_X1 _23619_ (.A(_11314_),
    .B1(_11358_),
    .B2(_11245_),
    .ZN(_13924_));
 AND4_X1 _23620_ (.A1(_12722_),
    .A2(_13922_),
    .A3(_13923_),
    .A4(_13924_),
    .ZN(_13925_));
 OAI211_X2 _23621_ (.A(_11153_),
    .B(_11319_),
    .C1(_11378_),
    .C2(_12262_),
    .ZN(_13926_));
 OAI211_X2 _23622_ (.A(_11153_),
    .B(_11319_),
    .C1(_11190_),
    .C2(_11230_),
    .ZN(_13927_));
 OAI211_X2 _23623_ (.A(_13926_),
    .B(_13927_),
    .C1(_11337_),
    .C2(_11357_),
    .ZN(_13928_));
 NAND3_X1 _23624_ (.A1(_11190_),
    .A2(_11319_),
    .A3(_11298_),
    .ZN(_13929_));
 NAND3_X1 _23625_ (.A1(_11379_),
    .A2(_11319_),
    .A3(_11298_),
    .ZN(_13930_));
 NAND2_X1 _23626_ (.A1(_13929_),
    .A2(_13930_),
    .ZN(_13931_));
 AND2_X1 _23627_ (.A1(_11309_),
    .A2(_12327_),
    .ZN(_13932_));
 NOR4_X2 _23628_ (.A1(_13928_),
    .A2(_13931_),
    .A3(_11307_),
    .A4(_13932_),
    .ZN(_13933_));
 NAND4_X2 _23629_ (.A1(_13912_),
    .A2(_13921_),
    .A3(_13925_),
    .A4(_13933_),
    .ZN(_13934_));
 AND4_X1 _23630_ (.A1(_12274_),
    .A2(_11242_),
    .A3(_11163_),
    .A4(_11348_),
    .ZN(_13935_));
 AND3_X1 _23631_ (.A1(_11242_),
    .A2(_11188_),
    .A3(_11186_),
    .ZN(_13936_));
 NOR3_X1 _23632_ (.A1(_13935_),
    .A2(_13936_),
    .A3(_12322_),
    .ZN(_13937_));
 NOR4_X2 _23633_ (.A1(_11287_),
    .A2(_13760_),
    .A3(_13054_),
    .A4(_11285_),
    .ZN(_13938_));
 OAI21_X1 _23634_ (.A(_11263_),
    .B1(_11345_),
    .B2(_11179_),
    .ZN(_13939_));
 OAI21_X1 _23635_ (.A(_11263_),
    .B1(_11377_),
    .B2(_11250_),
    .ZN(_13940_));
 OAI21_X1 _23636_ (.A(_11263_),
    .B1(_11207_),
    .B2(_11229_),
    .ZN(_13941_));
 AND4_X1 _23637_ (.A1(_13521_),
    .A2(_13939_),
    .A3(_13940_),
    .A4(_13941_),
    .ZN(_13942_));
 AOI21_X1 _23638_ (.A(_11290_),
    .B1(_11191_),
    .B2(_11278_),
    .ZN(_13943_));
 AND4_X1 _23639_ (.A1(_11213_),
    .A2(_11183_),
    .A3(_11241_),
    .A4(_11169_),
    .ZN(_13944_));
 NOR4_X1 _23640_ (.A1(_13943_),
    .A2(_12319_),
    .A3(_13765_),
    .A4(_13944_),
    .ZN(_13945_));
 AND4_X2 _23641_ (.A1(_13937_),
    .A2(_13938_),
    .A3(_13942_),
    .A4(_13945_),
    .ZN(_13946_));
 NAND3_X1 _23642_ (.A1(_11171_),
    .A2(_11164_),
    .A3(_11348_),
    .ZN(_13947_));
 AND4_X1 _23643_ (.A1(_12307_),
    .A2(_13334_),
    .A3(_12309_),
    .A4(_13947_),
    .ZN(_13948_));
 AOI21_X1 _23644_ (.A(_12295_),
    .B1(_12999_),
    .B2(_11180_),
    .ZN(_13949_));
 AOI21_X1 _23645_ (.A(_12295_),
    .B1(_11249_),
    .B2(_11280_),
    .ZN(_13950_));
 AOI211_X4 _23646_ (.A(_13949_),
    .B(_13950_),
    .C1(_12301_),
    .C2(_11157_),
    .ZN(_13951_));
 NAND4_X1 _23647_ (.A1(_11167_),
    .A2(_11326_),
    .A3(_11233_),
    .A4(_11322_),
    .ZN(_13952_));
 OAI21_X1 _23648_ (.A(_11222_),
    .B1(_12349_),
    .B2(_12301_),
    .ZN(_13953_));
 OAI21_X1 _23649_ (.A(_11222_),
    .B1(_11250_),
    .B2(_11364_),
    .ZN(_13954_));
 AND2_X1 _23650_ (.A1(_13953_),
    .A2(_13954_),
    .ZN(_13955_));
 OAI21_X1 _23651_ (.A(_12683_),
    .B1(_12704_),
    .B2(_11207_),
    .ZN(_13956_));
 OAI211_X2 _23652_ (.A(_11204_),
    .B(_12265_),
    .C1(_11244_),
    .C2(_11217_),
    .ZN(_13957_));
 AND4_X1 _23653_ (.A1(_13952_),
    .A2(_13955_),
    .A3(_13956_),
    .A4(_13957_),
    .ZN(_13958_));
 NAND4_X4 _23654_ (.A1(_13946_),
    .A2(_13948_),
    .A3(_13951_),
    .A4(_13958_),
    .ZN(_13959_));
 NOR2_X4 _23655_ (.A1(_13934_),
    .A2(_13959_),
    .ZN(_13960_));
 XOR2_X2 _23656_ (.A(_11958_),
    .B(_13960_),
    .Z(_13961_));
 NAND2_X1 _23657_ (.A1(_11573_),
    .A2(_11481_),
    .ZN(_13962_));
 OAI221_X1 _23658_ (.A(_13962_),
    .B1(_11523_),
    .B2(_11541_),
    .C1(_12423_),
    .C2(_11604_),
    .ZN(_13963_));
 AOI211_X2 _23659_ (.A(_13732_),
    .B(_13963_),
    .C1(_12972_),
    .C2(_11502_),
    .ZN(_13964_));
 NOR2_X1 _23660_ (.A1(_13417_),
    .A2(_11601_),
    .ZN(_13965_));
 AND2_X1 _23661_ (.A1(_11539_),
    .A2(_11561_),
    .ZN(_13966_));
 NOR4_X1 _23662_ (.A1(_13965_),
    .A2(_13966_),
    .A3(_13428_),
    .A4(_13429_),
    .ZN(_13967_));
 NOR4_X1 _23663_ (.A1(_12818_),
    .A2(_12819_),
    .A3(_12782_),
    .A4(_12795_),
    .ZN(_13968_));
 AND2_X1 _23664_ (.A1(_11482_),
    .A2(_11502_),
    .ZN(_13969_));
 NOR4_X2 _23665_ (.A1(_12376_),
    .A2(_13969_),
    .A3(_12769_),
    .A4(_12360_),
    .ZN(_13970_));
 NAND4_X1 _23666_ (.A1(_13964_),
    .A2(_13967_),
    .A3(_13968_),
    .A4(_13970_),
    .ZN(_13971_));
 OAI21_X1 _23667_ (.A(_12764_),
    .B1(_12423_),
    .B2(_12387_),
    .ZN(_13972_));
 AOI221_X1 _23668_ (.A(_13972_),
    .B1(_11519_),
    .B2(_11446_),
    .C1(_12379_),
    .C2(_11424_),
    .ZN(_13973_));
 AND2_X1 _23669_ (.A1(_11479_),
    .A2(_11519_),
    .ZN(_13974_));
 OAI21_X1 _23670_ (.A(_12925_),
    .B1(_11617_),
    .B2(_11489_),
    .ZN(_13975_));
 AOI211_X2 _23671_ (.A(_13974_),
    .B(_13975_),
    .C1(_12386_),
    .C2(_11501_),
    .ZN(_13976_));
 AND2_X1 _23672_ (.A1(_11510_),
    .A2(_11391_),
    .ZN(_13977_));
 AND2_X1 _23673_ (.A1(_11515_),
    .A2(_11433_),
    .ZN(_13978_));
 NOR4_X2 _23674_ (.A1(_12756_),
    .A2(_12978_),
    .A3(_13977_),
    .A4(_13978_),
    .ZN(_13979_));
 AND3_X1 _23675_ (.A1(_11459_),
    .A2(_11464_),
    .A3(_11478_),
    .ZN(_13980_));
 AOI211_X2 _23676_ (.A(_12777_),
    .B(_13980_),
    .C1(_11459_),
    .C2(_11606_),
    .ZN(_13981_));
 NAND4_X1 _23677_ (.A1(_13973_),
    .A2(_13976_),
    .A3(_13979_),
    .A4(_13981_),
    .ZN(_13982_));
 OAI21_X1 _23678_ (.A(_11567_),
    .B1(_12812_),
    .B2(_11434_),
    .ZN(_13983_));
 NAND4_X1 _23679_ (.A1(_11537_),
    .A2(_11445_),
    .A3(_11414_),
    .A4(_11599_),
    .ZN(_13984_));
 OAI211_X2 _23680_ (.A(_11567_),
    .B(_11411_),
    .C1(_11600_),
    .C2(_11601_),
    .ZN(_13985_));
 NAND4_X1 _23681_ (.A1(_13983_),
    .A2(_13736_),
    .A3(_13984_),
    .A4(_13985_),
    .ZN(_13986_));
 AND3_X2 _23682_ (.A1(_11585_),
    .A2(_12393_),
    .A3(_11391_),
    .ZN(_13987_));
 AOI211_X2 _23683_ (.A(_13691_),
    .B(_13987_),
    .C1(_11556_),
    .C2(_11515_),
    .ZN(_13988_));
 OAI21_X1 _23684_ (.A(_12456_),
    .B1(_11570_),
    .B2(_12379_),
    .ZN(_13989_));
 AND3_X2 _23685_ (.A1(_11597_),
    .A2(_12393_),
    .A3(_12430_),
    .ZN(_13990_));
 AOI21_X1 _23686_ (.A(_13990_),
    .B1(_12456_),
    .B2(_12812_),
    .ZN(_13991_));
 OAI21_X1 _23687_ (.A(_11554_),
    .B1(_11499_),
    .B2(_11548_),
    .ZN(_13992_));
 OAI21_X1 _23688_ (.A(_11554_),
    .B1(_12409_),
    .B2(_11496_),
    .ZN(_13993_));
 AND2_X1 _23689_ (.A1(_13992_),
    .A2(_13993_),
    .ZN(_13994_));
 NAND4_X1 _23690_ (.A1(_13988_),
    .A2(_13989_),
    .A3(_13991_),
    .A4(_13994_),
    .ZN(_13995_));
 NOR4_X1 _23691_ (.A1(_13971_),
    .A2(_13982_),
    .A3(_13986_),
    .A4(_13995_),
    .ZN(_13996_));
 AOI21_X1 _23692_ (.A(_11525_),
    .B1(_11617_),
    .B2(_12400_),
    .ZN(_13997_));
 AOI211_X2 _23693_ (.A(_12437_),
    .B(_13997_),
    .C1(_11447_),
    .C2(_11561_),
    .ZN(_13998_));
 NAND3_X1 _23694_ (.A1(_11442_),
    .A2(_11415_),
    .A3(_11412_),
    .ZN(_13999_));
 AOI22_X1 _23695_ (.A1(_11543_),
    .A2(_12463_),
    .B1(_11544_),
    .B2(_11396_),
    .ZN(_14000_));
 NAND4_X1 _23696_ (.A1(_13998_),
    .A2(_12411_),
    .A3(_13999_),
    .A4(_14000_),
    .ZN(_14001_));
 OR4_X2 _23697_ (.A1(_11471_),
    .A2(_11588_),
    .A3(_11473_),
    .A4(_13707_),
    .ZN(_14002_));
 AND3_X1 _23698_ (.A1(_12409_),
    .A2(_11591_),
    .A3(_11586_),
    .ZN(_14003_));
 INV_X1 _23699_ (.A(_14003_),
    .ZN(_14004_));
 OAI21_X1 _23700_ (.A(_11442_),
    .B1(_12417_),
    .B2(_12972_),
    .ZN(_14005_));
 NAND2_X1 _23701_ (.A1(_11470_),
    .A2(_11505_),
    .ZN(_14006_));
 NAND4_X1 _23702_ (.A1(_13668_),
    .A2(_14004_),
    .A3(_14005_),
    .A4(_14006_),
    .ZN(_14007_));
 AOI221_X2 _23703_ (.A(_13702_),
    .B1(_11510_),
    .B2(_11616_),
    .C1(_11529_),
    .C2(_12920_),
    .ZN(_14008_));
 INV_X1 _23704_ (.A(_11495_),
    .ZN(_14009_));
 NOR2_X1 _23705_ (.A1(_13398_),
    .A2(_12436_),
    .ZN(_14010_));
 NAND4_X1 _23706_ (.A1(_14008_),
    .A2(_14009_),
    .A3(_12794_),
    .A4(_14010_),
    .ZN(_14011_));
 NOR4_X1 _23707_ (.A1(_14001_),
    .A2(_14002_),
    .A3(_14007_),
    .A4(_14011_),
    .ZN(_14012_));
 AND2_X1 _23708_ (.A1(_13996_),
    .A2(_14012_),
    .ZN(_14013_));
 BUF_X4 _23709_ (.A(_14013_),
    .Z(_14014_));
 XNOR2_X1 _23710_ (.A(_14014_),
    .B(_13846_),
    .ZN(_14015_));
 XNOR2_X1 _23711_ (.A(_13961_),
    .B(_14015_),
    .ZN(_14016_));
 AND3_X1 _23712_ (.A1(_12826_),
    .A2(_12121_),
    .A3(_13592_),
    .ZN(_14017_));
 OAI211_X2 _23713_ (.A(_14017_),
    .B(_13255_),
    .C1(_12092_),
    .C2(_12138_),
    .ZN(_14018_));
 AND2_X1 _23714_ (.A1(_12162_),
    .A2(_12071_),
    .ZN(_14019_));
 OAI211_X2 _23715_ (.A(_13895_),
    .B(_13263_),
    .C1(_12144_),
    .C2(_12839_),
    .ZN(_14020_));
 AOI21_X1 _23716_ (.A(_12853_),
    .B1(_12153_),
    .B2(_12073_),
    .ZN(_14021_));
 AOI21_X1 _23717_ (.A(_12853_),
    .B1(_12155_),
    .B2(_12130_),
    .ZN(_14022_));
 OR4_X2 _23718_ (.A1(_14019_),
    .A2(_14020_),
    .A3(_14021_),
    .A4(_14022_),
    .ZN(_14023_));
 NOR2_X1 _23719_ (.A1(_12131_),
    .A2(_12580_),
    .ZN(_14024_));
 NOR4_X2 _23720_ (.A1(_14018_),
    .A2(_14023_),
    .A3(_14024_),
    .A4(_13169_),
    .ZN(_14025_));
 NAND4_X1 _23721_ (.A1(_13213_),
    .A2(_12087_),
    .A3(_13855_),
    .A4(_12900_),
    .ZN(_14026_));
 OAI211_X2 _23722_ (.A(_12863_),
    .B(_12496_),
    .C1(_12050_),
    .C2(_12484_),
    .ZN(_14027_));
 OAI221_X1 _23723_ (.A(_14027_),
    .B1(_13191_),
    .B2(_12063_),
    .C1(_12899_),
    .C2(_12031_),
    .ZN(_14028_));
 NAND4_X1 _23724_ (.A1(_12496_),
    .A2(_12089_),
    .A3(_12528_),
    .A4(_11962_),
    .ZN(_14029_));
 NAND4_X1 _23725_ (.A1(_12496_),
    .A2(_12089_),
    .A3(_12090_),
    .A4(_11962_),
    .ZN(_14030_));
 OAI21_X1 _23726_ (.A(_12056_),
    .B1(_12025_),
    .B2(_12119_),
    .ZN(_14031_));
 NAND4_X1 _23727_ (.A1(_12057_),
    .A2(_14029_),
    .A3(_14030_),
    .A4(_14031_),
    .ZN(_14032_));
 OAI21_X1 _23728_ (.A(_12487_),
    .B1(_12834_),
    .B2(_12019_),
    .ZN(_14033_));
 OAI21_X1 _23729_ (.A(_12487_),
    .B1(_12163_),
    .B2(_12075_),
    .ZN(_14034_));
 OAI211_X2 _23730_ (.A(_12035_),
    .B(_12496_),
    .C1(_13164_),
    .C2(_12015_),
    .ZN(_14035_));
 NAND4_X1 _23731_ (.A1(_14033_),
    .A2(_14034_),
    .A3(_13856_),
    .A4(_14035_),
    .ZN(_14036_));
 NOR4_X1 _23732_ (.A1(_14026_),
    .A2(_14028_),
    .A3(_14032_),
    .A4(_14036_),
    .ZN(_14037_));
 AND3_X1 _23733_ (.A1(_12142_),
    .A2(_11990_),
    .A3(_12532_),
    .ZN(_14038_));
 OR4_X1 _23734_ (.A1(_13269_),
    .A2(_14038_),
    .A3(_12879_),
    .A4(_13272_),
    .ZN(_14039_));
 OAI21_X1 _23735_ (.A(_12150_),
    .B1(_12168_),
    .B2(_13884_),
    .ZN(_14040_));
 OAI21_X1 _23736_ (.A(_14040_),
    .B1(_12508_),
    .B2(_12151_),
    .ZN(_14041_));
 OAI21_X1 _23737_ (.A(_12108_),
    .B1(_12541_),
    .B2(_12068_),
    .ZN(_14042_));
 OAI21_X1 _23738_ (.A(_12108_),
    .B1(_13164_),
    .B2(_12015_),
    .ZN(_14043_));
 OAI211_X2 _23739_ (.A(_14042_),
    .B(_14043_),
    .C1(_13177_),
    .C2(_12045_),
    .ZN(_14044_));
 INV_X1 _23740_ (.A(_13581_),
    .ZN(_14045_));
 NAND2_X1 _23741_ (.A1(_12109_),
    .A2(_12544_),
    .ZN(_14046_));
 NAND4_X1 _23742_ (.A1(_14045_),
    .A2(_14046_),
    .A3(_12859_),
    .A4(_13583_),
    .ZN(_14047_));
 NOR4_X1 _23743_ (.A1(_14039_),
    .A2(_14041_),
    .A3(_14044_),
    .A4(_14047_),
    .ZN(_14048_));
 AND2_X1 _23744_ (.A1(_12005_),
    .A2(_12012_),
    .ZN(_14049_));
 NOR3_X1 _23745_ (.A1(_12023_),
    .A2(_14049_),
    .A3(_12563_),
    .ZN(_14050_));
 OAI211_X2 _23746_ (.A(_14050_),
    .B(_12017_),
    .C1(_12561_),
    .C2(_12045_),
    .ZN(_14051_));
 OAI21_X1 _23747_ (.A(_13144_),
    .B1(_12168_),
    .B2(_13884_),
    .ZN(_14052_));
 OAI211_X2 _23748_ (.A(_12863_),
    .B(_11985_),
    .C1(_13164_),
    .C2(_12050_),
    .ZN(_14053_));
 NAND4_X1 _23749_ (.A1(_12863_),
    .A2(_12528_),
    .A3(_12089_),
    .A4(_11985_),
    .ZN(_14054_));
 NAND3_X1 _23750_ (.A1(_14052_),
    .A2(_14053_),
    .A3(_14054_),
    .ZN(_14055_));
 INV_X1 _23751_ (.A(_11979_),
    .ZN(_14056_));
 OAI21_X1 _23752_ (.A(_11964_),
    .B1(_12109_),
    .B2(_12152_),
    .ZN(_14057_));
 NAND4_X1 _23753_ (.A1(_14056_),
    .A2(_12848_),
    .A3(_13150_),
    .A4(_14057_),
    .ZN(_14058_));
 OAI21_X1 _23754_ (.A(_13132_),
    .B1(_12168_),
    .B2(_12122_),
    .ZN(_14059_));
 OAI211_X2 _23755_ (.A(_13132_),
    .B(_12528_),
    .C1(_12024_),
    .C2(_12031_),
    .ZN(_14060_));
 OAI211_X2 _23756_ (.A(_14059_),
    .B(_14060_),
    .C1(_12043_),
    .C2(_12059_),
    .ZN(_14061_));
 NOR4_X1 _23757_ (.A1(_14051_),
    .A2(_14055_),
    .A3(_14058_),
    .A4(_14061_),
    .ZN(_14062_));
 AND4_X1 _23758_ (.A1(_14025_),
    .A2(_14037_),
    .A3(_14048_),
    .A4(_14062_),
    .ZN(_14063_));
 NAND2_X2 _23759_ (.A1(_14063_),
    .A2(_12883_),
    .ZN(_14064_));
 XNOR2_X1 _23760_ (.A(_14016_),
    .B(_14064_),
    .ZN(_14065_));
 XOR2_X1 _23761_ (.A(_14065_),
    .B(_17269_),
    .Z(_14066_));
 MUX2_X1 _23762_ (.A(_13907_),
    .B(_14066_),
    .S(_11149_),
    .Z(_00723_));
 NOR2_X1 _23763_ (.A1(_11127_),
    .A2(_17162_),
    .ZN(_14067_));
 BUF_X2 _23764_ (.A(_14067_),
    .Z(_14068_));
 NOR2_X2 _23765_ (.A1(_11103_),
    .A2(_17161_),
    .ZN(_14069_));
 AND2_X2 _23766_ (.A1(_14068_),
    .A2(_14069_),
    .ZN(_14070_));
 AND2_X1 _23767_ (.A1(_17164_),
    .A2(_17165_),
    .ZN(_14071_));
 BUF_X4 _23768_ (.A(_14071_),
    .Z(_14072_));
 NOR2_X1 _23769_ (.A1(_17167_),
    .A2(_17168_),
    .ZN(_14073_));
 AND2_X2 _23770_ (.A1(_14072_),
    .A2(_14073_),
    .ZN(_14074_));
 BUF_X4 _23771_ (.A(_14074_),
    .Z(_14075_));
 AND2_X1 _23772_ (.A1(_14070_),
    .A2(_14075_),
    .ZN(_14076_));
 AND2_X2 _23773_ (.A1(_17162_),
    .A2(_17163_),
    .ZN(_14077_));
 BUF_X4 _23774_ (.A(_14077_),
    .Z(_14078_));
 INV_X1 _23775_ (.A(_14078_),
    .ZN(_14079_));
 INV_X1 _23776_ (.A(_14074_),
    .ZN(_14080_));
 INV_X32 _23777_ (.A(_17160_),
    .ZN(_14081_));
 AOI211_X4 _23778_ (.A(_14079_),
    .B(_14080_),
    .C1(_14081_),
    .C2(_11111_),
    .ZN(_14082_));
 INV_X2 _23779_ (.A(_14069_),
    .ZN(_14083_));
 NOR2_X1 _23780_ (.A1(_17162_),
    .A2(_17163_),
    .ZN(_14084_));
 BUF_X2 _23781_ (.A(_14084_),
    .Z(_14085_));
 NAND2_X1 _23782_ (.A1(_14083_),
    .A2(_14085_),
    .ZN(_14086_));
 NOR2_X1 _23783_ (.A1(_14080_),
    .A2(_14086_),
    .ZN(_14087_));
 INV_X1 _23784_ (.A(_17162_),
    .ZN(_14088_));
 NOR2_X2 _23785_ (.A1(_14088_),
    .A2(_17163_),
    .ZN(_14089_));
 BUF_X4 _23786_ (.A(_14089_),
    .Z(_14090_));
 INV_X2 _23787_ (.A(_17161_),
    .ZN(_14091_));
 NOR2_X4 _23788_ (.A1(_14091_),
    .A2(_11103_),
    .ZN(_14092_));
 BUF_X2 _23789_ (.A(_14092_),
    .Z(_14093_));
 AND3_X1 _23790_ (.A1(_14074_),
    .A2(_14090_),
    .A3(_14093_),
    .ZN(_14094_));
 OR4_X1 _23791_ (.A1(_14076_),
    .A2(_14082_),
    .A3(_14087_),
    .A4(_14094_),
    .ZN(_14095_));
 NOR2_X1 _23792_ (.A1(_14081_),
    .A2(_17161_),
    .ZN(_14096_));
 AND2_X1 _23793_ (.A1(_14089_),
    .A2(_14096_),
    .ZN(_14097_));
 NOR2_X1 _23794_ (.A1(_17164_),
    .A2(_17165_),
    .ZN(_14098_));
 AND2_X1 _23795_ (.A1(_14073_),
    .A2(_14098_),
    .ZN(_14099_));
 CLKBUF_X2 _23796_ (.A(_14099_),
    .Z(_14100_));
 AND2_X1 _23797_ (.A1(_14097_),
    .A2(_14100_),
    .ZN(_14101_));
 AND2_X2 _23798_ (.A1(_14089_),
    .A2(_11111_),
    .ZN(_14102_));
 BUF_X2 _23799_ (.A(_14100_),
    .Z(_14103_));
 AND2_X1 _23800_ (.A1(_14102_),
    .A2(_14103_),
    .ZN(_14104_));
 AND2_X2 _23801_ (.A1(_14084_),
    .A2(_11111_),
    .ZN(_14105_));
 AND2_X1 _23802_ (.A1(_14100_),
    .A2(_14105_),
    .ZN(_14106_));
 NOR3_X1 _23803_ (.A1(_14101_),
    .A2(_14104_),
    .A3(_14106_),
    .ZN(_14107_));
 BUF_X4 _23804_ (.A(_14068_),
    .Z(_14108_));
 BUF_X4 _23805_ (.A(_14108_),
    .Z(_14109_));
 NAND3_X1 _23806_ (.A1(_14103_),
    .A2(_14083_),
    .A3(_14109_),
    .ZN(_14110_));
 INV_X1 _23807_ (.A(_14099_),
    .ZN(_14111_));
 NAND2_X1 _23808_ (.A1(_14083_),
    .A2(_14078_),
    .ZN(_14112_));
 AND2_X1 _23809_ (.A1(_17160_),
    .A2(_17161_),
    .ZN(_14113_));
 BUF_X4 _23810_ (.A(_14113_),
    .Z(_14114_));
 NOR2_X1 _23811_ (.A1(_14112_),
    .A2(_14114_),
    .ZN(_14115_));
 INV_X1 _23812_ (.A(_14115_),
    .ZN(_14116_));
 OAI211_X2 _23813_ (.A(_14107_),
    .B(_14110_),
    .C1(_14111_),
    .C2(_14116_),
    .ZN(_14117_));
 INV_X16 _23814_ (.A(_17165_),
    .ZN(_14118_));
 AND2_X2 _23815_ (.A1(_14118_),
    .A2(_17164_),
    .ZN(_14119_));
 AND2_X1 _23816_ (.A1(_14119_),
    .A2(_14073_),
    .ZN(_14120_));
 BUF_X2 _23817_ (.A(_14120_),
    .Z(_14121_));
 BUF_X4 _23818_ (.A(_14121_),
    .Z(_14122_));
 AND2_X2 _23819_ (.A1(_14092_),
    .A2(_14085_),
    .ZN(_14123_));
 AND2_X1 _23820_ (.A1(_14114_),
    .A2(_14084_),
    .ZN(_14124_));
 BUF_X4 _23821_ (.A(_14124_),
    .Z(_14125_));
 OAI21_X1 _23822_ (.A(_14122_),
    .B1(_14123_),
    .B2(_14125_),
    .ZN(_14126_));
 AND2_X1 _23823_ (.A1(_14068_),
    .A2(_14114_),
    .ZN(_14127_));
 BUF_X2 _23824_ (.A(_14127_),
    .Z(_14128_));
 OAI21_X1 _23825_ (.A(_14122_),
    .B1(_14070_),
    .B2(_14128_),
    .ZN(_14129_));
 INV_X1 _23826_ (.A(_14114_),
    .ZN(_14130_));
 NAND2_X1 _23827_ (.A1(_14130_),
    .A2(_14089_),
    .ZN(_14131_));
 NOR2_X1 _23828_ (.A1(_14131_),
    .A2(_14069_),
    .ZN(_14132_));
 INV_X1 _23829_ (.A(_14132_),
    .ZN(_14133_));
 INV_X1 _23830_ (.A(_14120_),
    .ZN(_14134_));
 OAI211_X2 _23831_ (.A(_14126_),
    .B(_14129_),
    .C1(_14133_),
    .C2(_14134_),
    .ZN(_14135_));
 NOR2_X1 _23832_ (.A1(_14118_),
    .A2(_17164_),
    .ZN(_14136_));
 AND2_X1 _23833_ (.A1(_14136_),
    .A2(_14073_),
    .ZN(_14137_));
 AND2_X1 _23834_ (.A1(_17161_),
    .A2(_17163_),
    .ZN(_14138_));
 AND2_X1 _23835_ (.A1(_14138_),
    .A2(_14088_),
    .ZN(_14139_));
 BUF_X2 _23836_ (.A(_14139_),
    .Z(_14140_));
 AND2_X1 _23837_ (.A1(_14137_),
    .A2(_14140_),
    .ZN(_14141_));
 BUF_X4 _23838_ (.A(_14096_),
    .Z(_14142_));
 AND4_X1 _23839_ (.A1(_14073_),
    .A2(_14136_),
    .A3(_14108_),
    .A4(_14142_),
    .ZN(_14143_));
 NOR2_X1 _23840_ (.A1(_14141_),
    .A2(_14143_),
    .ZN(_14144_));
 INV_X1 _23841_ (.A(_14085_),
    .ZN(_14145_));
 NOR2_X1 _23842_ (.A1(_14145_),
    .A2(_14114_),
    .ZN(_14146_));
 AND2_X1 _23843_ (.A1(_14137_),
    .A2(_14146_),
    .ZN(_14147_));
 INV_X1 _23844_ (.A(_14147_),
    .ZN(_14148_));
 BUF_X2 _23845_ (.A(_14137_),
    .Z(_14149_));
 BUF_X4 _23846_ (.A(_14090_),
    .Z(_14150_));
 NAND4_X1 _23847_ (.A1(_14149_),
    .A2(_14083_),
    .A3(_14130_),
    .A4(_14150_),
    .ZN(_14151_));
 AND2_X4 _23848_ (.A1(_14077_),
    .A2(_14069_),
    .ZN(_14152_));
 BUF_X2 _23849_ (.A(_14152_),
    .Z(_14153_));
 AND2_X2 _23850_ (.A1(_14138_),
    .A2(_17162_),
    .ZN(_14154_));
 BUF_X4 _23851_ (.A(_14154_),
    .Z(_14155_));
 OAI21_X1 _23852_ (.A(_14149_),
    .B1(_14153_),
    .B2(_14155_),
    .ZN(_14156_));
 NAND4_X1 _23853_ (.A1(_14144_),
    .A2(_14148_),
    .A3(_14151_),
    .A4(_14156_),
    .ZN(_14157_));
 NOR4_X1 _23854_ (.A1(_14095_),
    .A2(_14117_),
    .A3(_14135_),
    .A4(_14157_),
    .ZN(_14158_));
 BUF_X4 _23855_ (.A(_14119_),
    .Z(_14159_));
 INV_X1 _23856_ (.A(_17167_),
    .ZN(_14160_));
 NOR2_X1 _23857_ (.A1(_14160_),
    .A2(_17168_),
    .ZN(_14161_));
 BUF_X4 _23858_ (.A(_14161_),
    .Z(_14162_));
 NAND4_X1 _23859_ (.A1(_14159_),
    .A2(_14108_),
    .A3(_14162_),
    .A4(_11104_),
    .ZN(_14163_));
 AND2_X2 _23860_ (.A1(_14119_),
    .A2(_14162_),
    .ZN(_14164_));
 INV_X1 _23861_ (.A(_14164_),
    .ZN(_14165_));
 AND2_X2 _23862_ (.A1(_14077_),
    .A2(_14113_),
    .ZN(_14166_));
 INV_X1 _23863_ (.A(_14166_),
    .ZN(_14167_));
 OAI21_X1 _23864_ (.A(_14163_),
    .B1(_14165_),
    .B2(_14167_),
    .ZN(_14168_));
 INV_X1 _23865_ (.A(_14102_),
    .ZN(_14169_));
 INV_X1 _23866_ (.A(_14092_),
    .ZN(_14170_));
 NAND2_X1 _23867_ (.A1(_14170_),
    .A2(_14085_),
    .ZN(_14171_));
 AOI21_X1 _23868_ (.A(_14165_),
    .B1(_14169_),
    .B2(_14171_),
    .ZN(_14172_));
 BUF_X2 _23869_ (.A(_14098_),
    .Z(_14173_));
 AND2_X1 _23870_ (.A1(_14162_),
    .A2(_14173_),
    .ZN(_14174_));
 INV_X1 _23871_ (.A(_14174_),
    .ZN(_14175_));
 AND2_X2 _23872_ (.A1(_14089_),
    .A2(_14069_),
    .ZN(_14176_));
 INV_X1 _23873_ (.A(_14176_),
    .ZN(_14177_));
 AND2_X1 _23874_ (.A1(_14084_),
    .A2(_14091_),
    .ZN(_14178_));
 BUF_X2 _23875_ (.A(_14178_),
    .Z(_14179_));
 INV_X1 _23876_ (.A(_14179_),
    .ZN(_14180_));
 AOI21_X1 _23877_ (.A(_14175_),
    .B1(_14177_),
    .B2(_14180_),
    .ZN(_14181_));
 BUF_X4 _23878_ (.A(_14174_),
    .Z(_14182_));
 AND2_X1 _23879_ (.A1(_14092_),
    .A2(_14077_),
    .ZN(_14183_));
 BUF_X2 _23880_ (.A(_14183_),
    .Z(_14184_));
 AND2_X2 _23881_ (.A1(_14077_),
    .A2(_14091_),
    .ZN(_14185_));
 OAI21_X1 _23882_ (.A(_14182_),
    .B1(_14184_),
    .B2(_14185_),
    .ZN(_14186_));
 NAND4_X1 _23883_ (.A1(_14108_),
    .A2(_14162_),
    .A3(_11104_),
    .A4(_14173_),
    .ZN(_14187_));
 NAND2_X1 _23884_ (.A1(_14186_),
    .A2(_14187_),
    .ZN(_14188_));
 OR4_X1 _23885_ (.A1(_14168_),
    .A2(_14172_),
    .A3(_14181_),
    .A4(_14188_),
    .ZN(_14189_));
 AND2_X1 _23886_ (.A1(_14136_),
    .A2(_14161_),
    .ZN(_14190_));
 BUF_X4 _23887_ (.A(_14190_),
    .Z(_14191_));
 AND2_X2 _23888_ (.A1(_14089_),
    .A2(_14091_),
    .ZN(_14192_));
 AND2_X1 _23889_ (.A1(_14191_),
    .A2(_14192_),
    .ZN(_14193_));
 NAND2_X1 _23890_ (.A1(_14191_),
    .A2(_14184_),
    .ZN(_14194_));
 INV_X1 _23891_ (.A(_14190_),
    .ZN(_14195_));
 OAI21_X1 _23892_ (.A(_14068_),
    .B1(_11103_),
    .B2(_14091_),
    .ZN(_14196_));
 OAI21_X1 _23893_ (.A(_14194_),
    .B1(_14195_),
    .B2(_14196_),
    .ZN(_14197_));
 AND2_X2 _23894_ (.A1(_14089_),
    .A2(_14092_),
    .ZN(_14198_));
 NAND2_X1 _23895_ (.A1(_14198_),
    .A2(_14191_),
    .ZN(_14199_));
 AND2_X2 _23896_ (.A1(_14089_),
    .A2(_14114_),
    .ZN(_14200_));
 INV_X1 _23897_ (.A(_14200_),
    .ZN(_14201_));
 OAI21_X1 _23898_ (.A(_14199_),
    .B1(_14195_),
    .B2(_14201_),
    .ZN(_14202_));
 AND2_X2 _23899_ (.A1(_14096_),
    .A2(_14084_),
    .ZN(_14203_));
 NAND2_X1 _23900_ (.A1(_14191_),
    .A2(_14203_),
    .ZN(_14204_));
 INV_X1 _23901_ (.A(_14124_),
    .ZN(_14205_));
 OAI21_X1 _23902_ (.A(_14204_),
    .B1(_14195_),
    .B2(_14205_),
    .ZN(_14206_));
 OR4_X1 _23903_ (.A1(_14193_),
    .A2(_14197_),
    .A3(_14202_),
    .A4(_14206_),
    .ZN(_14207_));
 INV_X2 _23904_ (.A(_14112_),
    .ZN(_14208_));
 AND2_X2 _23905_ (.A1(_14161_),
    .A2(_14072_),
    .ZN(_14209_));
 BUF_X4 _23906_ (.A(_14209_),
    .Z(_14210_));
 NAND3_X1 _23907_ (.A1(_14208_),
    .A2(_14130_),
    .A3(_14210_),
    .ZN(_14211_));
 NAND2_X1 _23908_ (.A1(_14128_),
    .A2(_14210_),
    .ZN(_14212_));
 NAND2_X1 _23909_ (.A1(_14211_),
    .A2(_14212_),
    .ZN(_14213_));
 AND2_X1 _23910_ (.A1(_14069_),
    .A2(_14084_),
    .ZN(_14214_));
 BUF_X4 _23911_ (.A(_14214_),
    .Z(_14215_));
 OAI21_X1 _23912_ (.A(_14210_),
    .B1(_14203_),
    .B2(_14215_),
    .ZN(_14216_));
 AND2_X2 _23913_ (.A1(_14090_),
    .A2(_11103_),
    .ZN(_14217_));
 NAND2_X1 _23914_ (.A1(_14217_),
    .A2(_14210_),
    .ZN(_14218_));
 INV_X1 _23915_ (.A(_14209_),
    .ZN(_14219_));
 OAI211_X2 _23916_ (.A(_14216_),
    .B(_14218_),
    .C1(_14219_),
    .C2(_14205_),
    .ZN(_14220_));
 NOR4_X1 _23917_ (.A1(_14189_),
    .A2(_14207_),
    .A3(_14213_),
    .A4(_14220_),
    .ZN(_14221_));
 AND2_X2 _23918_ (.A1(_14160_),
    .A2(_17168_),
    .ZN(_14222_));
 AND2_X2 _23919_ (.A1(_14119_),
    .A2(_14222_),
    .ZN(_14223_));
 AND3_X1 _23920_ (.A1(_14223_),
    .A2(_14083_),
    .A3(_14146_),
    .ZN(_14224_));
 AOI21_X1 _23921_ (.A(_14224_),
    .B1(_14155_),
    .B2(_14223_),
    .ZN(_14225_));
 INV_X1 _23922_ (.A(_14089_),
    .ZN(_14226_));
 NOR2_X1 _23923_ (.A1(_14226_),
    .A2(_14092_),
    .ZN(_14227_));
 AND2_X1 _23924_ (.A1(_14222_),
    .A2(_14098_),
    .ZN(_14228_));
 NAND2_X1 _23925_ (.A1(_14227_),
    .A2(_14228_),
    .ZN(_14229_));
 BUF_X4 _23926_ (.A(_14222_),
    .Z(_14230_));
 BUF_X4 _23927_ (.A(_14081_),
    .Z(_14231_));
 BUF_X4 _23928_ (.A(_14085_),
    .Z(_14232_));
 NAND4_X1 _23929_ (.A1(_14230_),
    .A2(_14231_),
    .A3(_14173_),
    .A4(_14232_),
    .ZN(_14233_));
 BUF_X4 _23930_ (.A(_14228_),
    .Z(_14234_));
 AND2_X1 _23931_ (.A1(_14068_),
    .A2(_11103_),
    .ZN(_14235_));
 OAI21_X1 _23932_ (.A(_14234_),
    .B1(_14208_),
    .B2(_14235_),
    .ZN(_14236_));
 NAND4_X1 _23933_ (.A1(_14225_),
    .A2(_14229_),
    .A3(_14233_),
    .A4(_14236_),
    .ZN(_14237_));
 AND2_X1 _23934_ (.A1(_14222_),
    .A2(_14136_),
    .ZN(_14238_));
 BUF_X2 _23935_ (.A(_14238_),
    .Z(_14239_));
 BUF_X4 _23936_ (.A(_14185_),
    .Z(_14240_));
 OAI21_X1 _23937_ (.A(_14239_),
    .B1(_14240_),
    .B2(_14166_),
    .ZN(_14241_));
 NAND4_X1 _23938_ (.A1(_14230_),
    .A2(_14136_),
    .A3(_14108_),
    .A4(_14142_),
    .ZN(_14242_));
 NAND2_X1 _23939_ (.A1(_14241_),
    .A2(_14242_),
    .ZN(_14243_));
 AND2_X2 _23940_ (.A1(_14222_),
    .A2(_14071_),
    .ZN(_14244_));
 BUF_X4 _23941_ (.A(_14244_),
    .Z(_14245_));
 AND2_X1 _23942_ (.A1(_14227_),
    .A2(_14245_),
    .ZN(_14246_));
 NOR2_X1 _23943_ (.A1(_14145_),
    .A2(_14142_),
    .ZN(_14247_));
 AND2_X1 _23944_ (.A1(_14244_),
    .A2(_14247_),
    .ZN(_14248_));
 AND2_X1 _23945_ (.A1(_14244_),
    .A2(_14153_),
    .ZN(_14249_));
 OR3_X1 _23946_ (.A1(_14246_),
    .A2(_14248_),
    .A3(_14249_),
    .ZN(_14250_));
 AND2_X1 _23947_ (.A1(_14238_),
    .A2(_14176_),
    .ZN(_14251_));
 NOR4_X1 _23948_ (.A1(_14237_),
    .A2(_14243_),
    .A3(_14250_),
    .A4(_14251_),
    .ZN(_14252_));
 AND2_X4 _23949_ (.A1(_17167_),
    .A2(_17168_),
    .ZN(_14253_));
 BUF_X2 _23950_ (.A(_14253_),
    .Z(_14254_));
 AND2_X1 _23951_ (.A1(_14072_),
    .A2(_14254_),
    .ZN(_14255_));
 BUF_X4 _23952_ (.A(_14255_),
    .Z(_14256_));
 BUF_X4 _23953_ (.A(_14256_),
    .Z(_14257_));
 OAI21_X1 _23954_ (.A(_14257_),
    .B1(_14184_),
    .B2(_14109_),
    .ZN(_14258_));
 AND2_X1 _23955_ (.A1(_14254_),
    .A2(_14098_),
    .ZN(_14259_));
 BUF_X4 _23956_ (.A(_14259_),
    .Z(_14260_));
 BUF_X4 _23957_ (.A(_14078_),
    .Z(_14261_));
 BUF_X8 _23958_ (.A(_14091_),
    .Z(_14262_));
 OAI211_X2 _23959_ (.A(_14260_),
    .B(_14261_),
    .C1(_14231_),
    .C2(_14262_),
    .ZN(_14263_));
 NAND3_X1 _23960_ (.A1(_14260_),
    .A2(_14108_),
    .A3(_14142_),
    .ZN(_14264_));
 INV_X1 _23961_ (.A(_14260_),
    .ZN(_14265_));
 INV_X1 _23962_ (.A(_14127_),
    .ZN(_14266_));
 OAI211_X2 _23963_ (.A(_14263_),
    .B(_14264_),
    .C1(_14265_),
    .C2(_14266_),
    .ZN(_14267_));
 AND2_X2 _23964_ (.A1(_14119_),
    .A2(_14253_),
    .ZN(_14268_));
 INV_X1 _23965_ (.A(_14268_),
    .ZN(_14269_));
 INV_X1 _23966_ (.A(_14097_),
    .ZN(_14270_));
 INV_X1 _23967_ (.A(_14123_),
    .ZN(_14271_));
 AOI21_X1 _23968_ (.A(_14269_),
    .B1(_14270_),
    .B2(_14271_),
    .ZN(_14272_));
 INV_X1 _23969_ (.A(_14068_),
    .ZN(_14273_));
 OAI21_X1 _23970_ (.A(_14273_),
    .B1(_14112_),
    .B2(_14114_),
    .ZN(_14274_));
 BUF_X2 _23971_ (.A(_14268_),
    .Z(_14275_));
 AND2_X1 _23972_ (.A1(_14274_),
    .A2(_14275_),
    .ZN(_14276_));
 AND3_X1 _23973_ (.A1(_14259_),
    .A2(_14093_),
    .A3(_14085_),
    .ZN(_14277_));
 NOR4_X1 _23974_ (.A1(_14267_),
    .A2(_14272_),
    .A3(_14276_),
    .A4(_14277_),
    .ZN(_14278_));
 AND2_X2 _23975_ (.A1(_14136_),
    .A2(_14253_),
    .ZN(_14279_));
 BUF_X4 _23976_ (.A(_14279_),
    .Z(_14280_));
 INV_X1 _23977_ (.A(_14142_),
    .ZN(_14281_));
 AND4_X1 _23978_ (.A1(_14170_),
    .A2(_14280_),
    .A3(_14281_),
    .A4(_14232_),
    .ZN(_14282_));
 INV_X1 _23979_ (.A(_14280_),
    .ZN(_14283_));
 NAND2_X1 _23980_ (.A1(_14281_),
    .A2(_14068_),
    .ZN(_14284_));
 NOR2_X1 _23981_ (.A1(_14283_),
    .A2(_14284_),
    .ZN(_14285_));
 AND2_X1 _23982_ (.A1(_14192_),
    .A2(_14280_),
    .ZN(_14286_));
 AND2_X2 _23983_ (.A1(_14078_),
    .A2(_11103_),
    .ZN(_14287_));
 AND2_X1 _23984_ (.A1(_14280_),
    .A2(_14287_),
    .ZN(_14288_));
 NOR4_X1 _23985_ (.A1(_14282_),
    .A2(_14285_),
    .A3(_14286_),
    .A4(_14288_),
    .ZN(_14289_));
 AND2_X1 _23986_ (.A1(_14176_),
    .A2(_14255_),
    .ZN(_14290_));
 AND2_X2 _23987_ (.A1(_14203_),
    .A2(_14255_),
    .ZN(_14291_));
 AOI211_X4 _23988_ (.A(_14290_),
    .B(_14291_),
    .C1(_14105_),
    .C2(_14256_),
    .ZN(_14292_));
 AND4_X1 _23989_ (.A1(_14258_),
    .A2(_14278_),
    .A3(_14289_),
    .A4(_14292_),
    .ZN(_14293_));
 NAND4_X1 _23990_ (.A1(_14158_),
    .A2(_14221_),
    .A3(_14252_),
    .A4(_14293_),
    .ZN(_14294_));
 AND2_X1 _23991_ (.A1(_14103_),
    .A2(_14215_),
    .ZN(_14295_));
 NOR2_X1 _23992_ (.A1(_14294_),
    .A2(_14295_),
    .ZN(_14296_));
 INV_X1 _23993_ (.A(_00988_),
    .ZN(_14297_));
 XNOR2_X1 _23994_ (.A(_14296_),
    .B(_14297_),
    .ZN(_14298_));
 MUX2_X1 _23995_ (.A(_01325_),
    .B(_14298_),
    .S(_03749_),
    .Z(_01058_));
 AND2_X1 _23996_ (.A1(_14090_),
    .A2(_14081_),
    .ZN(_14299_));
 OAI21_X1 _23997_ (.A(_14121_),
    .B1(_14299_),
    .B2(_14179_),
    .ZN(_14300_));
 AND2_X1 _23998_ (.A1(_14139_),
    .A2(_14099_),
    .ZN(_14301_));
 INV_X1 _23999_ (.A(_14183_),
    .ZN(_14302_));
 AOI21_X1 _24000_ (.A(_14111_),
    .B1(_14302_),
    .B2(_14167_),
    .ZN(_14303_));
 AOI211_X4 _24001_ (.A(_14301_),
    .B(_14303_),
    .C1(_14185_),
    .C2(_14100_),
    .ZN(_14304_));
 AND3_X1 _24002_ (.A1(_14100_),
    .A2(_14069_),
    .A3(_14090_),
    .ZN(_14305_));
 AND3_X1 _24003_ (.A1(_14100_),
    .A2(_14090_),
    .A3(_14093_),
    .ZN(_14306_));
 NOR4_X1 _24004_ (.A1(_14101_),
    .A2(_14305_),
    .A3(_14306_),
    .A4(_14106_),
    .ZN(_14307_));
 OAI21_X1 _24005_ (.A(_14121_),
    .B1(_14184_),
    .B2(_14140_),
    .ZN(_14308_));
 AND4_X1 _24006_ (.A1(_14300_),
    .A2(_14304_),
    .A3(_14307_),
    .A4(_14308_),
    .ZN(_14309_));
 NOR3_X1 _24007_ (.A1(_17164_),
    .A2(_17167_),
    .A3(_17168_),
    .ZN(_14310_));
 NAND3_X1 _24008_ (.A1(_14130_),
    .A2(_14310_),
    .A3(_14090_),
    .ZN(_14311_));
 NOR2_X1 _24009_ (.A1(_14311_),
    .A2(_14118_),
    .ZN(_14312_));
 INV_X1 _24010_ (.A(_14312_),
    .ZN(_14313_));
 NAND2_X1 _24011_ (.A1(_14149_),
    .A2(_14247_),
    .ZN(_14314_));
 AOI211_X4 _24012_ (.A(_14079_),
    .B(_14080_),
    .C1(_11104_),
    .C2(_11111_),
    .ZN(_14315_));
 OAI211_X2 _24013_ (.A(_14075_),
    .B(_14108_),
    .C1(_11104_),
    .C2(_14262_),
    .ZN(_14316_));
 INV_X1 _24014_ (.A(_14316_),
    .ZN(_14317_));
 AND3_X1 _24015_ (.A1(_14075_),
    .A2(_11104_),
    .A3(_14090_),
    .ZN(_14318_));
 NOR4_X1 _24016_ (.A1(_14315_),
    .A2(_14317_),
    .A3(_14087_),
    .A4(_14318_),
    .ZN(_14319_));
 NAND4_X1 _24017_ (.A1(_14309_),
    .A2(_14313_),
    .A3(_14314_),
    .A4(_14319_),
    .ZN(_14320_));
 INV_X1 _24018_ (.A(_14215_),
    .ZN(_14321_));
 NAND2_X1 _24019_ (.A1(_14205_),
    .A2(_14321_),
    .ZN(_14322_));
 OAI21_X1 _24020_ (.A(_14260_),
    .B1(_14322_),
    .B2(_14217_),
    .ZN(_14323_));
 OAI211_X2 _24021_ (.A(_14260_),
    .B(_14078_),
    .C1(_14231_),
    .C2(_11111_),
    .ZN(_14324_));
 OAI211_X2 _24022_ (.A(_14323_),
    .B(_14324_),
    .C1(_14265_),
    .C2(_14266_),
    .ZN(_14325_));
 AND2_X1 _24023_ (.A1(_14067_),
    .A2(_14092_),
    .ZN(_14326_));
 BUF_X2 _24024_ (.A(_14326_),
    .Z(_14327_));
 AND2_X1 _24025_ (.A1(_14327_),
    .A2(_14279_),
    .ZN(_14328_));
 AND2_X1 _24026_ (.A1(_14279_),
    .A2(_14152_),
    .ZN(_14329_));
 AND3_X1 _24027_ (.A1(_14166_),
    .A2(_14136_),
    .A3(_14254_),
    .ZN(_14330_));
 OR2_X4 _24028_ (.A1(_14329_),
    .A2(_14330_),
    .ZN(_14331_));
 AND2_X2 _24029_ (.A1(_14067_),
    .A2(_14091_),
    .ZN(_14332_));
 AND2_X1 _24030_ (.A1(_14332_),
    .A2(_14279_),
    .ZN(_14333_));
 AND2_X1 _24031_ (.A1(_14198_),
    .A2(_14279_),
    .ZN(_14334_));
 OR4_X2 _24032_ (.A1(_14328_),
    .A2(_14331_),
    .A3(_14333_),
    .A4(_14334_),
    .ZN(_14335_));
 AND2_X1 _24033_ (.A1(_14268_),
    .A2(_14326_),
    .ZN(_14336_));
 NAND2_X1 _24034_ (.A1(_14268_),
    .A2(_14102_),
    .ZN(_14337_));
 OAI21_X1 _24035_ (.A(_14337_),
    .B1(_14269_),
    .B2(_14270_),
    .ZN(_14338_));
 NAND2_X1 _24036_ (.A1(_14268_),
    .A2(_14166_),
    .ZN(_14339_));
 NAND2_X1 _24037_ (.A1(_14268_),
    .A2(_14152_),
    .ZN(_14340_));
 NAND2_X1 _24038_ (.A1(_14339_),
    .A2(_14340_),
    .ZN(_14341_));
 AND4_X1 _24039_ (.A1(_11103_),
    .A2(_14119_),
    .A3(_14254_),
    .A4(_14085_),
    .ZN(_14342_));
 OR4_X1 _24040_ (.A1(_14336_),
    .A2(_14338_),
    .A3(_14341_),
    .A4(_14342_),
    .ZN(_14343_));
 NAND2_X1 _24041_ (.A1(_14128_),
    .A2(_14256_),
    .ZN(_14344_));
 NAND2_X1 _24042_ (.A1(_14198_),
    .A2(_14256_),
    .ZN(_14345_));
 NAND2_X1 _24043_ (.A1(_14192_),
    .A2(_14256_),
    .ZN(_14346_));
 NAND2_X1 _24044_ (.A1(_14256_),
    .A2(_14154_),
    .ZN(_14347_));
 NAND4_X1 _24045_ (.A1(_14344_),
    .A2(_14345_),
    .A3(_14346_),
    .A4(_14347_),
    .ZN(_14348_));
 OR4_X1 _24046_ (.A1(_14325_),
    .A2(_14335_),
    .A3(_14343_),
    .A4(_14348_),
    .ZN(_14349_));
 INV_X1 _24047_ (.A(_14131_),
    .ZN(_14350_));
 AND2_X1 _24048_ (.A1(_14085_),
    .A2(_11103_),
    .ZN(_14351_));
 OAI21_X1 _24049_ (.A(_14182_),
    .B1(_14350_),
    .B2(_14351_),
    .ZN(_14352_));
 OAI211_X2 _24050_ (.A(_14182_),
    .B(_14078_),
    .C1(_14093_),
    .C2(_14142_),
    .ZN(_14353_));
 OAI211_X2 _24051_ (.A(_14352_),
    .B(_14353_),
    .C1(_14273_),
    .C2(_14175_),
    .ZN(_14354_));
 BUF_X4 _24052_ (.A(_14164_),
    .Z(_14355_));
 OAI21_X1 _24053_ (.A(_14355_),
    .B1(_14200_),
    .B2(_14215_),
    .ZN(_14356_));
 OAI21_X1 _24054_ (.A(_14355_),
    .B1(_14153_),
    .B2(_14166_),
    .ZN(_14357_));
 NAND2_X1 _24055_ (.A1(_14164_),
    .A2(_14332_),
    .ZN(_14358_));
 NAND3_X1 _24056_ (.A1(_14327_),
    .A2(_14159_),
    .A3(_14162_),
    .ZN(_14359_));
 NAND4_X1 _24057_ (.A1(_14356_),
    .A2(_14357_),
    .A3(_14358_),
    .A4(_14359_),
    .ZN(_14360_));
 OAI21_X1 _24058_ (.A(_14191_),
    .B1(_14184_),
    .B2(_14140_),
    .ZN(_14361_));
 INV_X1 _24059_ (.A(_14086_),
    .ZN(_14362_));
 NAND2_X1 _24060_ (.A1(_14362_),
    .A2(_14191_),
    .ZN(_14363_));
 INV_X1 _24061_ (.A(_14299_),
    .ZN(_14364_));
 OAI211_X2 _24062_ (.A(_14361_),
    .B(_14363_),
    .C1(_14364_),
    .C2(_14195_),
    .ZN(_14365_));
 OAI21_X1 _24063_ (.A(_14209_),
    .B1(_14203_),
    .B2(_14125_),
    .ZN(_14366_));
 NAND4_X1 _24064_ (.A1(_14209_),
    .A2(_14083_),
    .A3(_14130_),
    .A4(_14068_),
    .ZN(_14367_));
 NAND2_X1 _24065_ (.A1(_14208_),
    .A2(_14209_),
    .ZN(_14368_));
 NAND4_X1 _24066_ (.A1(_14090_),
    .A2(_14162_),
    .A3(_14069_),
    .A4(_14072_),
    .ZN(_14369_));
 NAND4_X1 _24067_ (.A1(_14366_),
    .A2(_14367_),
    .A3(_14368_),
    .A4(_14369_),
    .ZN(_14370_));
 OR4_X1 _24068_ (.A1(_14354_),
    .A2(_14360_),
    .A3(_14365_),
    .A4(_14370_),
    .ZN(_14371_));
 AND2_X1 _24069_ (.A1(_14244_),
    .A2(_14183_),
    .ZN(_14372_));
 AND2_X1 _24070_ (.A1(_14244_),
    .A2(_14185_),
    .ZN(_14373_));
 AOI221_X4 _24071_ (.A(_14372_),
    .B1(_14244_),
    .B2(_14235_),
    .C1(_11104_),
    .C2(_14373_),
    .ZN(_14374_));
 AND2_X1 _24072_ (.A1(_14232_),
    .A2(_14081_),
    .ZN(_14375_));
 OAI21_X1 _24073_ (.A(_14245_),
    .B1(_14198_),
    .B2(_14375_),
    .ZN(_14376_));
 AND2_X1 _24074_ (.A1(_14374_),
    .A2(_14376_),
    .ZN(_14377_));
 AND2_X1 _24075_ (.A1(_14228_),
    .A2(_14166_),
    .ZN(_14378_));
 NAND4_X1 _24076_ (.A1(_14222_),
    .A2(_14173_),
    .A3(_14092_),
    .A4(_14085_),
    .ZN(_14379_));
 NAND2_X1 _24077_ (.A1(_14229_),
    .A2(_14379_),
    .ZN(_14380_));
 INV_X2 _24078_ (.A(_14326_),
    .ZN(_14381_));
 AND2_X1 _24079_ (.A1(_14068_),
    .A2(_14096_),
    .ZN(_14382_));
 INV_X1 _24080_ (.A(_14382_),
    .ZN(_14383_));
 NAND2_X1 _24081_ (.A1(_14381_),
    .A2(_14383_),
    .ZN(_14384_));
 AOI211_X4 _24082_ (.A(_14378_),
    .B(_14380_),
    .C1(_14228_),
    .C2(_14384_),
    .ZN(_14385_));
 AND2_X1 _24083_ (.A1(_14223_),
    .A2(_14332_),
    .ZN(_14386_));
 INV_X1 _24084_ (.A(_14223_),
    .ZN(_14387_));
 INV_X1 _24085_ (.A(_14192_),
    .ZN(_14388_));
 AOI21_X1 _24086_ (.A(_14387_),
    .B1(_14388_),
    .B2(_14271_),
    .ZN(_14389_));
 AOI211_X4 _24087_ (.A(_14386_),
    .B(_14389_),
    .C1(_14261_),
    .C2(_14223_),
    .ZN(_14390_));
 AND2_X1 _24088_ (.A1(_14239_),
    .A2(_14105_),
    .ZN(_14391_));
 INV_X1 _24089_ (.A(_14196_),
    .ZN(_14392_));
 AND2_X1 _24090_ (.A1(_14392_),
    .A2(_14239_),
    .ZN(_14393_));
 BUF_X2 _24091_ (.A(_14097_),
    .Z(_14394_));
 AND2_X1 _24092_ (.A1(_14238_),
    .A2(_14394_),
    .ZN(_14395_));
 AND2_X1 _24093_ (.A1(_14238_),
    .A2(_14203_),
    .ZN(_14396_));
 NOR4_X1 _24094_ (.A1(_14391_),
    .A2(_14393_),
    .A3(_14395_),
    .A4(_14396_),
    .ZN(_14397_));
 NAND4_X1 _24095_ (.A1(_14377_),
    .A2(_14385_),
    .A3(_14390_),
    .A4(_14397_),
    .ZN(_14398_));
 OR4_X2 _24096_ (.A1(_14320_),
    .A2(_14349_),
    .A3(_14371_),
    .A4(_14398_),
    .ZN(_14399_));
 NOR2_X2 _24097_ (.A1(_14399_),
    .A2(_14295_),
    .ZN(_14400_));
 INV_X1 _24098_ (.A(_00989_),
    .ZN(_14401_));
 XNOR2_X1 _24099_ (.A(_14400_),
    .B(_14401_),
    .ZN(_14402_));
 BUF_X4 _24100_ (.A(_03738_),
    .Z(_14403_));
 MUX2_X1 _24101_ (.A(_01326_),
    .B(_14402_),
    .S(_14403_),
    .Z(_01069_));
 XOR2_X1 _24102_ (.A(_17270_),
    .B(_17074_),
    .Z(_14404_));
 XNOR2_X1 _24103_ (.A(_11387_),
    .B(_11857_),
    .ZN(_14405_));
 XOR2_X1 _24104_ (.A(_14014_),
    .B(_00990_),
    .Z(_14406_));
 XOR2_X1 _24105_ (.A(_14405_),
    .B(_14406_),
    .Z(_14407_));
 XNOR2_X1 _24106_ (.A(_14407_),
    .B(_12584_),
    .ZN(_14408_));
 MUX2_X1 _24107_ (.A(_14404_),
    .B(_14408_),
    .S(_11149_),
    .Z(_00684_));
 AND2_X1 _24108_ (.A1(_14223_),
    .A2(_14105_),
    .ZN(_14409_));
 INV_X1 _24109_ (.A(_14409_),
    .ZN(_14410_));
 AND3_X1 _24110_ (.A1(_14127_),
    .A2(_14159_),
    .A3(_14230_),
    .ZN(_14411_));
 AOI211_X4 _24111_ (.A(_14411_),
    .B(_14386_),
    .C1(_14240_),
    .C2(_14223_),
    .ZN(_14412_));
 OAI211_X2 _24112_ (.A(_14234_),
    .B(_11127_),
    .C1(_17162_),
    .C2(_14170_),
    .ZN(_14413_));
 OAI211_X2 _24113_ (.A(_14173_),
    .B(_14230_),
    .C1(_14240_),
    .C2(_14109_),
    .ZN(_14414_));
 AND4_X1 _24114_ (.A1(_14410_),
    .A2(_14412_),
    .A3(_14413_),
    .A4(_14414_),
    .ZN(_14415_));
 OAI21_X1 _24115_ (.A(_14260_),
    .B1(_14327_),
    .B2(_14235_),
    .ZN(_14416_));
 NAND3_X1 _24116_ (.A1(_14240_),
    .A2(_14260_),
    .A3(_11105_),
    .ZN(_14417_));
 AND2_X1 _24117_ (.A1(_14416_),
    .A2(_14417_),
    .ZN(_14418_));
 INV_X1 _24118_ (.A(_14336_),
    .ZN(_14419_));
 AND2_X1 _24119_ (.A1(_14268_),
    .A2(_14154_),
    .ZN(_14420_));
 INV_X1 _24120_ (.A(_14420_),
    .ZN(_14421_));
 AND2_X1 _24121_ (.A1(_14268_),
    .A2(_14382_),
    .ZN(_14422_));
 INV_X1 _24122_ (.A(_14422_),
    .ZN(_14423_));
 AND4_X1 _24123_ (.A1(_14419_),
    .A2(_14421_),
    .A3(_14423_),
    .A4(_14340_),
    .ZN(_14424_));
 AND2_X1 _24124_ (.A1(_14259_),
    .A2(_14124_),
    .ZN(_14425_));
 AND3_X1 _24125_ (.A1(_14150_),
    .A2(_14173_),
    .A3(_14254_),
    .ZN(_14426_));
 NOR3_X1 _24126_ (.A1(_14277_),
    .A2(_14425_),
    .A3(_14426_),
    .ZN(_14427_));
 NAND2_X1 _24127_ (.A1(_14275_),
    .A2(_14105_),
    .ZN(_14428_));
 NAND3_X1 _24128_ (.A1(_14203_),
    .A2(_14159_),
    .A3(_14254_),
    .ZN(_14429_));
 AND3_X1 _24129_ (.A1(_14428_),
    .A2(_14337_),
    .A3(_14429_),
    .ZN(_14430_));
 AND4_X1 _24130_ (.A1(_14418_),
    .A2(_14424_),
    .A3(_14427_),
    .A4(_14430_),
    .ZN(_14431_));
 OAI21_X1 _24131_ (.A(_14239_),
    .B1(_14394_),
    .B2(_14102_),
    .ZN(_14432_));
 INV_X1 _24132_ (.A(_14245_),
    .ZN(_14433_));
 INV_X1 _24133_ (.A(_14332_),
    .ZN(_14434_));
 AOI21_X1 _24134_ (.A(_14433_),
    .B1(_14381_),
    .B2(_14434_),
    .ZN(_14435_));
 NOR3_X1 _24135_ (.A1(_14435_),
    .A2(_14249_),
    .A3(_14372_),
    .ZN(_14436_));
 OAI21_X1 _24136_ (.A(_14239_),
    .B1(_14115_),
    .B2(_14327_),
    .ZN(_14437_));
 OAI21_X1 _24137_ (.A(_14245_),
    .B1(_14350_),
    .B2(_14247_),
    .ZN(_14438_));
 AND4_X1 _24138_ (.A1(_14432_),
    .A2(_14436_),
    .A3(_14437_),
    .A4(_14438_),
    .ZN(_14439_));
 OAI21_X1 _24139_ (.A(_14257_),
    .B1(_14327_),
    .B2(_14128_),
    .ZN(_14440_));
 NAND4_X1 _24140_ (.A1(_14257_),
    .A2(_14170_),
    .A3(_14281_),
    .A4(_14232_),
    .ZN(_14441_));
 NAND4_X1 _24141_ (.A1(_14261_),
    .A2(_14072_),
    .A3(_14254_),
    .A4(_11105_),
    .ZN(_14442_));
 NAND4_X1 _24142_ (.A1(_14440_),
    .A2(_14346_),
    .A3(_14441_),
    .A4(_14442_),
    .ZN(_14443_));
 AOI21_X1 _24143_ (.A(_14283_),
    .B1(_14381_),
    .B2(_14383_),
    .ZN(_14444_));
 NAND2_X1 _24144_ (.A1(_14170_),
    .A2(_14078_),
    .ZN(_14445_));
 NOR2_X1 _24145_ (.A1(_14283_),
    .A2(_14445_),
    .ZN(_14446_));
 AND2_X1 _24146_ (.A1(_14102_),
    .A2(_14279_),
    .ZN(_14447_));
 NOR4_X1 _24147_ (.A1(_14443_),
    .A2(_14444_),
    .A3(_14446_),
    .A4(_14447_),
    .ZN(_14448_));
 NAND4_X1 _24148_ (.A1(_14415_),
    .A2(_14431_),
    .A3(_14439_),
    .A4(_14448_),
    .ZN(_14449_));
 BUF_X4 _24149_ (.A(_14191_),
    .Z(_14450_));
 NOR2_X1 _24150_ (.A1(_14284_),
    .A2(_14093_),
    .ZN(_14451_));
 OAI21_X1 _24151_ (.A(_14450_),
    .B1(_14451_),
    .B2(_14115_),
    .ZN(_14452_));
 AND2_X1 _24152_ (.A1(_14191_),
    .A2(_14200_),
    .ZN(_14453_));
 AOI221_X4 _24153_ (.A(_14453_),
    .B1(_14450_),
    .B2(_14203_),
    .C1(_11105_),
    .C2(_14193_),
    .ZN(_14454_));
 OAI21_X1 _24154_ (.A(_14210_),
    .B1(_14217_),
    .B2(_14125_),
    .ZN(_14455_));
 OAI211_X2 _24155_ (.A(_14210_),
    .B(_14262_),
    .C1(_14287_),
    .C2(_14109_),
    .ZN(_14456_));
 AND4_X1 _24156_ (.A1(_14452_),
    .A2(_14454_),
    .A3(_14455_),
    .A4(_14456_),
    .ZN(_14457_));
 AND3_X1 _24157_ (.A1(_14103_),
    .A2(_14108_),
    .A3(_14093_),
    .ZN(_14458_));
 AND3_X1 _24158_ (.A1(_14100_),
    .A2(_14078_),
    .A3(_14170_),
    .ZN(_14459_));
 OR2_X1 _24159_ (.A1(_14458_),
    .A2(_14459_),
    .ZN(_14460_));
 OAI21_X1 _24160_ (.A(_14122_),
    .B1(_14198_),
    .B2(_14125_),
    .ZN(_14461_));
 NAND2_X1 _24161_ (.A1(_14122_),
    .A2(_14128_),
    .ZN(_14462_));
 NAND2_X1 _24162_ (.A1(_14122_),
    .A2(_14332_),
    .ZN(_14463_));
 NAND2_X1 _24163_ (.A1(_14122_),
    .A2(_14240_),
    .ZN(_14464_));
 NAND4_X1 _24164_ (.A1(_14461_),
    .A2(_14462_),
    .A3(_14463_),
    .A4(_14464_),
    .ZN(_14465_));
 AND3_X1 _24165_ (.A1(_14146_),
    .A2(_14083_),
    .A3(_14103_),
    .ZN(_14466_));
 NOR4_X1 _24166_ (.A1(_14460_),
    .A2(_14465_),
    .A3(_14104_),
    .A4(_14466_),
    .ZN(_14467_));
 OAI21_X1 _24167_ (.A(_14075_),
    .B1(_14070_),
    .B2(_14287_),
    .ZN(_14468_));
 NAND4_X1 _24168_ (.A1(_14075_),
    .A2(_14083_),
    .A3(_14130_),
    .A4(_14150_),
    .ZN(_14469_));
 OAI211_X2 _24169_ (.A(_14468_),
    .B(_14469_),
    .C1(_14080_),
    .C2(_14180_),
    .ZN(_14470_));
 NAND4_X1 _24170_ (.A1(_14136_),
    .A2(_14109_),
    .A3(_14093_),
    .A4(_14073_),
    .ZN(_14471_));
 NAND4_X1 _24171_ (.A1(_14136_),
    .A2(_14261_),
    .A3(_14114_),
    .A4(_14073_),
    .ZN(_14472_));
 INV_X1 _24172_ (.A(_14149_),
    .ZN(_14473_));
 OAI211_X2 _24173_ (.A(_14471_),
    .B(_14472_),
    .C1(_14473_),
    .C2(_14434_),
    .ZN(_14474_));
 AOI21_X1 _24174_ (.A(_14473_),
    .B1(_14169_),
    .B2(_14388_),
    .ZN(_14475_));
 NOR2_X1 _24175_ (.A1(_14473_),
    .A2(_14171_),
    .ZN(_14476_));
 NOR4_X1 _24176_ (.A1(_14470_),
    .A2(_14474_),
    .A3(_14475_),
    .A4(_14476_),
    .ZN(_14477_));
 OAI21_X1 _24177_ (.A(_14182_),
    .B1(_14394_),
    .B2(_14123_),
    .ZN(_14478_));
 OAI21_X1 _24178_ (.A(_14355_),
    .B1(_14394_),
    .B2(_14125_),
    .ZN(_14479_));
 OAI21_X1 _24179_ (.A(_14355_),
    .B1(_14327_),
    .B2(_14287_),
    .ZN(_14480_));
 OAI21_X1 _24180_ (.A(_14182_),
    .B1(_14327_),
    .B2(_14155_),
    .ZN(_14481_));
 AND4_X1 _24181_ (.A1(_14478_),
    .A2(_14479_),
    .A3(_14480_),
    .A4(_14481_),
    .ZN(_14482_));
 NAND4_X1 _24182_ (.A1(_14457_),
    .A2(_14467_),
    .A3(_14477_),
    .A4(_14482_),
    .ZN(_14483_));
 NOR2_X1 _24183_ (.A1(_14449_),
    .A2(_14483_),
    .ZN(_14484_));
 XOR2_X1 _24184_ (.A(_14484_),
    .B(_00991_),
    .Z(_14485_));
 MUX2_X1 _24185_ (.A(_01327_),
    .B(_14485_),
    .S(_14403_),
    .Z(_01080_));
 NAND4_X1 _24186_ (.A1(_14230_),
    .A2(_11105_),
    .A3(_14072_),
    .A4(_14232_),
    .ZN(_14486_));
 AND4_X1 _24187_ (.A1(_14068_),
    .A2(_14244_),
    .A3(_14170_),
    .A4(_14281_),
    .ZN(_14487_));
 AOI221_X4 _24188_ (.A(_14487_),
    .B1(_11105_),
    .B2(_14373_),
    .C1(_14155_),
    .C2(_14245_),
    .ZN(_14488_));
 OAI211_X2 _24189_ (.A(_14245_),
    .B(_14150_),
    .C1(_14231_),
    .C2(_11111_),
    .ZN(_14489_));
 INV_X1 _24190_ (.A(_14238_),
    .ZN(_14490_));
 AOI21_X1 _24191_ (.A(_14490_),
    .B1(_14167_),
    .B2(_14381_),
    .ZN(_14491_));
 AND2_X1 _24192_ (.A1(_14238_),
    .A2(_14200_),
    .ZN(_14492_));
 NOR4_X1 _24193_ (.A1(_14491_),
    .A2(_14251_),
    .A3(_14391_),
    .A4(_14492_),
    .ZN(_14493_));
 AND4_X1 _24194_ (.A1(_14486_),
    .A2(_14488_),
    .A3(_14489_),
    .A4(_14493_),
    .ZN(_14494_));
 AND2_X1 _24195_ (.A1(_14234_),
    .A2(_14140_),
    .ZN(_14495_));
 INV_X1 _24196_ (.A(_14495_),
    .ZN(_14496_));
 AND2_X1 _24197_ (.A1(_14142_),
    .A2(_14078_),
    .ZN(_14497_));
 BUF_X4 _24198_ (.A(_14497_),
    .Z(_14498_));
 OAI21_X1 _24199_ (.A(_14234_),
    .B1(_14184_),
    .B2(_14498_),
    .ZN(_14499_));
 INV_X1 _24200_ (.A(_14171_),
    .ZN(_14500_));
 OAI21_X1 _24201_ (.A(_14234_),
    .B1(_14500_),
    .B2(_14176_),
    .ZN(_14501_));
 AND3_X1 _24202_ (.A1(_14496_),
    .A2(_14499_),
    .A3(_14501_),
    .ZN(_14502_));
 INV_X1 _24203_ (.A(_14384_),
    .ZN(_14503_));
 AOI21_X1 _24204_ (.A(_14387_),
    .B1(_14503_),
    .B2(_14079_),
    .ZN(_14504_));
 AOI211_X4 _24205_ (.A(_14409_),
    .B(_14504_),
    .C1(_14217_),
    .C2(_14223_),
    .ZN(_14505_));
 NAND2_X1 _24206_ (.A1(_14275_),
    .A2(_14128_),
    .ZN(_14506_));
 OAI21_X1 _24207_ (.A(_14275_),
    .B1(_14176_),
    .B2(_14200_),
    .ZN(_14507_));
 NAND4_X1 _24208_ (.A1(_14421_),
    .A2(_14506_),
    .A3(_14429_),
    .A4(_14507_),
    .ZN(_14508_));
 OAI211_X2 _24209_ (.A(_14280_),
    .B(_14150_),
    .C1(_14231_),
    .C2(_14262_),
    .ZN(_14509_));
 OAI211_X2 _24210_ (.A(_14280_),
    .B(_14232_),
    .C1(_14093_),
    .C2(_14142_),
    .ZN(_14510_));
 OAI211_X2 _24211_ (.A(_14280_),
    .B(_14109_),
    .C1(_11105_),
    .C2(_14262_),
    .ZN(_14511_));
 OAI21_X1 _24212_ (.A(_14280_),
    .B1(_14153_),
    .B2(_14155_),
    .ZN(_14512_));
 NAND4_X1 _24213_ (.A1(_14509_),
    .A2(_14510_),
    .A3(_14511_),
    .A4(_14512_),
    .ZN(_14513_));
 BUF_X4 _24214_ (.A(_14260_),
    .Z(_14514_));
 OAI21_X1 _24215_ (.A(_14514_),
    .B1(_14240_),
    .B2(_14155_),
    .ZN(_14515_));
 OAI211_X2 _24216_ (.A(_14514_),
    .B(_14109_),
    .C1(_11105_),
    .C2(_14262_),
    .ZN(_14516_));
 OAI21_X1 _24217_ (.A(_14514_),
    .B1(_14125_),
    .B2(_14179_),
    .ZN(_14517_));
 NAND2_X1 _24218_ (.A1(_14176_),
    .A2(_14514_),
    .ZN(_14518_));
 NAND4_X1 _24219_ (.A1(_14515_),
    .A2(_14516_),
    .A3(_14517_),
    .A4(_14518_),
    .ZN(_14519_));
 OAI211_X2 _24220_ (.A(_14257_),
    .B(_14109_),
    .C1(_11105_),
    .C2(_11111_),
    .ZN(_14520_));
 OAI211_X2 _24221_ (.A(_14257_),
    .B(_14150_),
    .C1(_14069_),
    .C2(_14114_),
    .ZN(_14521_));
 NAND3_X1 _24222_ (.A1(_14257_),
    .A2(_14261_),
    .A3(_14093_),
    .ZN(_14522_));
 OAI21_X1 _24223_ (.A(_14257_),
    .B1(_14215_),
    .B2(_14105_),
    .ZN(_14523_));
 NAND4_X1 _24224_ (.A1(_14520_),
    .A2(_14521_),
    .A3(_14522_),
    .A4(_14523_),
    .ZN(_14524_));
 NOR4_X1 _24225_ (.A1(_14508_),
    .A2(_14513_),
    .A3(_14519_),
    .A4(_14524_),
    .ZN(_14525_));
 NAND4_X1 _24226_ (.A1(_14494_),
    .A2(_14502_),
    .A3(_14505_),
    .A4(_14525_),
    .ZN(_14526_));
 OAI21_X1 _24227_ (.A(_14103_),
    .B1(_14132_),
    .B2(_14351_),
    .ZN(_14527_));
 AND2_X1 _24228_ (.A1(_14152_),
    .A2(_14100_),
    .ZN(_14528_));
 AND2_X1 _24229_ (.A1(_14184_),
    .A2(_14100_),
    .ZN(_14529_));
 AOI211_X4 _24230_ (.A(_14528_),
    .B(_14529_),
    .C1(_14103_),
    .C2(_14128_),
    .ZN(_14530_));
 OAI21_X1 _24231_ (.A(_14122_),
    .B1(_14192_),
    .B2(_14247_),
    .ZN(_14531_));
 NAND2_X1 _24232_ (.A1(_14122_),
    .A2(_14153_),
    .ZN(_14532_));
 AND2_X1 _24233_ (.A1(_14129_),
    .A2(_14532_),
    .ZN(_14533_));
 AND4_X1 _24234_ (.A1(_14527_),
    .A2(_14530_),
    .A3(_14531_),
    .A4(_14533_),
    .ZN(_14534_));
 OAI21_X1 _24235_ (.A(_14450_),
    .B1(_14362_),
    .B2(_14394_),
    .ZN(_14535_));
 OAI21_X1 _24236_ (.A(_14450_),
    .B1(_14498_),
    .B2(_14155_),
    .ZN(_14536_));
 NAND2_X1 _24237_ (.A1(_14450_),
    .A2(_14235_),
    .ZN(_14537_));
 AND2_X1 _24238_ (.A1(_14536_),
    .A2(_14537_),
    .ZN(_14538_));
 OAI21_X1 _24239_ (.A(_14210_),
    .B1(_14132_),
    .B2(_14125_),
    .ZN(_14539_));
 AND2_X1 _24240_ (.A1(_14108_),
    .A2(_14231_),
    .ZN(_14540_));
 OAI21_X1 _24241_ (.A(_14210_),
    .B1(_14498_),
    .B2(_14540_),
    .ZN(_14541_));
 AND4_X1 _24242_ (.A1(_14535_),
    .A2(_14538_),
    .A3(_14539_),
    .A4(_14541_),
    .ZN(_14542_));
 NAND2_X1 _24243_ (.A1(_14355_),
    .A2(_14261_),
    .ZN(_14543_));
 INV_X1 _24244_ (.A(_14140_),
    .ZN(_14544_));
 OAI211_X2 _24245_ (.A(_14358_),
    .B(_14543_),
    .C1(_14165_),
    .C2(_14544_),
    .ZN(_14545_));
 OAI211_X2 _24246_ (.A(_14182_),
    .B(_14232_),
    .C1(_14231_),
    .C2(_11111_),
    .ZN(_14546_));
 OAI21_X1 _24247_ (.A(_14546_),
    .B1(_14131_),
    .B2(_14175_),
    .ZN(_14547_));
 NAND2_X1 _24248_ (.A1(_14355_),
    .A2(_14217_),
    .ZN(_14548_));
 OAI21_X1 _24249_ (.A(_14548_),
    .B1(_14165_),
    .B2(_14205_),
    .ZN(_14549_));
 AND2_X1 _24250_ (.A1(_14077_),
    .A2(_14081_),
    .ZN(_14550_));
 INV_X1 _24251_ (.A(_14550_),
    .ZN(_14551_));
 AOI21_X1 _24252_ (.A(_14175_),
    .B1(_14383_),
    .B2(_14551_),
    .ZN(_14552_));
 NOR4_X1 _24253_ (.A1(_14545_),
    .A2(_14547_),
    .A3(_14549_),
    .A4(_14552_),
    .ZN(_14553_));
 NAND2_X1 _24254_ (.A1(_14149_),
    .A2(_14498_),
    .ZN(_14554_));
 OAI21_X1 _24255_ (.A(_14149_),
    .B1(_14203_),
    .B2(_14217_),
    .ZN(_14555_));
 NAND3_X1 _24256_ (.A1(_14227_),
    .A2(_14075_),
    .A3(_14281_),
    .ZN(_14556_));
 NAND2_X1 _24257_ (.A1(_14153_),
    .A2(_14074_),
    .ZN(_14557_));
 AND4_X1 _24258_ (.A1(_14554_),
    .A2(_14555_),
    .A3(_14556_),
    .A4(_14557_),
    .ZN(_14558_));
 NAND4_X1 _24259_ (.A1(_14534_),
    .A2(_14542_),
    .A3(_14553_),
    .A4(_14558_),
    .ZN(_14559_));
 NOR2_X1 _24260_ (.A1(_14526_),
    .A2(_14559_),
    .ZN(_14560_));
 INV_X1 _24261_ (.A(_00992_),
    .ZN(_14561_));
 XNOR2_X1 _24262_ (.A(_14560_),
    .B(_14561_),
    .ZN(_14562_));
 MUX2_X1 _24263_ (.A(_01328_),
    .B(_14562_),
    .S(_14403_),
    .Z(_01083_));
 NAND2_X1 _24264_ (.A1(_14362_),
    .A2(_14103_),
    .ZN(_14563_));
 INV_X1 _24265_ (.A(_14563_),
    .ZN(_14564_));
 AND2_X1 _24266_ (.A1(_14070_),
    .A2(_14100_),
    .ZN(_14565_));
 NOR4_X1 _24267_ (.A1(_14564_),
    .A2(_14565_),
    .A3(_14305_),
    .A4(_14459_),
    .ZN(_14566_));
 AND2_X1 _24268_ (.A1(_14227_),
    .A2(_14120_),
    .ZN(_14567_));
 AOI21_X1 _24269_ (.A(_14134_),
    .B1(_14383_),
    .B2(_14551_),
    .ZN(_14568_));
 AOI211_X4 _24270_ (.A(_14567_),
    .B(_14568_),
    .C1(_14121_),
    .C2(_14125_),
    .ZN(_14569_));
 OAI21_X1 _24271_ (.A(_14149_),
    .B1(_14451_),
    .B2(_14261_),
    .ZN(_14570_));
 AND3_X1 _24272_ (.A1(_14570_),
    .A2(_14148_),
    .A3(_14313_),
    .ZN(_14571_));
 AND2_X1 _24273_ (.A1(_14074_),
    .A2(_14154_),
    .ZN(_14572_));
 AND2_X1 _24274_ (.A1(_14382_),
    .A2(_14074_),
    .ZN(_14573_));
 AOI211_X4 _24275_ (.A(_14572_),
    .B(_14573_),
    .C1(_14075_),
    .C2(_14227_),
    .ZN(_14574_));
 AND4_X1 _24276_ (.A1(_14566_),
    .A2(_14569_),
    .A3(_14571_),
    .A4(_14574_),
    .ZN(_14575_));
 AOI21_X1 _24277_ (.A(_14175_),
    .B1(_14364_),
    .B2(_14205_),
    .ZN(_14576_));
 OAI21_X1 _24278_ (.A(_14164_),
    .B1(_14394_),
    .B2(_14102_),
    .ZN(_14577_));
 OAI21_X1 _24279_ (.A(_14164_),
    .B1(_14184_),
    .B2(_14140_),
    .ZN(_14578_));
 OAI211_X2 _24280_ (.A(_14577_),
    .B(_14578_),
    .C1(_14180_),
    .C2(_14165_),
    .ZN(_14579_));
 AOI211_X4 _24281_ (.A(_14576_),
    .B(_14579_),
    .C1(_14109_),
    .C2(_14182_),
    .ZN(_14580_));
 OAI21_X1 _24282_ (.A(_14450_),
    .B1(_14322_),
    .B2(_14198_),
    .ZN(_14581_));
 OAI21_X1 _24283_ (.A(_14450_),
    .B1(_14498_),
    .B2(_14153_),
    .ZN(_14582_));
 AND4_X1 _24284_ (.A1(_14194_),
    .A2(_14581_),
    .A3(_14537_),
    .A4(_14582_),
    .ZN(_14583_));
 AND2_X1 _24285_ (.A1(_14332_),
    .A2(_14209_),
    .ZN(_14584_));
 AND2_X1 _24286_ (.A1(_14327_),
    .A2(_14209_),
    .ZN(_14585_));
 NOR2_X1 _24287_ (.A1(_14584_),
    .A2(_14585_),
    .ZN(_14586_));
 NAND2_X1 _24288_ (.A1(_14210_),
    .A2(_14261_),
    .ZN(_14587_));
 OAI211_X2 _24289_ (.A(_14072_),
    .B(_14162_),
    .C1(_14215_),
    .C2(_14150_),
    .ZN(_14588_));
 AND3_X1 _24290_ (.A1(_14586_),
    .A2(_14587_),
    .A3(_14588_),
    .ZN(_14589_));
 AND4_X1 _24291_ (.A1(_14575_),
    .A2(_14580_),
    .A3(_14583_),
    .A4(_14589_),
    .ZN(_14590_));
 NAND2_X1 _24292_ (.A1(_14208_),
    .A2(_14234_),
    .ZN(_14591_));
 NAND2_X1 _24293_ (.A1(_14496_),
    .A2(_14591_),
    .ZN(_14592_));
 INV_X1 _24294_ (.A(_14198_),
    .ZN(_14593_));
 AOI21_X1 _24295_ (.A(_14387_),
    .B1(_14593_),
    .B2(_14205_),
    .ZN(_14594_));
 AOI21_X1 _24296_ (.A(_14387_),
    .B1(_14544_),
    .B2(_14445_),
    .ZN(_14595_));
 NOR4_X1 _24297_ (.A1(_14592_),
    .A2(_14594_),
    .A3(_14595_),
    .A4(_14380_),
    .ZN(_14596_));
 AND4_X1 _24298_ (.A1(_14419_),
    .A2(_14421_),
    .A3(_14423_),
    .A4(_14506_),
    .ZN(_14597_));
 OAI21_X1 _24299_ (.A(_14514_),
    .B1(_14299_),
    .B2(_14179_),
    .ZN(_14598_));
 AND2_X1 _24300_ (.A1(_14275_),
    .A2(_14123_),
    .ZN(_14599_));
 AND2_X1 _24301_ (.A1(_14275_),
    .A2(_14198_),
    .ZN(_14600_));
 AND2_X1 _24302_ (.A1(_14275_),
    .A2(_14179_),
    .ZN(_14601_));
 NOR3_X1 _24303_ (.A1(_14599_),
    .A2(_14600_),
    .A3(_14601_),
    .ZN(_14602_));
 AND4_X1 _24304_ (.A1(_14418_),
    .A2(_14597_),
    .A3(_14598_),
    .A4(_14602_),
    .ZN(_14603_));
 NAND2_X1 _24305_ (.A1(_14245_),
    .A2(_14498_),
    .ZN(_14604_));
 OAI21_X1 _24306_ (.A(_14245_),
    .B1(_14394_),
    .B2(_14123_),
    .ZN(_14605_));
 OAI211_X2 _24307_ (.A(_14604_),
    .B(_14605_),
    .C1(_14503_),
    .C2(_14433_),
    .ZN(_14606_));
 AND4_X1 _24308_ (.A1(_14081_),
    .A2(_14105_),
    .A3(_14136_),
    .A4(_14222_),
    .ZN(_14607_));
 OR2_X1 _24309_ (.A1(_14396_),
    .A2(_14607_),
    .ZN(_14608_));
 NOR4_X1 _24310_ (.A1(_14606_),
    .A2(_14608_),
    .A3(_14243_),
    .A4(_14492_),
    .ZN(_14609_));
 AND2_X1 _24311_ (.A1(_14382_),
    .A2(_14256_),
    .ZN(_14610_));
 INV_X1 _24312_ (.A(_14610_),
    .ZN(_14611_));
 INV_X1 _24313_ (.A(_14290_),
    .ZN(_14612_));
 NAND4_X1 _24314_ (.A1(_14261_),
    .A2(_14072_),
    .A3(_14254_),
    .A4(_14262_),
    .ZN(_14613_));
 NAND4_X1 _24315_ (.A1(_14611_),
    .A2(_14612_),
    .A3(_14347_),
    .A4(_14613_),
    .ZN(_14614_));
 INV_X1 _24316_ (.A(_14217_),
    .ZN(_14615_));
 AOI21_X1 _24317_ (.A(_14283_),
    .B1(_14615_),
    .B2(_14086_),
    .ZN(_14616_));
 NOR4_X1 _24318_ (.A1(_14614_),
    .A2(_14288_),
    .A3(_14333_),
    .A4(_14616_),
    .ZN(_14617_));
 AND4_X1 _24319_ (.A1(_14596_),
    .A2(_14603_),
    .A3(_14609_),
    .A4(_14617_),
    .ZN(_14618_));
 AND3_X1 _24320_ (.A1(_14590_),
    .A2(_00993_),
    .A3(_14618_),
    .ZN(_14619_));
 AOI21_X1 _24321_ (.A(_00993_),
    .B1(_14590_),
    .B2(_14618_),
    .ZN(_14620_));
 NOR2_X1 _24322_ (.A1(_14619_),
    .A2(_14620_),
    .ZN(_14621_));
 MUX2_X1 _24323_ (.A(_01203_),
    .B(_14621_),
    .S(_14403_),
    .Z(_01084_));
 NAND2_X1 _24324_ (.A1(_14075_),
    .A2(_14155_),
    .ZN(_14622_));
 OAI221_X1 _24325_ (.A(_14622_),
    .B1(_14169_),
    .B2(_14219_),
    .C1(_14180_),
    .C2(_14269_),
    .ZN(_14623_));
 AND2_X1 _24326_ (.A1(_14567_),
    .A2(_14281_),
    .ZN(_14624_));
 AND3_X1 _24327_ (.A1(_14208_),
    .A2(_14121_),
    .A3(_14130_),
    .ZN(_14625_));
 NOR4_X1 _24328_ (.A1(_14623_),
    .A2(_14608_),
    .A3(_14624_),
    .A4(_14625_),
    .ZN(_14626_));
 AND2_X1 _24329_ (.A1(_14121_),
    .A2(_14140_),
    .ZN(_14627_));
 INV_X1 _24330_ (.A(_14627_),
    .ZN(_14628_));
 NAND3_X1 _24331_ (.A1(_14138_),
    .A2(_14073_),
    .A3(_14173_),
    .ZN(_14629_));
 AND3_X1 _24332_ (.A1(_14628_),
    .A2(_14346_),
    .A3(_14629_),
    .ZN(_14630_));
 OAI22_X1 _24333_ (.A1(_14387_),
    .A2(_14388_),
    .B1(_14434_),
    .B2(_14219_),
    .ZN(_14631_));
 AOI221_X4 _24334_ (.A(_14631_),
    .B1(_14240_),
    .B2(_14074_),
    .C1(_14332_),
    .C2(_14275_),
    .ZN(_14632_));
 INV_X1 _24335_ (.A(_14203_),
    .ZN(_14633_));
 OAI22_X1 _24336_ (.A1(_14433_),
    .A2(_14201_),
    .B1(_14219_),
    .B2(_14633_),
    .ZN(_14634_));
 AND2_X1 _24337_ (.A1(_14268_),
    .A2(_14127_),
    .ZN(_14635_));
 AND2_X1 _24338_ (.A1(_14121_),
    .A2(_14070_),
    .ZN(_14636_));
 NOR4_X1 _24339_ (.A1(_14634_),
    .A2(_14248_),
    .A3(_14635_),
    .A4(_14636_),
    .ZN(_14637_));
 AND4_X1 _24340_ (.A1(_14626_),
    .A2(_14630_),
    .A3(_14632_),
    .A4(_14637_),
    .ZN(_14638_));
 AOI21_X1 _24341_ (.A(_14321_),
    .B1(_14387_),
    .B2(_14490_),
    .ZN(_14639_));
 AND3_X1 _24342_ (.A1(_14075_),
    .A2(_14093_),
    .A3(_14232_),
    .ZN(_14640_));
 OR2_X1 _24343_ (.A1(_14639_),
    .A2(_14640_),
    .ZN(_14641_));
 AND3_X1 _24344_ (.A1(_14275_),
    .A2(_14231_),
    .A3(_14102_),
    .ZN(_14642_));
 AND2_X1 _24345_ (.A1(_14327_),
    .A2(_14256_),
    .ZN(_14643_));
 OR2_X1 _24346_ (.A1(_14642_),
    .A2(_14643_),
    .ZN(_14644_));
 NOR4_X1 _24347_ (.A1(_14641_),
    .A2(_14644_),
    .A3(_14213_),
    .A4(_14564_),
    .ZN(_14645_));
 NOR2_X1 _24348_ (.A1(_14445_),
    .A2(_14142_),
    .ZN(_14646_));
 OAI21_X1 _24349_ (.A(_14234_),
    .B1(_14646_),
    .B2(_14382_),
    .ZN(_14647_));
 OAI21_X1 _24350_ (.A(_14182_),
    .B1(_14123_),
    .B2(_14217_),
    .ZN(_14648_));
 OAI21_X1 _24351_ (.A(_14149_),
    .B1(_14550_),
    .B2(_14109_),
    .ZN(_14649_));
 NAND3_X1 _24352_ (.A1(_14647_),
    .A2(_14648_),
    .A3(_14649_),
    .ZN(_14650_));
 AND3_X1 _24353_ (.A1(_14140_),
    .A2(_14072_),
    .A3(_14230_),
    .ZN(_14651_));
 OR2_X1 _24354_ (.A1(_14372_),
    .A2(_14651_),
    .ZN(_14652_));
 AND2_X1 _24355_ (.A1(_14200_),
    .A2(_14256_),
    .ZN(_14653_));
 OR2_X1 _24356_ (.A1(_14653_),
    .A2(_14528_),
    .ZN(_14654_));
 OAI211_X2 _24357_ (.A(_14363_),
    .B(_14311_),
    .C1(_14473_),
    .C2(_14171_),
    .ZN(_14655_));
 NOR4_X1 _24358_ (.A1(_14650_),
    .A2(_14652_),
    .A3(_14654_),
    .A4(_14655_),
    .ZN(_14656_));
 AND2_X1 _24359_ (.A1(_14186_),
    .A2(_14187_),
    .ZN(_14657_));
 AOI211_X4 _24360_ (.A(_14425_),
    .B(_14277_),
    .C1(_14514_),
    .C2(_14179_),
    .ZN(_14658_));
 NAND4_X1 _24361_ (.A1(_14514_),
    .A2(_14083_),
    .A3(_14130_),
    .A4(_14150_),
    .ZN(_14659_));
 OAI21_X1 _24362_ (.A(_14514_),
    .B1(_14498_),
    .B2(_14540_),
    .ZN(_14660_));
 AND4_X1 _24363_ (.A1(_14657_),
    .A2(_14658_),
    .A3(_14659_),
    .A4(_14660_),
    .ZN(_14661_));
 NAND4_X1 _24364_ (.A1(_14638_),
    .A2(_14645_),
    .A3(_14656_),
    .A4(_14661_),
    .ZN(_14662_));
 OAI21_X1 _24365_ (.A(_14199_),
    .B1(_14134_),
    .B2(_14205_),
    .ZN(_14663_));
 OR2_X1 _24366_ (.A1(_14663_),
    .A2(_14565_),
    .ZN(_14664_));
 AOI21_X1 _24367_ (.A(_14490_),
    .B1(_14593_),
    .B2(_14381_),
    .ZN(_14665_));
 AND2_X1 _24368_ (.A1(_14176_),
    .A2(_14279_),
    .ZN(_14666_));
 OR3_X1 _24369_ (.A1(_14665_),
    .A2(_14666_),
    .A3(_14291_),
    .ZN(_14667_));
 AND2_X1 _24370_ (.A1(_14244_),
    .A2(_14070_),
    .ZN(_14668_));
 AND2_X1 _24371_ (.A1(_14228_),
    .A2(_14124_),
    .ZN(_14669_));
 OR2_X1 _24372_ (.A1(_14668_),
    .A2(_14669_),
    .ZN(_14670_));
 AOI21_X1 _24373_ (.A(_14266_),
    .B1(_14490_),
    .B2(_14080_),
    .ZN(_14671_));
 OR4_X2 _24374_ (.A1(_14664_),
    .A2(_14667_),
    .A3(_14670_),
    .A4(_14671_),
    .ZN(_14672_));
 NAND2_X1 _24375_ (.A1(_14384_),
    .A2(_14223_),
    .ZN(_14673_));
 NAND4_X1 _24376_ (.A1(_14673_),
    .A2(_14496_),
    .A3(_14428_),
    .A4(_14537_),
    .ZN(_14674_));
 AND2_X1 _24377_ (.A1(_14279_),
    .A2(_14179_),
    .ZN(_14675_));
 NOR2_X1 _24378_ (.A1(_14373_),
    .A2(_14675_),
    .ZN(_14676_));
 NAND2_X1 _24379_ (.A1(_14256_),
    .A2(_14550_),
    .ZN(_14677_));
 OAI21_X1 _24380_ (.A(_14280_),
    .B1(_14184_),
    .B2(_14128_),
    .ZN(_14678_));
 AOI22_X1 _24381_ (.A1(_14239_),
    .A2(_14155_),
    .B1(_14450_),
    .B2(_14287_),
    .ZN(_14679_));
 NAND4_X1 _24382_ (.A1(_14676_),
    .A2(_14677_),
    .A3(_14678_),
    .A4(_14679_),
    .ZN(_14680_));
 AND3_X1 _24383_ (.A1(_14198_),
    .A2(_14119_),
    .A3(_14162_),
    .ZN(_14681_));
 AND2_X1 _24384_ (.A1(_14164_),
    .A2(_14124_),
    .ZN(_14682_));
 AOI211_X4 _24385_ (.A(_14681_),
    .B(_14682_),
    .C1(_14192_),
    .C2(_14164_),
    .ZN(_14683_));
 OAI21_X1 _24386_ (.A(_14355_),
    .B1(_14070_),
    .B2(_14140_),
    .ZN(_14684_));
 OAI211_X2 _24387_ (.A(_14683_),
    .B(_14684_),
    .C1(_14111_),
    .C2(_14321_),
    .ZN(_14685_));
 OR4_X1 _24388_ (.A1(_14672_),
    .A2(_14674_),
    .A3(_14680_),
    .A4(_14685_),
    .ZN(_14686_));
 NOR2_X2 _24389_ (.A1(_14662_),
    .A2(_14686_),
    .ZN(_14687_));
 XOR2_X1 _24390_ (.A(_14687_),
    .B(_00994_),
    .Z(_14688_));
 MUX2_X1 _24391_ (.A(_01204_),
    .B(_14688_),
    .S(_14403_),
    .Z(_01085_));
 OR3_X1 _24392_ (.A1(_14101_),
    .A2(_14104_),
    .A3(_14305_),
    .ZN(_14689_));
 NOR3_X1 _24393_ (.A1(_14689_),
    .A2(_14564_),
    .A3(_14460_),
    .ZN(_14690_));
 AND2_X1 _24394_ (.A1(_14120_),
    .A2(_14183_),
    .ZN(_14691_));
 AND2_X1 _24395_ (.A1(_14121_),
    .A2(_14382_),
    .ZN(_14692_));
 AOI211_X4 _24396_ (.A(_14691_),
    .B(_14692_),
    .C1(_14166_),
    .C2(_14121_),
    .ZN(_14693_));
 NAND4_X1 _24397_ (.A1(_14159_),
    .A2(_14073_),
    .A3(_14069_),
    .A4(_14232_),
    .ZN(_14694_));
 AOI21_X1 _24398_ (.A(_14134_),
    .B1(_14593_),
    .B2(_14201_),
    .ZN(_14695_));
 AOI21_X1 _24399_ (.A(_14695_),
    .B1(_14122_),
    .B2(_14192_),
    .ZN(_14696_));
 AND4_X1 _24400_ (.A1(_14126_),
    .A2(_14693_),
    .A3(_14694_),
    .A4(_14696_),
    .ZN(_14697_));
 AND2_X1 _24401_ (.A1(_14149_),
    .A2(_14153_),
    .ZN(_14698_));
 INV_X1 _24402_ (.A(_14698_),
    .ZN(_14699_));
 NAND2_X1 _24403_ (.A1(_14699_),
    .A2(_14554_),
    .ZN(_14700_));
 AND2_X1 _24404_ (.A1(_14149_),
    .A2(_14203_),
    .ZN(_14701_));
 AND2_X1 _24405_ (.A1(_14137_),
    .A2(_14102_),
    .ZN(_14702_));
 NOR4_X1 _24406_ (.A1(_14700_),
    .A2(_14701_),
    .A3(_14702_),
    .A4(_14141_),
    .ZN(_14703_));
 AND2_X1 _24407_ (.A1(_14074_),
    .A2(_14351_),
    .ZN(_14704_));
 OAI21_X1 _24408_ (.A(_14557_),
    .B1(_14167_),
    .B2(_14080_),
    .ZN(_14705_));
 AOI211_X4 _24409_ (.A(_14704_),
    .B(_14705_),
    .C1(_14075_),
    .C2(_14128_),
    .ZN(_14706_));
 AND4_X1 _24410_ (.A1(_14690_),
    .A2(_14697_),
    .A3(_14703_),
    .A4(_14706_),
    .ZN(_14707_));
 OAI21_X1 _24411_ (.A(_14234_),
    .B1(_14322_),
    .B2(_14299_),
    .ZN(_14708_));
 AOI211_X4 _24412_ (.A(_14251_),
    .B(_14492_),
    .C1(_14239_),
    .C2(_14215_),
    .ZN(_14709_));
 AND4_X1 _24413_ (.A1(_14114_),
    .A2(_14222_),
    .A3(_14072_),
    .A4(_14085_),
    .ZN(_14710_));
 AND2_X1 _24414_ (.A1(_14244_),
    .A2(_14179_),
    .ZN(_14711_));
 AOI211_X4 _24415_ (.A(_14710_),
    .B(_14711_),
    .C1(_14132_),
    .C2(_14245_),
    .ZN(_14712_));
 OAI21_X1 _24416_ (.A(_14239_),
    .B1(_14392_),
    .B2(_14155_),
    .ZN(_14713_));
 OAI211_X2 _24417_ (.A(_14245_),
    .B(_17163_),
    .C1(_14262_),
    .C2(_14088_),
    .ZN(_14714_));
 AND4_X1 _24418_ (.A1(_14709_),
    .A2(_14712_),
    .A3(_14713_),
    .A4(_14714_),
    .ZN(_14715_));
 AND4_X1 _24419_ (.A1(_14081_),
    .A2(_14230_),
    .A3(_14173_),
    .A4(_14108_),
    .ZN(_14716_));
 AOI211_X4 _24420_ (.A(_14716_),
    .B(_14378_),
    .C1(_14240_),
    .C2(_14234_),
    .ZN(_14717_));
 NOR2_X1 _24421_ (.A1(_14387_),
    .A2(_14445_),
    .ZN(_14718_));
 AND3_X1 _24422_ (.A1(_14215_),
    .A2(_14159_),
    .A3(_14230_),
    .ZN(_14719_));
 NOR4_X1 _24423_ (.A1(_14718_),
    .A2(_14409_),
    .A3(_14386_),
    .A4(_14719_),
    .ZN(_14720_));
 AND4_X1 _24424_ (.A1(_14708_),
    .A2(_14715_),
    .A3(_14717_),
    .A4(_14720_),
    .ZN(_14721_));
 OAI21_X1 _24425_ (.A(_14450_),
    .B1(_14392_),
    .B2(_14153_),
    .ZN(_14722_));
 OAI21_X1 _24426_ (.A(_14450_),
    .B1(_14179_),
    .B2(_14125_),
    .ZN(_14723_));
 OAI211_X2 _24427_ (.A(_14722_),
    .B(_14723_),
    .C1(_14388_),
    .C2(_14195_),
    .ZN(_14724_));
 NAND2_X1 _24428_ (.A1(_14500_),
    .A2(_14355_),
    .ZN(_14725_));
 NAND4_X1 _24429_ (.A1(_14725_),
    .A2(_14358_),
    .A3(_14548_),
    .A4(_14543_),
    .ZN(_14726_));
 OAI21_X1 _24430_ (.A(_14182_),
    .B1(_14498_),
    .B2(_14540_),
    .ZN(_14727_));
 OAI21_X1 _24431_ (.A(_14727_),
    .B1(_14133_),
    .B2(_14175_),
    .ZN(_14728_));
 OAI21_X1 _24432_ (.A(_14210_),
    .B1(_14200_),
    .B2(_14375_),
    .ZN(_14729_));
 OAI211_X2 _24433_ (.A(_14729_),
    .B(_14368_),
    .C1(_14219_),
    .C2(_14381_),
    .ZN(_14730_));
 NOR4_X1 _24434_ (.A1(_14724_),
    .A2(_14726_),
    .A3(_14728_),
    .A4(_14730_),
    .ZN(_14731_));
 OAI21_X1 _24435_ (.A(_14275_),
    .B1(_14498_),
    .B2(_14540_),
    .ZN(_14732_));
 OAI211_X2 _24436_ (.A(_14159_),
    .B(_14254_),
    .C1(_14125_),
    .C2(_14215_),
    .ZN(_14733_));
 NAND4_X1 _24437_ (.A1(_14159_),
    .A2(_14231_),
    .A3(_14150_),
    .A4(_14254_),
    .ZN(_14734_));
 AND3_X1 _24438_ (.A1(_14732_),
    .A2(_14733_),
    .A3(_14734_),
    .ZN(_14735_));
 AND2_X1 _24439_ (.A1(_14153_),
    .A2(_14260_),
    .ZN(_14736_));
 AOI21_X1 _24440_ (.A(_14265_),
    .B1(_14381_),
    .B2(_14434_),
    .ZN(_14737_));
 NAND2_X1 _24441_ (.A1(_14633_),
    .A2(_14201_),
    .ZN(_14738_));
 AOI211_X4 _24442_ (.A(_14736_),
    .B(_14737_),
    .C1(_14514_),
    .C2(_14738_),
    .ZN(_14739_));
 AND2_X1 _24443_ (.A1(_14128_),
    .A2(_14280_),
    .ZN(_14740_));
 NOR4_X1 _24444_ (.A1(_14286_),
    .A2(_14446_),
    .A3(_14740_),
    .A4(_14675_),
    .ZN(_14741_));
 INV_X1 _24445_ (.A(_14653_),
    .ZN(_14742_));
 OAI21_X1 _24446_ (.A(_14257_),
    .B1(_14498_),
    .B2(_14070_),
    .ZN(_14743_));
 NAND3_X1 _24447_ (.A1(_14257_),
    .A2(_14150_),
    .A3(_14142_),
    .ZN(_14744_));
 AND4_X1 _24448_ (.A1(_14345_),
    .A2(_14742_),
    .A3(_14743_),
    .A4(_14744_),
    .ZN(_14745_));
 AND4_X1 _24449_ (.A1(_14735_),
    .A2(_14739_),
    .A3(_14741_),
    .A4(_14745_),
    .ZN(_14746_));
 NAND4_X1 _24450_ (.A1(_14707_),
    .A2(_14721_),
    .A3(_14731_),
    .A4(_14746_),
    .ZN(_14747_));
 NOR2_X1 _24451_ (.A1(_14747_),
    .A2(_14295_),
    .ZN(_14748_));
 XOR2_X1 _24452_ (.A(_14748_),
    .B(_00995_),
    .Z(_14749_));
 MUX2_X1 _24453_ (.A(_01205_),
    .B(_14749_),
    .S(_14403_),
    .Z(_01086_));
 NAND3_X1 _24454_ (.A1(_14227_),
    .A2(_14103_),
    .A3(_14281_),
    .ZN(_14750_));
 OAI211_X2 _24455_ (.A(_14103_),
    .B(_14261_),
    .C1(_14231_),
    .C2(_14262_),
    .ZN(_14751_));
 AND2_X1 _24456_ (.A1(_14750_),
    .A2(_14751_),
    .ZN(_14752_));
 OAI21_X1 _24457_ (.A(_14355_),
    .B1(_14384_),
    .B2(_14166_),
    .ZN(_14753_));
 NAND4_X1 _24458_ (.A1(_14159_),
    .A2(_11104_),
    .A3(_14162_),
    .A4(_14232_),
    .ZN(_14754_));
 OAI21_X1 _24459_ (.A(_14355_),
    .B1(_14198_),
    .B2(_14394_),
    .ZN(_14755_));
 AND3_X1 _24460_ (.A1(_14753_),
    .A2(_14754_),
    .A3(_14755_),
    .ZN(_14756_));
 AND2_X1 _24461_ (.A1(_14191_),
    .A2(_14382_),
    .ZN(_14757_));
 OAI21_X1 _24462_ (.A(_14190_),
    .B1(_14105_),
    .B2(_14178_),
    .ZN(_14758_));
 OAI21_X1 _24463_ (.A(_14758_),
    .B1(_14195_),
    .B2(_14201_),
    .ZN(_14759_));
 AOI211_X4 _24464_ (.A(_14757_),
    .B(_14759_),
    .C1(_14154_),
    .C2(_14191_),
    .ZN(_14760_));
 AND4_X1 _24465_ (.A1(_11103_),
    .A2(_14162_),
    .A3(_14078_),
    .A4(_14173_),
    .ZN(_14761_));
 AND2_X1 _24466_ (.A1(_14174_),
    .A2(_14140_),
    .ZN(_14762_));
 AOI211_X4 _24467_ (.A(_14761_),
    .B(_14762_),
    .C1(_14738_),
    .C2(_14182_),
    .ZN(_14763_));
 OAI211_X2 _24468_ (.A(_14209_),
    .B(_14090_),
    .C1(_11104_),
    .C2(_14262_),
    .ZN(_14764_));
 AND4_X1 _24469_ (.A1(_14368_),
    .A2(_14586_),
    .A3(_14366_),
    .A4(_14764_),
    .ZN(_14765_));
 AND4_X1 _24470_ (.A1(_14756_),
    .A2(_14760_),
    .A3(_14763_),
    .A4(_14765_),
    .ZN(_14766_));
 AND2_X1 _24471_ (.A1(_14120_),
    .A2(_14123_),
    .ZN(_14767_));
 AOI221_X4 _24472_ (.A(_14767_),
    .B1(_14121_),
    .B2(_14179_),
    .C1(_14281_),
    .C2(_14567_),
    .ZN(_14768_));
 OAI21_X1 _24473_ (.A(_14122_),
    .B1(_14240_),
    .B2(_14166_),
    .ZN(_14769_));
 AND4_X1 _24474_ (.A1(_14628_),
    .A2(_14768_),
    .A3(_14463_),
    .A4(_14769_),
    .ZN(_14770_));
 INV_X1 _24475_ (.A(_14702_),
    .ZN(_14771_));
 NAND4_X1 _24476_ (.A1(_14144_),
    .A2(_14148_),
    .A3(_14771_),
    .A4(_14554_),
    .ZN(_14772_));
 AOI21_X1 _24477_ (.A(_14080_),
    .B1(_14551_),
    .B2(_14544_),
    .ZN(_14773_));
 NOR4_X1 _24478_ (.A1(_14772_),
    .A2(_14318_),
    .A3(_14704_),
    .A4(_14773_),
    .ZN(_14774_));
 AND4_X1 _24479_ (.A1(_14752_),
    .A2(_14766_),
    .A3(_14770_),
    .A4(_14774_),
    .ZN(_14775_));
 NAND3_X1 _24480_ (.A1(_14332_),
    .A2(_14173_),
    .A3(_14230_),
    .ZN(_14776_));
 OAI21_X1 _24481_ (.A(_14223_),
    .B1(_14384_),
    .B2(_14646_),
    .ZN(_14777_));
 OAI211_X2 _24482_ (.A(_14159_),
    .B(_14230_),
    .C1(_14102_),
    .C2(_14351_),
    .ZN(_14778_));
 OAI21_X1 _24483_ (.A(_14234_),
    .B1(_14322_),
    .B2(_14394_),
    .ZN(_14779_));
 AND4_X1 _24484_ (.A1(_14776_),
    .A2(_14777_),
    .A3(_14778_),
    .A4(_14779_),
    .ZN(_14780_));
 NOR2_X1 _24485_ (.A1(_14599_),
    .A2(_14600_),
    .ZN(_14781_));
 AOI221_X4 _24486_ (.A(_14635_),
    .B1(_14185_),
    .B2(_14268_),
    .C1(_11104_),
    .C2(_14420_),
    .ZN(_14782_));
 AOI22_X1 _24487_ (.A1(_14426_),
    .A2(_14083_),
    .B1(_14514_),
    .B2(_14215_),
    .ZN(_14783_));
 AND2_X1 _24488_ (.A1(_14154_),
    .A2(_14259_),
    .ZN(_14784_));
 AND2_X1 _24489_ (.A1(_14497_),
    .A2(_14259_),
    .ZN(_14785_));
 AOI211_X4 _24490_ (.A(_14784_),
    .B(_14785_),
    .C1(_14332_),
    .C2(_14260_),
    .ZN(_14786_));
 AND4_X1 _24491_ (.A1(_14781_),
    .A2(_14782_),
    .A3(_14783_),
    .A4(_14786_),
    .ZN(_14787_));
 AND2_X1 _24492_ (.A1(_14394_),
    .A2(_14279_),
    .ZN(_14788_));
 AND2_X1 _24493_ (.A1(_14123_),
    .A2(_14279_),
    .ZN(_14789_));
 OR4_X1 _24494_ (.A1(_14788_),
    .A2(_14447_),
    .A3(_14789_),
    .A4(_14675_),
    .ZN(_14790_));
 NAND2_X1 _24495_ (.A1(_14146_),
    .A2(_14257_),
    .ZN(_14791_));
 NAND4_X1 _24496_ (.A1(_14611_),
    .A2(_14346_),
    .A3(_14677_),
    .A4(_14791_),
    .ZN(_14792_));
 NOR4_X1 _24497_ (.A1(_14790_),
    .A2(_14792_),
    .A3(_14331_),
    .A4(_14285_),
    .ZN(_14793_));
 OAI21_X1 _24498_ (.A(_14239_),
    .B1(_14327_),
    .B2(_14332_),
    .ZN(_14794_));
 OAI21_X1 _24499_ (.A(_14239_),
    .B1(_14184_),
    .B2(_14240_),
    .ZN(_14795_));
 OAI211_X2 _24500_ (.A(_14794_),
    .B(_14795_),
    .C1(_14490_),
    .C2(_14321_),
    .ZN(_14796_));
 NOR4_X1 _24501_ (.A1(_14652_),
    .A2(_14796_),
    .A3(_14246_),
    .A4(_14711_),
    .ZN(_14797_));
 AND4_X1 _24502_ (.A1(_14780_),
    .A2(_14787_),
    .A3(_14793_),
    .A4(_14797_),
    .ZN(_14798_));
 AND2_X1 _24503_ (.A1(_14775_),
    .A2(_14798_),
    .ZN(_14799_));
 XOR2_X1 _24504_ (.A(_14799_),
    .B(_00996_),
    .Z(_14800_));
 MUX2_X1 _24505_ (.A(_01206_),
    .B(_14800_),
    .S(_14403_),
    .Z(_01087_));
 AND2_X1 _24506_ (.A1(_17170_),
    .A2(_17171_),
    .ZN(_14801_));
 AND2_X2 _24507_ (.A1(_17172_),
    .A2(_17173_),
    .ZN(_14802_));
 AND2_X2 _24508_ (.A1(_14801_),
    .A2(_14802_),
    .ZN(_14803_));
 NOR2_X1 _24509_ (.A1(_09531_),
    .A2(_04121_),
    .ZN(_14804_));
 BUF_X4 _24510_ (.A(_14804_),
    .Z(_14805_));
 AND2_X2 _24511_ (.A1(_17166_),
    .A2(_17169_),
    .ZN(_14806_));
 BUF_X2 _24512_ (.A(_14806_),
    .Z(_14807_));
 AND3_X1 _24513_ (.A1(_14803_),
    .A2(_14805_),
    .A3(_14807_),
    .ZN(_14808_));
 INV_X1 _24514_ (.A(_17166_),
    .ZN(_14809_));
 NOR2_X1 _24515_ (.A1(_14809_),
    .A2(_17169_),
    .ZN(_14810_));
 NOR2_X4 _24516_ (.A1(_17144_),
    .A2(_17155_),
    .ZN(_14811_));
 AND2_X2 _24517_ (.A1(_14810_),
    .A2(_14811_),
    .ZN(_14812_));
 AND2_X1 _24518_ (.A1(_14812_),
    .A2(_14803_),
    .ZN(_14813_));
 INV_X1 _24519_ (.A(_14813_),
    .ZN(_14814_));
 NOR2_X1 _24520_ (.A1(_09095_),
    .A2(_17155_),
    .ZN(_14815_));
 BUF_X4 _24521_ (.A(_14815_),
    .Z(_14816_));
 NOR2_X1 _24522_ (.A1(_17166_),
    .A2(_17169_),
    .ZN(_14817_));
 BUF_X2 _24523_ (.A(_14817_),
    .Z(_14818_));
 AND2_X1 _24524_ (.A1(_14816_),
    .A2(_14818_),
    .ZN(_14819_));
 BUF_X2 _24525_ (.A(_14803_),
    .Z(_14820_));
 NAND2_X1 _24526_ (.A1(_14819_),
    .A2(_14820_),
    .ZN(_14821_));
 INV_X1 _24527_ (.A(_14820_),
    .ZN(_14822_));
 AND2_X2 _24528_ (.A1(_14818_),
    .A2(_17155_),
    .ZN(_14823_));
 INV_X1 _24529_ (.A(_14823_),
    .ZN(_14824_));
 OAI211_X2 _24530_ (.A(_14814_),
    .B(_14821_),
    .C1(_14822_),
    .C2(_14824_),
    .ZN(_14825_));
 INV_X1 _24531_ (.A(_17169_),
    .ZN(_14826_));
 NOR2_X1 _24532_ (.A1(_14826_),
    .A2(_17166_),
    .ZN(_14827_));
 BUF_X2 _24533_ (.A(_14827_),
    .Z(_14828_));
 BUF_X4 _24534_ (.A(_14828_),
    .Z(_14829_));
 CLKBUF_X2 _24535_ (.A(_14801_),
    .Z(_14830_));
 AND4_X1 _24536_ (.A1(_09531_),
    .A2(_14829_),
    .A3(_14830_),
    .A4(_14802_),
    .ZN(_14831_));
 AND2_X1 _24537_ (.A1(_14828_),
    .A2(_17155_),
    .ZN(_14832_));
 BUF_X2 _24538_ (.A(_14832_),
    .Z(_14833_));
 AND2_X1 _24539_ (.A1(_14833_),
    .A2(_14820_),
    .ZN(_14834_));
 OR4_X1 _24540_ (.A1(_14808_),
    .A2(_14825_),
    .A3(_14831_),
    .A4(_14834_),
    .ZN(_14835_));
 AND2_X2 _24541_ (.A1(_14804_),
    .A2(_14817_),
    .ZN(_14836_));
 NOR2_X1 _24542_ (.A1(_17170_),
    .A2(_17171_),
    .ZN(_14837_));
 AND2_X1 _24543_ (.A1(_14802_),
    .A2(_14837_),
    .ZN(_14838_));
 BUF_X2 _24544_ (.A(_14838_),
    .Z(_14839_));
 AND2_X1 _24545_ (.A1(_14836_),
    .A2(_14839_),
    .ZN(_14840_));
 BUF_X4 _24546_ (.A(_14807_),
    .Z(_14841_));
 AND3_X1 _24547_ (.A1(_14839_),
    .A2(_14805_),
    .A3(_14841_),
    .ZN(_14842_));
 AND3_X1 _24548_ (.A1(_14839_),
    .A2(_04121_),
    .A3(_14829_),
    .ZN(_14843_));
 AND2_X1 _24549_ (.A1(_14806_),
    .A2(_09531_),
    .ZN(_14844_));
 BUF_X2 _24550_ (.A(_14844_),
    .Z(_14845_));
 AND2_X1 _24551_ (.A1(_14845_),
    .A2(_14839_),
    .ZN(_14846_));
 OR4_X1 _24552_ (.A1(_14840_),
    .A2(_14842_),
    .A3(_14843_),
    .A4(_14846_),
    .ZN(_14847_));
 INV_X1 _24553_ (.A(_14811_),
    .ZN(_14848_));
 NAND2_X2 _24554_ (.A1(_14848_),
    .A2(_14807_),
    .ZN(_14849_));
 INV_X1 _24555_ (.A(_14849_),
    .ZN(_14850_));
 INV_X1 _24556_ (.A(_17171_),
    .ZN(_14851_));
 AND2_X2 _24557_ (.A1(_14851_),
    .A2(_17170_),
    .ZN(_14852_));
 AND2_X1 _24558_ (.A1(_14852_),
    .A2(_14802_),
    .ZN(_14853_));
 CLKBUF_X2 _24559_ (.A(_14853_),
    .Z(_14854_));
 AND2_X2 _24560_ (.A1(_04121_),
    .A2(_17155_),
    .ZN(_14855_));
 INV_X1 _24561_ (.A(_14855_),
    .ZN(_14856_));
 AND3_X1 _24562_ (.A1(_14850_),
    .A2(_14854_),
    .A3(_14856_),
    .ZN(_14857_));
 AND2_X1 _24563_ (.A1(_14854_),
    .A2(_14836_),
    .ZN(_14858_));
 BUF_X2 _24564_ (.A(_14810_),
    .Z(_14859_));
 AND2_X1 _24565_ (.A1(_14859_),
    .A2(_14815_),
    .ZN(_14860_));
 BUF_X2 _24566_ (.A(_14860_),
    .Z(_14861_));
 AND2_X1 _24567_ (.A1(_14854_),
    .A2(_14861_),
    .ZN(_14862_));
 AND2_X1 _24568_ (.A1(_14854_),
    .A2(_14829_),
    .ZN(_14863_));
 OR4_X1 _24569_ (.A1(_14857_),
    .A2(_14858_),
    .A3(_14862_),
    .A4(_14863_),
    .ZN(_14864_));
 NOR2_X1 _24570_ (.A1(_14851_),
    .A2(_17170_),
    .ZN(_14865_));
 BUF_X2 _24571_ (.A(_14865_),
    .Z(_14866_));
 AND2_X2 _24572_ (.A1(_14866_),
    .A2(_14802_),
    .ZN(_14867_));
 INV_X1 _24573_ (.A(_14867_),
    .ZN(_14868_));
 INV_X1 _24574_ (.A(_14828_),
    .ZN(_14869_));
 OR3_X1 _24575_ (.A1(_14868_),
    .A2(_14816_),
    .A3(_14869_),
    .ZN(_14870_));
 BUF_X4 _24576_ (.A(_14867_),
    .Z(_14871_));
 AND2_X1 _24577_ (.A1(_14855_),
    .A2(_14818_),
    .ZN(_14872_));
 INV_X1 _24578_ (.A(_14872_),
    .ZN(_14873_));
 AND2_X1 _24579_ (.A1(_14811_),
    .A2(_14817_),
    .ZN(_14874_));
 INV_X1 _24580_ (.A(_14874_),
    .ZN(_14875_));
 NAND2_X1 _24581_ (.A1(_14873_),
    .A2(_14875_),
    .ZN(_14876_));
 AND2_X2 _24582_ (.A1(_14810_),
    .A2(_09531_),
    .ZN(_14877_));
 OAI21_X1 _24583_ (.A(_14871_),
    .B1(_14876_),
    .B2(_14877_),
    .ZN(_14878_));
 AND2_X1 _24584_ (.A1(_14807_),
    .A2(_04121_),
    .ZN(_14879_));
 INV_X1 _24585_ (.A(_14879_),
    .ZN(_14880_));
 OAI211_X2 _24586_ (.A(_14870_),
    .B(_14878_),
    .C1(_14880_),
    .C2(_14868_),
    .ZN(_14881_));
 NOR4_X1 _24587_ (.A1(_14835_),
    .A2(_14847_),
    .A3(_14864_),
    .A4(_14881_),
    .ZN(_14882_));
 NOR2_X1 _24588_ (.A1(_17172_),
    .A2(_17173_),
    .ZN(_14883_));
 AND2_X2 _24589_ (.A1(_14883_),
    .A2(_14837_),
    .ZN(_14884_));
 AND3_X1 _24590_ (.A1(_14884_),
    .A2(_14816_),
    .A3(_14828_),
    .ZN(_14885_));
 NOR2_X1 _24591_ (.A1(_14849_),
    .A2(_14855_),
    .ZN(_14886_));
 BUF_X2 _24592_ (.A(_14884_),
    .Z(_14887_));
 AND3_X1 _24593_ (.A1(_14884_),
    .A2(_09101_),
    .A3(_14809_),
    .ZN(_14888_));
 AOI221_X4 _24594_ (.A(_14885_),
    .B1(_14886_),
    .B2(_14887_),
    .C1(_17169_),
    .C2(_14888_),
    .ZN(_14889_));
 AND2_X2 _24595_ (.A1(_14810_),
    .A2(_17155_),
    .ZN(_14890_));
 AND2_X1 _24596_ (.A1(_14890_),
    .A2(_14884_),
    .ZN(_14891_));
 INV_X1 _24597_ (.A(_14891_),
    .ZN(_14892_));
 NAND2_X1 _24598_ (.A1(_14884_),
    .A2(_14823_),
    .ZN(_14893_));
 NAND3_X1 _24599_ (.A1(_14884_),
    .A2(_14859_),
    .A3(_14816_),
    .ZN(_14894_));
 NAND4_X1 _24600_ (.A1(_14889_),
    .A2(_14892_),
    .A3(_14893_),
    .A4(_14894_),
    .ZN(_14895_));
 AND2_X2 _24601_ (.A1(_14807_),
    .A2(_14855_),
    .ZN(_14896_));
 BUF_X2 _24602_ (.A(_14883_),
    .Z(_14897_));
 AND2_X2 _24603_ (.A1(_14801_),
    .A2(_14897_),
    .ZN(_14898_));
 AND2_X1 _24604_ (.A1(_14896_),
    .A2(_14898_),
    .ZN(_14899_));
 INV_X1 _24605_ (.A(_14899_),
    .ZN(_14900_));
 AND2_X2 _24606_ (.A1(_14828_),
    .A2(_14811_),
    .ZN(_14901_));
 BUF_X4 _24607_ (.A(_14898_),
    .Z(_14902_));
 NAND2_X1 _24608_ (.A1(_14901_),
    .A2(_14902_),
    .ZN(_14903_));
 NAND2_X1 _24609_ (.A1(_14898_),
    .A2(_14845_),
    .ZN(_14904_));
 AND3_X1 _24610_ (.A1(_14900_),
    .A2(_14903_),
    .A3(_14904_),
    .ZN(_14905_));
 BUF_X4 _24611_ (.A(_14818_),
    .Z(_14906_));
 NAND3_X1 _24612_ (.A1(_14902_),
    .A2(_14848_),
    .A3(_14906_),
    .ZN(_14907_));
 INV_X1 _24613_ (.A(_14898_),
    .ZN(_14908_));
 AND2_X1 _24614_ (.A1(_14810_),
    .A2(_14804_),
    .ZN(_14909_));
 BUF_X2 _24615_ (.A(_14909_),
    .Z(_14910_));
 INV_X1 _24616_ (.A(_14910_),
    .ZN(_14911_));
 OAI211_X2 _24617_ (.A(_14905_),
    .B(_14907_),
    .C1(_14908_),
    .C2(_14911_),
    .ZN(_14912_));
 AND2_X2 _24618_ (.A1(_14827_),
    .A2(_14855_),
    .ZN(_14913_));
 INV_X1 _24619_ (.A(_14913_),
    .ZN(_14914_));
 INV_X1 _24620_ (.A(_14901_),
    .ZN(_14915_));
 NAND2_X1 _24621_ (.A1(_14914_),
    .A2(_14915_),
    .ZN(_14916_));
 AND2_X2 _24622_ (.A1(_14852_),
    .A2(_14883_),
    .ZN(_14917_));
 BUF_X4 _24623_ (.A(_14917_),
    .Z(_14918_));
 NAND2_X1 _24624_ (.A1(_14916_),
    .A2(_14918_),
    .ZN(_14919_));
 OAI21_X1 _24625_ (.A(_14918_),
    .B1(_14836_),
    .B2(_14872_),
    .ZN(_14920_));
 INV_X1 _24626_ (.A(_14917_),
    .ZN(_14921_));
 NAND2_X1 _24627_ (.A1(_14856_),
    .A2(_14859_),
    .ZN(_14922_));
 NOR2_X1 _24628_ (.A1(_14922_),
    .A2(_14811_),
    .ZN(_14923_));
 INV_X1 _24629_ (.A(_14923_),
    .ZN(_14924_));
 OAI211_X2 _24630_ (.A(_14919_),
    .B(_14920_),
    .C1(_14921_),
    .C2(_14924_),
    .ZN(_14925_));
 AND2_X1 _24631_ (.A1(_14866_),
    .A2(_14897_),
    .ZN(_14926_));
 BUF_X2 _24632_ (.A(_14926_),
    .Z(_14927_));
 INV_X1 _24633_ (.A(_14818_),
    .ZN(_14928_));
 NOR2_X1 _24634_ (.A1(_14928_),
    .A2(_14855_),
    .ZN(_14929_));
 AND2_X1 _24635_ (.A1(_14927_),
    .A2(_14929_),
    .ZN(_14930_));
 INV_X1 _24636_ (.A(_14930_),
    .ZN(_14931_));
 AND2_X1 _24637_ (.A1(_14848_),
    .A2(_14828_),
    .ZN(_14932_));
 NAND2_X1 _24638_ (.A1(_14932_),
    .A2(_14927_),
    .ZN(_14933_));
 BUF_X4 _24639_ (.A(_14859_),
    .Z(_14934_));
 NAND4_X1 _24640_ (.A1(_14927_),
    .A2(_14934_),
    .A3(_14848_),
    .A4(_14856_),
    .ZN(_14935_));
 AND2_X2 _24641_ (.A1(_14806_),
    .A2(_14811_),
    .ZN(_14936_));
 BUF_X4 _24642_ (.A(_14936_),
    .Z(_14937_));
 AND2_X2 _24643_ (.A1(_14806_),
    .A2(_17155_),
    .ZN(_14938_));
 OAI21_X1 _24644_ (.A(_14927_),
    .B1(_14937_),
    .B2(_14938_),
    .ZN(_14939_));
 NAND4_X1 _24645_ (.A1(_14931_),
    .A2(_14933_),
    .A3(_14935_),
    .A4(_14939_),
    .ZN(_14940_));
 NOR4_X1 _24646_ (.A1(_14895_),
    .A2(_14912_),
    .A3(_14925_),
    .A4(_14940_),
    .ZN(_14941_));
 INV_X1 _24647_ (.A(_17173_),
    .ZN(_14942_));
 AND2_X2 _24648_ (.A1(_14942_),
    .A2(_17172_),
    .ZN(_14943_));
 AND2_X1 _24649_ (.A1(_14943_),
    .A2(_14837_),
    .ZN(_14944_));
 BUF_X4 _24650_ (.A(_14944_),
    .Z(_14945_));
 AND2_X1 _24651_ (.A1(_14804_),
    .A2(_14806_),
    .ZN(_14946_));
 BUF_X2 _24652_ (.A(_14946_),
    .Z(_14947_));
 OAI21_X1 _24653_ (.A(_14945_),
    .B1(_14947_),
    .B2(_14845_),
    .ZN(_14948_));
 AND2_X1 _24654_ (.A1(_14818_),
    .A2(_09531_),
    .ZN(_14949_));
 BUF_X4 _24655_ (.A(_14949_),
    .Z(_14950_));
 OAI21_X1 _24656_ (.A(_14945_),
    .B1(_14812_),
    .B2(_14950_),
    .ZN(_14951_));
 BUF_X4 _24657_ (.A(_14943_),
    .Z(_14952_));
 BUF_X4 _24658_ (.A(_14829_),
    .Z(_14953_));
 BUF_X2 _24659_ (.A(_14837_),
    .Z(_14954_));
 NAND4_X1 _24660_ (.A1(_14952_),
    .A2(_04132_),
    .A3(_14953_),
    .A4(_14954_),
    .ZN(_14955_));
 NAND3_X1 _24661_ (.A1(_14948_),
    .A2(_14951_),
    .A3(_14955_),
    .ZN(_14956_));
 BUF_X4 _24662_ (.A(_14896_),
    .Z(_14957_));
 BUF_X4 _24663_ (.A(_14852_),
    .Z(_14958_));
 NAND3_X1 _24664_ (.A1(_14957_),
    .A2(_14958_),
    .A3(_14952_),
    .ZN(_14959_));
 BUF_X4 _24665_ (.A(_04121_),
    .Z(_14960_));
 NAND4_X1 _24666_ (.A1(_14952_),
    .A2(_14958_),
    .A3(_14829_),
    .A4(_14960_),
    .ZN(_14961_));
 NAND2_X1 _24667_ (.A1(_14959_),
    .A2(_14961_),
    .ZN(_14962_));
 AND2_X1 _24668_ (.A1(_14943_),
    .A2(_14852_),
    .ZN(_14963_));
 INV_X1 _24669_ (.A(_14963_),
    .ZN(_14964_));
 INV_X1 _24670_ (.A(_14805_),
    .ZN(_14965_));
 NAND2_X1 _24671_ (.A1(_14965_),
    .A2(_14906_),
    .ZN(_14966_));
 NOR2_X1 _24672_ (.A1(_14964_),
    .A2(_14966_),
    .ZN(_14967_));
 AND2_X1 _24673_ (.A1(_14963_),
    .A2(_14890_),
    .ZN(_14968_));
 OR3_X1 _24674_ (.A1(_14962_),
    .A2(_14967_),
    .A3(_14968_),
    .ZN(_14969_));
 AND2_X2 _24675_ (.A1(_14943_),
    .A2(_14801_),
    .ZN(_14970_));
 AND2_X1 _24676_ (.A1(_14815_),
    .A2(_14806_),
    .ZN(_14971_));
 BUF_X2 _24677_ (.A(_14971_),
    .Z(_14972_));
 OAI21_X1 _24678_ (.A(_14970_),
    .B1(_14947_),
    .B2(_14972_),
    .ZN(_14973_));
 NAND3_X1 _24679_ (.A1(_14913_),
    .A2(_14830_),
    .A3(_14952_),
    .ZN(_14974_));
 NAND2_X1 _24680_ (.A1(_14973_),
    .A2(_14974_),
    .ZN(_14975_));
 INV_X1 _24681_ (.A(_14975_),
    .ZN(_14976_));
 BUF_X4 _24682_ (.A(_14970_),
    .Z(_14977_));
 OAI211_X2 _24683_ (.A(_14977_),
    .B(_14906_),
    .C1(_04132_),
    .C2(_09532_),
    .ZN(_14978_));
 AND2_X2 _24684_ (.A1(_14859_),
    .A2(_04121_),
    .ZN(_14979_));
 INV_X1 _24685_ (.A(_14979_),
    .ZN(_14980_));
 INV_X1 _24686_ (.A(_14970_),
    .ZN(_14981_));
 OAI211_X2 _24687_ (.A(_14976_),
    .B(_14978_),
    .C1(_14980_),
    .C2(_14981_),
    .ZN(_14982_));
 AND2_X1 _24688_ (.A1(_14943_),
    .A2(_14865_),
    .ZN(_14983_));
 BUF_X2 _24689_ (.A(_14983_),
    .Z(_14984_));
 BUF_X2 _24690_ (.A(_14984_),
    .Z(_14985_));
 OAI21_X1 _24691_ (.A(_14985_),
    .B1(_14877_),
    .B2(_14890_),
    .ZN(_14986_));
 NOR3_X1 _24692_ (.A1(_14805_),
    .A2(_17166_),
    .A3(_14826_),
    .ZN(_14987_));
 OAI21_X1 _24693_ (.A(_14985_),
    .B1(_14987_),
    .B2(_14947_),
    .ZN(_14988_));
 BUF_X4 _24694_ (.A(_14872_),
    .Z(_14989_));
 NAND2_X1 _24695_ (.A1(_14985_),
    .A2(_14989_),
    .ZN(_14990_));
 BUF_X2 _24696_ (.A(_14819_),
    .Z(_14991_));
 NAND2_X1 _24697_ (.A1(_14985_),
    .A2(_14991_),
    .ZN(_14992_));
 NAND4_X1 _24698_ (.A1(_14986_),
    .A2(_14988_),
    .A3(_14990_),
    .A4(_14992_),
    .ZN(_14993_));
 NOR4_X1 _24699_ (.A1(_14956_),
    .A2(_14969_),
    .A3(_14982_),
    .A4(_14993_),
    .ZN(_14994_));
 NOR2_X1 _24700_ (.A1(_14942_),
    .A2(_17172_),
    .ZN(_14995_));
 AND2_X1 _24701_ (.A1(_14852_),
    .A2(_14995_),
    .ZN(_14996_));
 BUF_X2 _24702_ (.A(_14996_),
    .Z(_14997_));
 AND3_X1 _24703_ (.A1(_14997_),
    .A2(_14848_),
    .A3(_14929_),
    .ZN(_14998_));
 AOI21_X1 _24704_ (.A(_14998_),
    .B1(_14938_),
    .B2(_14997_),
    .ZN(_14999_));
 AND2_X1 _24705_ (.A1(_14995_),
    .A2(_14801_),
    .ZN(_15000_));
 BUF_X4 _24706_ (.A(_15000_),
    .Z(_15001_));
 AND2_X1 _24707_ (.A1(_15001_),
    .A2(_14936_),
    .ZN(_15002_));
 AND2_X1 _24708_ (.A1(_14810_),
    .A2(_14855_),
    .ZN(_15003_));
 BUF_X2 _24709_ (.A(_15003_),
    .Z(_15004_));
 NAND2_X1 _24710_ (.A1(_15000_),
    .A2(_15004_),
    .ZN(_15005_));
 INV_X1 _24711_ (.A(_14877_),
    .ZN(_15006_));
 INV_X1 _24712_ (.A(_15000_),
    .ZN(_15007_));
 OAI21_X1 _24713_ (.A(_15005_),
    .B1(_15006_),
    .B2(_15007_),
    .ZN(_15008_));
 NOR2_X1 _24714_ (.A1(_14928_),
    .A2(_14816_),
    .ZN(_15009_));
 AOI211_X4 _24715_ (.A(_15002_),
    .B(_15008_),
    .C1(_15001_),
    .C2(_15009_),
    .ZN(_15010_));
 AND2_X2 _24716_ (.A1(_14995_),
    .A2(_14954_),
    .ZN(_15011_));
 BUF_X2 _24717_ (.A(_15011_),
    .Z(_15012_));
 AND2_X1 _24718_ (.A1(_14828_),
    .A2(_04121_),
    .ZN(_15013_));
 OAI21_X1 _24719_ (.A(_15012_),
    .B1(_14850_),
    .B2(_15013_),
    .ZN(_15014_));
 NAND3_X1 _24720_ (.A1(_15011_),
    .A2(_14859_),
    .A3(_14965_),
    .ZN(_15015_));
 BUF_X4 _24721_ (.A(_14995_),
    .Z(_15016_));
 NAND4_X1 _24722_ (.A1(_15016_),
    .A2(_09095_),
    .A3(_14954_),
    .A4(_14906_),
    .ZN(_15017_));
 AND3_X1 _24723_ (.A1(_15014_),
    .A2(_15015_),
    .A3(_15017_),
    .ZN(_15018_));
 AND2_X2 _24724_ (.A1(_14866_),
    .A2(_14995_),
    .ZN(_15019_));
 AND2_X1 _24725_ (.A1(_15019_),
    .A2(_14812_),
    .ZN(_15020_));
 INV_X1 _24726_ (.A(_15020_),
    .ZN(_15021_));
 BUF_X2 _24727_ (.A(_15019_),
    .Z(_15022_));
 NAND2_X1 _24728_ (.A1(_15022_),
    .A2(_14957_),
    .ZN(_15023_));
 AND2_X2 _24729_ (.A1(_14816_),
    .A2(_14828_),
    .ZN(_15024_));
 OAI21_X1 _24730_ (.A(_15022_),
    .B1(_15024_),
    .B2(_14845_),
    .ZN(_15025_));
 AND3_X1 _24731_ (.A1(_15021_),
    .A2(_15023_),
    .A3(_15025_),
    .ZN(_15026_));
 AND4_X1 _24732_ (.A1(_14999_),
    .A2(_15010_),
    .A3(_15018_),
    .A4(_15026_),
    .ZN(_15027_));
 NAND4_X1 _24733_ (.A1(_14882_),
    .A2(_14941_),
    .A3(_14994_),
    .A4(_15027_),
    .ZN(_15028_));
 BUF_X4 _24734_ (.A(_14874_),
    .Z(_15029_));
 AND2_X1 _24735_ (.A1(_14887_),
    .A2(_15029_),
    .ZN(_15030_));
 NOR2_X1 _24736_ (.A1(_15028_),
    .A2(_15030_),
    .ZN(_15031_));
 XOR2_X1 _24737_ (.A(_15031_),
    .B(_00997_),
    .Z(_15032_));
 MUX2_X1 _24738_ (.A(_01207_),
    .B(_15032_),
    .S(_14403_),
    .Z(_01088_));
 AND2_X1 _24739_ (.A1(_14853_),
    .A2(_14936_),
    .ZN(_15033_));
 AND2_X1 _24740_ (.A1(_14804_),
    .A2(_14827_),
    .ZN(_15034_));
 BUF_X2 _24741_ (.A(_15034_),
    .Z(_15035_));
 AND2_X1 _24742_ (.A1(_14854_),
    .A2(_15035_),
    .ZN(_15036_));
 AOI211_X4 _24743_ (.A(_15033_),
    .B(_15036_),
    .C1(_14854_),
    .C2(_14957_),
    .ZN(_15037_));
 BUF_X4 _24744_ (.A(_14854_),
    .Z(_15038_));
 OAI21_X1 _24745_ (.A(_15038_),
    .B1(_14861_),
    .B2(_14890_),
    .ZN(_15039_));
 INV_X1 _24746_ (.A(_14853_),
    .ZN(_15040_));
 AND2_X1 _24747_ (.A1(_14818_),
    .A2(_04121_),
    .ZN(_15041_));
 INV_X1 _24748_ (.A(_15041_),
    .ZN(_15042_));
 OAI211_X2 _24749_ (.A(_15037_),
    .B(_15039_),
    .C1(_15040_),
    .C2(_15042_),
    .ZN(_15043_));
 BUF_X4 _24750_ (.A(_14839_),
    .Z(_15044_));
 OAI21_X1 _24751_ (.A(_15044_),
    .B1(_14876_),
    .B2(_14979_),
    .ZN(_15045_));
 AND2_X1 _24752_ (.A1(_14913_),
    .A2(_14838_),
    .ZN(_15046_));
 INV_X1 _24753_ (.A(_15046_),
    .ZN(_15047_));
 OAI211_X2 _24754_ (.A(_15044_),
    .B(_14841_),
    .C1(_09096_),
    .C2(_09101_),
    .ZN(_15048_));
 NAND3_X1 _24755_ (.A1(_15045_),
    .A2(_15047_),
    .A3(_15048_),
    .ZN(_15049_));
 AND2_X2 _24756_ (.A1(_14828_),
    .A2(_09531_),
    .ZN(_15050_));
 AND2_X1 _24757_ (.A1(_14867_),
    .A2(_15050_),
    .ZN(_15051_));
 INV_X1 _24758_ (.A(_15051_),
    .ZN(_15052_));
 AND2_X1 _24759_ (.A1(_14910_),
    .A2(_14871_),
    .ZN(_15053_));
 INV_X1 _24760_ (.A(_15053_),
    .ZN(_15054_));
 NAND2_X1 _24761_ (.A1(_15035_),
    .A2(_14871_),
    .ZN(_15055_));
 OAI21_X1 _24762_ (.A(_14867_),
    .B1(_14896_),
    .B2(_14937_),
    .ZN(_15056_));
 NAND4_X1 _24763_ (.A1(_15052_),
    .A2(_15054_),
    .A3(_15055_),
    .A4(_15056_),
    .ZN(_15057_));
 AND2_X1 _24764_ (.A1(_14877_),
    .A2(_14803_),
    .ZN(_15058_));
 INV_X1 _24765_ (.A(_15058_),
    .ZN(_15059_));
 NAND2_X1 _24766_ (.A1(_14820_),
    .A2(_14938_),
    .ZN(_15060_));
 NAND2_X1 _24767_ (.A1(_14913_),
    .A2(_14820_),
    .ZN(_15061_));
 NAND2_X1 _24768_ (.A1(_14909_),
    .A2(_14820_),
    .ZN(_15062_));
 NAND4_X1 _24769_ (.A1(_15059_),
    .A2(_15060_),
    .A3(_15061_),
    .A4(_15062_),
    .ZN(_15063_));
 NOR4_X1 _24770_ (.A1(_15043_),
    .A2(_15049_),
    .A3(_15057_),
    .A4(_15063_),
    .ZN(_15064_));
 AND2_X1 _24771_ (.A1(_14833_),
    .A2(_14884_),
    .ZN(_15065_));
 INV_X1 _24772_ (.A(_14884_),
    .ZN(_15066_));
 OAI21_X1 _24773_ (.A(_14893_),
    .B1(_15066_),
    .B2(_14922_),
    .ZN(_15067_));
 AOI211_X4 _24774_ (.A(_15065_),
    .B(_15067_),
    .C1(_14841_),
    .C2(_14887_),
    .ZN(_15068_));
 INV_X1 _24775_ (.A(_14950_),
    .ZN(_15069_));
 AND2_X1 _24776_ (.A1(_14859_),
    .A2(_09095_),
    .ZN(_15070_));
 INV_X1 _24777_ (.A(_15070_),
    .ZN(_15071_));
 AOI21_X1 _24778_ (.A(_14921_),
    .B1(_15069_),
    .B2(_15071_),
    .ZN(_15072_));
 AND2_X1 _24779_ (.A1(_14917_),
    .A2(_14946_),
    .ZN(_15073_));
 AND2_X1 _24780_ (.A1(_14917_),
    .A2(_14833_),
    .ZN(_15074_));
 NOR3_X1 _24781_ (.A1(_15072_),
    .A2(_15073_),
    .A3(_15074_),
    .ZN(_15075_));
 INV_X1 _24782_ (.A(_14927_),
    .ZN(_15076_));
 NOR2_X1 _24783_ (.A1(_15076_),
    .A2(_14922_),
    .ZN(_15077_));
 AOI21_X1 _24784_ (.A(_15077_),
    .B1(_14927_),
    .B2(_15009_),
    .ZN(_15078_));
 NAND2_X1 _24785_ (.A1(_14848_),
    .A2(_14818_),
    .ZN(_15079_));
 INV_X1 _24786_ (.A(_15079_),
    .ZN(_15080_));
 OAI21_X1 _24787_ (.A(_14902_),
    .B1(_15080_),
    .B2(_14979_),
    .ZN(_15081_));
 NAND2_X1 _24788_ (.A1(_14947_),
    .A2(_14902_),
    .ZN(_15082_));
 OAI211_X2 _24789_ (.A(_14902_),
    .B(_14829_),
    .C1(_14960_),
    .C2(_09532_),
    .ZN(_15083_));
 AND4_X1 _24790_ (.A1(_14904_),
    .A2(_15081_),
    .A3(_15082_),
    .A4(_15083_),
    .ZN(_15084_));
 AND4_X1 _24791_ (.A1(_15068_),
    .A2(_15075_),
    .A3(_15078_),
    .A4(_15084_),
    .ZN(_15085_));
 NAND3_X1 _24792_ (.A1(_14946_),
    .A2(_14954_),
    .A3(_14943_),
    .ZN(_15086_));
 NAND3_X1 _24793_ (.A1(_14972_),
    .A2(_14954_),
    .A3(_14943_),
    .ZN(_15087_));
 NAND2_X1 _24794_ (.A1(_15086_),
    .A2(_15087_),
    .ZN(_15088_));
 INV_X1 _24795_ (.A(_14944_),
    .ZN(_15089_));
 AOI21_X1 _24796_ (.A(_15089_),
    .B1(_15042_),
    .B2(_14922_),
    .ZN(_15090_));
 AOI211_X4 _24797_ (.A(_15088_),
    .B(_15090_),
    .C1(_14953_),
    .C2(_14944_),
    .ZN(_15091_));
 AND2_X1 _24798_ (.A1(_15080_),
    .A2(_14984_),
    .ZN(_15092_));
 NAND2_X1 _24799_ (.A1(_14984_),
    .A2(_14946_),
    .ZN(_15093_));
 INV_X1 _24800_ (.A(_14983_),
    .ZN(_15094_));
 INV_X1 _24801_ (.A(_14832_),
    .ZN(_15095_));
 OAI21_X1 _24802_ (.A(_15093_),
    .B1(_15094_),
    .B2(_15095_),
    .ZN(_15096_));
 AOI211_X4 _24803_ (.A(_15092_),
    .B(_15096_),
    .C1(_15070_),
    .C2(_14985_),
    .ZN(_15097_));
 BUF_X4 _24804_ (.A(_14963_),
    .Z(_15098_));
 AND2_X1 _24805_ (.A1(_15098_),
    .A2(_15050_),
    .ZN(_15099_));
 INV_X1 _24806_ (.A(_15099_),
    .ZN(_15100_));
 OAI211_X2 _24807_ (.A(_14958_),
    .B(_14952_),
    .C1(_15004_),
    .C2(_15029_),
    .ZN(_15101_));
 OAI211_X2 _24808_ (.A(_14958_),
    .B(_14952_),
    .C1(_14957_),
    .C2(_14937_),
    .ZN(_15102_));
 NAND3_X1 _24809_ (.A1(_15035_),
    .A2(_14958_),
    .A3(_14952_),
    .ZN(_15103_));
 AND4_X1 _24810_ (.A1(_15100_),
    .A2(_15101_),
    .A3(_15102_),
    .A4(_15103_),
    .ZN(_15104_));
 AND2_X1 _24811_ (.A1(_14850_),
    .A2(_14970_),
    .ZN(_15105_));
 AND3_X1 _24812_ (.A1(_14970_),
    .A2(_14932_),
    .A3(_14856_),
    .ZN(_15106_));
 AND2_X1 _24813_ (.A1(_14970_),
    .A2(_15041_),
    .ZN(_15107_));
 AND4_X1 _24814_ (.A1(_14859_),
    .A2(_14943_),
    .A3(_14830_),
    .A4(_14811_),
    .ZN(_15108_));
 NOR4_X1 _24815_ (.A1(_15105_),
    .A2(_15106_),
    .A3(_15107_),
    .A4(_15108_),
    .ZN(_15109_));
 AND4_X1 _24816_ (.A1(_15091_),
    .A2(_15097_),
    .A3(_15104_),
    .A4(_15109_),
    .ZN(_15110_));
 BUF_X4 _24817_ (.A(_15001_),
    .Z(_15111_));
 OAI211_X2 _24818_ (.A(_15111_),
    .B(_14841_),
    .C1(_14805_),
    .C2(_14816_),
    .ZN(_15112_));
 AND2_X1 _24819_ (.A1(_14818_),
    .A2(_09095_),
    .ZN(_15113_));
 OAI21_X1 _24820_ (.A(_15111_),
    .B1(_14910_),
    .B2(_15113_),
    .ZN(_15114_));
 NAND4_X1 _24821_ (.A1(_14953_),
    .A2(_15016_),
    .A3(_04132_),
    .A4(_14830_),
    .ZN(_15115_));
 AND3_X1 _24822_ (.A1(_15112_),
    .A2(_15114_),
    .A3(_15115_),
    .ZN(_15116_));
 AND2_X1 _24823_ (.A1(_14997_),
    .A2(_14807_),
    .ZN(_15117_));
 NAND3_X1 _24824_ (.A1(_14836_),
    .A2(_14852_),
    .A3(_15016_),
    .ZN(_15118_));
 INV_X2 _24825_ (.A(_14996_),
    .ZN(_15119_));
 OAI21_X1 _24826_ (.A(_15118_),
    .B1(_15119_),
    .B2(_15006_),
    .ZN(_15120_));
 AOI211_X4 _24827_ (.A(_15117_),
    .B(_15120_),
    .C1(_15050_),
    .C2(_14997_),
    .ZN(_15121_));
 AND3_X1 _24828_ (.A1(_14932_),
    .A2(_14856_),
    .A3(_15011_),
    .ZN(_15122_));
 NAND4_X1 _24829_ (.A1(_14805_),
    .A2(_15016_),
    .A3(_14954_),
    .A4(_14818_),
    .ZN(_15123_));
 NAND2_X1 _24830_ (.A1(_15015_),
    .A2(_15123_),
    .ZN(_15124_));
 AOI211_X4 _24831_ (.A(_15122_),
    .B(_15124_),
    .C1(_15012_),
    .C2(_14957_),
    .ZN(_15125_));
 AND2_X1 _24832_ (.A1(_15022_),
    .A2(_14823_),
    .ZN(_15126_));
 AND2_X1 _24833_ (.A1(_14861_),
    .A2(_15022_),
    .ZN(_15127_));
 AND2_X1 _24834_ (.A1(_14987_),
    .A2(_15019_),
    .ZN(_15128_));
 AND2_X1 _24835_ (.A1(_15022_),
    .A2(_14991_),
    .ZN(_15129_));
 NOR4_X1 _24836_ (.A1(_15126_),
    .A2(_15127_),
    .A3(_15128_),
    .A4(_15129_),
    .ZN(_15130_));
 AND4_X1 _24837_ (.A1(_15116_),
    .A2(_15121_),
    .A3(_15125_),
    .A4(_15130_),
    .ZN(_15131_));
 NAND4_X1 _24838_ (.A1(_15064_),
    .A2(_15085_),
    .A3(_15110_),
    .A4(_15131_),
    .ZN(_15132_));
 NOR2_X1 _24839_ (.A1(_15132_),
    .A2(_15030_),
    .ZN(_15133_));
 XOR2_X1 _24840_ (.A(_15133_),
    .B(_00998_),
    .Z(_15134_));
 MUX2_X1 _24841_ (.A(_01208_),
    .B(_15134_),
    .S(_14403_),
    .Z(_01089_));
 INV_X1 _24842_ (.A(_14838_),
    .ZN(_15135_));
 AOI211_X4 _24843_ (.A(_14869_),
    .B(_15135_),
    .C1(_09095_),
    .C2(_09531_),
    .ZN(_15136_));
 AND2_X1 _24844_ (.A1(_14972_),
    .A2(_15044_),
    .ZN(_15137_));
 OR2_X1 _24845_ (.A1(_15136_),
    .A2(_15137_),
    .ZN(_15138_));
 OAI21_X1 _24846_ (.A(_15038_),
    .B1(_15035_),
    .B2(_15024_),
    .ZN(_15139_));
 OAI21_X1 _24847_ (.A(_15038_),
    .B1(_14991_),
    .B2(_14823_),
    .ZN(_15140_));
 OAI21_X1 _24848_ (.A(_15038_),
    .B1(_14938_),
    .B2(_14937_),
    .ZN(_15141_));
 NAND2_X1 _24849_ (.A1(_15038_),
    .A2(_14890_),
    .ZN(_15142_));
 NAND4_X1 _24850_ (.A1(_15139_),
    .A2(_15140_),
    .A3(_15141_),
    .A4(_15142_),
    .ZN(_15143_));
 AND3_X1 _24851_ (.A1(_14859_),
    .A2(_14802_),
    .A3(_14954_),
    .ZN(_15144_));
 INV_X1 _24852_ (.A(_14836_),
    .ZN(_15145_));
 AOI21_X1 _24853_ (.A(_15135_),
    .B1(_15145_),
    .B2(_14873_),
    .ZN(_15146_));
 NOR4_X1 _24854_ (.A1(_15138_),
    .A2(_15143_),
    .A3(_15144_),
    .A4(_15146_),
    .ZN(_15147_));
 OAI21_X1 _24855_ (.A(_14997_),
    .B1(_14913_),
    .B2(_15050_),
    .ZN(_15148_));
 NAND2_X1 _24856_ (.A1(_14997_),
    .A2(_14823_),
    .ZN(_15149_));
 INV_X1 _24857_ (.A(_14844_),
    .ZN(_15150_));
 OAI211_X2 _24858_ (.A(_15148_),
    .B(_15149_),
    .C1(_15150_),
    .C2(_15119_),
    .ZN(_15151_));
 INV_X1 _24859_ (.A(_15012_),
    .ZN(_15152_));
 NOR2_X1 _24860_ (.A1(_15152_),
    .A2(_14966_),
    .ZN(_15153_));
 NAND2_X1 _24861_ (.A1(_15012_),
    .A2(_14845_),
    .ZN(_15154_));
 OAI21_X1 _24862_ (.A(_15154_),
    .B1(_15152_),
    .B2(_14869_),
    .ZN(_15155_));
 AND2_X1 _24863_ (.A1(_15012_),
    .A2(_14934_),
    .ZN(_15156_));
 NOR4_X1 _24864_ (.A1(_15151_),
    .A2(_15153_),
    .A3(_15155_),
    .A4(_15156_),
    .ZN(_15157_));
 NAND2_X1 _24865_ (.A1(_15111_),
    .A2(_15009_),
    .ZN(_15158_));
 OAI21_X1 _24866_ (.A(_15022_),
    .B1(_14886_),
    .B2(_15035_),
    .ZN(_15159_));
 NAND2_X1 _24867_ (.A1(_14861_),
    .A2(_15022_),
    .ZN(_15160_));
 NAND2_X1 _24868_ (.A1(_15022_),
    .A2(_14890_),
    .ZN(_15161_));
 AND3_X1 _24869_ (.A1(_15159_),
    .A2(_15160_),
    .A3(_15161_),
    .ZN(_15162_));
 OAI211_X2 _24870_ (.A(_15111_),
    .B(_14934_),
    .C1(_09096_),
    .C2(_09532_),
    .ZN(_15163_));
 OAI211_X2 _24871_ (.A(_15001_),
    .B(_14953_),
    .C1(_09096_),
    .C2(_09532_),
    .ZN(_15164_));
 OAI21_X1 _24872_ (.A(_15001_),
    .B1(_14947_),
    .B2(_14937_),
    .ZN(_15165_));
 AND2_X1 _24873_ (.A1(_15164_),
    .A2(_15165_),
    .ZN(_15166_));
 AND4_X1 _24874_ (.A1(_15158_),
    .A2(_15162_),
    .A3(_15163_),
    .A4(_15166_),
    .ZN(_15167_));
 NAND2_X1 _24875_ (.A1(_14867_),
    .A2(_14890_),
    .ZN(_15168_));
 NOR3_X1 _24876_ (.A1(_14822_),
    .A2(_14966_),
    .A3(_14816_),
    .ZN(_15169_));
 AND4_X1 _24877_ (.A1(_14960_),
    .A2(_14830_),
    .A3(_14802_),
    .A4(_14807_),
    .ZN(_15170_));
 NOR4_X1 _24878_ (.A1(_15169_),
    .A2(_15058_),
    .A3(_14834_),
    .A4(_15170_),
    .ZN(_15171_));
 AND2_X1 _24879_ (.A1(_14867_),
    .A2(_14879_),
    .ZN(_15172_));
 AND2_X1 _24880_ (.A1(_14867_),
    .A2(_14936_),
    .ZN(_15173_));
 NOR2_X1 _24881_ (.A1(_15172_),
    .A2(_15173_),
    .ZN(_15174_));
 NAND3_X1 _24882_ (.A1(_14932_),
    .A2(_14871_),
    .A3(_14856_),
    .ZN(_15175_));
 AND4_X1 _24883_ (.A1(_15168_),
    .A2(_15171_),
    .A3(_15174_),
    .A4(_15175_),
    .ZN(_15176_));
 NAND4_X1 _24884_ (.A1(_15147_),
    .A2(_15157_),
    .A3(_15167_),
    .A4(_15176_),
    .ZN(_15177_));
 OAI21_X1 _24885_ (.A(_14985_),
    .B1(_14916_),
    .B2(_14886_),
    .ZN(_15178_));
 AND2_X1 _24886_ (.A1(_14983_),
    .A2(_15004_),
    .ZN(_15179_));
 AND2_X1 _24887_ (.A1(_14983_),
    .A2(_14949_),
    .ZN(_15180_));
 AOI221_X4 _24888_ (.A(_15179_),
    .B1(_14861_),
    .B2(_14984_),
    .C1(_14960_),
    .C2(_15180_),
    .ZN(_15181_));
 OAI21_X1 _24889_ (.A(_14977_),
    .B1(_14979_),
    .B2(_14989_),
    .ZN(_15182_));
 OAI21_X1 _24890_ (.A(_14977_),
    .B1(_14972_),
    .B2(_15050_),
    .ZN(_15183_));
 AND4_X1 _24891_ (.A1(_15178_),
    .A2(_15181_),
    .A3(_15182_),
    .A4(_15183_),
    .ZN(_15184_));
 NAND2_X1 _24892_ (.A1(_14965_),
    .A2(_14807_),
    .ZN(_15185_));
 INV_X1 _24893_ (.A(_15185_),
    .ZN(_15186_));
 NAND2_X1 _24894_ (.A1(_15186_),
    .A2(_14887_),
    .ZN(_15187_));
 NAND3_X1 _24895_ (.A1(_14887_),
    .A2(_14805_),
    .A3(_14829_),
    .ZN(_15188_));
 AND2_X1 _24896_ (.A1(_15187_),
    .A2(_15188_),
    .ZN(_15189_));
 NAND2_X1 _24897_ (.A1(_15080_),
    .A2(_14887_),
    .ZN(_15190_));
 INV_X1 _24898_ (.A(_15190_),
    .ZN(_15191_));
 AOI21_X1 _24899_ (.A(_14891_),
    .B1(_15191_),
    .B2(_14856_),
    .ZN(_15192_));
 OAI211_X2 _24900_ (.A(_14918_),
    .B(_14953_),
    .C1(_04132_),
    .C2(_09532_),
    .ZN(_15193_));
 NAND3_X1 _24901_ (.A1(_14845_),
    .A2(_14958_),
    .A3(_14897_),
    .ZN(_15194_));
 AND2_X1 _24902_ (.A1(_15193_),
    .A2(_15194_),
    .ZN(_15195_));
 OAI21_X1 _24903_ (.A(_14918_),
    .B1(_14910_),
    .B2(_14989_),
    .ZN(_15196_));
 AND4_X1 _24904_ (.A1(_15189_),
    .A2(_15192_),
    .A3(_15195_),
    .A4(_15196_),
    .ZN(_15197_));
 AOI21_X1 _24905_ (.A(_14908_),
    .B1(_14924_),
    .B2(_15069_),
    .ZN(_15198_));
 OAI21_X1 _24906_ (.A(_14927_),
    .B1(_14991_),
    .B2(_15029_),
    .ZN(_15199_));
 NAND2_X1 _24907_ (.A1(_14927_),
    .A2(_14877_),
    .ZN(_15200_));
 NAND3_X1 _24908_ (.A1(_14989_),
    .A2(_14866_),
    .A3(_14897_),
    .ZN(_15201_));
 NAND2_X1 _24909_ (.A1(_14926_),
    .A2(_14890_),
    .ZN(_15202_));
 NAND4_X1 _24910_ (.A1(_15199_),
    .A2(_15200_),
    .A3(_15201_),
    .A4(_15202_),
    .ZN(_15203_));
 NAND4_X1 _24911_ (.A1(_14805_),
    .A2(_14953_),
    .A3(_14866_),
    .A4(_14897_),
    .ZN(_15204_));
 NAND4_X1 _24912_ (.A1(_14866_),
    .A2(_14841_),
    .A3(_14855_),
    .A4(_14897_),
    .ZN(_15205_));
 INV_X1 _24913_ (.A(_15050_),
    .ZN(_15206_));
 OAI211_X2 _24914_ (.A(_15204_),
    .B(_15205_),
    .C1(_15206_),
    .C2(_15076_),
    .ZN(_15207_));
 AOI21_X1 _24915_ (.A(_14908_),
    .B1(_14915_),
    .B2(_14880_),
    .ZN(_15208_));
 NOR4_X1 _24916_ (.A1(_15198_),
    .A2(_15203_),
    .A3(_15207_),
    .A4(_15208_),
    .ZN(_15209_));
 OAI21_X1 _24917_ (.A(_14945_),
    .B1(_14861_),
    .B2(_14836_),
    .ZN(_15210_));
 OAI21_X1 _24918_ (.A(_15098_),
    .B1(_14861_),
    .B2(_14989_),
    .ZN(_15211_));
 OAI21_X1 _24919_ (.A(_15098_),
    .B1(_15035_),
    .B2(_14879_),
    .ZN(_15212_));
 OAI21_X1 _24920_ (.A(_14945_),
    .B1(_15035_),
    .B2(_14938_),
    .ZN(_15213_));
 AND4_X1 _24921_ (.A1(_15210_),
    .A2(_15211_),
    .A3(_15212_),
    .A4(_15213_),
    .ZN(_15214_));
 NAND4_X1 _24922_ (.A1(_15184_),
    .A2(_15197_),
    .A3(_15209_),
    .A4(_15214_),
    .ZN(_15215_));
 NOR2_X1 _24923_ (.A1(_15177_),
    .A2(_15215_),
    .ZN(_15216_));
 XOR2_X1 _24924_ (.A(_15216_),
    .B(_00999_),
    .Z(_15217_));
 MUX2_X1 _24925_ (.A(_01209_),
    .B(_15217_),
    .S(_14403_),
    .Z(_01059_));
 NAND3_X1 _24926_ (.A1(_15044_),
    .A2(_14934_),
    .A3(_14811_),
    .ZN(_15218_));
 AND3_X1 _24927_ (.A1(_14819_),
    .A2(_14802_),
    .A3(_14852_),
    .ZN(_15219_));
 INV_X1 _24928_ (.A(_14938_),
    .ZN(_15220_));
 AOI21_X1 _24929_ (.A(_15040_),
    .B1(_15220_),
    .B2(_14914_),
    .ZN(_15221_));
 INV_X1 _24930_ (.A(_14812_),
    .ZN(_15222_));
 INV_X1 _24931_ (.A(_15003_),
    .ZN(_15223_));
 NAND2_X1 _24932_ (.A1(_15222_),
    .A2(_15223_),
    .ZN(_15224_));
 AOI211_X4 _24933_ (.A(_15219_),
    .B(_15221_),
    .C1(_15038_),
    .C2(_15224_),
    .ZN(_15225_));
 AND2_X1 _24934_ (.A1(_15050_),
    .A2(_14839_),
    .ZN(_15226_));
 AOI211_X4 _24935_ (.A(_15046_),
    .B(_15226_),
    .C1(_14841_),
    .C2(_14839_),
    .ZN(_15227_));
 OAI21_X1 _24936_ (.A(_15044_),
    .B1(_14989_),
    .B2(_14950_),
    .ZN(_15228_));
 AND4_X1 _24937_ (.A1(_15218_),
    .A2(_15225_),
    .A3(_15227_),
    .A4(_15228_),
    .ZN(_15229_));
 OAI211_X2 _24938_ (.A(_14871_),
    .B(_14906_),
    .C1(_14805_),
    .C2(_14816_),
    .ZN(_15230_));
 AND2_X1 _24939_ (.A1(_15024_),
    .A2(_14803_),
    .ZN(_15231_));
 NOR3_X1 _24940_ (.A1(_14834_),
    .A2(_15231_),
    .A3(_14808_),
    .ZN(_15232_));
 AND2_X1 _24941_ (.A1(_15003_),
    .A2(_14803_),
    .ZN(_15233_));
 INV_X1 _24942_ (.A(_15233_),
    .ZN(_15234_));
 OAI21_X1 _24943_ (.A(_14820_),
    .B1(_15029_),
    .B2(_14823_),
    .ZN(_15235_));
 AND4_X1 _24944_ (.A1(_14814_),
    .A2(_15232_),
    .A3(_15234_),
    .A4(_15235_),
    .ZN(_15236_));
 OAI211_X2 _24945_ (.A(_14871_),
    .B(_14934_),
    .C1(_09096_),
    .C2(_09532_),
    .ZN(_15237_));
 NAND2_X1 _24946_ (.A1(_14871_),
    .A2(_14913_),
    .ZN(_15238_));
 OAI21_X1 _24947_ (.A(_14871_),
    .B1(_14937_),
    .B2(_14938_),
    .ZN(_15239_));
 AND3_X1 _24948_ (.A1(_15052_),
    .A2(_15238_),
    .A3(_15239_),
    .ZN(_15240_));
 AND4_X1 _24949_ (.A1(_15230_),
    .A2(_15236_),
    .A3(_15237_),
    .A4(_15240_),
    .ZN(_15241_));
 OAI21_X1 _24950_ (.A(_15012_),
    .B1(_14886_),
    .B2(_14833_),
    .ZN(_15242_));
 NAND2_X1 _24951_ (.A1(_14812_),
    .A2(_15012_),
    .ZN(_15243_));
 OAI211_X2 _24952_ (.A(_15242_),
    .B(_15243_),
    .C1(_15152_),
    .C2(_14966_),
    .ZN(_15244_));
 AND2_X1 _24953_ (.A1(_14932_),
    .A2(_14856_),
    .ZN(_15245_));
 AND2_X1 _24954_ (.A1(_15245_),
    .A2(_14997_),
    .ZN(_15246_));
 OAI21_X1 _24955_ (.A(_15149_),
    .B1(_15119_),
    .B2(_14980_),
    .ZN(_15247_));
 NOR4_X1 _24956_ (.A1(_15244_),
    .A2(_15246_),
    .A3(_15117_),
    .A4(_15247_),
    .ZN(_15248_));
 NAND4_X1 _24957_ (.A1(_15016_),
    .A2(_04132_),
    .A3(_14830_),
    .A4(_14906_),
    .ZN(_15249_));
 AND2_X1 _24958_ (.A1(_15034_),
    .A2(_15019_),
    .ZN(_15250_));
 INV_X1 _24959_ (.A(_15250_),
    .ZN(_15251_));
 NAND2_X1 _24960_ (.A1(_15251_),
    .A2(_15023_),
    .ZN(_15252_));
 AND2_X1 _24961_ (.A1(_15019_),
    .A2(_15004_),
    .ZN(_15253_));
 NOR4_X1 _24962_ (.A1(_15252_),
    .A2(_15020_),
    .A3(_15126_),
    .A4(_15253_),
    .ZN(_15254_));
 OAI211_X2 _24963_ (.A(_15111_),
    .B(_14934_),
    .C1(_09096_),
    .C2(_09101_),
    .ZN(_15255_));
 AND4_X1 _24964_ (.A1(_17155_),
    .A2(_14995_),
    .A3(_14801_),
    .A4(_14807_),
    .ZN(_15256_));
 AND2_X1 _24965_ (.A1(_14972_),
    .A2(_15000_),
    .ZN(_15257_));
 AOI211_X4 _24966_ (.A(_15256_),
    .B(_15257_),
    .C1(_15001_),
    .C2(_14916_),
    .ZN(_15258_));
 AND4_X1 _24967_ (.A1(_15249_),
    .A2(_15254_),
    .A3(_15255_),
    .A4(_15258_),
    .ZN(_15259_));
 NAND4_X1 _24968_ (.A1(_15229_),
    .A2(_15241_),
    .A3(_15248_),
    .A4(_15259_),
    .ZN(_15260_));
 OAI21_X1 _24969_ (.A(_14985_),
    .B1(_15080_),
    .B2(_14861_),
    .ZN(_15261_));
 AND3_X1 _24970_ (.A1(_14971_),
    .A2(_14866_),
    .A3(_14943_),
    .ZN(_15262_));
 AND2_X1 _24971_ (.A1(_14983_),
    .A2(_15013_),
    .ZN(_15263_));
 AOI211_X4 _24972_ (.A(_15262_),
    .B(_15263_),
    .C1(_14938_),
    .C2(_14984_),
    .ZN(_15264_));
 OAI21_X1 _24973_ (.A(_14977_),
    .B1(_14923_),
    .B2(_14989_),
    .ZN(_15265_));
 AND2_X1 _24974_ (.A1(_14828_),
    .A2(_09095_),
    .ZN(_15266_));
 OAI21_X1 _24975_ (.A(_14977_),
    .B1(_14972_),
    .B2(_15266_),
    .ZN(_15267_));
 AND4_X1 _24976_ (.A1(_15261_),
    .A2(_15264_),
    .A3(_15265_),
    .A4(_15267_),
    .ZN(_15268_));
 INV_X1 _24977_ (.A(_14916_),
    .ZN(_15269_));
 INV_X1 _24978_ (.A(_14937_),
    .ZN(_15270_));
 AOI21_X1 _24979_ (.A(_14921_),
    .B1(_15269_),
    .B2(_15270_),
    .ZN(_15271_));
 AND2_X1 _24980_ (.A1(_14946_),
    .A2(_14884_),
    .ZN(_15272_));
 AND3_X1 _24981_ (.A1(_14887_),
    .A2(_14855_),
    .A3(_14829_),
    .ZN(_15273_));
 AND2_X1 _24982_ (.A1(_14937_),
    .A2(_14887_),
    .ZN(_15274_));
 OR3_X1 _24983_ (.A1(_15272_),
    .A2(_15273_),
    .A3(_15274_),
    .ZN(_15275_));
 AOI21_X1 _24984_ (.A(_15066_),
    .B1(_14924_),
    .B2(_15042_),
    .ZN(_15276_));
 NAND4_X1 _24985_ (.A1(_14958_),
    .A2(_14811_),
    .A3(_14897_),
    .A4(_14906_),
    .ZN(_15277_));
 OAI211_X2 _24986_ (.A(_14920_),
    .B(_15277_),
    .C1(_15006_),
    .C2(_14921_),
    .ZN(_15278_));
 NOR4_X1 _24987_ (.A1(_15271_),
    .A2(_15275_),
    .A3(_15276_),
    .A4(_15278_),
    .ZN(_15279_));
 NAND2_X1 _24988_ (.A1(_14972_),
    .A2(_14926_),
    .ZN(_15280_));
 OAI21_X1 _24989_ (.A(_14902_),
    .B1(_14812_),
    .B2(_15004_),
    .ZN(_15281_));
 OAI21_X1 _24990_ (.A(_14927_),
    .B1(_14991_),
    .B2(_14979_),
    .ZN(_15282_));
 NAND2_X1 _24991_ (.A1(_14937_),
    .A2(_14898_),
    .ZN(_15283_));
 AND4_X1 _24992_ (.A1(_15280_),
    .A2(_15281_),
    .A3(_15282_),
    .A4(_15283_),
    .ZN(_15284_));
 OAI211_X2 _24993_ (.A(_14945_),
    .B(_14906_),
    .C1(_09096_),
    .C2(_09101_),
    .ZN(_15285_));
 AND2_X1 _24994_ (.A1(_14806_),
    .A2(_09095_),
    .ZN(_15286_));
 OAI21_X1 _24995_ (.A(_14945_),
    .B1(_15024_),
    .B2(_15286_),
    .ZN(_15287_));
 OAI211_X2 _24996_ (.A(_15285_),
    .B(_15287_),
    .C1(_15089_),
    .C2(_14922_),
    .ZN(_15288_));
 OAI21_X1 _24997_ (.A(_14963_),
    .B1(_14946_),
    .B2(_14896_),
    .ZN(_15289_));
 OAI21_X1 _24998_ (.A(_15289_),
    .B1(_15150_),
    .B2(_14964_),
    .ZN(_15290_));
 AOI21_X1 _24999_ (.A(_14964_),
    .B1(_15206_),
    .B2(_15095_),
    .ZN(_15291_));
 NAND2_X1 _25000_ (.A1(_15098_),
    .A2(_14979_),
    .ZN(_15292_));
 OAI21_X1 _25001_ (.A(_15292_),
    .B1(_14964_),
    .B2(_14873_),
    .ZN(_15293_));
 NOR4_X1 _25002_ (.A1(_15288_),
    .A2(_15290_),
    .A3(_15291_),
    .A4(_15293_),
    .ZN(_15294_));
 NAND4_X1 _25003_ (.A1(_15268_),
    .A2(_15279_),
    .A3(_15284_),
    .A4(_15294_),
    .ZN(_15295_));
 NOR2_X1 _25004_ (.A1(_15260_),
    .A2(_15295_),
    .ZN(_15296_));
 XOR2_X1 _25005_ (.A(_15296_),
    .B(_01000_),
    .Z(_15297_));
 BUF_X4 _25006_ (.A(_03738_),
    .Z(_15298_));
 MUX2_X1 _25007_ (.A(_01210_),
    .B(_15297_),
    .S(_15298_),
    .Z(_01060_));
 XOR2_X1 _25008_ (.A(_17271_),
    .B(_17075_),
    .Z(_15299_));
 XOR2_X2 _25009_ (.A(_11624_),
    .B(_14014_),
    .Z(_15300_));
 XNOR2_X1 _25010_ (.A(_12358_),
    .B(_15300_),
    .ZN(_15301_));
 XOR2_X1 _25011_ (.A(_12584_),
    .B(_12904_),
    .Z(_15302_));
 XNOR2_X1 _25012_ (.A(_15301_),
    .B(_15302_),
    .ZN(_15303_));
 INV_X1 _25013_ (.A(_17271_),
    .ZN(_15304_));
 XNOR2_X1 _25014_ (.A(_15303_),
    .B(_15304_),
    .ZN(_15305_));
 BUF_X4 _25015_ (.A(_09099_),
    .Z(_15306_));
 MUX2_X1 _25016_ (.A(_15299_),
    .B(_15305_),
    .S(_15306_),
    .Z(_00685_));
 AOI211_X4 _25017_ (.A(_14960_),
    .B(_14921_),
    .C1(_15220_),
    .C2(_15150_),
    .ZN(_15307_));
 AND2_X1 _25018_ (.A1(_14918_),
    .A2(_14872_),
    .ZN(_15308_));
 AND2_X1 _25019_ (.A1(_14917_),
    .A2(_15024_),
    .ZN(_15309_));
 AOI21_X1 _25020_ (.A(_14921_),
    .B1(_15006_),
    .B2(_15223_),
    .ZN(_15310_));
 NOR4_X1 _25021_ (.A1(_15307_),
    .A2(_15308_),
    .A3(_15309_),
    .A4(_15310_),
    .ZN(_15311_));
 NAND2_X1 _25022_ (.A1(_14812_),
    .A2(_14884_),
    .ZN(_15312_));
 OAI21_X1 _25023_ (.A(_14887_),
    .B1(_15186_),
    .B2(_14901_),
    .ZN(_15313_));
 AND4_X1 _25024_ (.A1(_15190_),
    .A2(_15311_),
    .A3(_15312_),
    .A4(_15313_),
    .ZN(_15314_));
 INV_X1 _25025_ (.A(_14807_),
    .ZN(_15315_));
 AOI21_X1 _25026_ (.A(_15076_),
    .B1(_15269_),
    .B2(_15315_),
    .ZN(_15316_));
 NAND2_X1 _25027_ (.A1(_15024_),
    .A2(_14902_),
    .ZN(_15317_));
 OAI211_X2 _25028_ (.A(_14902_),
    .B(_14934_),
    .C1(_04132_),
    .C2(_09532_),
    .ZN(_15318_));
 NAND4_X1 _25029_ (.A1(_14900_),
    .A2(_15082_),
    .A3(_15317_),
    .A4(_15318_),
    .ZN(_15319_));
 NOR4_X1 _25030_ (.A1(_15316_),
    .A2(_15319_),
    .A3(_14930_),
    .A4(_15077_),
    .ZN(_15320_));
 NAND2_X1 _25031_ (.A1(_14945_),
    .A2(_14953_),
    .ZN(_15321_));
 AND2_X1 _25032_ (.A1(_14963_),
    .A2(_14860_),
    .ZN(_15322_));
 AOI211_X4 _25033_ (.A(_14968_),
    .B(_15322_),
    .C1(_14950_),
    .C2(_15098_),
    .ZN(_15323_));
 OAI21_X1 _25034_ (.A(_14945_),
    .B1(_15070_),
    .B2(_14989_),
    .ZN(_15324_));
 OAI21_X1 _25035_ (.A(_15098_),
    .B1(_14947_),
    .B2(_14833_),
    .ZN(_15325_));
 AND4_X1 _25036_ (.A1(_15321_),
    .A2(_15323_),
    .A3(_15324_),
    .A4(_15325_),
    .ZN(_15326_));
 NOR3_X1 _25037_ (.A1(_14855_),
    .A2(_17166_),
    .A3(_14826_),
    .ZN(_15327_));
 OAI21_X1 _25038_ (.A(_14977_),
    .B1(_14841_),
    .B2(_15327_),
    .ZN(_15328_));
 AND2_X1 _25039_ (.A1(_14985_),
    .A2(_14947_),
    .ZN(_15329_));
 AND2_X1 _25040_ (.A1(_14984_),
    .A2(_14937_),
    .ZN(_15330_));
 NOR4_X1 _25041_ (.A1(_15329_),
    .A2(_15263_),
    .A3(_15330_),
    .A4(_15262_),
    .ZN(_15331_));
 OAI21_X1 _25042_ (.A(_14985_),
    .B1(_14876_),
    .B2(_14910_),
    .ZN(_15332_));
 NAND2_X1 _25043_ (.A1(_14977_),
    .A2(_15029_),
    .ZN(_15333_));
 NAND2_X1 _25044_ (.A1(_14970_),
    .A2(_14877_),
    .ZN(_15334_));
 NAND2_X1 _25045_ (.A1(_14970_),
    .A2(_14890_),
    .ZN(_15335_));
 AND3_X1 _25046_ (.A1(_15333_),
    .A2(_15334_),
    .A3(_15335_),
    .ZN(_15336_));
 AND4_X1 _25047_ (.A1(_15328_),
    .A2(_15331_),
    .A3(_15332_),
    .A4(_15336_),
    .ZN(_15337_));
 NAND4_X1 _25048_ (.A1(_15314_),
    .A2(_15320_),
    .A3(_15326_),
    .A4(_15337_),
    .ZN(_15338_));
 INV_X1 _25049_ (.A(_14860_),
    .ZN(_15339_));
 AOI21_X1 _25050_ (.A(_15007_),
    .B1(_15339_),
    .B2(_15145_),
    .ZN(_15340_));
 AOI211_X4 _25051_ (.A(_15257_),
    .B(_15340_),
    .C1(_15111_),
    .C2(_15245_),
    .ZN(_15341_));
 AND2_X1 _25052_ (.A1(_15019_),
    .A2(_14836_),
    .ZN(_15342_));
 NOR3_X1 _25053_ (.A1(_15129_),
    .A2(_15253_),
    .A3(_15342_),
    .ZN(_15343_));
 AND4_X1 _25054_ (.A1(_15023_),
    .A2(_15341_),
    .A3(_15025_),
    .A4(_15343_),
    .ZN(_15344_));
 AOI21_X1 _25055_ (.A(_15119_),
    .B1(_14873_),
    .B2(_14911_),
    .ZN(_15345_));
 AOI21_X1 _25056_ (.A(_15119_),
    .B1(_15095_),
    .B2(_15185_),
    .ZN(_15346_));
 AOI21_X1 _25057_ (.A(_15152_),
    .B1(_14849_),
    .B2(_15095_),
    .ZN(_15347_));
 NOR4_X1 _25058_ (.A1(_15345_),
    .A2(_15346_),
    .A3(_15347_),
    .A4(_15124_),
    .ZN(_15348_));
 OAI21_X1 _25059_ (.A(_15038_),
    .B1(_15024_),
    .B2(_14833_),
    .ZN(_15349_));
 OAI21_X1 _25060_ (.A(_15349_),
    .B1(_15220_),
    .B2(_15040_),
    .ZN(_15350_));
 NAND2_X1 _25061_ (.A1(_15038_),
    .A2(_14836_),
    .ZN(_15351_));
 OAI221_X1 _25062_ (.A(_15351_),
    .B1(_15040_),
    .B2(_15069_),
    .C1(_15142_),
    .C2(_04132_),
    .ZN(_15352_));
 AOI21_X1 _25063_ (.A(_15135_),
    .B1(_15071_),
    .B2(_15069_),
    .ZN(_15353_));
 NOR4_X1 _25064_ (.A1(_15138_),
    .A2(_15350_),
    .A3(_15352_),
    .A4(_15353_),
    .ZN(_15354_));
 INV_X1 _25065_ (.A(_15231_),
    .ZN(_15355_));
 OAI211_X2 _25066_ (.A(_15355_),
    .B(_14814_),
    .C1(_14822_),
    .C2(_15315_),
    .ZN(_15356_));
 AOI21_X1 _25067_ (.A(_14868_),
    .B1(_14980_),
    .B2(_15079_),
    .ZN(_15357_));
 NOR4_X1 _25068_ (.A1(_15356_),
    .A2(_15172_),
    .A3(_15051_),
    .A4(_15357_),
    .ZN(_15358_));
 NAND4_X1 _25069_ (.A1(_15344_),
    .A2(_15348_),
    .A3(_15354_),
    .A4(_15358_),
    .ZN(_15359_));
 NOR2_X1 _25070_ (.A1(_15338_),
    .A2(_15359_),
    .ZN(_15360_));
 XOR2_X1 _25071_ (.A(_15360_),
    .B(_01001_),
    .Z(_15361_));
 MUX2_X1 _25072_ (.A(_01211_),
    .B(_15361_),
    .S(_15298_),
    .Z(_01061_));
 AND3_X1 _25073_ (.A1(_14872_),
    .A2(_15016_),
    .A3(_14954_),
    .ZN(_15362_));
 OAI211_X2 _25074_ (.A(_15011_),
    .B(_14829_),
    .C1(_14960_),
    .C2(_09101_),
    .ZN(_15363_));
 OAI21_X1 _25075_ (.A(_15011_),
    .B1(_14896_),
    .B2(_14936_),
    .ZN(_15364_));
 NAND2_X1 _25076_ (.A1(_15363_),
    .A2(_15364_),
    .ZN(_15365_));
 AOI21_X1 _25077_ (.A(_15119_),
    .B1(_15006_),
    .B2(_14875_),
    .ZN(_15366_));
 OR4_X1 _25078_ (.A1(_15362_),
    .A2(_15246_),
    .A3(_15365_),
    .A4(_15366_),
    .ZN(_15367_));
 AOI21_X1 _25079_ (.A(_15040_),
    .B1(_14914_),
    .B2(_15206_),
    .ZN(_15368_));
 AND2_X1 _25080_ (.A1(_14854_),
    .A2(_14823_),
    .ZN(_15369_));
 AND2_X1 _25081_ (.A1(_14854_),
    .A2(_14949_),
    .ZN(_15370_));
 AND2_X1 _25082_ (.A1(_14854_),
    .A2(_14910_),
    .ZN(_15371_));
 NOR4_X1 _25083_ (.A1(_15368_),
    .A2(_15369_),
    .A3(_15370_),
    .A4(_15371_),
    .ZN(_15372_));
 AOI21_X1 _25084_ (.A(_15146_),
    .B1(_14950_),
    .B2(_15044_),
    .ZN(_15373_));
 NAND4_X1 _25085_ (.A1(_15044_),
    .A2(_14934_),
    .A3(_14848_),
    .A4(_14856_),
    .ZN(_15374_));
 OAI21_X1 _25086_ (.A(_15044_),
    .B1(_14972_),
    .B2(_15266_),
    .ZN(_15375_));
 NAND4_X1 _25087_ (.A1(_15372_),
    .A2(_15373_),
    .A3(_15374_),
    .A4(_15375_),
    .ZN(_15376_));
 AND2_X1 _25088_ (.A1(_15019_),
    .A2(_14938_),
    .ZN(_15377_));
 AOI211_X4 _25089_ (.A(_15377_),
    .B(_15250_),
    .C1(_14913_),
    .C2(_15019_),
    .ZN(_15378_));
 AND2_X1 _25090_ (.A1(_14947_),
    .A2(_15001_),
    .ZN(_15379_));
 AND2_X1 _25091_ (.A1(_14901_),
    .A2(_15001_),
    .ZN(_15380_));
 AND2_X1 _25092_ (.A1(_15001_),
    .A2(_14833_),
    .ZN(_15381_));
 AND2_X1 _25093_ (.A1(_15001_),
    .A2(_14845_),
    .ZN(_15382_));
 NOR4_X1 _25094_ (.A1(_15379_),
    .A2(_15380_),
    .A3(_15381_),
    .A4(_15382_),
    .ZN(_15383_));
 NAND2_X1 _25095_ (.A1(_15022_),
    .A2(_14819_),
    .ZN(_15384_));
 INV_X1 _25096_ (.A(_15342_),
    .ZN(_15385_));
 NAND2_X1 _25097_ (.A1(_14910_),
    .A2(_15019_),
    .ZN(_15386_));
 NAND3_X1 _25098_ (.A1(_15029_),
    .A2(_14866_),
    .A3(_15016_),
    .ZN(_15387_));
 AND4_X1 _25099_ (.A1(_15384_),
    .A2(_15385_),
    .A3(_15386_),
    .A4(_15387_),
    .ZN(_15388_));
 OAI21_X1 _25100_ (.A(_15111_),
    .B1(_15004_),
    .B2(_15009_),
    .ZN(_15389_));
 NAND4_X1 _25101_ (.A1(_15378_),
    .A2(_15383_),
    .A3(_15388_),
    .A4(_15389_),
    .ZN(_15390_));
 AND2_X1 _25102_ (.A1(_14991_),
    .A2(_14820_),
    .ZN(_15391_));
 NOR3_X1 _25103_ (.A1(_15391_),
    .A2(_15233_),
    .A3(_15058_),
    .ZN(_15392_));
 OAI21_X1 _25104_ (.A(_14871_),
    .B1(_14947_),
    .B2(_14913_),
    .ZN(_15393_));
 OAI21_X1 _25105_ (.A(_14871_),
    .B1(_14812_),
    .B2(_14950_),
    .ZN(_15394_));
 OAI21_X1 _25106_ (.A(_14820_),
    .B1(_15035_),
    .B2(_15286_),
    .ZN(_15395_));
 NAND4_X1 _25107_ (.A1(_15392_),
    .A2(_15393_),
    .A3(_15394_),
    .A4(_15395_),
    .ZN(_15396_));
 NOR4_X1 _25108_ (.A1(_15367_),
    .A2(_15376_),
    .A3(_15390_),
    .A4(_15396_),
    .ZN(_15397_));
 AND2_X1 _25109_ (.A1(_15224_),
    .A2(_14917_),
    .ZN(_15398_));
 AND3_X1 _25110_ (.A1(_14850_),
    .A2(_14917_),
    .A3(_14856_),
    .ZN(_15399_));
 AOI21_X1 _25111_ (.A(_14921_),
    .B1(_14915_),
    .B2(_15095_),
    .ZN(_15400_));
 OR4_X1 _25112_ (.A1(_15308_),
    .A2(_15398_),
    .A3(_15399_),
    .A4(_15400_),
    .ZN(_15401_));
 NOR2_X1 _25113_ (.A1(_15066_),
    .A2(_14922_),
    .ZN(_15402_));
 AOI221_X4 _25114_ (.A(_15066_),
    .B1(_14960_),
    .B2(_09531_),
    .C1(_15315_),
    .C2(_14869_),
    .ZN(_15403_));
 NOR4_X1 _25115_ (.A1(_15401_),
    .A2(_15191_),
    .A3(_15402_),
    .A4(_15403_),
    .ZN(_15404_));
 OAI21_X1 _25116_ (.A(_14902_),
    .B1(_14947_),
    .B2(_14957_),
    .ZN(_15405_));
 OAI211_X2 _25117_ (.A(_15405_),
    .B(_14904_),
    .C1(_14914_),
    .C2(_14908_),
    .ZN(_15406_));
 OAI211_X2 _25118_ (.A(_15199_),
    .B(_15201_),
    .C1(_14922_),
    .C2(_15076_),
    .ZN(_15407_));
 NAND2_X1 _25119_ (.A1(_14926_),
    .A2(_14833_),
    .ZN(_15408_));
 NAND4_X1 _25120_ (.A1(_14866_),
    .A2(_09096_),
    .A3(_14841_),
    .A4(_14897_),
    .ZN(_15409_));
 OAI211_X2 _25121_ (.A(_15408_),
    .B(_15409_),
    .C1(_15206_),
    .C2(_15076_),
    .ZN(_15410_));
 AND4_X1 _25122_ (.A1(_14830_),
    .A2(_14805_),
    .A3(_14897_),
    .A4(_14906_),
    .ZN(_15411_));
 NOR4_X1 _25123_ (.A1(_15406_),
    .A2(_15407_),
    .A3(_15410_),
    .A4(_15411_),
    .ZN(_15412_));
 NAND2_X1 _25124_ (.A1(_14984_),
    .A2(_15013_),
    .ZN(_15413_));
 OAI21_X1 _25125_ (.A(_15413_),
    .B1(_15094_),
    .B2(_14880_),
    .ZN(_15414_));
 AND2_X1 _25126_ (.A1(_14984_),
    .A2(_14910_),
    .ZN(_15415_));
 OR3_X1 _25127_ (.A1(_15414_),
    .A2(_15415_),
    .A3(_15092_),
    .ZN(_15416_));
 OAI21_X1 _25128_ (.A(_14945_),
    .B1(_14836_),
    .B2(_14979_),
    .ZN(_15417_));
 NAND3_X1 _25129_ (.A1(_15417_),
    .A2(_14948_),
    .A3(_14955_),
    .ZN(_15418_));
 OAI21_X1 _25130_ (.A(_15098_),
    .B1(_14910_),
    .B2(_14877_),
    .ZN(_15419_));
 OAI21_X1 _25131_ (.A(_15098_),
    .B1(_14901_),
    .B2(_14833_),
    .ZN(_15420_));
 OAI211_X2 _25132_ (.A(_15419_),
    .B(_15420_),
    .C1(_14873_),
    .C2(_14964_),
    .ZN(_15421_));
 OAI21_X1 _25133_ (.A(_14977_),
    .B1(_14913_),
    .B2(_15050_),
    .ZN(_15422_));
 NAND2_X1 _25134_ (.A1(_14977_),
    .A2(_14991_),
    .ZN(_15423_));
 NAND4_X1 _25135_ (.A1(_14973_),
    .A2(_15422_),
    .A3(_15423_),
    .A4(_15335_),
    .ZN(_15424_));
 NOR4_X1 _25136_ (.A1(_15416_),
    .A2(_15418_),
    .A3(_15421_),
    .A4(_15424_),
    .ZN(_15425_));
 NAND4_X1 _25137_ (.A1(_15397_),
    .A2(_15404_),
    .A3(_15412_),
    .A4(_15425_),
    .ZN(_15426_));
 NOR2_X1 _25138_ (.A1(_15426_),
    .A2(_15030_),
    .ZN(_15427_));
 INV_X1 _25139_ (.A(_01002_),
    .ZN(_15428_));
 XNOR2_X1 _25140_ (.A(_15427_),
    .B(_15428_),
    .ZN(_15429_));
 MUX2_X1 _25141_ (.A(_01212_),
    .B(_15429_),
    .S(_15298_),
    .Z(_01062_));
 OAI21_X1 _25142_ (.A(_15044_),
    .B1(_15004_),
    .B2(_14991_),
    .ZN(_15430_));
 OAI21_X1 _25143_ (.A(_14803_),
    .B1(_14972_),
    .B2(_14901_),
    .ZN(_15431_));
 NAND3_X1 _25144_ (.A1(_14820_),
    .A2(_14859_),
    .A3(_14816_),
    .ZN(_15432_));
 AND4_X1 _25145_ (.A1(_15062_),
    .A2(_15234_),
    .A3(_15431_),
    .A4(_15432_),
    .ZN(_15433_));
 OAI21_X1 _25146_ (.A(_14867_),
    .B1(_14877_),
    .B2(_14950_),
    .ZN(_15434_));
 AND4_X1 _25147_ (.A1(_15238_),
    .A2(_15433_),
    .A3(_15174_),
    .A4(_15434_),
    .ZN(_15435_));
 OAI21_X1 _25148_ (.A(_15038_),
    .B1(_14972_),
    .B2(_15266_),
    .ZN(_15436_));
 OAI211_X2 _25149_ (.A(_14802_),
    .B(_14958_),
    .C1(_14989_),
    .C2(_15029_),
    .ZN(_15437_));
 NAND4_X1 _25150_ (.A1(_14958_),
    .A2(_09095_),
    .A3(_14934_),
    .A4(_14802_),
    .ZN(_15438_));
 AND3_X1 _25151_ (.A1(_15436_),
    .A2(_15437_),
    .A3(_15438_),
    .ZN(_15439_));
 AND2_X1 _25152_ (.A1(_14936_),
    .A2(_14839_),
    .ZN(_15440_));
 AOI211_X4 _25153_ (.A(_15440_),
    .B(_15226_),
    .C1(_15035_),
    .C2(_14839_),
    .ZN(_15441_));
 AND4_X1 _25154_ (.A1(_15430_),
    .A2(_15435_),
    .A3(_15439_),
    .A4(_15441_),
    .ZN(_15442_));
 AND2_X1 _25155_ (.A1(_14983_),
    .A2(_14823_),
    .ZN(_15443_));
 AOI221_X4 _25156_ (.A(_15180_),
    .B1(_14877_),
    .B2(_14984_),
    .C1(_14960_),
    .C2(_15443_),
    .ZN(_15444_));
 NAND2_X1 _25157_ (.A1(_14985_),
    .A2(_14987_),
    .ZN(_15445_));
 OAI211_X2 _25158_ (.A(_15444_),
    .B(_15445_),
    .C1(_15270_),
    .C2(_15094_),
    .ZN(_15446_));
 NOR2_X1 _25159_ (.A1(_15290_),
    .A2(_15099_),
    .ZN(_15447_));
 OAI211_X2 _25160_ (.A(_15447_),
    .B(_15292_),
    .C1(_14966_),
    .C2(_14964_),
    .ZN(_15448_));
 NAND4_X1 _25161_ (.A1(_14952_),
    .A2(_09096_),
    .A3(_14953_),
    .A4(_14954_),
    .ZN(_15449_));
 OAI211_X2 _25162_ (.A(_15087_),
    .B(_15449_),
    .C1(_14924_),
    .C2(_15089_),
    .ZN(_15450_));
 AND2_X1 _25163_ (.A1(_14970_),
    .A2(_15113_),
    .ZN(_15451_));
 AND2_X1 _25164_ (.A1(_14970_),
    .A2(_15035_),
    .ZN(_15452_));
 AND3_X1 _25165_ (.A1(_15004_),
    .A2(_14830_),
    .A3(_14943_),
    .ZN(_15453_));
 OR4_X4 _25166_ (.A1(_15451_),
    .A2(_15105_),
    .A3(_15452_),
    .A4(_15453_),
    .ZN(_15454_));
 NOR4_X1 _25167_ (.A1(_15446_),
    .A2(_15448_),
    .A3(_15450_),
    .A4(_15454_),
    .ZN(_15455_));
 INV_X1 _25168_ (.A(_15253_),
    .ZN(_15456_));
 NAND2_X1 _25169_ (.A1(_15021_),
    .A2(_15456_),
    .ZN(_15457_));
 AND3_X1 _25170_ (.A1(_15029_),
    .A2(_14866_),
    .A3(_15016_),
    .ZN(_15458_));
 OR4_X1 _25171_ (.A1(_15377_),
    .A2(_15457_),
    .A3(_15128_),
    .A4(_15458_),
    .ZN(_15459_));
 OAI21_X1 _25172_ (.A(_15012_),
    .B1(_14876_),
    .B2(_15070_),
    .ZN(_15460_));
 NAND2_X1 _25173_ (.A1(_15012_),
    .A2(_14957_),
    .ZN(_15461_));
 NAND4_X1 _25174_ (.A1(_14953_),
    .A2(_15016_),
    .A3(_09096_),
    .A4(_14954_),
    .ZN(_15462_));
 NAND4_X1 _25175_ (.A1(_15460_),
    .A2(_15461_),
    .A3(_15154_),
    .A4(_15462_),
    .ZN(_15463_));
 NAND2_X1 _25176_ (.A1(_15186_),
    .A2(_14997_),
    .ZN(_15464_));
 OAI211_X2 _25177_ (.A(_14958_),
    .B(_15016_),
    .C1(_15029_),
    .C2(_14823_),
    .ZN(_15465_));
 OAI211_X2 _25178_ (.A(_15464_),
    .B(_15465_),
    .C1(_15206_),
    .C2(_15119_),
    .ZN(_15466_));
 OAI21_X1 _25179_ (.A(_15111_),
    .B1(_14989_),
    .B2(_14950_),
    .ZN(_15467_));
 OAI211_X2 _25180_ (.A(_15111_),
    .B(_17169_),
    .C1(_09532_),
    .C2(_14809_),
    .ZN(_15468_));
 OAI211_X2 _25181_ (.A(_15467_),
    .B(_15468_),
    .C1(_14924_),
    .C2(_15007_),
    .ZN(_15469_));
 NOR4_X1 _25182_ (.A1(_15459_),
    .A2(_15463_),
    .A3(_15466_),
    .A4(_15469_),
    .ZN(_15470_));
 OAI21_X1 _25183_ (.A(_14918_),
    .B1(_15009_),
    .B2(_14934_),
    .ZN(_15471_));
 AND3_X1 _25184_ (.A1(_14892_),
    .A2(_15312_),
    .A3(_14894_),
    .ZN(_15472_));
 AND3_X1 _25185_ (.A1(_15472_),
    .A2(_15190_),
    .A3(_15189_),
    .ZN(_15473_));
 OAI211_X2 _25186_ (.A(_14900_),
    .B(_15283_),
    .C1(_14914_),
    .C2(_14908_),
    .ZN(_15474_));
 AND2_X1 _25187_ (.A1(_14902_),
    .A2(_15041_),
    .ZN(_15475_));
 NAND2_X1 _25188_ (.A1(_14926_),
    .A2(_14936_),
    .ZN(_15476_));
 NAND3_X1 _25189_ (.A1(_15408_),
    .A2(_15280_),
    .A3(_15476_),
    .ZN(_15477_));
 NAND2_X1 _25190_ (.A1(_14991_),
    .A2(_14927_),
    .ZN(_15478_));
 NAND2_X1 _25191_ (.A1(_15478_),
    .A2(_15202_),
    .ZN(_15479_));
 NOR4_X1 _25192_ (.A1(_15474_),
    .A2(_15475_),
    .A3(_15477_),
    .A4(_15479_),
    .ZN(_15480_));
 AOI211_X4 _25193_ (.A(_15073_),
    .B(_15309_),
    .C1(_14918_),
    .C2(_14896_),
    .ZN(_15481_));
 AND4_X1 _25194_ (.A1(_15471_),
    .A2(_15473_),
    .A3(_15480_),
    .A4(_15481_),
    .ZN(_15482_));
 NAND4_X1 _25195_ (.A1(_15442_),
    .A2(_15455_),
    .A3(_15470_),
    .A4(_15482_),
    .ZN(_15483_));
 NOR2_X2 _25196_ (.A1(_15483_),
    .A2(_15030_),
    .ZN(_15484_));
 INV_X1 _25197_ (.A(_01003_),
    .ZN(_15485_));
 XNOR2_X1 _25198_ (.A(_15484_),
    .B(_15485_),
    .ZN(_15486_));
 MUX2_X1 _25199_ (.A(_01214_),
    .B(_15486_),
    .S(_15298_),
    .Z(_01063_));
 AOI21_X1 _25200_ (.A(_15066_),
    .B1(_15222_),
    .B2(_15223_),
    .ZN(_15487_));
 AOI211_X4 _25201_ (.A(_15272_),
    .B(_15487_),
    .C1(_14845_),
    .C2(_14887_),
    .ZN(_15488_));
 AND2_X1 _25202_ (.A1(_14917_),
    .A2(_14836_),
    .ZN(_15489_));
 AOI211_X4 _25203_ (.A(_15489_),
    .B(_15398_),
    .C1(_14918_),
    .C2(_14950_),
    .ZN(_15490_));
 AND2_X1 _25204_ (.A1(_14918_),
    .A2(_14901_),
    .ZN(_15491_));
 NOR3_X1 _25205_ (.A1(_15491_),
    .A2(_15074_),
    .A3(_15309_),
    .ZN(_15492_));
 OAI21_X1 _25206_ (.A(_14918_),
    .B1(_14957_),
    .B2(_14845_),
    .ZN(_15493_));
 AND4_X1 _25207_ (.A1(_15488_),
    .A2(_15490_),
    .A3(_15492_),
    .A4(_15493_),
    .ZN(_15494_));
 NAND2_X1 _25208_ (.A1(_14984_),
    .A2(_15024_),
    .ZN(_15495_));
 OAI21_X1 _25209_ (.A(_15495_),
    .B1(_15094_),
    .B2(_15220_),
    .ZN(_15496_));
 OR4_X1 _25210_ (.A1(_15179_),
    .A2(_15496_),
    .A3(_15443_),
    .A4(_15180_),
    .ZN(_15497_));
 AND2_X1 _25211_ (.A1(_14977_),
    .A2(_15327_),
    .ZN(_15498_));
 NAND3_X1 _25212_ (.A1(_15004_),
    .A2(_14830_),
    .A3(_14952_),
    .ZN(_15499_));
 OAI211_X2 _25213_ (.A(_15334_),
    .B(_15499_),
    .C1(_14981_),
    .C2(_15042_),
    .ZN(_15500_));
 NOR4_X1 _25214_ (.A1(_15497_),
    .A2(_15105_),
    .A3(_15498_),
    .A4(_15500_),
    .ZN(_15501_));
 NAND4_X1 _25215_ (.A1(_14931_),
    .A2(_14933_),
    .A3(_15202_),
    .A4(_15280_),
    .ZN(_15502_));
 AND4_X1 _25216_ (.A1(_09101_),
    .A2(_14829_),
    .A3(_14830_),
    .A4(_14897_),
    .ZN(_15503_));
 NAND2_X1 _25217_ (.A1(_15082_),
    .A2(_15283_),
    .ZN(_15504_));
 AOI21_X1 _25218_ (.A(_14908_),
    .B1(_14980_),
    .B2(_15042_),
    .ZN(_15505_));
 NOR4_X1 _25219_ (.A1(_15502_),
    .A2(_15503_),
    .A3(_15504_),
    .A4(_15505_),
    .ZN(_15506_));
 OAI21_X1 _25220_ (.A(_15098_),
    .B1(_14861_),
    .B2(_14910_),
    .ZN(_15507_));
 NAND4_X1 _25221_ (.A1(_14852_),
    .A2(_14952_),
    .A3(_14960_),
    .A4(_14906_),
    .ZN(_15508_));
 AND2_X1 _25222_ (.A1(_15507_),
    .A2(_15508_),
    .ZN(_15509_));
 OAI21_X1 _25223_ (.A(_15098_),
    .B1(_15245_),
    .B2(_14957_),
    .ZN(_15510_));
 OAI21_X1 _25224_ (.A(_14945_),
    .B1(_14991_),
    .B2(_15004_),
    .ZN(_15511_));
 OAI21_X1 _25225_ (.A(_14944_),
    .B1(_14833_),
    .B2(_14879_),
    .ZN(_15512_));
 AND4_X1 _25226_ (.A1(_15509_),
    .A2(_15510_),
    .A3(_15511_),
    .A4(_15512_),
    .ZN(_15513_));
 AND4_X1 _25227_ (.A1(_15494_),
    .A2(_15501_),
    .A3(_15506_),
    .A4(_15513_),
    .ZN(_15514_));
 AND2_X1 _25228_ (.A1(_15050_),
    .A2(_15011_),
    .ZN(_15515_));
 INV_X1 _25229_ (.A(_15515_),
    .ZN(_15516_));
 NOR2_X1 _25230_ (.A1(_14896_),
    .A2(_14936_),
    .ZN(_15517_));
 NOR2_X1 _25231_ (.A1(_15119_),
    .A2(_15517_),
    .ZN(_15518_));
 AOI21_X1 _25232_ (.A(_15518_),
    .B1(_14997_),
    .B2(_15245_),
    .ZN(_15519_));
 OAI21_X1 _25233_ (.A(_14997_),
    .B1(_14890_),
    .B2(_15041_),
    .ZN(_15520_));
 OAI21_X1 _25234_ (.A(_15012_),
    .B1(_14876_),
    .B2(_14861_),
    .ZN(_15521_));
 AND4_X1 _25235_ (.A1(_15516_),
    .A2(_15519_),
    .A3(_15520_),
    .A4(_15521_),
    .ZN(_15522_));
 NOR2_X1 _25236_ (.A1(_15371_),
    .A2(_14858_),
    .ZN(_15523_));
 OAI21_X1 _25237_ (.A(_15038_),
    .B1(_14957_),
    .B2(_14845_),
    .ZN(_15524_));
 OAI211_X2 _25238_ (.A(_15523_),
    .B(_15524_),
    .C1(_15040_),
    .C2(_14914_),
    .ZN(_15525_));
 AND2_X1 _25239_ (.A1(_15044_),
    .A2(_15029_),
    .ZN(_15526_));
 AND2_X1 _25240_ (.A1(_15144_),
    .A2(_14848_),
    .ZN(_15527_));
 OAI211_X2 _25241_ (.A(_14839_),
    .B(_14841_),
    .C1(_14960_),
    .C2(_09101_),
    .ZN(_15528_));
 OAI21_X1 _25242_ (.A(_15528_),
    .B1(_15206_),
    .B2(_15135_),
    .ZN(_15529_));
 NOR4_X1 _25243_ (.A1(_15525_),
    .A2(_15526_),
    .A3(_15527_),
    .A4(_15529_),
    .ZN(_15530_));
 NOR2_X1 _25244_ (.A1(_15379_),
    .A2(_15381_),
    .ZN(_15531_));
 AOI21_X1 _25245_ (.A(_15008_),
    .B1(_15111_),
    .B2(_14950_),
    .ZN(_15532_));
 OAI221_X1 _25246_ (.A(_15022_),
    .B1(_09095_),
    .B2(_09532_),
    .C1(_14841_),
    .C2(_14953_),
    .ZN(_15533_));
 AND4_X1 _25247_ (.A1(_15531_),
    .A2(_15532_),
    .A3(_15387_),
    .A4(_15533_),
    .ZN(_15534_));
 AND2_X1 _25248_ (.A1(_14929_),
    .A2(_14803_),
    .ZN(_15535_));
 AND2_X1 _25249_ (.A1(_14803_),
    .A2(_15286_),
    .ZN(_15536_));
 OR4_X1 _25250_ (.A1(_15058_),
    .A2(_15231_),
    .A3(_15535_),
    .A4(_15536_),
    .ZN(_15537_));
 AOI21_X1 _25251_ (.A(_14868_),
    .B1(_15145_),
    .B2(_15069_),
    .ZN(_15538_));
 NAND2_X1 _25252_ (.A1(_14870_),
    .A2(_15056_),
    .ZN(_15539_));
 OAI21_X1 _25253_ (.A(_15168_),
    .B1(_15339_),
    .B2(_14868_),
    .ZN(_15540_));
 NOR4_X1 _25254_ (.A1(_15537_),
    .A2(_15538_),
    .A3(_15539_),
    .A4(_15540_),
    .ZN(_15541_));
 AND4_X1 _25255_ (.A1(_15522_),
    .A2(_15530_),
    .A3(_15534_),
    .A4(_15541_),
    .ZN(_15542_));
 AND2_X1 _25256_ (.A1(_15514_),
    .A2(_15542_),
    .ZN(_15543_));
 INV_X1 _25257_ (.A(_01004_),
    .ZN(_15544_));
 XNOR2_X1 _25258_ (.A(_15543_),
    .B(_15544_),
    .ZN(_15545_));
 MUX2_X1 _25259_ (.A(_01215_),
    .B(_15545_),
    .S(_15298_),
    .Z(_01064_));
 INV_X1 _25260_ (.A(_17146_),
    .ZN(_15546_));
 NOR2_X1 _25261_ (.A1(_15546_),
    .A2(_17145_),
    .ZN(_15547_));
 NOR2_X1 _25262_ (.A1(_17174_),
    .A2(_17175_),
    .ZN(_15548_));
 AND2_X1 _25263_ (.A1(_15547_),
    .A2(_15548_),
    .ZN(_15549_));
 AND2_X1 _25264_ (.A1(_17147_),
    .A2(_17148_),
    .ZN(_15550_));
 CLKBUF_X2 _25265_ (.A(_15550_),
    .Z(_15551_));
 NOR2_X1 _25266_ (.A1(_17149_),
    .A2(_17150_),
    .ZN(_15552_));
 AND2_X1 _25267_ (.A1(_15551_),
    .A2(_15552_),
    .ZN(_15553_));
 BUF_X4 _25268_ (.A(_15553_),
    .Z(_15554_));
 AND2_X1 _25269_ (.A1(_15549_),
    .A2(_15554_),
    .ZN(_15555_));
 NOR2_X1 _25270_ (.A1(_17145_),
    .A2(_17146_),
    .ZN(_15556_));
 BUF_X2 _25271_ (.A(_15556_),
    .Z(_15557_));
 INV_X1 _25272_ (.A(_15557_),
    .ZN(_15558_));
 NOR2_X1 _25273_ (.A1(_15558_),
    .A2(_15548_),
    .ZN(_15559_));
 AND2_X1 _25274_ (.A1(_15559_),
    .A2(_15554_),
    .ZN(_15560_));
 NOR2_X1 _25275_ (.A1(_15555_),
    .A2(_15560_),
    .ZN(_15561_));
 AND2_X2 _25276_ (.A1(_11041_),
    .A2(_17150_),
    .ZN(_15562_));
 NOR2_X1 _25277_ (.A1(_17147_),
    .A2(_17148_),
    .ZN(_15563_));
 AND2_X2 _25278_ (.A1(_15562_),
    .A2(_15563_),
    .ZN(_15564_));
 AND2_X1 _25279_ (.A1(_17145_),
    .A2(_17146_),
    .ZN(_15565_));
 INV_X1 _25280_ (.A(_15565_),
    .ZN(_15566_));
 NOR2_X1 _25281_ (.A1(_15566_),
    .A2(_15548_),
    .ZN(_15567_));
 AND2_X1 _25282_ (.A1(_15564_),
    .A2(_15567_),
    .ZN(_15568_));
 INV_X1 _25283_ (.A(_17145_),
    .ZN(_15569_));
 NOR2_X1 _25284_ (.A1(_15569_),
    .A2(_17146_),
    .ZN(_15570_));
 CLKBUF_X2 _25285_ (.A(_15570_),
    .Z(_15571_));
 AND2_X1 _25286_ (.A1(_15571_),
    .A2(_15548_),
    .ZN(_15572_));
 BUF_X2 _25287_ (.A(_15572_),
    .Z(_15573_));
 NOR2_X1 _25288_ (.A1(_11035_),
    .A2(_17147_),
    .ZN(_15574_));
 AND2_X1 _25289_ (.A1(_15562_),
    .A2(_15574_),
    .ZN(_15575_));
 BUF_X2 _25290_ (.A(_15575_),
    .Z(_15576_));
 AND2_X1 _25291_ (.A1(_15562_),
    .A2(_15551_),
    .ZN(_15577_));
 BUF_X4 _25292_ (.A(_15577_),
    .Z(_15578_));
 INV_X1 _25293_ (.A(_17174_),
    .ZN(_15579_));
 NOR2_X1 _25294_ (.A1(_15579_),
    .A2(_11003_),
    .ZN(_15580_));
 BUF_X4 _25295_ (.A(_15580_),
    .Z(_15581_));
 NOR2_X1 _25296_ (.A1(_15558_),
    .A2(_15581_),
    .ZN(_15582_));
 AND2_X1 _25297_ (.A1(_15565_),
    .A2(_15548_),
    .ZN(_15583_));
 BUF_X2 _25298_ (.A(_15583_),
    .Z(_15584_));
 NOR2_X1 _25299_ (.A1(_15582_),
    .A2(_15584_),
    .ZN(_15585_));
 INV_X1 _25300_ (.A(_15585_),
    .ZN(_15586_));
 AOI221_X4 _25301_ (.A(_15568_),
    .B1(_15573_),
    .B2(_15576_),
    .C1(_15578_),
    .C2(_15586_),
    .ZN(_15587_));
 BUF_X2 _25302_ (.A(_15565_),
    .Z(_15588_));
 AND2_X1 _25303_ (.A1(_17174_),
    .A2(_17175_),
    .ZN(_15589_));
 BUF_X4 _25304_ (.A(_15589_),
    .Z(_15590_));
 AND2_X2 _25305_ (.A1(_15588_),
    .A2(_15590_),
    .ZN(_15591_));
 AND2_X1 _25306_ (.A1(_15591_),
    .A2(_15553_),
    .ZN(_15592_));
 NOR2_X1 _25307_ (.A1(_11041_),
    .A2(_17150_),
    .ZN(_15593_));
 AND2_X2 _25308_ (.A1(_15593_),
    .A2(_15563_),
    .ZN(_15594_));
 AND2_X2 _25309_ (.A1(_15571_),
    .A2(_11003_),
    .ZN(_15595_));
 BUF_X2 _25310_ (.A(_15574_),
    .Z(_15596_));
 AND2_X1 _25311_ (.A1(_15596_),
    .A2(_15593_),
    .ZN(_15597_));
 BUF_X4 _25312_ (.A(_15597_),
    .Z(_15598_));
 AOI221_X4 _25313_ (.A(_15592_),
    .B1(_15573_),
    .B2(_15594_),
    .C1(_15595_),
    .C2(_15598_),
    .ZN(_15599_));
 NOR2_X2 _25314_ (.A1(_11010_),
    .A2(_17174_),
    .ZN(_15600_));
 AND2_X1 _25315_ (.A1(_15600_),
    .A2(_15571_),
    .ZN(_15601_));
 BUF_X2 _25316_ (.A(_15601_),
    .Z(_15602_));
 BUF_X4 _25317_ (.A(_15554_),
    .Z(_15603_));
 AND2_X1 _25318_ (.A1(_15574_),
    .A2(_15552_),
    .ZN(_15604_));
 BUF_X2 _25319_ (.A(_15604_),
    .Z(_15605_));
 AOI22_X1 _25320_ (.A1(_15602_),
    .A2(_15603_),
    .B1(_15605_),
    .B2(_15584_),
    .ZN(_15606_));
 AND4_X1 _25321_ (.A1(_15561_),
    .A2(_15587_),
    .A3(_15599_),
    .A4(_15606_),
    .ZN(_15607_));
 AND2_X1 _25322_ (.A1(_15581_),
    .A2(_15571_),
    .ZN(_15608_));
 INV_X1 _25323_ (.A(_15608_),
    .ZN(_15609_));
 NOR2_X1 _25324_ (.A1(_11029_),
    .A2(_17148_),
    .ZN(_15610_));
 AND2_X2 _25325_ (.A1(_17149_),
    .A2(_17150_),
    .ZN(_15611_));
 AND2_X2 _25326_ (.A1(_15610_),
    .A2(_15611_),
    .ZN(_15612_));
 INV_X1 _25327_ (.A(_15612_),
    .ZN(_15613_));
 AND2_X2 _25328_ (.A1(_15600_),
    .A2(_15557_),
    .ZN(_15614_));
 INV_X1 _25329_ (.A(_15614_),
    .ZN(_15615_));
 AND2_X2 _25330_ (.A1(_15611_),
    .A2(_15563_),
    .ZN(_15616_));
 INV_X1 _25331_ (.A(_15616_),
    .ZN(_15617_));
 OAI22_X1 _25332_ (.A1(_15609_),
    .A2(_15613_),
    .B1(_15615_),
    .B2(_15617_),
    .ZN(_15618_));
 AND2_X1 _25333_ (.A1(_15596_),
    .A2(_15611_),
    .ZN(_15619_));
 BUF_X2 _25334_ (.A(_15619_),
    .Z(_15620_));
 BUF_X4 _25335_ (.A(_15620_),
    .Z(_15621_));
 BUF_X4 _25336_ (.A(_15547_),
    .Z(_15622_));
 BUF_X4 _25337_ (.A(_15622_),
    .Z(_15623_));
 BUF_X4 _25338_ (.A(_15600_),
    .Z(_15624_));
 OAI211_X2 _25339_ (.A(_15621_),
    .B(_15623_),
    .C1(_15624_),
    .C2(_15590_),
    .ZN(_15625_));
 BUF_X4 _25340_ (.A(_15548_),
    .Z(_15626_));
 NAND4_X1 _25341_ (.A1(_15596_),
    .A2(_15623_),
    .A3(_15626_),
    .A4(_15611_),
    .ZN(_15627_));
 NAND2_X1 _25342_ (.A1(_15625_),
    .A2(_15627_),
    .ZN(_15628_));
 AND2_X1 _25343_ (.A1(_15550_),
    .A2(_15611_),
    .ZN(_15629_));
 BUF_X2 _25344_ (.A(_15629_),
    .Z(_15630_));
 AND2_X1 _25345_ (.A1(_15573_),
    .A2(_15630_),
    .ZN(_15631_));
 AND2_X2 _25346_ (.A1(_15581_),
    .A2(_15557_),
    .ZN(_15632_));
 AND2_X1 _25347_ (.A1(_15632_),
    .A2(_15629_),
    .ZN(_15633_));
 NOR4_X1 _25348_ (.A1(_15618_),
    .A2(_15628_),
    .A3(_15631_),
    .A4(_15633_),
    .ZN(_15634_));
 BUF_X4 _25349_ (.A(_15612_),
    .Z(_15635_));
 BUF_X4 _25350_ (.A(_15557_),
    .Z(_15636_));
 AND2_X2 _25351_ (.A1(_15636_),
    .A2(_11003_),
    .ZN(_15637_));
 AND2_X1 _25352_ (.A1(_15635_),
    .A2(_15637_),
    .ZN(_15638_));
 BUF_X4 _25353_ (.A(_15579_),
    .Z(_15639_));
 BUF_X4 _25354_ (.A(_15639_),
    .Z(_15640_));
 AND2_X1 _25355_ (.A1(_15638_),
    .A2(_15640_),
    .ZN(_15641_));
 BUF_X2 _25356_ (.A(_15605_),
    .Z(_15642_));
 NOR2_X1 _25357_ (.A1(_15558_),
    .A2(_15590_),
    .ZN(_15643_));
 AND2_X1 _25358_ (.A1(_15642_),
    .A2(_15643_),
    .ZN(_15644_));
 INV_X1 _25359_ (.A(_15548_),
    .ZN(_15645_));
 NAND2_X1 _25360_ (.A1(_15645_),
    .A2(_15623_),
    .ZN(_15646_));
 INV_X1 _25361_ (.A(_15596_),
    .ZN(_15647_));
 BUF_X2 _25362_ (.A(_15552_),
    .Z(_15648_));
 INV_X1 _25363_ (.A(_15648_),
    .ZN(_15649_));
 NOR3_X1 _25364_ (.A1(_15646_),
    .A2(_15647_),
    .A3(_15649_),
    .ZN(_15650_));
 BUF_X2 _25365_ (.A(_15616_),
    .Z(_15651_));
 BUF_X4 _25366_ (.A(_15588_),
    .Z(_15652_));
 AND3_X1 _25367_ (.A1(_15651_),
    .A2(_15652_),
    .A3(_15624_),
    .ZN(_15653_));
 NOR4_X1 _25368_ (.A1(_15641_),
    .A2(_15644_),
    .A3(_15650_),
    .A4(_15653_),
    .ZN(_15654_));
 AND2_X1 _25369_ (.A1(_15589_),
    .A2(_15556_),
    .ZN(_15655_));
 BUF_X2 _25370_ (.A(_15655_),
    .Z(_15656_));
 AND2_X1 _25371_ (.A1(_15598_),
    .A2(_15656_),
    .ZN(_15657_));
 INV_X1 _25372_ (.A(_15657_),
    .ZN(_15658_));
 BUF_X4 _25373_ (.A(_15598_),
    .Z(_15659_));
 AND2_X1 _25374_ (.A1(_15659_),
    .A2(_15632_),
    .ZN(_15660_));
 INV_X1 _25375_ (.A(_15660_),
    .ZN(_15661_));
 AND2_X2 _25376_ (.A1(_15593_),
    .A2(_15551_),
    .ZN(_15662_));
 BUF_X2 _25377_ (.A(_15662_),
    .Z(_15663_));
 AND2_X1 _25378_ (.A1(_15548_),
    .A2(_15557_),
    .ZN(_15664_));
 BUF_X2 _25379_ (.A(_15664_),
    .Z(_15665_));
 NAND2_X1 _25380_ (.A1(_15663_),
    .A2(_15665_),
    .ZN(_15666_));
 AND2_X1 _25381_ (.A1(_15565_),
    .A2(_11003_),
    .ZN(_15667_));
 BUF_X2 _25382_ (.A(_15667_),
    .Z(_15668_));
 NAND3_X1 _25383_ (.A1(_15659_),
    .A2(_15640_),
    .A3(_15668_),
    .ZN(_15669_));
 AND4_X1 _25384_ (.A1(_15658_),
    .A2(_15661_),
    .A3(_15666_),
    .A4(_15669_),
    .ZN(_15670_));
 AND4_X1 _25385_ (.A1(_15607_),
    .A2(_15634_),
    .A3(_15654_),
    .A4(_15670_),
    .ZN(_15671_));
 AND2_X2 _25386_ (.A1(_15552_),
    .A2(_15563_),
    .ZN(_15672_));
 BUF_X4 _25387_ (.A(_15672_),
    .Z(_15673_));
 AND2_X1 _25388_ (.A1(_15595_),
    .A2(_15673_),
    .ZN(_15674_));
 INV_X1 _25389_ (.A(_15674_),
    .ZN(_15675_));
 NAND3_X1 _25390_ (.A1(_15637_),
    .A2(_11035_),
    .A3(_15648_),
    .ZN(_15676_));
 BUF_X4 _25391_ (.A(_15673_),
    .Z(_15677_));
 BUF_X4 _25392_ (.A(_15623_),
    .Z(_15678_));
 BUF_X2 _25393_ (.A(_15570_),
    .Z(_15679_));
 BUF_X4 _25394_ (.A(_15679_),
    .Z(_15680_));
 OAI211_X2 _25395_ (.A(_15677_),
    .B(_15581_),
    .C1(_15678_),
    .C2(_15680_),
    .ZN(_15681_));
 AND3_X1 _25396_ (.A1(_15675_),
    .A2(_15676_),
    .A3(_15681_),
    .ZN(_15682_));
 AND2_X2 _25397_ (.A1(_15557_),
    .A2(_10996_),
    .ZN(_15683_));
 NAND2_X1 _25398_ (.A1(_15663_),
    .A2(_15683_),
    .ZN(_15684_));
 AND2_X1 _25399_ (.A1(_15557_),
    .A2(_11010_),
    .ZN(_15685_));
 BUF_X4 _25400_ (.A(_15685_),
    .Z(_15686_));
 BUF_X4 _25401_ (.A(_15594_),
    .Z(_15687_));
 AND2_X1 _25402_ (.A1(_15565_),
    .A2(_11010_),
    .ZN(_15688_));
 BUF_X2 _25403_ (.A(_15688_),
    .Z(_15689_));
 AOI22_X1 _25404_ (.A1(_15686_),
    .A2(_15687_),
    .B1(_15689_),
    .B2(_15603_),
    .ZN(_15690_));
 AND2_X1 _25405_ (.A1(_15571_),
    .A2(_11010_),
    .ZN(_15691_));
 BUF_X2 _25406_ (.A(_15691_),
    .Z(_15692_));
 NAND2_X1 _25407_ (.A1(_15598_),
    .A2(_15692_),
    .ZN(_15693_));
 AND2_X2 _25408_ (.A1(_15610_),
    .A2(_15593_),
    .ZN(_15694_));
 BUF_X2 _25409_ (.A(_15694_),
    .Z(_15695_));
 NAND2_X1 _25410_ (.A1(_15695_),
    .A2(_15595_),
    .ZN(_15696_));
 AND4_X1 _25411_ (.A1(_15684_),
    .A2(_15690_),
    .A3(_15693_),
    .A4(_15696_),
    .ZN(_15697_));
 INV_X1 _25412_ (.A(_15589_),
    .ZN(_15698_));
 BUF_X2 _25413_ (.A(_15698_),
    .Z(_15699_));
 AND2_X1 _25414_ (.A1(_15567_),
    .A2(_15699_),
    .ZN(_15700_));
 AND2_X1 _25415_ (.A1(_15547_),
    .A2(_11003_),
    .ZN(_15701_));
 BUF_X2 _25416_ (.A(_15701_),
    .Z(_15702_));
 OAI21_X1 _25417_ (.A(_15677_),
    .B1(_15700_),
    .B2(_15702_),
    .ZN(_15703_));
 AND2_X1 _25418_ (.A1(_15622_),
    .A2(_15590_),
    .ZN(_15704_));
 BUF_X2 _25419_ (.A(_15704_),
    .Z(_15705_));
 OR2_X1 _25420_ (.A1(_15705_),
    .A2(_15549_),
    .ZN(_15706_));
 AND2_X1 _25421_ (.A1(_15610_),
    .A2(_15648_),
    .ZN(_15707_));
 BUF_X4 _25422_ (.A(_15707_),
    .Z(_15708_));
 BUF_X4 _25423_ (.A(_15708_),
    .Z(_15709_));
 NAND2_X1 _25424_ (.A1(_15706_),
    .A2(_15709_),
    .ZN(_15710_));
 BUF_X2 _25425_ (.A(_15608_),
    .Z(_15711_));
 OAI21_X1 _25426_ (.A(_15709_),
    .B1(_15602_),
    .B2(_15711_),
    .ZN(_15712_));
 AND3_X1 _25427_ (.A1(_15703_),
    .A2(_15710_),
    .A3(_15712_),
    .ZN(_15713_));
 AND2_X1 _25428_ (.A1(_15665_),
    .A2(_15677_),
    .ZN(_15714_));
 INV_X1 _25429_ (.A(_15714_),
    .ZN(_15715_));
 AND2_X1 _25430_ (.A1(_15605_),
    .A2(_15668_),
    .ZN(_15716_));
 NAND2_X1 _25431_ (.A1(_15699_),
    .A2(_15679_),
    .ZN(_15717_));
 NOR2_X1 _25432_ (.A1(_15717_),
    .A2(_15626_),
    .ZN(_15718_));
 AND2_X2 _25433_ (.A1(_15679_),
    .A2(_10996_),
    .ZN(_15719_));
 AOI221_X4 _25434_ (.A(_15716_),
    .B1(_15605_),
    .B2(_15718_),
    .C1(_15719_),
    .C2(_15663_),
    .ZN(_15720_));
 AND3_X1 _25435_ (.A1(_15713_),
    .A2(_15715_),
    .A3(_15720_),
    .ZN(_15721_));
 NAND4_X1 _25436_ (.A1(_15671_),
    .A2(_15682_),
    .A3(_15697_),
    .A4(_15721_),
    .ZN(_15722_));
 AND2_X1 _25437_ (.A1(_15622_),
    .A2(_10996_),
    .ZN(_15723_));
 OAI21_X1 _25438_ (.A(_15695_),
    .B1(_15723_),
    .B2(_15591_),
    .ZN(_15724_));
 AND2_X1 _25439_ (.A1(_15576_),
    .A2(_15591_),
    .ZN(_15725_));
 INV_X1 _25440_ (.A(_15725_),
    .ZN(_15726_));
 AND2_X2 _25441_ (.A1(_15581_),
    .A2(_15547_),
    .ZN(_15727_));
 OAI21_X1 _25442_ (.A(_15576_),
    .B1(_15727_),
    .B2(_15689_),
    .ZN(_15728_));
 AND2_X1 _25443_ (.A1(_15726_),
    .A2(_15728_),
    .ZN(_15729_));
 INV_X1 _25444_ (.A(_15729_),
    .ZN(_15730_));
 INV_X1 _25445_ (.A(_15570_),
    .ZN(_15731_));
 NOR2_X1 _25446_ (.A1(_15731_),
    .A2(_15600_),
    .ZN(_15732_));
 BUF_X4 _25447_ (.A(_15578_),
    .Z(_15733_));
 AND2_X1 _25448_ (.A1(_15732_),
    .A2(_15733_),
    .ZN(_15734_));
 NOR2_X1 _25449_ (.A1(_15730_),
    .A2(_15734_),
    .ZN(_15735_));
 INV_X1 _25450_ (.A(_15600_),
    .ZN(_15736_));
 AND3_X1 _25451_ (.A1(_15694_),
    .A2(_15636_),
    .A3(_15736_),
    .ZN(_15737_));
 OAI21_X1 _25452_ (.A(_15622_),
    .B1(_10996_),
    .B2(_11010_),
    .ZN(_15738_));
 INV_X1 _25453_ (.A(_15738_),
    .ZN(_15739_));
 AOI21_X1 _25454_ (.A(_15737_),
    .B1(_15659_),
    .B2(_15739_),
    .ZN(_15740_));
 BUF_X4 _25455_ (.A(_15564_),
    .Z(_15741_));
 AND2_X1 _25456_ (.A1(_15557_),
    .A2(_15639_),
    .ZN(_15742_));
 OAI21_X1 _25457_ (.A(_15741_),
    .B1(_15723_),
    .B2(_15742_),
    .ZN(_15743_));
 NAND2_X1 _25458_ (.A1(_15732_),
    .A2(_15564_),
    .ZN(_15744_));
 AND2_X1 _25459_ (.A1(_15743_),
    .A2(_15744_),
    .ZN(_15745_));
 AND4_X1 _25460_ (.A1(_15724_),
    .A2(_15735_),
    .A3(_15740_),
    .A4(_15745_),
    .ZN(_15746_));
 NAND3_X1 _25461_ (.A1(_15567_),
    .A2(_15663_),
    .A3(_15699_),
    .ZN(_15747_));
 NAND2_X1 _25462_ (.A1(_15705_),
    .A2(_15663_),
    .ZN(_15748_));
 AND2_X1 _25463_ (.A1(_15747_),
    .A2(_15748_),
    .ZN(_15749_));
 INV_X1 _25464_ (.A(_15700_),
    .ZN(_15750_));
 INV_X1 _25465_ (.A(_15622_),
    .ZN(_15751_));
 AOI21_X1 _25466_ (.A(_15613_),
    .B1(_15750_),
    .B2(_15751_),
    .ZN(_15752_));
 AND2_X1 _25467_ (.A1(_15723_),
    .A2(_15651_),
    .ZN(_15753_));
 CLKBUF_X2 _25468_ (.A(_15562_),
    .Z(_15754_));
 BUF_X2 _25469_ (.A(_15610_),
    .Z(_15755_));
 AND3_X1 _25470_ (.A1(_15668_),
    .A2(_15754_),
    .A3(_15755_),
    .ZN(_15756_));
 AND2_X1 _25471_ (.A1(_15689_),
    .A2(_15651_),
    .ZN(_15757_));
 OR3_X1 _25472_ (.A1(_15753_),
    .A2(_15756_),
    .A3(_15757_),
    .ZN(_15758_));
 AND2_X1 _25473_ (.A1(_15562_),
    .A2(_15610_),
    .ZN(_15759_));
 BUF_X2 _25474_ (.A(_15759_),
    .Z(_15760_));
 AND3_X1 _25475_ (.A1(_15760_),
    .A2(_15645_),
    .A3(_15643_),
    .ZN(_15761_));
 AND2_X1 _25476_ (.A1(_15692_),
    .A2(_15621_),
    .ZN(_15762_));
 NOR4_X1 _25477_ (.A1(_15752_),
    .A2(_15758_),
    .A3(_15761_),
    .A4(_15762_),
    .ZN(_15763_));
 AND2_X1 _25478_ (.A1(_15600_),
    .A2(_15588_),
    .ZN(_15764_));
 BUF_X2 _25479_ (.A(_15764_),
    .Z(_15765_));
 OAI21_X1 _25480_ (.A(_15594_),
    .B1(_15765_),
    .B2(_15689_),
    .ZN(_15766_));
 NAND4_X1 _25481_ (.A1(_15623_),
    .A2(_15593_),
    .A3(_10996_),
    .A4(_15563_),
    .ZN(_15767_));
 AND2_X1 _25482_ (.A1(_15766_),
    .A2(_15767_),
    .ZN(_15768_));
 INV_X1 _25483_ (.A(_15655_),
    .ZN(_15769_));
 INV_X1 _25484_ (.A(_15664_),
    .ZN(_15770_));
 NAND2_X1 _25485_ (.A1(_15769_),
    .A2(_15770_),
    .ZN(_15771_));
 AND2_X2 _25486_ (.A1(_15588_),
    .A2(_10996_),
    .ZN(_15772_));
 OAI21_X1 _25487_ (.A(_15621_),
    .B1(_15771_),
    .B2(_15772_),
    .ZN(_15773_));
 BUF_X4 _25488_ (.A(_15630_),
    .Z(_15774_));
 OAI21_X1 _25489_ (.A(_15774_),
    .B1(_15765_),
    .B2(_15678_),
    .ZN(_15775_));
 NAND2_X1 _25490_ (.A1(_15774_),
    .A2(_15637_),
    .ZN(_15776_));
 AND4_X1 _25491_ (.A1(_15768_),
    .A2(_15773_),
    .A3(_15775_),
    .A4(_15776_),
    .ZN(_15777_));
 NAND4_X1 _25492_ (.A1(_15746_),
    .A2(_15749_),
    .A3(_15763_),
    .A4(_15777_),
    .ZN(_15778_));
 NOR2_X1 _25493_ (.A1(_15722_),
    .A2(_15778_),
    .ZN(_15779_));
 XOR2_X1 _25494_ (.A(_15779_),
    .B(_01005_),
    .Z(_15780_));
 MUX2_X1 _25495_ (.A(_01216_),
    .B(_15780_),
    .S(_15298_),
    .Z(_01065_));
 AND2_X1 _25496_ (.A1(_15679_),
    .A2(_15639_),
    .ZN(_15781_));
 OAI21_X1 _25497_ (.A(_15708_),
    .B1(_15781_),
    .B2(_15686_),
    .ZN(_15782_));
 AND3_X1 _25498_ (.A1(_15672_),
    .A2(_15626_),
    .A3(_15571_),
    .ZN(_15783_));
 AND3_X1 _25499_ (.A1(_15672_),
    .A2(_15581_),
    .A3(_15571_),
    .ZN(_15784_));
 AND3_X1 _25500_ (.A1(_15672_),
    .A2(_15600_),
    .A3(_15571_),
    .ZN(_15785_));
 OR3_X1 _25501_ (.A1(_15783_),
    .A2(_15784_),
    .A3(_15785_),
    .ZN(_15786_));
 AOI21_X1 _25502_ (.A(_15786_),
    .B1(_15637_),
    .B2(_15673_),
    .ZN(_15787_));
 AND2_X1 _25503_ (.A1(_15688_),
    .A2(_15672_),
    .ZN(_15788_));
 NAND3_X1 _25504_ (.A1(_15672_),
    .A2(_15600_),
    .A3(_15622_),
    .ZN(_15789_));
 NAND3_X1 _25505_ (.A1(_15672_),
    .A2(_15590_),
    .A3(_15622_),
    .ZN(_15790_));
 NAND2_X1 _25506_ (.A1(_15789_),
    .A2(_15790_),
    .ZN(_15791_));
 AOI211_X4 _25507_ (.A(_15788_),
    .B(_15791_),
    .C1(_15667_),
    .C2(_15673_),
    .ZN(_15792_));
 OAI21_X1 _25508_ (.A(_15708_),
    .B1(_15765_),
    .B2(_15702_),
    .ZN(_15793_));
 AND4_X1 _25509_ (.A1(_15782_),
    .A2(_15787_),
    .A3(_15792_),
    .A4(_15793_),
    .ZN(_15794_));
 INV_X1 _25510_ (.A(_15717_),
    .ZN(_15795_));
 OAI21_X1 _25511_ (.A(_15642_),
    .B1(_15795_),
    .B2(_15582_),
    .ZN(_15796_));
 OAI21_X1 _25512_ (.A(_15603_),
    .B1(_15719_),
    .B2(_15559_),
    .ZN(_15797_));
 AND2_X1 _25513_ (.A1(_15689_),
    .A2(_15554_),
    .ZN(_15798_));
 INV_X1 _25514_ (.A(_15798_),
    .ZN(_15799_));
 NAND2_X1 _25515_ (.A1(_15705_),
    .A2(_15554_),
    .ZN(_15800_));
 NAND2_X1 _25516_ (.A1(_15764_),
    .A2(_15554_),
    .ZN(_15801_));
 OAI211_X2 _25517_ (.A(_15554_),
    .B(_15623_),
    .C1(_15626_),
    .C2(_15581_),
    .ZN(_15802_));
 AND4_X1 _25518_ (.A1(_15799_),
    .A2(_15800_),
    .A3(_15801_),
    .A4(_15802_),
    .ZN(_15803_));
 AND4_X1 _25519_ (.A1(_15794_),
    .A2(_15796_),
    .A3(_15797_),
    .A4(_15803_),
    .ZN(_15804_));
 AND2_X1 _25520_ (.A1(_15594_),
    .A2(_15622_),
    .ZN(_15805_));
 AND2_X1 _25521_ (.A1(_15594_),
    .A2(_15764_),
    .ZN(_15806_));
 AND2_X2 _25522_ (.A1(_15580_),
    .A2(_15588_),
    .ZN(_15807_));
 AOI211_X4 _25523_ (.A(_15805_),
    .B(_15806_),
    .C1(_15594_),
    .C2(_15807_),
    .ZN(_15808_));
 NAND2_X1 _25524_ (.A1(_15795_),
    .A2(_15687_),
    .ZN(_15809_));
 INV_X1 _25525_ (.A(_15683_),
    .ZN(_15810_));
 INV_X1 _25526_ (.A(_15687_),
    .ZN(_15811_));
 OAI211_X2 _25527_ (.A(_15808_),
    .B(_15809_),
    .C1(_15810_),
    .C2(_15811_),
    .ZN(_15812_));
 AND2_X2 _25528_ (.A1(_15547_),
    .A2(_11010_),
    .ZN(_15813_));
 AND2_X1 _25529_ (.A1(_15694_),
    .A2(_15813_),
    .ZN(_15814_));
 AND2_X1 _25530_ (.A1(_15571_),
    .A2(_15589_),
    .ZN(_15815_));
 BUF_X2 _25531_ (.A(_15815_),
    .Z(_15816_));
 NOR2_X1 _25532_ (.A1(_15816_),
    .A2(_15665_),
    .ZN(_15817_));
 INV_X1 _25533_ (.A(_15694_),
    .ZN(_15818_));
 NOR2_X1 _25534_ (.A1(_15817_),
    .A2(_15818_),
    .ZN(_15819_));
 NOR2_X1 _25535_ (.A1(_15591_),
    .A2(_15583_),
    .ZN(_15820_));
 NOR2_X1 _25536_ (.A1(_15820_),
    .A2(_15818_),
    .ZN(_15821_));
 AND2_X2 _25537_ (.A1(_15600_),
    .A2(_15547_),
    .ZN(_15822_));
 AND2_X1 _25538_ (.A1(_15822_),
    .A2(_15694_),
    .ZN(_15823_));
 OR4_X1 _25539_ (.A1(_15814_),
    .A2(_15819_),
    .A3(_15821_),
    .A4(_15823_),
    .ZN(_15824_));
 AND2_X1 _25540_ (.A1(_15662_),
    .A2(_15683_),
    .ZN(_15825_));
 INV_X1 _25541_ (.A(_15662_),
    .ZN(_15826_));
 INV_X1 _25542_ (.A(_15822_),
    .ZN(_15827_));
 INV_X1 _25543_ (.A(_15727_),
    .ZN(_15828_));
 AOI21_X1 _25544_ (.A(_15826_),
    .B1(_15827_),
    .B2(_15828_),
    .ZN(_15829_));
 AND4_X1 _25545_ (.A1(_15551_),
    .A2(_15679_),
    .A3(_15593_),
    .A4(_15626_),
    .ZN(_15830_));
 AND2_X1 _25546_ (.A1(_15567_),
    .A2(_15662_),
    .ZN(_15831_));
 OR4_X1 _25547_ (.A1(_15825_),
    .A2(_15829_),
    .A3(_15830_),
    .A4(_15831_),
    .ZN(_15832_));
 AND2_X1 _25548_ (.A1(_15597_),
    .A2(_15559_),
    .ZN(_15833_));
 INV_X1 _25549_ (.A(_15833_),
    .ZN(_15834_));
 OAI21_X1 _25550_ (.A(_15659_),
    .B1(_15765_),
    .B2(_15702_),
    .ZN(_15835_));
 INV_X1 _25551_ (.A(_15781_),
    .ZN(_15836_));
 INV_X1 _25552_ (.A(_15597_),
    .ZN(_15837_));
 OAI211_X2 _25553_ (.A(_15834_),
    .B(_15835_),
    .C1(_15836_),
    .C2(_15837_),
    .ZN(_15838_));
 NOR4_X1 _25554_ (.A1(_15812_),
    .A2(_15824_),
    .A3(_15832_),
    .A4(_15838_),
    .ZN(_15839_));
 OAI21_X1 _25555_ (.A(_15733_),
    .B1(_15765_),
    .B2(_15807_),
    .ZN(_15840_));
 OAI21_X1 _25556_ (.A(_15578_),
    .B1(_15602_),
    .B2(_15742_),
    .ZN(_15841_));
 NAND4_X1 _25557_ (.A1(_15754_),
    .A2(_15623_),
    .A3(_10997_),
    .A4(_15551_),
    .ZN(_15842_));
 AND3_X1 _25558_ (.A1(_15840_),
    .A2(_15841_),
    .A3(_15842_),
    .ZN(_15843_));
 AND2_X1 _25559_ (.A1(_15739_),
    .A2(_15576_),
    .ZN(_15844_));
 AND2_X1 _25560_ (.A1(_15576_),
    .A2(_15637_),
    .ZN(_15845_));
 AND2_X1 _25561_ (.A1(_15575_),
    .A2(_15632_),
    .ZN(_15846_));
 AND3_X1 _25562_ (.A1(_15608_),
    .A2(_15754_),
    .A3(_15596_),
    .ZN(_15847_));
 NOR4_X1 _25563_ (.A1(_15844_),
    .A2(_15845_),
    .A3(_15846_),
    .A4(_15847_),
    .ZN(_15848_));
 OAI21_X1 _25564_ (.A(_15564_),
    .B1(_15822_),
    .B2(_15727_),
    .ZN(_15849_));
 NAND4_X1 _25565_ (.A1(_15754_),
    .A2(_15624_),
    .A3(_15636_),
    .A4(_15563_),
    .ZN(_15850_));
 NAND2_X1 _25566_ (.A1(_15564_),
    .A2(_15591_),
    .ZN(_15851_));
 AND4_X1 _25567_ (.A1(_15744_),
    .A2(_15849_),
    .A3(_15850_),
    .A4(_15851_),
    .ZN(_15852_));
 NAND2_X1 _25568_ (.A1(_15760_),
    .A2(_15692_),
    .ZN(_15853_));
 INV_X1 _25569_ (.A(_15759_),
    .ZN(_15854_));
 OAI21_X1 _25570_ (.A(_15853_),
    .B1(_15854_),
    .B2(_15615_),
    .ZN(_15855_));
 AND2_X1 _25571_ (.A1(_15760_),
    .A2(_15652_),
    .ZN(_15856_));
 AND2_X1 _25572_ (.A1(_15759_),
    .A2(_15813_),
    .ZN(_15857_));
 NOR3_X1 _25573_ (.A1(_15855_),
    .A2(_15856_),
    .A3(_15857_),
    .ZN(_15858_));
 AND4_X1 _25574_ (.A1(_15843_),
    .A2(_15848_),
    .A3(_15852_),
    .A4(_15858_),
    .ZN(_15859_));
 AND2_X1 _25575_ (.A1(_15584_),
    .A2(_15616_),
    .ZN(_15860_));
 AND2_X1 _25576_ (.A1(_15668_),
    .A2(_15616_),
    .ZN(_15861_));
 OR2_X1 _25577_ (.A1(_15860_),
    .A2(_15861_),
    .ZN(_15862_));
 AND2_X1 _25578_ (.A1(_15705_),
    .A2(_15651_),
    .ZN(_15863_));
 AOI21_X1 _25579_ (.A(_15617_),
    .B1(_15769_),
    .B2(_15770_),
    .ZN(_15864_));
 AND4_X1 _25580_ (.A1(_10996_),
    .A2(_15679_),
    .A3(_15563_),
    .A4(_15611_),
    .ZN(_15865_));
 NOR4_X1 _25581_ (.A1(_15862_),
    .A2(_15863_),
    .A3(_15864_),
    .A4(_15865_),
    .ZN(_15866_));
 INV_X1 _25582_ (.A(_15595_),
    .ZN(_15867_));
 AOI21_X1 _25583_ (.A(_15613_),
    .B1(_15609_),
    .B2(_15867_),
    .ZN(_15868_));
 NAND3_X1 _25584_ (.A1(_15583_),
    .A2(_15755_),
    .A3(_15611_),
    .ZN(_15869_));
 NAND2_X1 _25585_ (.A1(_15612_),
    .A2(_15667_),
    .ZN(_15870_));
 OAI221_X1 _25586_ (.A(_15869_),
    .B1(_15827_),
    .B2(_15613_),
    .C1(_15639_),
    .C2(_15870_),
    .ZN(_15871_));
 AOI211_X4 _25587_ (.A(_15868_),
    .B(_15871_),
    .C1(_15683_),
    .C2(_15612_),
    .ZN(_15872_));
 AND2_X1 _25588_ (.A1(_15619_),
    .A2(_15583_),
    .ZN(_15873_));
 AND3_X1 _25589_ (.A1(_15591_),
    .A2(_15596_),
    .A3(_15611_),
    .ZN(_15874_));
 OR2_X1 _25590_ (.A1(_15873_),
    .A2(_15874_),
    .ZN(_15875_));
 AND2_X1 _25591_ (.A1(_15822_),
    .A2(_15620_),
    .ZN(_15876_));
 AND2_X1 _25592_ (.A1(_15813_),
    .A2(_15620_),
    .ZN(_15877_));
 AND2_X1 _25593_ (.A1(_15602_),
    .A2(_15620_),
    .ZN(_15878_));
 NOR4_X1 _25594_ (.A1(_15875_),
    .A2(_15876_),
    .A3(_15877_),
    .A4(_15878_),
    .ZN(_15879_));
 AND2_X1 _25595_ (.A1(_15704_),
    .A2(_15629_),
    .ZN(_15880_));
 INV_X1 _25596_ (.A(_15629_),
    .ZN(_15881_));
 AOI211_X4 _25597_ (.A(_15731_),
    .B(_15881_),
    .C1(_10996_),
    .C2(_11003_),
    .ZN(_15882_));
 AOI211_X4 _25598_ (.A(_15880_),
    .B(_15882_),
    .C1(_15668_),
    .C2(_15630_),
    .ZN(_15883_));
 AND4_X1 _25599_ (.A1(_15866_),
    .A2(_15872_),
    .A3(_15879_),
    .A4(_15883_),
    .ZN(_15884_));
 NAND4_X1 _25600_ (.A1(_15804_),
    .A2(_15839_),
    .A3(_15859_),
    .A4(_15884_),
    .ZN(_15885_));
 NOR2_X1 _25601_ (.A1(_15885_),
    .A2(_15714_),
    .ZN(_15886_));
 INV_X1 _25602_ (.A(_01006_),
    .ZN(_15887_));
 XNOR2_X1 _25603_ (.A(_15886_),
    .B(_15887_),
    .ZN(_15888_));
 MUX2_X1 _25604_ (.A(_01217_),
    .B(_15888_),
    .S(_15298_),
    .Z(_01066_));
 AND2_X1 _25605_ (.A1(_15760_),
    .A2(_15689_),
    .ZN(_15889_));
 AND2_X1 _25606_ (.A1(_15760_),
    .A2(_15637_),
    .ZN(_15890_));
 AND3_X1 _25607_ (.A1(_15705_),
    .A2(_15754_),
    .A3(_15755_),
    .ZN(_15891_));
 NOR4_X1 _25608_ (.A1(_15889_),
    .A2(_15890_),
    .A3(_15857_),
    .A4(_15891_),
    .ZN(_15892_));
 OAI21_X1 _25609_ (.A(_15741_),
    .B1(_15689_),
    .B2(_15678_),
    .ZN(_15893_));
 OAI211_X2 _25610_ (.A(_15741_),
    .B(_15546_),
    .C1(_17145_),
    .C2(_15736_),
    .ZN(_15894_));
 AND3_X1 _25611_ (.A1(_15892_),
    .A2(_15893_),
    .A3(_15894_),
    .ZN(_15895_));
 OAI21_X1 _25612_ (.A(_15578_),
    .B1(_15665_),
    .B2(_15637_),
    .ZN(_15896_));
 INV_X1 _25613_ (.A(_15575_),
    .ZN(_15897_));
 AOI21_X1 _25614_ (.A(_15897_),
    .B1(_15750_),
    .B2(_15827_),
    .ZN(_15898_));
 AOI211_X4 _25615_ (.A(_15847_),
    .B(_15898_),
    .C1(_15595_),
    .C2(_15576_),
    .ZN(_15899_));
 OAI21_X1 _25616_ (.A(_15733_),
    .B1(_15602_),
    .B2(_15692_),
    .ZN(_15900_));
 AND2_X1 _25617_ (.A1(_15578_),
    .A2(_15764_),
    .ZN(_15901_));
 INV_X1 _25618_ (.A(_15578_),
    .ZN(_15902_));
 INV_X1 _25619_ (.A(_15813_),
    .ZN(_15903_));
 AOI21_X1 _25620_ (.A(_15902_),
    .B1(_15827_),
    .B2(_15903_),
    .ZN(_15904_));
 AOI211_X4 _25621_ (.A(_15901_),
    .B(_15904_),
    .C1(_15733_),
    .C2(_15584_),
    .ZN(_15905_));
 AND4_X1 _25622_ (.A1(_15896_),
    .A2(_15899_),
    .A3(_15900_),
    .A4(_15905_),
    .ZN(_15906_));
 INV_X1 _25623_ (.A(_15638_),
    .ZN(_15907_));
 NAND2_X1 _25624_ (.A1(_15632_),
    .A2(_15635_),
    .ZN(_15908_));
 OAI211_X2 _25625_ (.A(_15907_),
    .B(_15908_),
    .C1(_15867_),
    .C2(_15613_),
    .ZN(_15909_));
 AOI21_X1 _25626_ (.A(_15613_),
    .B1(_15827_),
    .B2(_15828_),
    .ZN(_15910_));
 NAND2_X1 _25627_ (.A1(_15870_),
    .A2(_15869_),
    .ZN(_15911_));
 OR2_X1 _25628_ (.A1(_15910_),
    .A2(_15911_),
    .ZN(_15912_));
 AOI21_X1 _25629_ (.A(_15617_),
    .B1(_15615_),
    .B2(_15769_),
    .ZN(_15913_));
 AND3_X1 _25630_ (.A1(_15679_),
    .A2(_15563_),
    .A3(_15611_),
    .ZN(_15914_));
 OR2_X1 _25631_ (.A1(_15913_),
    .A2(_15914_),
    .ZN(_15915_));
 AND2_X1 _25632_ (.A1(_15807_),
    .A2(_15651_),
    .ZN(_15916_));
 INV_X1 _25633_ (.A(_15916_),
    .ZN(_15917_));
 OAI211_X2 _25634_ (.A(_15651_),
    .B(_15623_),
    .C1(_10997_),
    .C2(_11004_),
    .ZN(_15918_));
 NAND2_X1 _25635_ (.A1(_15917_),
    .A2(_15918_),
    .ZN(_15919_));
 NOR4_X1 _25636_ (.A1(_15909_),
    .A2(_15912_),
    .A3(_15915_),
    .A4(_15919_),
    .ZN(_15920_));
 NAND2_X1 _25637_ (.A1(_15691_),
    .A2(_15630_),
    .ZN(_15921_));
 INV_X1 _25638_ (.A(_15620_),
    .ZN(_15922_));
 AOI21_X1 _25639_ (.A(_15922_),
    .B1(_15827_),
    .B2(_15828_),
    .ZN(_15923_));
 AND2_X1 _25640_ (.A1(_15619_),
    .A2(_15772_),
    .ZN(_15924_));
 AND2_X1 _25641_ (.A1(_15595_),
    .A2(_15620_),
    .ZN(_15925_));
 NOR4_X1 _25642_ (.A1(_15923_),
    .A2(_15924_),
    .A3(_15925_),
    .A4(_15873_),
    .ZN(_15926_));
 OAI21_X1 _25643_ (.A(_15774_),
    .B1(_15656_),
    .B2(_15665_),
    .ZN(_15927_));
 OAI21_X1 _25644_ (.A(_15774_),
    .B1(_15702_),
    .B2(_15772_),
    .ZN(_15928_));
 AND4_X1 _25645_ (.A1(_15921_),
    .A2(_15926_),
    .A3(_15927_),
    .A4(_15928_),
    .ZN(_15929_));
 AND4_X1 _25646_ (.A1(_15895_),
    .A2(_15906_),
    .A3(_15920_),
    .A4(_15929_),
    .ZN(_15930_));
 AND2_X1 _25647_ (.A1(_15708_),
    .A2(_15656_),
    .ZN(_15931_));
 INV_X1 _25648_ (.A(_15931_),
    .ZN(_15932_));
 NAND2_X1 _25649_ (.A1(_15602_),
    .A2(_15709_),
    .ZN(_15933_));
 NAND3_X1 _25650_ (.A1(_15689_),
    .A2(_15648_),
    .A3(_15755_),
    .ZN(_15934_));
 OAI211_X2 _25651_ (.A(_15709_),
    .B(_15678_),
    .C1(_10997_),
    .C2(_11011_),
    .ZN(_15935_));
 NAND4_X1 _25652_ (.A1(_15932_),
    .A2(_15933_),
    .A3(_15934_),
    .A4(_15935_),
    .ZN(_15936_));
 NOR2_X1 _25653_ (.A1(_15566_),
    .A2(_15600_),
    .ZN(_15937_));
 NAND2_X1 _25654_ (.A1(_15937_),
    .A2(_15677_),
    .ZN(_15938_));
 NAND2_X1 _25655_ (.A1(_15938_),
    .A2(_15789_),
    .ZN(_15939_));
 AND3_X1 _25656_ (.A1(_15559_),
    .A2(_15699_),
    .A3(_15677_),
    .ZN(_15940_));
 NOR4_X1 _25657_ (.A1(_15936_),
    .A2(_15674_),
    .A3(_15939_),
    .A4(_15940_),
    .ZN(_15941_));
 OAI21_X1 _25658_ (.A(_15659_),
    .B1(_15706_),
    .B2(_15700_),
    .ZN(_15942_));
 AND2_X1 _25659_ (.A1(_15662_),
    .A2(_15656_),
    .ZN(_15943_));
 INV_X1 _25660_ (.A(_15807_),
    .ZN(_15944_));
 AOI21_X1 _25661_ (.A(_15826_),
    .B1(_15903_),
    .B2(_15944_),
    .ZN(_15945_));
 AOI211_X4 _25662_ (.A(_15943_),
    .B(_15945_),
    .C1(_15719_),
    .C2(_15663_),
    .ZN(_15946_));
 OAI21_X1 _25663_ (.A(_15687_),
    .B1(_15711_),
    .B2(_15614_),
    .ZN(_15947_));
 OAI21_X1 _25664_ (.A(_15687_),
    .B1(_15822_),
    .B2(_15668_),
    .ZN(_15948_));
 OAI21_X1 _25665_ (.A(_15695_),
    .B1(_15711_),
    .B2(_15656_),
    .ZN(_15949_));
 OAI21_X1 _25666_ (.A(_15695_),
    .B1(_15822_),
    .B2(_15772_),
    .ZN(_15950_));
 AND4_X1 _25667_ (.A1(_15947_),
    .A2(_15948_),
    .A3(_15949_),
    .A4(_15950_),
    .ZN(_15951_));
 AND2_X1 _25668_ (.A1(_15659_),
    .A2(_15816_),
    .ZN(_15952_));
 AND2_X1 _25669_ (.A1(_15711_),
    .A2(_15598_),
    .ZN(_15953_));
 NOR3_X1 _25670_ (.A1(_15952_),
    .A2(_15953_),
    .A3(_15660_),
    .ZN(_15954_));
 AND4_X1 _25671_ (.A1(_15942_),
    .A2(_15946_),
    .A3(_15951_),
    .A4(_15954_),
    .ZN(_15955_));
 NAND4_X1 _25672_ (.A1(_15624_),
    .A2(_15596_),
    .A3(_15678_),
    .A4(_15648_),
    .ZN(_15956_));
 NAND4_X1 _25673_ (.A1(_15596_),
    .A2(_15652_),
    .A3(_15590_),
    .A4(_15648_),
    .ZN(_15957_));
 INV_X1 _25674_ (.A(_15604_),
    .ZN(_15958_));
 OAI211_X2 _25675_ (.A(_15956_),
    .B(_15957_),
    .C1(_15958_),
    .C2(_15903_),
    .ZN(_15959_));
 NAND2_X1 _25676_ (.A1(_15736_),
    .A2(_15557_),
    .ZN(_15960_));
 NOR2_X1 _25677_ (.A1(_15958_),
    .A2(_15960_),
    .ZN(_15961_));
 AND2_X1 _25678_ (.A1(_15642_),
    .A2(_15692_),
    .ZN(_15962_));
 AND2_X1 _25679_ (.A1(_15605_),
    .A2(_15595_),
    .ZN(_15963_));
 NOR4_X1 _25680_ (.A1(_15959_),
    .A2(_15961_),
    .A3(_15962_),
    .A4(_15963_),
    .ZN(_15964_));
 OAI21_X1 _25681_ (.A(_15603_),
    .B1(_15718_),
    .B2(_15686_),
    .ZN(_15965_));
 OAI21_X1 _25682_ (.A(_15603_),
    .B1(_15549_),
    .B2(_15772_),
    .ZN(_15966_));
 AND2_X1 _25683_ (.A1(_15965_),
    .A2(_15966_),
    .ZN(_15967_));
 AND4_X1 _25684_ (.A1(_15941_),
    .A2(_15955_),
    .A3(_15964_),
    .A4(_15967_),
    .ZN(_15968_));
 AND2_X2 _25685_ (.A1(_15930_),
    .A2(_15968_),
    .ZN(_15969_));
 XOR2_X1 _25686_ (.A(_15969_),
    .B(_01007_),
    .Z(_15970_));
 MUX2_X1 _25687_ (.A(_01218_),
    .B(_15970_),
    .S(_15298_),
    .Z(_01067_));
 OAI21_X1 _25688_ (.A(_15677_),
    .B1(_15718_),
    .B2(_15683_),
    .ZN(_15971_));
 AND2_X1 _25689_ (.A1(_15765_),
    .A2(_15673_),
    .ZN(_15972_));
 AOI221_X4 _25690_ (.A(_15972_),
    .B1(_15705_),
    .B2(_15677_),
    .C1(_15640_),
    .C2(_15788_),
    .ZN(_15973_));
 NAND2_X1 _25691_ (.A1(_15614_),
    .A2(_15708_),
    .ZN(_15974_));
 NAND2_X1 _25692_ (.A1(_15709_),
    .A2(_15692_),
    .ZN(_15975_));
 NAND4_X1 _25693_ (.A1(_15755_),
    .A2(_15626_),
    .A3(_15636_),
    .A4(_15648_),
    .ZN(_15976_));
 AND4_X1 _25694_ (.A1(_15974_),
    .A2(_15932_),
    .A3(_15975_),
    .A4(_15976_),
    .ZN(_15977_));
 OAI21_X1 _25695_ (.A(_15709_),
    .B1(_15706_),
    .B2(_15584_),
    .ZN(_15978_));
 AND4_X1 _25696_ (.A1(_15971_),
    .A2(_15973_),
    .A3(_15977_),
    .A4(_15978_),
    .ZN(_15979_));
 AOI211_X4 _25697_ (.A(_15566_),
    .B(_15837_),
    .C1(_15639_),
    .C2(_11011_),
    .ZN(_15980_));
 AND2_X1 _25698_ (.A1(_15598_),
    .A2(_15723_),
    .ZN(_15981_));
 OR4_X1 _25699_ (.A1(_15833_),
    .A2(_15980_),
    .A3(_15953_),
    .A4(_15981_),
    .ZN(_15982_));
 AND4_X1 _25700_ (.A1(_15645_),
    .A2(_15663_),
    .A3(_15699_),
    .A4(_15680_),
    .ZN(_15983_));
 AND2_X1 _25701_ (.A1(_15547_),
    .A2(_15639_),
    .ZN(_15984_));
 INV_X1 _25702_ (.A(_15984_),
    .ZN(_15985_));
 AOI21_X1 _25703_ (.A(_15826_),
    .B1(_15985_),
    .B2(_15944_),
    .ZN(_15986_));
 NOR4_X1 _25704_ (.A1(_15982_),
    .A2(_15943_),
    .A3(_15983_),
    .A4(_15986_),
    .ZN(_15987_));
 OAI21_X1 _25705_ (.A(_15603_),
    .B1(_15573_),
    .B2(_15816_),
    .ZN(_15988_));
 OAI21_X1 _25706_ (.A(_15642_),
    .B1(_15632_),
    .B2(_15719_),
    .ZN(_15989_));
 NAND2_X1 _25707_ (.A1(_15584_),
    .A2(_15603_),
    .ZN(_15990_));
 NAND2_X1 _25708_ (.A1(_15807_),
    .A2(_15642_),
    .ZN(_15991_));
 AND4_X1 _25709_ (.A1(_15988_),
    .A2(_15989_),
    .A3(_15990_),
    .A4(_15991_),
    .ZN(_15992_));
 INV_X1 _25710_ (.A(_15719_),
    .ZN(_15993_));
 AOI21_X1 _25711_ (.A(_15818_),
    .B1(_15769_),
    .B2(_15993_),
    .ZN(_15994_));
 AND2_X1 _25712_ (.A1(_15695_),
    .A2(_15702_),
    .ZN(_15995_));
 AND2_X1 _25713_ (.A1(_15694_),
    .A2(_15588_),
    .ZN(_15996_));
 NOR4_X1 _25714_ (.A1(_15994_),
    .A2(_15814_),
    .A3(_15995_),
    .A4(_15996_),
    .ZN(_15997_));
 OAI211_X2 _25715_ (.A(_15687_),
    .B(_15636_),
    .C1(_15640_),
    .C2(_11004_),
    .ZN(_15998_));
 AND2_X1 _25716_ (.A1(_15588_),
    .A2(_15639_),
    .ZN(_15999_));
 OAI21_X1 _25717_ (.A(_15687_),
    .B1(_15727_),
    .B2(_15999_),
    .ZN(_16000_));
 AND4_X1 _25718_ (.A1(_15809_),
    .A2(_15997_),
    .A3(_15998_),
    .A4(_16000_),
    .ZN(_16001_));
 AND4_X1 _25719_ (.A1(_15979_),
    .A2(_15987_),
    .A3(_15992_),
    .A4(_16001_),
    .ZN(_16002_));
 AND4_X1 _25720_ (.A1(_11004_),
    .A2(_15754_),
    .A3(_15551_),
    .A4(_15588_),
    .ZN(_16003_));
 AND2_X1 _25721_ (.A1(_15733_),
    .A2(_15807_),
    .ZN(_16004_));
 AOI211_X4 _25722_ (.A(_16003_),
    .B(_16004_),
    .C1(_15733_),
    .C2(_15706_),
    .ZN(_16005_));
 INV_X1 _25723_ (.A(_15591_),
    .ZN(_16006_));
 AOI21_X1 _25724_ (.A(_15897_),
    .B1(_15827_),
    .B2(_16006_),
    .ZN(_16007_));
 AND2_X1 _25725_ (.A1(_15576_),
    .A2(_15572_),
    .ZN(_16008_));
 AND2_X1 _25726_ (.A1(_15575_),
    .A2(_15816_),
    .ZN(_16009_));
 NOR4_X1 _25727_ (.A1(_16007_),
    .A2(_16008_),
    .A3(_15845_),
    .A4(_16009_),
    .ZN(_16010_));
 NAND4_X1 _25728_ (.A1(_15754_),
    .A2(_10997_),
    .A3(_15551_),
    .A4(_15636_),
    .ZN(_16011_));
 OAI211_X2 _25729_ (.A(_15733_),
    .B(_15680_),
    .C1(_15640_),
    .C2(_11004_),
    .ZN(_16012_));
 NAND4_X1 _25730_ (.A1(_16005_),
    .A2(_16010_),
    .A3(_16011_),
    .A4(_16012_),
    .ZN(_16013_));
 AND2_X1 _25731_ (.A1(_15813_),
    .A2(_15616_),
    .ZN(_16014_));
 OR2_X1 _25732_ (.A1(_15863_),
    .A2(_16014_),
    .ZN(_16015_));
 NAND3_X1 _25733_ (.A1(_15651_),
    .A2(_15626_),
    .A3(_15680_),
    .ZN(_16016_));
 NAND2_X1 _25734_ (.A1(_15651_),
    .A2(_15686_),
    .ZN(_16017_));
 OAI211_X2 _25735_ (.A(_16016_),
    .B(_16017_),
    .C1(_15769_),
    .C2(_15617_),
    .ZN(_16018_));
 NOR4_X1 _25736_ (.A1(_16015_),
    .A2(_16018_),
    .A3(_15757_),
    .A4(_15861_),
    .ZN(_16019_));
 AND2_X1 _25737_ (.A1(_15705_),
    .A2(_15612_),
    .ZN(_16020_));
 INV_X1 _25738_ (.A(_16020_),
    .ZN(_16021_));
 OAI21_X1 _25739_ (.A(_15635_),
    .B1(_15573_),
    .B2(_15816_),
    .ZN(_16022_));
 AND4_X1 _25740_ (.A1(_16021_),
    .A2(_15870_),
    .A3(_15908_),
    .A4(_16022_),
    .ZN(_16023_));
 OAI211_X2 _25741_ (.A(_15621_),
    .B(_15636_),
    .C1(_15581_),
    .C2(_15624_),
    .ZN(_16024_));
 OAI211_X2 _25742_ (.A(_15621_),
    .B(_15680_),
    .C1(_15640_),
    .C2(_11011_),
    .ZN(_16025_));
 OAI211_X2 _25743_ (.A(_15621_),
    .B(_15623_),
    .C1(_10997_),
    .C2(_11011_),
    .ZN(_16026_));
 OAI21_X1 _25744_ (.A(_15621_),
    .B1(_15584_),
    .B2(_15668_),
    .ZN(_16027_));
 AND4_X1 _25745_ (.A1(_16024_),
    .A2(_16025_),
    .A3(_16026_),
    .A4(_16027_),
    .ZN(_16028_));
 NAND3_X1 _25746_ (.A1(_15774_),
    .A2(_15652_),
    .A3(_15624_),
    .ZN(_16029_));
 OAI211_X2 _25747_ (.A(_15774_),
    .B(_15680_),
    .C1(_15626_),
    .C2(_15590_),
    .ZN(_16030_));
 OAI211_X2 _25748_ (.A(_15774_),
    .B(_15623_),
    .C1(_11004_),
    .C2(_15581_),
    .ZN(_16031_));
 OAI21_X1 _25749_ (.A(_15774_),
    .B1(_15665_),
    .B2(_15637_),
    .ZN(_16032_));
 AND4_X1 _25750_ (.A1(_16029_),
    .A2(_16030_),
    .A3(_16031_),
    .A4(_16032_),
    .ZN(_16033_));
 NAND4_X1 _25751_ (.A1(_16019_),
    .A2(_16023_),
    .A3(_16028_),
    .A4(_16033_),
    .ZN(_16034_));
 AND2_X1 _25752_ (.A1(_15741_),
    .A2(_15573_),
    .ZN(_16035_));
 INV_X1 _25753_ (.A(_15564_),
    .ZN(_16036_));
 NOR2_X1 _25754_ (.A1(_16036_),
    .A2(_15960_),
    .ZN(_16037_));
 AND3_X1 _25755_ (.A1(_15741_),
    .A2(_15699_),
    .A3(_15567_),
    .ZN(_16038_));
 AND2_X1 _25756_ (.A1(_15741_),
    .A2(_15702_),
    .ZN(_16039_));
 OR4_X1 _25757_ (.A1(_16035_),
    .A2(_16037_),
    .A3(_16038_),
    .A4(_16039_),
    .ZN(_16040_));
 NOR2_X1 _25758_ (.A1(_15822_),
    .A2(_15727_),
    .ZN(_16041_));
 NOR2_X1 _25759_ (.A1(_16041_),
    .A2(_15854_),
    .ZN(_16042_));
 AND3_X1 _25760_ (.A1(_15719_),
    .A2(_15754_),
    .A3(_15755_),
    .ZN(_16043_));
 OR4_X1 _25761_ (.A1(_15856_),
    .A2(_16042_),
    .A3(_15890_),
    .A4(_16043_),
    .ZN(_16044_));
 NOR4_X1 _25762_ (.A1(_16013_),
    .A2(_16034_),
    .A3(_16040_),
    .A4(_16044_),
    .ZN(_16045_));
 AND3_X1 _25763_ (.A1(_16002_),
    .A2(_01008_),
    .A3(_16045_),
    .ZN(_16046_));
 AOI21_X1 _25764_ (.A(_01008_),
    .B1(_16002_),
    .B2(_16045_),
    .ZN(_16047_));
 NOR2_X1 _25765_ (.A1(_16046_),
    .A2(_16047_),
    .ZN(_16048_));
 MUX2_X1 _25766_ (.A(_01219_),
    .B(_16048_),
    .S(_15298_),
    .Z(_01068_));
 OAI21_X1 _25767_ (.A(_15642_),
    .B1(_15705_),
    .B2(_15549_),
    .ZN(_16049_));
 AND2_X1 _25768_ (.A1(_15727_),
    .A2(_15554_),
    .ZN(_16050_));
 INV_X1 _25769_ (.A(_15554_),
    .ZN(_16051_));
 OAI21_X1 _25770_ (.A(_15801_),
    .B1(_16006_),
    .B2(_16051_),
    .ZN(_16052_));
 AOI211_X4 _25771_ (.A(_16050_),
    .B(_16052_),
    .C1(_15603_),
    .C2(_15732_),
    .ZN(_16053_));
 OAI21_X1 _25772_ (.A(_15642_),
    .B1(_15795_),
    .B2(_15643_),
    .ZN(_16054_));
 OAI21_X1 _25773_ (.A(_15642_),
    .B1(_15689_),
    .B2(_15668_),
    .ZN(_16055_));
 AND4_X1 _25774_ (.A1(_16049_),
    .A2(_16053_),
    .A3(_16054_),
    .A4(_16055_),
    .ZN(_16056_));
 NAND3_X1 _25775_ (.A1(_15677_),
    .A2(_15626_),
    .A3(_15678_),
    .ZN(_16057_));
 AND2_X1 _25776_ (.A1(_15727_),
    .A2(_15707_),
    .ZN(_16058_));
 INV_X1 _25777_ (.A(_16058_),
    .ZN(_16059_));
 OAI211_X2 _25778_ (.A(_15708_),
    .B(_15680_),
    .C1(_10997_),
    .C2(_11011_),
    .ZN(_16060_));
 OAI21_X1 _25779_ (.A(_15709_),
    .B1(_15765_),
    .B2(_15584_),
    .ZN(_16061_));
 AND4_X1 _25780_ (.A1(_15932_),
    .A2(_16059_),
    .A3(_16060_),
    .A4(_16061_),
    .ZN(_16062_));
 OAI21_X1 _25781_ (.A(_15677_),
    .B1(_15573_),
    .B2(_15559_),
    .ZN(_16063_));
 AND4_X1 _25782_ (.A1(_16057_),
    .A2(_16062_),
    .A3(_15938_),
    .A4(_16063_),
    .ZN(_16064_));
 NAND2_X1 _25783_ (.A1(_15711_),
    .A2(_15695_),
    .ZN(_16065_));
 INV_X1 _25784_ (.A(_15685_),
    .ZN(_16066_));
 OAI211_X2 _25785_ (.A(_16065_),
    .B(_15696_),
    .C1(_16066_),
    .C2(_15818_),
    .ZN(_16067_));
 AOI21_X1 _25786_ (.A(_15811_),
    .B1(_15769_),
    .B2(_15836_),
    .ZN(_16068_));
 NAND2_X1 _25787_ (.A1(_15695_),
    .A2(_15765_),
    .ZN(_16069_));
 INV_X1 _25788_ (.A(_15701_),
    .ZN(_16070_));
 OAI21_X1 _25789_ (.A(_16069_),
    .B1(_15818_),
    .B2(_16070_),
    .ZN(_16071_));
 NOR4_X1 _25790_ (.A1(_16067_),
    .A2(_16068_),
    .A3(_16071_),
    .A4(_15805_),
    .ZN(_16072_));
 INV_X1 _25791_ (.A(_15981_),
    .ZN(_16073_));
 NAND2_X1 _25792_ (.A1(_15602_),
    .A2(_15598_),
    .ZN(_16074_));
 OAI21_X1 _25793_ (.A(_15659_),
    .B1(_15656_),
    .B2(_15665_),
    .ZN(_16075_));
 OAI211_X2 _25794_ (.A(_15659_),
    .B(_15652_),
    .C1(_15640_),
    .C2(_11011_),
    .ZN(_16076_));
 NAND4_X1 _25795_ (.A1(_16073_),
    .A2(_16074_),
    .A3(_16075_),
    .A4(_16076_),
    .ZN(_16077_));
 AND2_X1 _25796_ (.A1(_15813_),
    .A2(_15662_),
    .ZN(_16078_));
 AND2_X1 _25797_ (.A1(_15822_),
    .A2(_15662_),
    .ZN(_16079_));
 OR2_X1 _25798_ (.A1(_16078_),
    .A2(_16079_),
    .ZN(_16080_));
 AND2_X1 _25799_ (.A1(_15663_),
    .A2(_15652_),
    .ZN(_16081_));
 NAND2_X1 _25800_ (.A1(_15692_),
    .A2(_15663_),
    .ZN(_16082_));
 OAI211_X2 _25801_ (.A(_16082_),
    .B(_15666_),
    .C1(_15867_),
    .C2(_15826_),
    .ZN(_16083_));
 NOR4_X1 _25802_ (.A1(_16077_),
    .A2(_16080_),
    .A3(_16081_),
    .A4(_16083_),
    .ZN(_16084_));
 NAND4_X1 _25803_ (.A1(_16056_),
    .A2(_16064_),
    .A3(_16072_),
    .A4(_16084_),
    .ZN(_16085_));
 AND3_X1 _25804_ (.A1(_15614_),
    .A2(_15562_),
    .A3(_15596_),
    .ZN(_16086_));
 OR3_X1 _25805_ (.A1(_15846_),
    .A2(_16009_),
    .A3(_16086_),
    .ZN(_16087_));
 AOI21_X1 _25806_ (.A(_15902_),
    .B1(_15615_),
    .B2(_15609_),
    .ZN(_16088_));
 AOI21_X1 _25807_ (.A(_15902_),
    .B1(_16041_),
    .B2(_15944_),
    .ZN(_16089_));
 NOR4_X1 _25808_ (.A1(_15730_),
    .A2(_16087_),
    .A3(_16088_),
    .A4(_16089_),
    .ZN(_16090_));
 OAI21_X1 _25809_ (.A(_15760_),
    .B1(_15602_),
    .B2(_15656_),
    .ZN(_16091_));
 NAND4_X1 _25810_ (.A1(_15754_),
    .A2(_15678_),
    .A3(_15755_),
    .A4(_11004_),
    .ZN(_16092_));
 NAND2_X1 _25811_ (.A1(_15760_),
    .A2(_15937_),
    .ZN(_16093_));
 NAND3_X1 _25812_ (.A1(_16091_),
    .A2(_16092_),
    .A3(_16093_),
    .ZN(_16094_));
 NAND2_X1 _25813_ (.A1(_15744_),
    .A2(_15850_),
    .ZN(_16095_));
 NOR4_X1 _25814_ (.A1(_16094_),
    .A2(_16095_),
    .A3(_15568_),
    .A4(_16039_),
    .ZN(_16096_));
 OAI211_X2 _25815_ (.A(_15635_),
    .B(_15678_),
    .C1(_11004_),
    .C2(_15581_),
    .ZN(_16097_));
 OAI21_X1 _25816_ (.A(_15635_),
    .B1(_15614_),
    .B2(_15686_),
    .ZN(_16098_));
 NAND2_X1 _25817_ (.A1(_15602_),
    .A2(_15635_),
    .ZN(_16099_));
 NAND4_X1 _25818_ (.A1(_16097_),
    .A2(_16098_),
    .A3(_15870_),
    .A4(_16099_),
    .ZN(_16100_));
 AOI21_X1 _25819_ (.A(_15617_),
    .B1(_15836_),
    .B2(_16066_),
    .ZN(_16101_));
 NOR3_X1 _25820_ (.A1(_15919_),
    .A2(_16100_),
    .A3(_16101_),
    .ZN(_16102_));
 AND2_X1 _25821_ (.A1(_15727_),
    .A2(_15630_),
    .ZN(_16103_));
 AOI211_X4 _25822_ (.A(_15631_),
    .B(_16103_),
    .C1(_15652_),
    .C2(_15630_),
    .ZN(_16104_));
 OAI21_X1 _25823_ (.A(_15621_),
    .B1(_15719_),
    .B2(_15559_),
    .ZN(_16105_));
 OAI21_X1 _25824_ (.A(_15621_),
    .B1(_15813_),
    .B2(_15772_),
    .ZN(_16106_));
 AND3_X1 _25825_ (.A1(_16104_),
    .A2(_16105_),
    .A3(_16106_),
    .ZN(_16107_));
 NAND4_X1 _25826_ (.A1(_16090_),
    .A2(_16096_),
    .A3(_16102_),
    .A4(_16107_),
    .ZN(_16108_));
 NOR2_X1 _25827_ (.A1(_16085_),
    .A2(_16108_),
    .ZN(_16109_));
 XOR2_X1 _25828_ (.A(_16109_),
    .B(_01009_),
    .Z(_16110_));
 MUX2_X1 _25829_ (.A(_01220_),
    .B(_16110_),
    .S(_15298_),
    .Z(_01070_));
 AND2_X1 _25830_ (.A1(_15564_),
    .A2(_15656_),
    .ZN(_16111_));
 AOI21_X1 _25831_ (.A(_16036_),
    .B1(_15828_),
    .B2(_16070_),
    .ZN(_16112_));
 INV_X1 _25832_ (.A(_15820_),
    .ZN(_16113_));
 AOI211_X4 _25833_ (.A(_16111_),
    .B(_16112_),
    .C1(_15741_),
    .C2(_16113_),
    .ZN(_16114_));
 AND2_X1 _25834_ (.A1(_15575_),
    .A2(_15601_),
    .ZN(_16115_));
 AND2_X1 _25835_ (.A1(_15575_),
    .A2(_15664_),
    .ZN(_16116_));
 OR4_X1 _25836_ (.A1(_15846_),
    .A2(_16115_),
    .A3(_16116_),
    .A4(_16086_),
    .ZN(_16117_));
 AND2_X1 _25837_ (.A1(_15576_),
    .A2(_15668_),
    .ZN(_16118_));
 AOI211_X4 _25838_ (.A(_15751_),
    .B(_15897_),
    .C1(_15736_),
    .C2(_15699_),
    .ZN(_16119_));
 NOR3_X1 _25839_ (.A1(_16117_),
    .A2(_16118_),
    .A3(_16119_),
    .ZN(_16120_));
 AND3_X1 _25840_ (.A1(_15664_),
    .A2(_15562_),
    .A3(_15755_),
    .ZN(_16121_));
 AOI211_X4 _25841_ (.A(_16121_),
    .B(_16042_),
    .C1(_15760_),
    .C2(_15692_),
    .ZN(_16122_));
 NAND2_X1 _25842_ (.A1(_15578_),
    .A2(_15816_),
    .ZN(_16123_));
 OAI211_X2 _25843_ (.A(_15578_),
    .B(_15652_),
    .C1(_15640_),
    .C2(_11011_),
    .ZN(_16124_));
 OAI21_X1 _25844_ (.A(_15578_),
    .B1(_15549_),
    .B2(_15701_),
    .ZN(_16125_));
 AND4_X1 _25845_ (.A1(_16123_),
    .A2(_16124_),
    .A3(_15896_),
    .A4(_16125_),
    .ZN(_16126_));
 AND4_X1 _25846_ (.A1(_16114_),
    .A2(_16120_),
    .A3(_16122_),
    .A4(_16126_),
    .ZN(_16127_));
 AND4_X1 _25847_ (.A1(_15645_),
    .A2(_15616_),
    .A3(_15699_),
    .A4(_15679_),
    .ZN(_16128_));
 AOI211_X4 _25848_ (.A(_16128_),
    .B(_15913_),
    .C1(_15686_),
    .C2(_15616_),
    .ZN(_16129_));
 OAI211_X2 _25849_ (.A(_16129_),
    .B(_15917_),
    .C1(_15985_),
    .C2(_15617_),
    .ZN(_16130_));
 NAND2_X1 _25850_ (.A1(_15813_),
    .A2(_15635_),
    .ZN(_16131_));
 OAI21_X1 _25851_ (.A(_15635_),
    .B1(_15637_),
    .B2(_15686_),
    .ZN(_16132_));
 NAND4_X1 _25852_ (.A1(_16021_),
    .A2(_16131_),
    .A3(_16099_),
    .A4(_16132_),
    .ZN(_16133_));
 AND2_X1 _25853_ (.A1(_15822_),
    .A2(_15630_),
    .ZN(_16134_));
 NAND2_X1 _25854_ (.A1(_15816_),
    .A2(_15630_),
    .ZN(_16135_));
 NAND2_X1 _25855_ (.A1(_15921_),
    .A2(_16135_),
    .ZN(_16136_));
 AND2_X1 _25856_ (.A1(_15630_),
    .A2(_15999_),
    .ZN(_16137_));
 OR4_X1 _25857_ (.A1(_16134_),
    .A2(_16136_),
    .A3(_15633_),
    .A4(_16137_),
    .ZN(_16138_));
 OAI21_X1 _25858_ (.A(_15620_),
    .B1(_15765_),
    .B2(_15705_),
    .ZN(_16139_));
 NAND2_X1 _25859_ (.A1(_15573_),
    .A2(_15620_),
    .ZN(_16140_));
 OAI211_X2 _25860_ (.A(_16139_),
    .B(_16140_),
    .C1(_16066_),
    .C2(_15922_),
    .ZN(_16141_));
 NOR4_X1 _25861_ (.A1(_16130_),
    .A2(_16133_),
    .A3(_16138_),
    .A4(_16141_),
    .ZN(_16142_));
 NOR2_X1 _25862_ (.A1(_16052_),
    .A2(_15798_),
    .ZN(_16143_));
 NAND4_X1 _25863_ (.A1(_15624_),
    .A2(_15551_),
    .A3(_15636_),
    .A4(_15648_),
    .ZN(_16144_));
 AND3_X1 _25864_ (.A1(_16143_),
    .A2(_15800_),
    .A3(_16144_),
    .ZN(_16145_));
 OR2_X1 _25865_ (.A1(_15572_),
    .A2(_15815_),
    .ZN(_16146_));
 AND2_X1 _25866_ (.A1(_16146_),
    .A2(_15708_),
    .ZN(_16147_));
 INV_X1 _25867_ (.A(_16147_),
    .ZN(_16148_));
 NAND3_X1 _25868_ (.A1(_15567_),
    .A2(_15708_),
    .A3(_15699_),
    .ZN(_16149_));
 OAI211_X2 _25869_ (.A(_15708_),
    .B(_15622_),
    .C1(_15639_),
    .C2(_11003_),
    .ZN(_16150_));
 AND4_X1 _25870_ (.A1(_15932_),
    .A2(_16148_),
    .A3(_16149_),
    .A4(_16150_),
    .ZN(_16151_));
 NAND2_X1 _25871_ (.A1(_15559_),
    .A2(_15673_),
    .ZN(_16152_));
 OAI21_X1 _25872_ (.A(_15673_),
    .B1(_15711_),
    .B2(_15573_),
    .ZN(_16153_));
 OAI221_X1 _25873_ (.A(_15673_),
    .B1(_15639_),
    .B2(_11003_),
    .C1(_15588_),
    .C2(_15622_),
    .ZN(_16154_));
 NAND3_X1 _25874_ (.A1(_15673_),
    .A2(_15624_),
    .A3(_15679_),
    .ZN(_16155_));
 AND4_X1 _25875_ (.A1(_16152_),
    .A2(_16153_),
    .A3(_16154_),
    .A4(_16155_),
    .ZN(_16156_));
 NAND2_X1 _25876_ (.A1(_15605_),
    .A2(_15701_),
    .ZN(_16157_));
 NAND4_X1 _25877_ (.A1(_15596_),
    .A2(_15639_),
    .A3(_15588_),
    .A4(_15648_),
    .ZN(_16158_));
 OAI211_X2 _25878_ (.A(_16157_),
    .B(_16158_),
    .C1(_15958_),
    .C2(_15903_),
    .ZN(_16159_));
 AOI211_X4 _25879_ (.A(_15961_),
    .B(_16159_),
    .C1(_15605_),
    .C2(_15795_),
    .ZN(_16160_));
 AND4_X1 _25880_ (.A1(_16145_),
    .A2(_16151_),
    .A3(_16156_),
    .A4(_16160_),
    .ZN(_16161_));
 AOI211_X4 _25881_ (.A(_15731_),
    .B(_15818_),
    .C1(_10996_),
    .C2(_11003_),
    .ZN(_16162_));
 AND2_X1 _25882_ (.A1(_15695_),
    .A2(_15656_),
    .ZN(_16163_));
 INV_X1 _25883_ (.A(_15549_),
    .ZN(_16164_));
 AOI21_X1 _25884_ (.A(_15818_),
    .B1(_16070_),
    .B2(_16164_),
    .ZN(_16165_));
 NOR3_X1 _25885_ (.A1(_16162_),
    .A2(_16163_),
    .A3(_16165_),
    .ZN(_16166_));
 OAI21_X1 _25886_ (.A(_15594_),
    .B1(_15614_),
    .B2(_15719_),
    .ZN(_16167_));
 AND3_X1 _25887_ (.A1(_16167_),
    .A2(_15767_),
    .A3(_15766_),
    .ZN(_16168_));
 NAND2_X1 _25888_ (.A1(_15598_),
    .A2(_15772_),
    .ZN(_16169_));
 AND4_X1 _25889_ (.A1(_16074_),
    .A2(_16073_),
    .A3(_15834_),
    .A4(_16169_),
    .ZN(_16170_));
 INV_X1 _25890_ (.A(_16078_),
    .ZN(_16171_));
 OAI21_X1 _25891_ (.A(_15663_),
    .B1(_15632_),
    .B2(_15595_),
    .ZN(_16172_));
 AND4_X1 _25892_ (.A1(_15748_),
    .A2(_16171_),
    .A3(_15747_),
    .A4(_16172_),
    .ZN(_16173_));
 AND4_X1 _25893_ (.A1(_16166_),
    .A2(_16168_),
    .A3(_16170_),
    .A4(_16173_),
    .ZN(_16174_));
 NAND4_X1 _25894_ (.A1(_16127_),
    .A2(_16142_),
    .A3(_16161_),
    .A4(_16174_),
    .ZN(_16175_));
 NOR2_X1 _25895_ (.A1(_16175_),
    .A2(_15714_),
    .ZN(_16176_));
 XOR2_X1 _25896_ (.A(_16176_),
    .B(_01010_),
    .Z(_16177_));
 BUF_X4 _25897_ (.A(_03738_),
    .Z(_16178_));
 MUX2_X1 _25898_ (.A(_01221_),
    .B(_16177_),
    .S(_16178_),
    .Z(_01071_));
 XOR2_X1 _25899_ (.A(_17241_),
    .B(_17076_),
    .Z(_16179_));
 XOR2_X2 _25900_ (.A(_12472_),
    .B(_12904_),
    .Z(_16180_));
 XNOR2_X2 _25901_ (.A(_16180_),
    .B(_12737_),
    .ZN(_16181_));
 XNOR2_X1 _25902_ (.A(_16181_),
    .B(_13199_),
    .ZN(_16182_));
 XOR2_X1 _25903_ (.A(_16182_),
    .B(_17241_),
    .Z(_16183_));
 MUX2_X1 _25904_ (.A(_16179_),
    .B(_16183_),
    .S(_15306_),
    .Z(_00686_));
 AND4_X1 _25905_ (.A1(_15551_),
    .A2(_15562_),
    .A3(_15557_),
    .A4(_15590_),
    .ZN(_16184_));
 AND4_X1 _25906_ (.A1(_15577_),
    .A2(_15645_),
    .A3(_15698_),
    .A4(_15571_),
    .ZN(_16185_));
 AOI211_X4 _25907_ (.A(_16184_),
    .B(_16185_),
    .C1(_15578_),
    .C2(_15685_),
    .ZN(_16186_));
 OAI21_X1 _25908_ (.A(_15733_),
    .B1(_15807_),
    .B2(_15584_),
    .ZN(_16187_));
 OAI21_X1 _25909_ (.A(_15733_),
    .B1(_15702_),
    .B2(_15813_),
    .ZN(_16188_));
 AND3_X1 _25910_ (.A1(_16186_),
    .A2(_16187_),
    .A3(_16188_),
    .ZN(_16189_));
 NAND2_X1 _25911_ (.A1(_15564_),
    .A2(_15688_),
    .ZN(_16190_));
 OAI211_X2 _25912_ (.A(_15851_),
    .B(_16190_),
    .C1(_16036_),
    .C2(_15985_),
    .ZN(_16191_));
 AND2_X1 _25913_ (.A1(_15771_),
    .A2(_15564_),
    .ZN(_16192_));
 AOI211_X4 _25914_ (.A(_16191_),
    .B(_16192_),
    .C1(_15781_),
    .C2(_15741_),
    .ZN(_16193_));
 AND2_X1 _25915_ (.A1(_15759_),
    .A2(_15937_),
    .ZN(_16194_));
 NOR4_X1 _25916_ (.A1(_15890_),
    .A2(_15857_),
    .A3(_16194_),
    .A4(_16121_),
    .ZN(_16195_));
 NOR2_X1 _25917_ (.A1(_16008_),
    .A2(_16009_),
    .ZN(_16196_));
 INV_X1 _25918_ (.A(_16196_),
    .ZN(_16197_));
 NOR4_X1 _25919_ (.A1(_16197_),
    .A2(_16118_),
    .A3(_15844_),
    .A4(_16116_),
    .ZN(_16198_));
 AND4_X1 _25920_ (.A1(_16189_),
    .A2(_16193_),
    .A3(_16195_),
    .A4(_16198_),
    .ZN(_16199_));
 AND3_X1 _25921_ (.A1(_15591_),
    .A2(_15648_),
    .A3(_15755_),
    .ZN(_16200_));
 AOI211_X4 _25922_ (.A(_16200_),
    .B(_16058_),
    .C1(_15708_),
    .C2(_15765_),
    .ZN(_16201_));
 AND3_X1 _25923_ (.A1(_15932_),
    .A2(_15974_),
    .A3(_15976_),
    .ZN(_16202_));
 OAI211_X2 _25924_ (.A(_15709_),
    .B(_15680_),
    .C1(_15624_),
    .C2(_15590_),
    .ZN(_16203_));
 NAND4_X1 _25925_ (.A1(_16201_),
    .A2(_15975_),
    .A3(_16202_),
    .A4(_16203_),
    .ZN(_16204_));
 AOI211_X4 _25926_ (.A(_15784_),
    .B(_15674_),
    .C1(_15573_),
    .C2(_15673_),
    .ZN(_16205_));
 NAND4_X1 _25927_ (.A1(_16205_),
    .A2(_16152_),
    .A3(_15789_),
    .A4(_15938_),
    .ZN(_16206_));
 AND2_X1 _25928_ (.A1(_15605_),
    .A2(_15632_),
    .ZN(_16207_));
 AND2_X1 _25929_ (.A1(_15605_),
    .A2(_15701_),
    .ZN(_16208_));
 AND2_X1 _25930_ (.A1(_15605_),
    .A2(_15688_),
    .ZN(_16209_));
 OR4_X1 _25931_ (.A1(_16207_),
    .A2(_16208_),
    .A3(_15963_),
    .A4(_16209_),
    .ZN(_16210_));
 OAI211_X2 _25932_ (.A(_15554_),
    .B(_15652_),
    .C1(_15626_),
    .C2(_15590_),
    .ZN(_16211_));
 OAI211_X2 _25933_ (.A(_16211_),
    .B(_15800_),
    .C1(_15810_),
    .C2(_16051_),
    .ZN(_16212_));
 NOR4_X1 _25934_ (.A1(_16204_),
    .A2(_16206_),
    .A3(_16210_),
    .A4(_16212_),
    .ZN(_16213_));
 OAI21_X1 _25935_ (.A(_15687_),
    .B1(_15602_),
    .B2(_15711_),
    .ZN(_16214_));
 OAI21_X1 _25936_ (.A(_15594_),
    .B1(_15984_),
    .B2(_15807_),
    .ZN(_16215_));
 AND2_X1 _25937_ (.A1(_16214_),
    .A2(_16215_),
    .ZN(_16216_));
 AND2_X1 _25938_ (.A1(_15694_),
    .A2(_15719_),
    .ZN(_16217_));
 NOR4_X1 _25939_ (.A1(_15737_),
    .A2(_15814_),
    .A3(_16217_),
    .A4(_15996_),
    .ZN(_16218_));
 AND2_X1 _25940_ (.A1(_15816_),
    .A2(_15662_),
    .ZN(_16219_));
 AND2_X1 _25941_ (.A1(_15662_),
    .A2(_15742_),
    .ZN(_16220_));
 NOR4_X1 _25942_ (.A1(_15831_),
    .A2(_16079_),
    .A3(_16219_),
    .A4(_16220_),
    .ZN(_16221_));
 NAND2_X1 _25943_ (.A1(_15598_),
    .A2(_15685_),
    .ZN(_16222_));
 OAI21_X1 _25944_ (.A(_15598_),
    .B1(_15739_),
    .B2(_15584_),
    .ZN(_16223_));
 AND4_X1 _25945_ (.A1(_15693_),
    .A2(_15658_),
    .A3(_16222_),
    .A4(_16223_),
    .ZN(_16224_));
 AND4_X1 _25946_ (.A1(_16216_),
    .A2(_16218_),
    .A3(_16221_),
    .A4(_16224_),
    .ZN(_16225_));
 OAI21_X1 _25947_ (.A(_15612_),
    .B1(_15984_),
    .B2(_15807_),
    .ZN(_16226_));
 OAI21_X1 _25948_ (.A(_15612_),
    .B1(_15656_),
    .B2(_15665_),
    .ZN(_16227_));
 NAND4_X1 _25949_ (.A1(_15755_),
    .A2(_15679_),
    .A3(_15640_),
    .A4(_15611_),
    .ZN(_16228_));
 AND3_X1 _25950_ (.A1(_16226_),
    .A2(_16227_),
    .A3(_16228_),
    .ZN(_16229_));
 AOI21_X1 _25951_ (.A(_15881_),
    .B1(_16164_),
    .B2(_15944_),
    .ZN(_16230_));
 AOI211_X4 _25952_ (.A(_15731_),
    .B(_15881_),
    .C1(_15736_),
    .C2(_15699_),
    .ZN(_16231_));
 AOI211_X4 _25953_ (.A(_16230_),
    .B(_16231_),
    .C1(_15711_),
    .C2(_15630_),
    .ZN(_16232_));
 INV_X1 _25954_ (.A(_15632_),
    .ZN(_16233_));
 INV_X1 _25955_ (.A(_15816_),
    .ZN(_16234_));
 AOI21_X1 _25956_ (.A(_15617_),
    .B1(_16233_),
    .B2(_16234_),
    .ZN(_16235_));
 AND2_X1 _25957_ (.A1(_15822_),
    .A2(_15651_),
    .ZN(_16236_));
 NOR4_X1 _25958_ (.A1(_16235_),
    .A2(_16236_),
    .A3(_16014_),
    .A4(_15860_),
    .ZN(_16237_));
 NOR2_X1 _25959_ (.A1(_15924_),
    .A2(_15873_),
    .ZN(_16238_));
 NAND2_X1 _25960_ (.A1(_15705_),
    .A2(_15620_),
    .ZN(_16239_));
 OAI21_X1 _25961_ (.A(_15620_),
    .B1(_15692_),
    .B2(_15686_),
    .ZN(_16240_));
 AND3_X1 _25962_ (.A1(_16238_),
    .A2(_16239_),
    .A3(_16240_),
    .ZN(_16241_));
 AND4_X1 _25963_ (.A1(_16229_),
    .A2(_16232_),
    .A3(_16237_),
    .A4(_16241_),
    .ZN(_16242_));
 NAND4_X1 _25964_ (.A1(_16199_),
    .A2(_16213_),
    .A3(_16225_),
    .A4(_16242_),
    .ZN(_16243_));
 NOR2_X1 _25965_ (.A1(_16243_),
    .A2(_15714_),
    .ZN(_16244_));
 INV_X1 _25966_ (.A(_01011_),
    .ZN(_16245_));
 XNOR2_X1 _25967_ (.A(_16244_),
    .B(_16245_),
    .ZN(_16246_));
 MUX2_X1 _25968_ (.A(_01222_),
    .B(_16246_),
    .S(_16178_),
    .Z(_01072_));
 AOI21_X1 _25969_ (.A(_15922_),
    .B1(_15615_),
    .B2(_16066_),
    .ZN(_16247_));
 AOI211_X4 _25970_ (.A(_15925_),
    .B(_16247_),
    .C1(_15711_),
    .C2(_15621_),
    .ZN(_16248_));
 NOR3_X1 _25971_ (.A1(_15628_),
    .A2(_15874_),
    .A3(_15873_),
    .ZN(_16249_));
 OAI21_X1 _25972_ (.A(_15774_),
    .B1(_15692_),
    .B2(_15643_),
    .ZN(_16250_));
 OAI21_X1 _25973_ (.A(_15774_),
    .B1(_15727_),
    .B2(_15999_),
    .ZN(_16251_));
 AND4_X1 _25974_ (.A1(_16248_),
    .A2(_16249_),
    .A3(_16250_),
    .A4(_16251_),
    .ZN(_16252_));
 NAND2_X1 _25975_ (.A1(_15741_),
    .A2(_15813_),
    .ZN(_16253_));
 AOI21_X1 _25976_ (.A(_16042_),
    .B1(_15760_),
    .B2(_16113_),
    .ZN(_16254_));
 OAI21_X1 _25977_ (.A(_15741_),
    .B1(_15771_),
    .B2(_15711_),
    .ZN(_16255_));
 OAI21_X1 _25978_ (.A(_15760_),
    .B1(_15595_),
    .B2(_15683_),
    .ZN(_16256_));
 AND4_X1 _25979_ (.A1(_16253_),
    .A2(_16254_),
    .A3(_16255_),
    .A4(_16256_),
    .ZN(_16257_));
 AND3_X1 _25980_ (.A1(_15702_),
    .A2(_15551_),
    .A3(_15754_),
    .ZN(_16258_));
 NOR2_X1 _25981_ (.A1(_15901_),
    .A2(_16258_),
    .ZN(_16259_));
 NAND2_X1 _25982_ (.A1(_15576_),
    .A2(_15665_),
    .ZN(_16260_));
 OAI221_X1 _25983_ (.A(_15576_),
    .B1(_15640_),
    .B2(_11011_),
    .C1(_15652_),
    .C2(_15678_),
    .ZN(_16261_));
 OAI21_X1 _25984_ (.A(_15733_),
    .B1(_15732_),
    .B2(_15686_),
    .ZN(_16262_));
 AND4_X1 _25985_ (.A1(_16259_),
    .A2(_16260_),
    .A3(_16261_),
    .A4(_16262_),
    .ZN(_16263_));
 AOI22_X1 _25986_ (.A1(_15914_),
    .A2(_15645_),
    .B1(_15665_),
    .B2(_15651_),
    .ZN(_16264_));
 AND2_X1 _25987_ (.A1(_15612_),
    .A2(_15591_),
    .ZN(_16265_));
 AOI211_X4 _25988_ (.A(_16265_),
    .B(_16020_),
    .C1(_15689_),
    .C2(_15635_),
    .ZN(_16266_));
 NOR3_X1 _25989_ (.A1(_15916_),
    .A2(_16014_),
    .A3(_15861_),
    .ZN(_16267_));
 OAI211_X2 _25990_ (.A(_15635_),
    .B(_15624_),
    .C1(_15636_),
    .C2(_15680_),
    .ZN(_16268_));
 AND4_X1 _25991_ (.A1(_16264_),
    .A2(_16266_),
    .A3(_16267_),
    .A4(_16268_),
    .ZN(_16269_));
 NAND4_X1 _25992_ (.A1(_16252_),
    .A2(_16257_),
    .A3(_16263_),
    .A4(_16269_),
    .ZN(_16270_));
 AOI211_X4 _25993_ (.A(_15788_),
    .B(_15972_),
    .C1(_15677_),
    .C2(_16146_),
    .ZN(_16271_));
 OAI21_X1 _25994_ (.A(_15709_),
    .B1(_15937_),
    .B2(_15678_),
    .ZN(_16272_));
 OAI21_X1 _25995_ (.A(_15709_),
    .B1(_15614_),
    .B2(_15686_),
    .ZN(_16273_));
 AND4_X1 _25996_ (.A1(_16148_),
    .A2(_16271_),
    .A3(_16272_),
    .A4(_16273_),
    .ZN(_16274_));
 AND2_X1 _25997_ (.A1(_15601_),
    .A2(_15694_),
    .ZN(_16275_));
 AOI221_X4 _25998_ (.A(_16275_),
    .B1(_15683_),
    .B2(_15695_),
    .C1(_11011_),
    .C2(_16217_),
    .ZN(_16276_));
 AOI21_X1 _25999_ (.A(_15818_),
    .B1(_15827_),
    .B2(_15828_),
    .ZN(_16277_));
 AOI21_X1 _26000_ (.A(_16277_),
    .B1(_15695_),
    .B2(_15591_),
    .ZN(_16278_));
 OAI21_X1 _26001_ (.A(_15687_),
    .B1(_15632_),
    .B2(_15816_),
    .ZN(_16279_));
 OAI21_X1 _26002_ (.A(_15687_),
    .B1(_15702_),
    .B2(_15772_),
    .ZN(_16280_));
 AND4_X1 _26003_ (.A1(_16276_),
    .A2(_16278_),
    .A3(_16279_),
    .A4(_16280_),
    .ZN(_16281_));
 OAI21_X1 _26004_ (.A(_15603_),
    .B1(_15702_),
    .B2(_15999_),
    .ZN(_16282_));
 AOI21_X1 _26005_ (.A(_15650_),
    .B1(_15642_),
    .B2(_15807_),
    .ZN(_16283_));
 OAI21_X1 _26006_ (.A(_15642_),
    .B1(_15595_),
    .B2(_15643_),
    .ZN(_16284_));
 OAI211_X2 _26007_ (.A(_15603_),
    .B(_10997_),
    .C1(_15636_),
    .C2(_15680_),
    .ZN(_16285_));
 AND4_X1 _26008_ (.A1(_16282_),
    .A2(_16283_),
    .A3(_16284_),
    .A4(_16285_),
    .ZN(_16286_));
 INV_X1 _26009_ (.A(_15952_),
    .ZN(_16287_));
 NAND2_X1 _26010_ (.A1(_15659_),
    .A2(_15637_),
    .ZN(_16288_));
 OAI21_X1 _26011_ (.A(_15659_),
    .B1(_15727_),
    .B2(_15668_),
    .ZN(_16289_));
 NAND4_X1 _26012_ (.A1(_16287_),
    .A2(_16288_),
    .A3(_16222_),
    .A4(_16289_),
    .ZN(_16290_));
 OAI211_X2 _26013_ (.A(_16082_),
    .B(_15684_),
    .C1(_16234_),
    .C2(_15826_),
    .ZN(_16291_));
 NOR4_X1 _26014_ (.A1(_16290_),
    .A2(_16080_),
    .A3(_15831_),
    .A4(_16291_),
    .ZN(_16292_));
 NAND4_X1 _26015_ (.A1(_16274_),
    .A2(_16281_),
    .A3(_16286_),
    .A4(_16292_),
    .ZN(_16293_));
 NOR2_X1 _26016_ (.A1(_16270_),
    .A2(_16293_),
    .ZN(_16294_));
 XOR2_X1 _26017_ (.A(_16294_),
    .B(_01012_),
    .Z(_16295_));
 MUX2_X1 _26018_ (.A(_01223_),
    .B(_16295_),
    .S(_16178_),
    .Z(_01073_));
 INV_X1 _26019_ (.A(_17151_),
    .ZN(_16296_));
 NOR2_X1 _26020_ (.A1(_16296_),
    .A2(_17152_),
    .ZN(_16297_));
 BUF_X4 _26021_ (.A(_16297_),
    .Z(_16298_));
 INV_X1 _26022_ (.A(_16298_),
    .ZN(_16299_));
 NOR2_X1 _26023_ (.A1(_11076_),
    .A2(_17153_),
    .ZN(_16300_));
 BUF_X4 _26024_ (.A(_16300_),
    .Z(_16301_));
 NAND2_X1 _26025_ (.A1(_16299_),
    .A2(_16301_),
    .ZN(_16302_));
 INV_X1 _26026_ (.A(_17152_),
    .ZN(_16303_));
 NOR2_X2 _26027_ (.A1(_16303_),
    .A2(_17151_),
    .ZN(_16304_));
 BUF_X4 _26028_ (.A(_16304_),
    .Z(_16305_));
 NOR2_X1 _26029_ (.A1(_16302_),
    .A2(_16305_),
    .ZN(_16306_));
 INV_X1 _26030_ (.A(_17157_),
    .ZN(_16307_));
 AND2_X2 _26031_ (.A1(_16307_),
    .A2(_17156_),
    .ZN(_16308_));
 NOR2_X1 _26032_ (.A1(_17158_),
    .A2(_17159_),
    .ZN(_16309_));
 AND2_X1 _26033_ (.A1(_16308_),
    .A2(_16309_),
    .ZN(_16310_));
 BUF_X4 _26034_ (.A(_16310_),
    .Z(_16311_));
 NAND2_X1 _26035_ (.A1(_16306_),
    .A2(_16311_),
    .ZN(_16312_));
 BUF_X4 _26036_ (.A(_16311_),
    .Z(_16313_));
 NOR2_X1 _26037_ (.A1(_17153_),
    .A2(_17154_),
    .ZN(_16314_));
 AND2_X2 _26038_ (.A1(_16314_),
    .A2(_17152_),
    .ZN(_16315_));
 NAND2_X1 _26039_ (.A1(_16313_),
    .A2(_16315_),
    .ZN(_16316_));
 INV_X1 _26040_ (.A(_16311_),
    .ZN(_16317_));
 NOR2_X4 _26041_ (.A1(_17151_),
    .A2(_17152_),
    .ZN(_16318_));
 INV_X1 _26042_ (.A(_16318_),
    .ZN(_16319_));
 NOR2_X1 _26043_ (.A1(_11068_),
    .A2(_17154_),
    .ZN(_16320_));
 BUF_X4 _26044_ (.A(_16320_),
    .Z(_16321_));
 NAND2_X1 _26045_ (.A1(_16319_),
    .A2(_16321_),
    .ZN(_16322_));
 AND2_X2 _26046_ (.A1(_17151_),
    .A2(_17152_),
    .ZN(_16323_));
 NOR2_X1 _26047_ (.A1(_16322_),
    .A2(_16323_),
    .ZN(_16324_));
 INV_X1 _26048_ (.A(_16324_),
    .ZN(_16325_));
 OAI211_X2 _26049_ (.A(_16312_),
    .B(_16316_),
    .C1(_16317_),
    .C2(_16325_),
    .ZN(_16326_));
 AND2_X1 _26050_ (.A1(_16321_),
    .A2(_17152_),
    .ZN(_16327_));
 BUF_X4 _26051_ (.A(_16327_),
    .Z(_16328_));
 NOR2_X1 _26052_ (.A1(_17156_),
    .A2(_17157_),
    .ZN(_16329_));
 BUF_X2 _26053_ (.A(_16309_),
    .Z(_16330_));
 AND2_X2 _26054_ (.A1(_16329_),
    .A2(_16330_),
    .ZN(_16331_));
 AND2_X1 _26055_ (.A1(_16328_),
    .A2(_16331_),
    .ZN(_16332_));
 INV_X1 _26056_ (.A(_16332_),
    .ZN(_16333_));
 BUF_X4 _26057_ (.A(_16321_),
    .Z(_16334_));
 NAND3_X1 _26058_ (.A1(_16331_),
    .A2(_16334_),
    .A3(_16298_),
    .ZN(_16335_));
 INV_X1 _26059_ (.A(_16315_),
    .ZN(_16336_));
 INV_X1 _26060_ (.A(_16331_),
    .ZN(_16337_));
 OAI211_X2 _26061_ (.A(_16333_),
    .B(_16335_),
    .C1(_16336_),
    .C2(_16337_),
    .ZN(_16338_));
 AND2_X1 _26062_ (.A1(_16300_),
    .A2(_17152_),
    .ZN(_16339_));
 BUF_X2 _26063_ (.A(_16339_),
    .Z(_16340_));
 NAND2_X1 _26064_ (.A1(_16340_),
    .A2(_16331_),
    .ZN(_16341_));
 NAND3_X1 _26065_ (.A1(_16331_),
    .A2(_16298_),
    .A3(_16301_),
    .ZN(_16342_));
 AND2_X2 _26066_ (.A1(_17153_),
    .A2(_17154_),
    .ZN(_16343_));
 AND2_X1 _26067_ (.A1(_16304_),
    .A2(_16343_),
    .ZN(_16344_));
 BUF_X4 _26068_ (.A(_16343_),
    .Z(_16345_));
 AND2_X4 _26069_ (.A1(_16297_),
    .A2(_16345_),
    .ZN(_16346_));
 NOR2_X4 _26070_ (.A1(_16344_),
    .A2(_16346_),
    .ZN(_16347_));
 OAI211_X2 _26071_ (.A(_16341_),
    .B(_16342_),
    .C1(_16347_),
    .C2(_16337_),
    .ZN(_16348_));
 NOR3_X1 _26072_ (.A1(_16326_),
    .A2(_16338_),
    .A3(_16348_),
    .ZN(_16349_));
 INV_X1 _26073_ (.A(_16345_),
    .ZN(_16350_));
 AND2_X1 _26074_ (.A1(_17156_),
    .A2(_17157_),
    .ZN(_16351_));
 AND2_X1 _26075_ (.A1(_16351_),
    .A2(_16330_),
    .ZN(_16352_));
 BUF_X4 _26076_ (.A(_16352_),
    .Z(_16353_));
 INV_X1 _26077_ (.A(_16353_),
    .ZN(_16354_));
 AOI211_X4 _26078_ (.A(_16350_),
    .B(_16354_),
    .C1(_16296_),
    .C2(_11056_),
    .ZN(_16355_));
 AND3_X1 _26079_ (.A1(_16353_),
    .A2(_16334_),
    .A3(_16305_),
    .ZN(_16356_));
 BUF_X4 _26080_ (.A(_16314_),
    .Z(_16357_));
 NAND2_X1 _26081_ (.A1(_16319_),
    .A2(_16357_),
    .ZN(_16358_));
 NOR2_X1 _26082_ (.A1(_16354_),
    .A2(_16358_),
    .ZN(_16359_));
 AND2_X2 _26083_ (.A1(_16300_),
    .A2(_16318_),
    .ZN(_16360_));
 AND2_X1 _26084_ (.A1(_16360_),
    .A2(_16353_),
    .ZN(_16361_));
 NOR4_X1 _26085_ (.A1(_16355_),
    .A2(_16356_),
    .A3(_16359_),
    .A4(_16361_),
    .ZN(_16362_));
 INV_X1 _26086_ (.A(_16323_),
    .ZN(_16363_));
 NOR2_X1 _26087_ (.A1(_16307_),
    .A2(_17156_),
    .ZN(_16364_));
 AND2_X1 _26088_ (.A1(_16364_),
    .A2(_16330_),
    .ZN(_16365_));
 BUF_X2 _26089_ (.A(_16365_),
    .Z(_16366_));
 BUF_X4 _26090_ (.A(_16366_),
    .Z(_16367_));
 INV_X1 _26091_ (.A(_16322_),
    .ZN(_16368_));
 OAI211_X2 _26092_ (.A(_16363_),
    .B(_16367_),
    .C1(_16368_),
    .C2(_16357_),
    .ZN(_16369_));
 AND2_X2 _26093_ (.A1(_16345_),
    .A2(_16318_),
    .ZN(_16370_));
 BUF_X2 _26094_ (.A(_16364_),
    .Z(_16371_));
 AND3_X1 _26095_ (.A1(_16370_),
    .A2(_16371_),
    .A3(_16330_),
    .ZN(_16372_));
 AND2_X1 _26096_ (.A1(_16345_),
    .A2(_17152_),
    .ZN(_16373_));
 AND2_X1 _26097_ (.A1(_16365_),
    .A2(_16373_),
    .ZN(_16374_));
 NAND2_X1 _26098_ (.A1(_16319_),
    .A2(_16301_),
    .ZN(_16375_));
 INV_X1 _26099_ (.A(_16375_),
    .ZN(_16376_));
 AOI211_X4 _26100_ (.A(_16372_),
    .B(_16374_),
    .C1(_16366_),
    .C2(_16376_),
    .ZN(_16377_));
 AND4_X1 _26101_ (.A1(_16349_),
    .A2(_16362_),
    .A3(_16369_),
    .A4(_16377_),
    .ZN(_16378_));
 AND2_X2 _26102_ (.A1(_17158_),
    .A2(_17159_),
    .ZN(_16379_));
 AND2_X2 _26103_ (.A1(_16364_),
    .A2(_16379_),
    .ZN(_16380_));
 BUF_X4 _26104_ (.A(_16380_),
    .Z(_16381_));
 AND2_X1 _26105_ (.A1(_16323_),
    .A2(_16314_),
    .ZN(_16382_));
 BUF_X4 _26106_ (.A(_16382_),
    .Z(_16383_));
 INV_X1 _26107_ (.A(_16383_),
    .ZN(_16384_));
 AND2_X1 _26108_ (.A1(_16314_),
    .A2(_16318_),
    .ZN(_16385_));
 INV_X1 _26109_ (.A(_16385_),
    .ZN(_16386_));
 NAND2_X1 _26110_ (.A1(_16384_),
    .A2(_16386_),
    .ZN(_16387_));
 BUF_X4 _26111_ (.A(_16303_),
    .Z(_16388_));
 AND2_X1 _26112_ (.A1(_16321_),
    .A2(_16388_),
    .ZN(_16389_));
 BUF_X2 _26113_ (.A(_16389_),
    .Z(_16390_));
 OAI21_X1 _26114_ (.A(_16381_),
    .B1(_16387_),
    .B2(_16390_),
    .ZN(_16391_));
 AND2_X1 _26115_ (.A1(_16308_),
    .A2(_16379_),
    .ZN(_16392_));
 BUF_X4 _26116_ (.A(_16392_),
    .Z(_16393_));
 AND2_X1 _26117_ (.A1(_16321_),
    .A2(_16298_),
    .ZN(_16394_));
 BUF_X2 _26118_ (.A(_16394_),
    .Z(_16395_));
 AND2_X1 _26119_ (.A1(_16304_),
    .A2(_16314_),
    .ZN(_16396_));
 BUF_X4 _26120_ (.A(_16396_),
    .Z(_16397_));
 OAI21_X1 _26121_ (.A(_16393_),
    .B1(_16395_),
    .B2(_16397_),
    .ZN(_16398_));
 AND2_X2 _26122_ (.A1(_16304_),
    .A2(_16300_),
    .ZN(_16399_));
 NAND2_X1 _26123_ (.A1(_16393_),
    .A2(_16399_),
    .ZN(_16400_));
 INV_X1 _26124_ (.A(_16392_),
    .ZN(_16401_));
 AND2_X1 _26125_ (.A1(_16300_),
    .A2(_16323_),
    .ZN(_16402_));
 INV_X1 _26126_ (.A(_16402_),
    .ZN(_16403_));
 OAI21_X1 _26127_ (.A(_16400_),
    .B1(_16401_),
    .B2(_16403_),
    .ZN(_16404_));
 NOR2_X1 _26128_ (.A1(_16347_),
    .A2(_16401_),
    .ZN(_16405_));
 AND2_X1 _26129_ (.A1(_16300_),
    .A2(_16388_),
    .ZN(_16406_));
 AOI211_X4 _26130_ (.A(_16404_),
    .B(_16405_),
    .C1(_16393_),
    .C2(_16406_),
    .ZN(_16407_));
 AND2_X1 _26131_ (.A1(_16379_),
    .A2(_16329_),
    .ZN(_16408_));
 BUF_X2 _26132_ (.A(_16408_),
    .Z(_16409_));
 BUF_X4 _26133_ (.A(_16409_),
    .Z(_16410_));
 NAND2_X1 _26134_ (.A1(_16397_),
    .A2(_16410_),
    .ZN(_16411_));
 AND2_X1 _26135_ (.A1(_16300_),
    .A2(_17151_),
    .ZN(_16412_));
 AND2_X1 _26136_ (.A1(_16412_),
    .A2(_16408_),
    .ZN(_16413_));
 NAND2_X1 _26137_ (.A1(_16346_),
    .A2(_16408_),
    .ZN(_16414_));
 NAND2_X1 _26138_ (.A1(_16370_),
    .A2(_16408_),
    .ZN(_16415_));
 NAND2_X1 _26139_ (.A1(_16414_),
    .A2(_16415_),
    .ZN(_16416_));
 AOI211_X4 _26140_ (.A(_16413_),
    .B(_16416_),
    .C1(_16344_),
    .C2(_16409_),
    .ZN(_16417_));
 AND4_X1 _26141_ (.A1(_16398_),
    .A2(_16407_),
    .A3(_16411_),
    .A4(_16417_),
    .ZN(_16418_));
 AND2_X2 _26142_ (.A1(_16345_),
    .A2(_17151_),
    .ZN(_16419_));
 AND2_X1 _26143_ (.A1(_16380_),
    .A2(_16419_),
    .ZN(_16420_));
 INV_X1 _26144_ (.A(_16380_),
    .ZN(_16421_));
 INV_X1 _26145_ (.A(_16399_),
    .ZN(_16422_));
 AOI21_X1 _26146_ (.A(_16421_),
    .B1(_16422_),
    .B2(_16403_),
    .ZN(_16423_));
 AOI211_X4 _26147_ (.A(_16420_),
    .B(_16423_),
    .C1(_16360_),
    .C2(_16380_),
    .ZN(_16424_));
 AND2_X1 _26148_ (.A1(_16379_),
    .A2(_16351_),
    .ZN(_16425_));
 CLKBUF_X2 _26149_ (.A(_16425_),
    .Z(_16426_));
 AND2_X1 _26150_ (.A1(_16344_),
    .A2(_16426_),
    .ZN(_16427_));
 AND2_X1 _26151_ (.A1(_16320_),
    .A2(_16318_),
    .ZN(_16428_));
 AND2_X1 _26152_ (.A1(_16428_),
    .A2(_16425_),
    .ZN(_16429_));
 INV_X1 _26153_ (.A(_16429_),
    .ZN(_16430_));
 AND2_X1 _26154_ (.A1(_16297_),
    .A2(_16314_),
    .ZN(_16431_));
 NAND2_X1 _26155_ (.A1(_16431_),
    .A2(_16426_),
    .ZN(_16432_));
 INV_X1 _26156_ (.A(_16426_),
    .ZN(_16433_));
 OAI211_X2 _26157_ (.A(_16430_),
    .B(_16432_),
    .C1(_16336_),
    .C2(_16433_),
    .ZN(_16434_));
 BUF_X4 _26158_ (.A(_16301_),
    .Z(_16435_));
 CLKBUF_X2 _26159_ (.A(_16426_),
    .Z(_16436_));
 AOI211_X4 _26160_ (.A(_16427_),
    .B(_16434_),
    .C1(_16435_),
    .C2(_16436_),
    .ZN(_16437_));
 AND4_X1 _26161_ (.A1(_16391_),
    .A2(_16418_),
    .A3(_16424_),
    .A4(_16437_),
    .ZN(_16438_));
 INV_X1 _26162_ (.A(_17158_),
    .ZN(_16439_));
 NOR2_X1 _26163_ (.A1(_16439_),
    .A2(_17159_),
    .ZN(_16440_));
 AND2_X1 _26164_ (.A1(_16364_),
    .A2(_16440_),
    .ZN(_16441_));
 BUF_X4 _26165_ (.A(_16441_),
    .Z(_16442_));
 BUF_X2 _26166_ (.A(_16344_),
    .Z(_16443_));
 AND2_X1 _26167_ (.A1(_16442_),
    .A2(_16443_),
    .ZN(_16444_));
 AND2_X2 _26168_ (.A1(_16320_),
    .A2(_16304_),
    .ZN(_16445_));
 AND2_X1 _26169_ (.A1(_16441_),
    .A2(_16445_),
    .ZN(_16446_));
 INV_X1 _26170_ (.A(_16446_),
    .ZN(_16447_));
 AND2_X1 _26171_ (.A1(_16320_),
    .A2(_16323_),
    .ZN(_16448_));
 BUF_X2 _26172_ (.A(_16448_),
    .Z(_16449_));
 AND2_X1 _26173_ (.A1(_16441_),
    .A2(_16449_),
    .ZN(_16450_));
 INV_X1 _26174_ (.A(_16450_),
    .ZN(_16451_));
 NAND2_X1 _26175_ (.A1(_16442_),
    .A2(_16390_),
    .ZN(_16452_));
 NAND3_X1 _26176_ (.A1(_16447_),
    .A2(_16451_),
    .A3(_16452_),
    .ZN(_16453_));
 BUF_X2 _26177_ (.A(_16431_),
    .Z(_16454_));
 NAND2_X1 _26178_ (.A1(_16442_),
    .A2(_16454_),
    .ZN(_16455_));
 NAND2_X1 _26179_ (.A1(_16442_),
    .A2(_16383_),
    .ZN(_16456_));
 NAND2_X1 _26180_ (.A1(_16455_),
    .A2(_16456_),
    .ZN(_16457_));
 BUF_X2 _26181_ (.A(_16440_),
    .Z(_16458_));
 NAND4_X1 _26182_ (.A1(_16301_),
    .A2(_16371_),
    .A3(_16458_),
    .A4(_16388_),
    .ZN(_16459_));
 INV_X1 _26183_ (.A(_16441_),
    .ZN(_16460_));
 OAI21_X1 _26184_ (.A(_16459_),
    .B1(_16460_),
    .B2(_16403_),
    .ZN(_16461_));
 OR4_X1 _26185_ (.A1(_16444_),
    .A2(_16453_),
    .A3(_16457_),
    .A4(_16461_),
    .ZN(_16462_));
 BUF_X2 _26186_ (.A(_16329_),
    .Z(_16463_));
 AND2_X2 _26187_ (.A1(_16458_),
    .A2(_16463_),
    .ZN(_16464_));
 AND2_X1 _26188_ (.A1(_16345_),
    .A2(_16388_),
    .ZN(_16465_));
 BUF_X2 _26189_ (.A(_16465_),
    .Z(_16466_));
 OAI21_X1 _26190_ (.A(_16464_),
    .B1(_16443_),
    .B2(_16466_),
    .ZN(_16467_));
 NAND4_X1 _26191_ (.A1(_16301_),
    .A2(_16458_),
    .A3(_11049_),
    .A4(_16463_),
    .ZN(_16468_));
 AND2_X1 _26192_ (.A1(_16467_),
    .A2(_16468_),
    .ZN(_16469_));
 BUF_X4 _26193_ (.A(_16464_),
    .Z(_16470_));
 NAND2_X1 _26194_ (.A1(_16428_),
    .A2(_16470_),
    .ZN(_16471_));
 AND2_X2 _26195_ (.A1(_16314_),
    .A2(_16303_),
    .ZN(_16472_));
 INV_X1 _26196_ (.A(_16472_),
    .ZN(_16473_));
 INV_X1 _26197_ (.A(_16464_),
    .ZN(_16474_));
 OAI211_X2 _26198_ (.A(_16469_),
    .B(_16471_),
    .C1(_16473_),
    .C2(_16474_),
    .ZN(_16475_));
 AND2_X1 _26199_ (.A1(_16308_),
    .A2(_16440_),
    .ZN(_16476_));
 BUF_X2 _26200_ (.A(_16476_),
    .Z(_16477_));
 AND2_X1 _26201_ (.A1(_16477_),
    .A2(_16382_),
    .ZN(_16478_));
 AND2_X1 _26202_ (.A1(_16477_),
    .A2(_16472_),
    .ZN(_16479_));
 NOR2_X1 _26203_ (.A1(_16478_),
    .A2(_16479_),
    .ZN(_16480_));
 BUF_X4 _26204_ (.A(_16477_),
    .Z(_16481_));
 NAND2_X1 _26205_ (.A1(_16481_),
    .A2(_16328_),
    .ZN(_16482_));
 AND2_X1 _26206_ (.A1(_16345_),
    .A2(_16323_),
    .ZN(_16483_));
 BUF_X4 _26207_ (.A(_16483_),
    .Z(_16484_));
 OAI21_X1 _26208_ (.A(_16481_),
    .B1(_16412_),
    .B2(_16484_),
    .ZN(_16485_));
 NAND3_X1 _26209_ (.A1(_16480_),
    .A2(_16482_),
    .A3(_16485_),
    .ZN(_16486_));
 BUF_X2 _26210_ (.A(_16351_),
    .Z(_16487_));
 AND2_X2 _26211_ (.A1(_16458_),
    .A2(_16487_),
    .ZN(_16488_));
 INV_X1 _26212_ (.A(_16488_),
    .ZN(_16489_));
 INV_X1 _26213_ (.A(_16344_),
    .ZN(_16490_));
 AOI21_X1 _26214_ (.A(_16489_),
    .B1(_16490_),
    .B2(_16403_),
    .ZN(_16491_));
 BUF_X2 _26215_ (.A(_16346_),
    .Z(_16492_));
 AND2_X1 _26216_ (.A1(_16492_),
    .A2(_16488_),
    .ZN(_16493_));
 NOR2_X1 _26217_ (.A1(_16491_),
    .A2(_16493_),
    .ZN(_16494_));
 NAND3_X1 _26218_ (.A1(_16472_),
    .A2(_16487_),
    .A3(_16458_),
    .ZN(_16495_));
 BUF_X2 _26219_ (.A(_16488_),
    .Z(_16496_));
 NAND2_X1 _26220_ (.A1(_16496_),
    .A2(_16383_),
    .ZN(_16497_));
 AND2_X2 _26221_ (.A1(_16321_),
    .A2(_17151_),
    .ZN(_16498_));
 NAND2_X1 _26222_ (.A1(_16498_),
    .A2(_16496_),
    .ZN(_16499_));
 NAND4_X1 _26223_ (.A1(_16494_),
    .A2(_16495_),
    .A3(_16497_),
    .A4(_16499_),
    .ZN(_16500_));
 NOR4_X1 _26224_ (.A1(_16462_),
    .A2(_16475_),
    .A3(_16486_),
    .A4(_16500_),
    .ZN(_16501_));
 AND2_X2 _26225_ (.A1(_16439_),
    .A2(_17159_),
    .ZN(_16502_));
 AND2_X2 _26226_ (.A1(_16502_),
    .A2(_16329_),
    .ZN(_16503_));
 INV_X1 _26227_ (.A(_16503_),
    .ZN(_16504_));
 OR2_X1 _26228_ (.A1(_16347_),
    .A2(_16504_),
    .ZN(_16505_));
 AND2_X1 _26229_ (.A1(_16503_),
    .A2(_16483_),
    .ZN(_16506_));
 INV_X1 _26230_ (.A(_16506_),
    .ZN(_16507_));
 NAND2_X1 _26231_ (.A1(_16505_),
    .A2(_16507_),
    .ZN(_16508_));
 BUF_X2 _26232_ (.A(_16503_),
    .Z(_16509_));
 AOI21_X1 _26233_ (.A(_16508_),
    .B1(_16412_),
    .B2(_16509_),
    .ZN(_16510_));
 INV_X1 _26234_ (.A(_16320_),
    .ZN(_16511_));
 NOR2_X1 _26235_ (.A1(_16511_),
    .A2(_16304_),
    .ZN(_16512_));
 NAND2_X1 _26236_ (.A1(_16512_),
    .A2(_16503_),
    .ZN(_16513_));
 AND2_X1 _26237_ (.A1(_16308_),
    .A2(_16502_),
    .ZN(_16514_));
 BUF_X2 _26238_ (.A(_16514_),
    .Z(_16515_));
 NOR3_X1 _26239_ (.A1(_16323_),
    .A2(_17153_),
    .A3(_17154_),
    .ZN(_16516_));
 AND3_X1 _26240_ (.A1(_16515_),
    .A2(_16319_),
    .A3(_16516_),
    .ZN(_16517_));
 BUF_X2 _26241_ (.A(_16373_),
    .Z(_16518_));
 AOI21_X1 _26242_ (.A(_16517_),
    .B1(_16518_),
    .B2(_16515_),
    .ZN(_16519_));
 BUF_X4 _26243_ (.A(_16502_),
    .Z(_16520_));
 BUF_X4 _26244_ (.A(_16520_),
    .Z(_16521_));
 BUF_X4 _26245_ (.A(_16296_),
    .Z(_16522_));
 NAND4_X1 _26246_ (.A1(_16521_),
    .A2(_16522_),
    .A3(_16357_),
    .A4(_16463_),
    .ZN(_16523_));
 NAND4_X1 _26247_ (.A1(_16510_),
    .A2(_16513_),
    .A3(_16519_),
    .A4(_16523_),
    .ZN(_16524_));
 AND3_X1 _26248_ (.A1(_16428_),
    .A2(_16371_),
    .A3(_16520_),
    .ZN(_16525_));
 AND2_X1 _26249_ (.A1(_16502_),
    .A2(_16364_),
    .ZN(_16526_));
 BUF_X2 _26250_ (.A(_16526_),
    .Z(_16527_));
 OAI21_X1 _26251_ (.A(_16527_),
    .B1(_16484_),
    .B2(_16466_),
    .ZN(_16528_));
 INV_X1 _26252_ (.A(_16527_),
    .ZN(_16529_));
 AND2_X2 _26253_ (.A1(_16297_),
    .A2(_16300_),
    .ZN(_16530_));
 INV_X1 _26254_ (.A(_16530_),
    .ZN(_16531_));
 OAI21_X1 _26255_ (.A(_16528_),
    .B1(_16529_),
    .B2(_16531_),
    .ZN(_16532_));
 AND2_X2 _26256_ (.A1(_16502_),
    .A2(_16351_),
    .ZN(_16533_));
 BUF_X4 _26257_ (.A(_16533_),
    .Z(_16534_));
 AND2_X1 _26258_ (.A1(_16512_),
    .A2(_16534_),
    .ZN(_16535_));
 AND2_X1 _26259_ (.A1(_16534_),
    .A2(_16370_),
    .ZN(_16536_));
 INV_X1 _26260_ (.A(_16314_),
    .ZN(_16537_));
 NOR2_X1 _26261_ (.A1(_16537_),
    .A2(_16298_),
    .ZN(_16538_));
 AND2_X1 _26262_ (.A1(_16534_),
    .A2(_16538_),
    .ZN(_16539_));
 OR3_X1 _26263_ (.A1(_16535_),
    .A2(_16536_),
    .A3(_16539_),
    .ZN(_16540_));
 NOR4_X1 _26264_ (.A1(_16524_),
    .A2(_16525_),
    .A3(_16532_),
    .A4(_16540_),
    .ZN(_16541_));
 AND4_X1 _26265_ (.A1(_16378_),
    .A2(_16438_),
    .A3(_16501_),
    .A4(_16541_),
    .ZN(_16542_));
 OAI21_X1 _26266_ (.A(_11076_),
    .B1(_16319_),
    .B2(_17153_),
    .ZN(_16543_));
 AND3_X1 _26267_ (.A1(_16463_),
    .A2(_16330_),
    .A3(_11076_),
    .ZN(_16544_));
 AND2_X1 _26268_ (.A1(_16543_),
    .A2(_16544_),
    .ZN(_16545_));
 INV_X1 _26269_ (.A(_16545_),
    .ZN(_16546_));
 NAND2_X1 _26270_ (.A1(_16542_),
    .A2(_16546_),
    .ZN(_16547_));
 XNOR2_X1 _26271_ (.A(_01014_),
    .B(_01013_),
    .ZN(_16548_));
 XNOR2_X1 _26272_ (.A(_16547_),
    .B(_16548_),
    .ZN(_16549_));
 MUX2_X1 _26273_ (.A(_01225_),
    .B(_16549_),
    .S(_16178_),
    .Z(_01074_));
 BUF_X2 _26274_ (.A(_16406_),
    .Z(_16550_));
 NAND2_X1 _26275_ (.A1(_16515_),
    .A2(_16550_),
    .ZN(_16551_));
 NAND4_X1 _26276_ (.A1(_16520_),
    .A2(_16357_),
    .A3(_16304_),
    .A4(_16463_),
    .ZN(_16552_));
 NAND2_X1 _26277_ (.A1(_16513_),
    .A2(_16552_),
    .ZN(_16553_));
 NOR2_X1 _26278_ (.A1(_16399_),
    .A2(_16530_),
    .ZN(_16554_));
 INV_X1 _26279_ (.A(_16554_),
    .ZN(_16555_));
 AOI211_X4 _26280_ (.A(_16506_),
    .B(_16553_),
    .C1(_16509_),
    .C2(_16555_),
    .ZN(_16556_));
 BUF_X4 _26281_ (.A(_16345_),
    .Z(_16557_));
 AND2_X1 _26282_ (.A1(_16514_),
    .A2(_16557_),
    .ZN(_16558_));
 INV_X1 _26283_ (.A(_16558_),
    .ZN(_16559_));
 OAI21_X1 _26284_ (.A(_16515_),
    .B1(_16397_),
    .B2(_16390_),
    .ZN(_16560_));
 AND4_X1 _26285_ (.A1(_16551_),
    .A2(_16556_),
    .A3(_16559_),
    .A4(_16560_),
    .ZN(_16561_));
 BUF_X4 _26286_ (.A(_16393_),
    .Z(_16562_));
 AND2_X2 _26287_ (.A1(_16314_),
    .A2(_11049_),
    .ZN(_16563_));
 OAI21_X1 _26288_ (.A(_16562_),
    .B1(_16368_),
    .B2(_16563_),
    .ZN(_16564_));
 AND2_X1 _26289_ (.A1(_16393_),
    .A2(_16399_),
    .ZN(_16565_));
 AND2_X1 _26290_ (.A1(_16393_),
    .A2(_16373_),
    .ZN(_16566_));
 AOI221_X4 _26291_ (.A(_16565_),
    .B1(_16393_),
    .B2(_16370_),
    .C1(_11049_),
    .C2(_16566_),
    .ZN(_16567_));
 AND2_X1 _26292_ (.A1(_16382_),
    .A2(_16408_),
    .ZN(_16568_));
 AND2_X1 _26293_ (.A1(_16409_),
    .A2(_16472_),
    .ZN(_16569_));
 AOI221_X4 _26294_ (.A(_16568_),
    .B1(_16498_),
    .B2(_16409_),
    .C1(_16296_),
    .C2(_16569_),
    .ZN(_16570_));
 AND2_X1 _26295_ (.A1(_16373_),
    .A2(_16409_),
    .ZN(_16571_));
 AND2_X1 _26296_ (.A1(_16402_),
    .A2(_16409_),
    .ZN(_16572_));
 AOI211_X4 _26297_ (.A(_16571_),
    .B(_16572_),
    .C1(_16409_),
    .C2(_16370_),
    .ZN(_16573_));
 AND4_X1 _26298_ (.A1(_16564_),
    .A2(_16567_),
    .A3(_16570_),
    .A4(_16573_),
    .ZN(_16574_));
 AND2_X1 _26299_ (.A1(_16526_),
    .A2(_16431_),
    .ZN(_16575_));
 INV_X1 _26300_ (.A(_16575_),
    .ZN(_16576_));
 NAND3_X1 _26301_ (.A1(_16395_),
    .A2(_16371_),
    .A3(_16520_),
    .ZN(_16577_));
 OAI211_X2 _26302_ (.A(_16576_),
    .B(_16577_),
    .C1(_16336_),
    .C2(_16529_),
    .ZN(_16578_));
 INV_X1 _26303_ (.A(_16533_),
    .ZN(_16579_));
 INV_X1 _26304_ (.A(_16328_),
    .ZN(_16580_));
 AOI211_X4 _26305_ (.A(_11049_),
    .B(_16579_),
    .C1(_16537_),
    .C2(_16580_),
    .ZN(_16581_));
 NAND2_X1 _26306_ (.A1(_16527_),
    .A2(_16406_),
    .ZN(_16582_));
 BUF_X2 _26307_ (.A(_16402_),
    .Z(_16583_));
 NAND2_X1 _26308_ (.A1(_16527_),
    .A2(_16583_),
    .ZN(_16584_));
 NAND2_X1 _26309_ (.A1(_16582_),
    .A2(_16584_),
    .ZN(_16585_));
 NAND2_X1 _26310_ (.A1(_16534_),
    .A2(_16443_),
    .ZN(_16586_));
 NAND4_X1 _26311_ (.A1(_16520_),
    .A2(_11049_),
    .A3(_16301_),
    .A4(_16487_),
    .ZN(_16587_));
 INV_X1 _26312_ (.A(_16492_),
    .ZN(_16588_));
 OAI211_X2 _26313_ (.A(_16586_),
    .B(_16587_),
    .C1(_16579_),
    .C2(_16588_),
    .ZN(_16589_));
 NOR4_X1 _26314_ (.A1(_16578_),
    .A2(_16581_),
    .A3(_16585_),
    .A4(_16589_),
    .ZN(_16590_));
 NAND2_X1 _26315_ (.A1(_16445_),
    .A2(_16381_),
    .ZN(_16591_));
 AND2_X1 _26316_ (.A1(_16583_),
    .A2(_16436_),
    .ZN(_16592_));
 AND2_X1 _26317_ (.A1(_16445_),
    .A2(_16426_),
    .ZN(_16593_));
 AND2_X1 _26318_ (.A1(_16389_),
    .A2(_16426_),
    .ZN(_16594_));
 AND2_X1 _26319_ (.A1(_16426_),
    .A2(_16518_),
    .ZN(_16595_));
 NOR4_X1 _26320_ (.A1(_16592_),
    .A2(_16593_),
    .A3(_16594_),
    .A4(_16595_),
    .ZN(_16596_));
 OAI211_X2 _26321_ (.A(_16381_),
    .B(_16435_),
    .C1(_16522_),
    .C2(_16388_),
    .ZN(_16597_));
 BUF_X4 _26322_ (.A(_16370_),
    .Z(_16598_));
 OAI21_X1 _26323_ (.A(_16380_),
    .B1(_16484_),
    .B2(_16598_),
    .ZN(_16599_));
 AND4_X1 _26324_ (.A1(_16591_),
    .A2(_16596_),
    .A3(_16597_),
    .A4(_16599_),
    .ZN(_16600_));
 AND4_X1 _26325_ (.A1(_16561_),
    .A2(_16574_),
    .A3(_16590_),
    .A4(_16600_),
    .ZN(_16601_));
 AND2_X1 _26326_ (.A1(_16311_),
    .A2(_16443_),
    .ZN(_16602_));
 INV_X1 _26327_ (.A(_16602_),
    .ZN(_16603_));
 AND2_X1 _26328_ (.A1(_16310_),
    .A2(_16339_),
    .ZN(_16604_));
 INV_X1 _26329_ (.A(_16604_),
    .ZN(_16605_));
 NAND3_X1 _26330_ (.A1(_16472_),
    .A2(_16308_),
    .A3(_16330_),
    .ZN(_16606_));
 AND2_X1 _26331_ (.A1(_16321_),
    .A2(_16296_),
    .ZN(_16607_));
 NAND2_X1 _26332_ (.A1(_16313_),
    .A2(_16607_),
    .ZN(_16608_));
 AND4_X1 _26333_ (.A1(_16603_),
    .A2(_16605_),
    .A3(_16606_),
    .A4(_16608_),
    .ZN(_16609_));
 BUF_X2 _26334_ (.A(_16331_),
    .Z(_16610_));
 NAND2_X1 _26335_ (.A1(_16610_),
    .A2(_16557_),
    .ZN(_16611_));
 NAND2_X1 _26336_ (.A1(_16363_),
    .A2(_16321_),
    .ZN(_16612_));
 INV_X1 _26337_ (.A(_16612_),
    .ZN(_16613_));
 OAI21_X1 _26338_ (.A(_16610_),
    .B1(_16613_),
    .B2(_16315_),
    .ZN(_16614_));
 AND4_X1 _26339_ (.A1(_16341_),
    .A2(_16609_),
    .A3(_16611_),
    .A4(_16614_),
    .ZN(_16615_));
 OAI21_X1 _26340_ (.A(_16367_),
    .B1(_16613_),
    .B2(_16538_),
    .ZN(_16616_));
 BUF_X4 _26341_ (.A(_16353_),
    .Z(_16617_));
 AOI21_X1 _26342_ (.A(_16359_),
    .B1(_16498_),
    .B2(_16617_),
    .ZN(_16618_));
 OAI211_X2 _26343_ (.A(_16617_),
    .B(_16435_),
    .C1(_11050_),
    .C2(_16388_),
    .ZN(_16619_));
 OAI211_X2 _26344_ (.A(_16617_),
    .B(_16557_),
    .C1(_16522_),
    .C2(_16388_),
    .ZN(_16620_));
 AND4_X1 _26345_ (.A1(_16616_),
    .A2(_16618_),
    .A3(_16619_),
    .A4(_16620_),
    .ZN(_16621_));
 NOR2_X1 _26346_ (.A1(_16474_),
    .A2(_16612_),
    .ZN(_16622_));
 INV_X1 _26347_ (.A(_16622_),
    .ZN(_16623_));
 NAND4_X1 _26348_ (.A1(_16458_),
    .A2(_11050_),
    .A3(_16357_),
    .A4(_16463_),
    .ZN(_16624_));
 OAI21_X1 _26349_ (.A(_16464_),
    .B1(_16550_),
    .B2(_16340_),
    .ZN(_16625_));
 OAI211_X2 _26350_ (.A(_16464_),
    .B(_16557_),
    .C1(_16298_),
    .C2(_16305_),
    .ZN(_16626_));
 AND4_X1 _26351_ (.A1(_16623_),
    .A2(_16624_),
    .A3(_16625_),
    .A4(_16626_),
    .ZN(_16627_));
 NOR2_X1 _26352_ (.A1(_16460_),
    .A2(_16358_),
    .ZN(_16628_));
 INV_X1 _26353_ (.A(_16339_),
    .ZN(_16629_));
 AOI21_X1 _26354_ (.A(_16460_),
    .B1(_16490_),
    .B2(_16629_),
    .ZN(_16630_));
 AOI211_X4 _26355_ (.A(_16628_),
    .B(_16630_),
    .C1(_16442_),
    .C2(_16607_),
    .ZN(_16631_));
 NAND2_X1 _26356_ (.A1(_16488_),
    .A2(_16563_),
    .ZN(_16632_));
 NAND4_X1 _26357_ (.A1(_16321_),
    .A2(_16458_),
    .A3(_16487_),
    .A4(_16318_),
    .ZN(_16633_));
 NAND2_X1 _26358_ (.A1(_16632_),
    .A2(_16633_),
    .ZN(_16634_));
 AND2_X1 _26359_ (.A1(_16488_),
    .A2(_16345_),
    .ZN(_16635_));
 AOI221_X4 _26360_ (.A(_16634_),
    .B1(_16635_),
    .B2(_16319_),
    .C1(_16496_),
    .C2(_16555_),
    .ZN(_16636_));
 AND2_X1 _26361_ (.A1(_16477_),
    .A2(_16406_),
    .ZN(_16637_));
 INV_X1 _26362_ (.A(_16637_),
    .ZN(_16638_));
 OAI21_X1 _26363_ (.A(_16477_),
    .B1(_16449_),
    .B2(_16385_),
    .ZN(_16639_));
 BUF_X4 _26364_ (.A(_16308_),
    .Z(_16640_));
 NAND3_X1 _26365_ (.A1(_16399_),
    .A2(_16640_),
    .A3(_16458_),
    .ZN(_16641_));
 OAI21_X1 _26366_ (.A(_16477_),
    .B1(_16484_),
    .B2(_16598_),
    .ZN(_16642_));
 AND4_X1 _26367_ (.A1(_16638_),
    .A2(_16639_),
    .A3(_16641_),
    .A4(_16642_),
    .ZN(_16643_));
 AND4_X1 _26368_ (.A1(_16627_),
    .A2(_16631_),
    .A3(_16636_),
    .A4(_16643_),
    .ZN(_16644_));
 NAND4_X1 _26369_ (.A1(_16601_),
    .A2(_16615_),
    .A3(_16621_),
    .A4(_16644_),
    .ZN(_16645_));
 NOR2_X1 _26370_ (.A1(_16645_),
    .A2(_16545_),
    .ZN(_16646_));
 XOR2_X1 _26371_ (.A(_01016_),
    .B(_01015_),
    .Z(_16647_));
 XNOR2_X1 _26372_ (.A(_16646_),
    .B(_16647_),
    .ZN(_16648_));
 MUX2_X1 _26373_ (.A(_01226_),
    .B(_16648_),
    .S(_16178_),
    .Z(_01075_));
 AND2_X1 _26374_ (.A1(_16340_),
    .A2(_16436_),
    .ZN(_16649_));
 INV_X1 _26375_ (.A(_16304_),
    .ZN(_16650_));
 AND3_X1 _26376_ (.A1(_16538_),
    .A2(_16436_),
    .A3(_16650_),
    .ZN(_16651_));
 AND4_X1 _26377_ (.A1(_11049_),
    .A2(_16379_),
    .A3(_16557_),
    .A4(_16487_),
    .ZN(_16652_));
 OR4_X1 _26378_ (.A1(_16649_),
    .A2(_16651_),
    .A3(_16594_),
    .A4(_16652_),
    .ZN(_16653_));
 AND2_X1 _26379_ (.A1(_16381_),
    .A2(_16328_),
    .ZN(_16654_));
 NOR2_X1 _26380_ (.A1(_16350_),
    .A2(_16304_),
    .ZN(_16655_));
 AND2_X1 _26381_ (.A1(_16655_),
    .A2(_16380_),
    .ZN(_16656_));
 AOI21_X1 _26382_ (.A(_16421_),
    .B1(_16422_),
    .B2(_16531_),
    .ZN(_16657_));
 NOR4_X1 _26383_ (.A1(_16653_),
    .A2(_16654_),
    .A3(_16656_),
    .A4(_16657_),
    .ZN(_16658_));
 NAND2_X1 _26384_ (.A1(_16393_),
    .A2(_16327_),
    .ZN(_16659_));
 NAND2_X1 _26385_ (.A1(_16562_),
    .A2(_16454_),
    .ZN(_16660_));
 NAND2_X1 _26386_ (.A1(_16393_),
    .A2(_16315_),
    .ZN(_16661_));
 AND3_X1 _26387_ (.A1(_16659_),
    .A2(_16660_),
    .A3(_16661_),
    .ZN(_16662_));
 NAND3_X1 _26388_ (.A1(_16598_),
    .A2(_16640_),
    .A3(_16379_),
    .ZN(_16663_));
 INV_X1 _26389_ (.A(_16566_),
    .ZN(_16664_));
 OAI21_X1 _26390_ (.A(_16562_),
    .B1(_16399_),
    .B2(_16530_),
    .ZN(_16665_));
 NAND4_X1 _26391_ (.A1(_16662_),
    .A2(_16663_),
    .A3(_16664_),
    .A4(_16665_),
    .ZN(_16666_));
 NAND3_X1 _26392_ (.A1(_16410_),
    .A2(_16435_),
    .A3(_16319_),
    .ZN(_16667_));
 NAND2_X1 _26393_ (.A1(_16414_),
    .A2(_16667_),
    .ZN(_16668_));
 OAI211_X2 _26394_ (.A(_16410_),
    .B(_16334_),
    .C1(_16298_),
    .C2(_16318_),
    .ZN(_16669_));
 INV_X1 _26395_ (.A(_16409_),
    .ZN(_16670_));
 OAI21_X1 _26396_ (.A(_16669_),
    .B1(_16670_),
    .B2(_16580_),
    .ZN(_16671_));
 INV_X1 _26397_ (.A(_16396_),
    .ZN(_16672_));
 AOI21_X1 _26398_ (.A(_16670_),
    .B1(_16672_),
    .B2(_16384_),
    .ZN(_16673_));
 NOR4_X1 _26399_ (.A1(_16666_),
    .A2(_16668_),
    .A3(_16671_),
    .A4(_16673_),
    .ZN(_16674_));
 AND2_X1 _26400_ (.A1(_16503_),
    .A2(_16339_),
    .ZN(_16675_));
 INV_X1 _26401_ (.A(_16675_),
    .ZN(_16676_));
 NAND3_X1 _26402_ (.A1(_16550_),
    .A2(_16521_),
    .A3(_16463_),
    .ZN(_16677_));
 NAND2_X1 _26403_ (.A1(_16503_),
    .A2(_16465_),
    .ZN(_16678_));
 NAND3_X1 _26404_ (.A1(_16676_),
    .A2(_16677_),
    .A3(_16678_),
    .ZN(_16679_));
 NAND2_X1 _26405_ (.A1(_16515_),
    .A2(_16315_),
    .ZN(_16680_));
 NAND2_X1 _26406_ (.A1(_16515_),
    .A2(_16466_),
    .ZN(_16681_));
 NAND3_X1 _26407_ (.A1(_16583_),
    .A2(_16640_),
    .A3(_16521_),
    .ZN(_16682_));
 NAND4_X1 _26408_ (.A1(_16680_),
    .A2(_16551_),
    .A3(_16681_),
    .A4(_16682_),
    .ZN(_16683_));
 OAI21_X1 _26409_ (.A(_16357_),
    .B1(_11049_),
    .B2(_16388_),
    .ZN(_16684_));
 INV_X1 _26410_ (.A(_16684_),
    .ZN(_16685_));
 AND2_X1 _26411_ (.A1(_16509_),
    .A2(_16685_),
    .ZN(_16686_));
 NAND2_X1 _26412_ (.A1(_16509_),
    .A2(_16428_),
    .ZN(_16687_));
 NAND2_X1 _26413_ (.A1(_16509_),
    .A2(_16395_),
    .ZN(_16688_));
 NAND4_X1 _26414_ (.A1(_16521_),
    .A2(_11056_),
    .A3(_16334_),
    .A4(_16463_),
    .ZN(_16689_));
 NAND3_X1 _26415_ (.A1(_16687_),
    .A2(_16688_),
    .A3(_16689_),
    .ZN(_16690_));
 NOR4_X1 _26416_ (.A1(_16679_),
    .A2(_16683_),
    .A3(_16686_),
    .A4(_16690_),
    .ZN(_16691_));
 AOI211_X4 _26417_ (.A(_16511_),
    .B(_16579_),
    .C1(_11050_),
    .C2(_11056_),
    .ZN(_16692_));
 OAI21_X1 _26418_ (.A(_16527_),
    .B1(_16395_),
    .B2(_16328_),
    .ZN(_16693_));
 NAND2_X1 _26419_ (.A1(_16527_),
    .A2(_16399_),
    .ZN(_16694_));
 OAI211_X2 _26420_ (.A(_16693_),
    .B(_16694_),
    .C1(_16347_),
    .C2(_16529_),
    .ZN(_16695_));
 NAND2_X1 _26421_ (.A1(_16534_),
    .A2(_16598_),
    .ZN(_16696_));
 NAND3_X1 _26422_ (.A1(_16550_),
    .A2(_16521_),
    .A3(_16487_),
    .ZN(_16697_));
 NAND4_X1 _26423_ (.A1(_16521_),
    .A2(_16305_),
    .A3(_16435_),
    .A4(_16487_),
    .ZN(_16698_));
 NAND4_X1 _26424_ (.A1(_16696_),
    .A2(_16586_),
    .A3(_16697_),
    .A4(_16698_),
    .ZN(_16699_));
 NOR4_X1 _26425_ (.A1(_16692_),
    .A2(_16695_),
    .A3(_16539_),
    .A4(_16699_),
    .ZN(_16700_));
 NAND4_X1 _26426_ (.A1(_16658_),
    .A2(_16674_),
    .A3(_16691_),
    .A4(_16700_),
    .ZN(_16701_));
 AND2_X1 _26427_ (.A1(_16366_),
    .A2(_16685_),
    .ZN(_16702_));
 AND2_X1 _26428_ (.A1(_16366_),
    .A2(_16328_),
    .ZN(_16703_));
 AOI211_X4 _26429_ (.A(_16702_),
    .B(_16703_),
    .C1(_16390_),
    .C2(_16366_),
    .ZN(_16704_));
 NAND2_X1 _26430_ (.A1(_16367_),
    .A2(_16550_),
    .ZN(_16705_));
 NAND4_X1 _26431_ (.A1(_16305_),
    .A2(_16435_),
    .A3(_16371_),
    .A4(_16330_),
    .ZN(_16706_));
 NAND4_X1 _26432_ (.A1(_16371_),
    .A2(_16557_),
    .A3(_16323_),
    .A4(_16330_),
    .ZN(_16707_));
 AND3_X1 _26433_ (.A1(_16705_),
    .A2(_16706_),
    .A3(_16707_),
    .ZN(_16708_));
 OAI21_X1 _26434_ (.A(_16617_),
    .B1(_16324_),
    .B2(_16472_),
    .ZN(_16709_));
 OAI21_X1 _26435_ (.A(_16617_),
    .B1(_16360_),
    .B2(_16419_),
    .ZN(_16710_));
 AND4_X1 _26436_ (.A1(_16704_),
    .A2(_16708_),
    .A3(_16709_),
    .A4(_16710_),
    .ZN(_16711_));
 BUF_X4 _26437_ (.A(_16442_),
    .Z(_16712_));
 NAND2_X1 _26438_ (.A1(_16306_),
    .A2(_16712_),
    .ZN(_16713_));
 OAI21_X1 _26439_ (.A(_16712_),
    .B1(_16443_),
    .B2(_16492_),
    .ZN(_16714_));
 OAI21_X1 _26440_ (.A(_16712_),
    .B1(_16395_),
    .B2(_16449_),
    .ZN(_16715_));
 NAND4_X1 _26441_ (.A1(_16713_),
    .A2(_16455_),
    .A3(_16714_),
    .A4(_16715_),
    .ZN(_16716_));
 NAND2_X1 _26442_ (.A1(_16499_),
    .A2(_16497_),
    .ZN(_16717_));
 AND2_X1 _26443_ (.A1(_16406_),
    .A2(_16488_),
    .ZN(_16718_));
 NOR4_X1 _26444_ (.A1(_16716_),
    .A2(_16493_),
    .A3(_16717_),
    .A4(_16718_),
    .ZN(_16719_));
 OAI21_X1 _26445_ (.A(_16470_),
    .B1(_16395_),
    .B2(_16397_),
    .ZN(_16720_));
 OAI21_X1 _26446_ (.A(_16481_),
    .B1(_16395_),
    .B2(_16383_),
    .ZN(_16721_));
 OAI21_X1 _26447_ (.A(_16481_),
    .B1(_16399_),
    .B2(_16419_),
    .ZN(_16722_));
 OAI21_X1 _26448_ (.A(_16470_),
    .B1(_16399_),
    .B2(_16518_),
    .ZN(_16723_));
 AND4_X1 _26449_ (.A1(_16720_),
    .A2(_16721_),
    .A3(_16722_),
    .A4(_16723_),
    .ZN(_16724_));
 NAND3_X1 _26450_ (.A1(_16583_),
    .A2(_16640_),
    .A3(_16330_),
    .ZN(_16725_));
 OAI21_X1 _26451_ (.A(_16311_),
    .B1(_16530_),
    .B2(_16360_),
    .ZN(_16726_));
 OAI21_X1 _26452_ (.A(_16311_),
    .B1(_16445_),
    .B2(_16383_),
    .ZN(_16727_));
 NAND3_X1 _26453_ (.A1(_16466_),
    .A2(_16308_),
    .A3(_16330_),
    .ZN(_16728_));
 AND4_X1 _26454_ (.A1(_16725_),
    .A2(_16726_),
    .A3(_16727_),
    .A4(_16728_),
    .ZN(_16729_));
 NAND3_X1 _26455_ (.A1(_16516_),
    .A2(_16319_),
    .A3(_16610_),
    .ZN(_16730_));
 AND2_X1 _26456_ (.A1(_16655_),
    .A2(_16610_),
    .ZN(_16731_));
 AND3_X1 _26457_ (.A1(_16331_),
    .A2(_16305_),
    .A3(_16301_),
    .ZN(_16732_));
 NOR2_X1 _26458_ (.A1(_16731_),
    .A2(_16732_),
    .ZN(_16733_));
 AND4_X1 _26459_ (.A1(_16333_),
    .A2(_16729_),
    .A3(_16730_),
    .A4(_16733_),
    .ZN(_16734_));
 NAND4_X1 _26460_ (.A1(_16711_),
    .A2(_16719_),
    .A3(_16724_),
    .A4(_16734_),
    .ZN(_16735_));
 NOR2_X1 _26461_ (.A1(_16701_),
    .A2(_16735_),
    .ZN(_16736_));
 XOR2_X1 _26462_ (.A(_01018_),
    .B(_01017_),
    .Z(_16737_));
 XNOR2_X1 _26463_ (.A(_16736_),
    .B(_16737_),
    .ZN(_16738_));
 MUX2_X1 _26464_ (.A(_01227_),
    .B(_16738_),
    .S(_16178_),
    .Z(_01076_));
 OAI21_X1 _26465_ (.A(_16610_),
    .B1(_16324_),
    .B2(_16563_),
    .ZN(_16739_));
 AND2_X1 _26466_ (.A1(_16533_),
    .A2(_16492_),
    .ZN(_16740_));
 AND4_X1 _26467_ (.A1(_16299_),
    .A2(_16533_),
    .A3(_16650_),
    .A4(_16300_),
    .ZN(_16741_));
 AOI211_X2 _26468_ (.A(_16740_),
    .B(_16741_),
    .C1(_16518_),
    .C2(_16534_),
    .ZN(_16742_));
 NAND4_X1 _26469_ (.A1(_16521_),
    .A2(_11050_),
    .A3(_16487_),
    .A4(_16357_),
    .ZN(_16743_));
 OAI211_X2 _26470_ (.A(_16534_),
    .B(_16334_),
    .C1(_16522_),
    .C2(_11056_),
    .ZN(_16744_));
 AND3_X1 _26471_ (.A1(_16742_),
    .A2(_16743_),
    .A3(_16744_),
    .ZN(_16745_));
 AND2_X1 _26472_ (.A1(_16443_),
    .A2(_16331_),
    .ZN(_16746_));
 NOR3_X1 _26473_ (.A1(_16298_),
    .A2(_11068_),
    .A3(_17154_),
    .ZN(_16747_));
 AND2_X1 _26474_ (.A1(_16747_),
    .A2(_16650_),
    .ZN(_16748_));
 AOI221_X4 _26475_ (.A(_16746_),
    .B1(_16583_),
    .B2(_16331_),
    .C1(_16562_),
    .C2(_16748_),
    .ZN(_16749_));
 AND2_X1 _26476_ (.A1(_16300_),
    .A2(_16296_),
    .ZN(_16750_));
 OAI21_X1 _26477_ (.A(_16496_),
    .B1(_16324_),
    .B2(_16750_),
    .ZN(_16751_));
 AND4_X2 _26478_ (.A1(_16739_),
    .A2(_16745_),
    .A3(_16749_),
    .A4(_16751_),
    .ZN(_16752_));
 NAND2_X1 _26479_ (.A1(_16313_),
    .A2(_16390_),
    .ZN(_16753_));
 AOI22_X1 _26480_ (.A1(_16313_),
    .A2(_16598_),
    .B1(_16428_),
    .B2(_16410_),
    .ZN(_16754_));
 NAND2_X1 _26481_ (.A1(_16481_),
    .A2(_16340_),
    .ZN(_01332_));
 NAND2_X1 _26482_ (.A1(_16598_),
    .A2(_16353_),
    .ZN(_01333_));
 AND4_X1 _26483_ (.A1(_16753_),
    .A2(_16754_),
    .A3(_01332_),
    .A4(_01333_),
    .ZN(_01334_));
 AOI21_X1 _26484_ (.A(_16433_),
    .B1(_16531_),
    .B2(_16386_),
    .ZN(_01335_));
 AND2_X1 _26485_ (.A1(_16442_),
    .A2(_16492_),
    .ZN(_01336_));
 NOR4_X1 _26486_ (.A1(_01335_),
    .A2(_01336_),
    .A3(_16493_),
    .A4(_16568_),
    .ZN(_01337_));
 OAI21_X1 _26487_ (.A(_16498_),
    .B1(_16515_),
    .B2(_16366_),
    .ZN(_01338_));
 NAND2_X1 _26488_ (.A1(_16492_),
    .A2(_16366_),
    .ZN(_01339_));
 NAND3_X1 _26489_ (.A1(_16747_),
    .A2(_16650_),
    .A3(_16353_),
    .ZN(_01340_));
 AND4_X1 _26490_ (.A1(_16687_),
    .A2(_01338_),
    .A3(_01339_),
    .A4(_01340_),
    .ZN(_01341_));
 NAND2_X1 _26491_ (.A1(_16454_),
    .A2(_16367_),
    .ZN(_01342_));
 NAND4_X1 _26492_ (.A1(_16518_),
    .A2(_11049_),
    .A3(_16371_),
    .A4(_16520_),
    .ZN(_01343_));
 NAND2_X1 _26493_ (.A1(_16397_),
    .A2(_16381_),
    .ZN(_01344_));
 AND4_X1 _26494_ (.A1(_01342_),
    .A2(_01343_),
    .A3(_01344_),
    .A4(_16497_),
    .ZN(_01345_));
 AND4_X1 _26495_ (.A1(_01334_),
    .A2(_01337_),
    .A3(_01341_),
    .A4(_01345_),
    .ZN(_01346_));
 AND2_X1 _26496_ (.A1(_16390_),
    .A2(_16380_),
    .ZN(_01347_));
 AND2_X1 _26497_ (.A1(_16345_),
    .A2(_16296_),
    .ZN(_01348_));
 AND2_X1 _26498_ (.A1(_16464_),
    .A2(_01348_),
    .ZN(_01349_));
 NOR4_X1 _26499_ (.A1(_16637_),
    .A2(_01347_),
    .A3(_01349_),
    .A4(_16569_),
    .ZN(_01350_));
 AOI221_X4 _26500_ (.A(_16478_),
    .B1(_16315_),
    .B2(_16436_),
    .C1(_16466_),
    .C2(_16410_),
    .ZN(_01351_));
 NAND2_X1 _26501_ (.A1(_16477_),
    .A2(_16557_),
    .ZN(_01352_));
 NAND2_X1 _26502_ (.A1(_16311_),
    .A2(_16538_),
    .ZN(_01353_));
 AND4_X1 _26503_ (.A1(_16680_),
    .A2(_16559_),
    .A3(_01352_),
    .A4(_01353_),
    .ZN(_01354_));
 NAND2_X1 _26504_ (.A1(_16481_),
    .A2(_16498_),
    .ZN(_01355_));
 AOI22_X1 _26505_ (.A1(_16518_),
    .A2(_16442_),
    .B1(_16550_),
    .B2(_16409_),
    .ZN(_01356_));
 AND3_X1 _26506_ (.A1(_16676_),
    .A2(_01355_),
    .A3(_01356_),
    .ZN(_01357_));
 AND4_X1 _26507_ (.A1(_01350_),
    .A2(_01351_),
    .A3(_01354_),
    .A4(_01357_),
    .ZN(_01358_));
 AND2_X1 _26508_ (.A1(_16380_),
    .A2(_16370_),
    .ZN(_01359_));
 NOR4_X1 _26509_ (.A1(_16628_),
    .A2(_16649_),
    .A3(_16427_),
    .A4(_01359_),
    .ZN(_01360_));
 AOI22_X1 _26510_ (.A1(_16413_),
    .A2(_11056_),
    .B1(_16509_),
    .B2(_16685_),
    .ZN(_01361_));
 AND4_X1 _26511_ (.A1(_16623_),
    .A2(_01360_),
    .A3(_16591_),
    .A4(_01361_),
    .ZN(_01362_));
 NAND4_X1 _26512_ (.A1(_16752_),
    .A2(_01346_),
    .A3(_01358_),
    .A4(_01362_),
    .ZN(_01363_));
 AND2_X1 _26513_ (.A1(_16393_),
    .A2(_16583_),
    .ZN(_01364_));
 INV_X1 _26514_ (.A(_01364_),
    .ZN(_01365_));
 OAI21_X1 _26515_ (.A(_16381_),
    .B1(_16454_),
    .B2(_16518_),
    .ZN(_01366_));
 AND3_X1 _26516_ (.A1(_01365_),
    .A2(_16664_),
    .A3(_01366_),
    .ZN(_01367_));
 NAND2_X1 _26517_ (.A1(_16712_),
    .A2(_16412_),
    .ZN(_01368_));
 OAI21_X1 _26518_ (.A(_16470_),
    .B1(_16530_),
    .B2(_16538_),
    .ZN(_01369_));
 AND4_X1 _26519_ (.A1(_16430_),
    .A2(_01367_),
    .A3(_01368_),
    .A4(_01369_),
    .ZN(_01370_));
 AND2_X1 _26520_ (.A1(_16527_),
    .A2(_16449_),
    .ZN(_01371_));
 NOR2_X1 _26521_ (.A1(_01371_),
    .A2(_16525_),
    .ZN(_01372_));
 INV_X1 _26522_ (.A(_16514_),
    .ZN(_01373_));
 OR2_X1 _26523_ (.A1(_16554_),
    .A2(_01373_),
    .ZN(_01374_));
 AND2_X1 _26524_ (.A1(_16583_),
    .A2(_16381_),
    .ZN(_01375_));
 AND2_X1 _26525_ (.A1(_16448_),
    .A2(_16426_),
    .ZN(_01376_));
 NOR2_X1 _26526_ (.A1(_01375_),
    .A2(_01376_),
    .ZN(_01377_));
 NAND2_X1 _26527_ (.A1(_16598_),
    .A2(_16610_),
    .ZN(_01378_));
 AND2_X1 _26528_ (.A1(_16694_),
    .A2(_01378_),
    .ZN(_01379_));
 AND4_X1 _26529_ (.A1(_01372_),
    .A2(_01374_),
    .A3(_01377_),
    .A4(_01379_),
    .ZN(_01380_));
 INV_X1 _26530_ (.A(_16347_),
    .ZN(_01381_));
 AOI22_X1 _26531_ (.A1(_01381_),
    .A2(_16509_),
    .B1(_16313_),
    .B2(_16306_),
    .ZN(_01382_));
 INV_X1 _26532_ (.A(_16395_),
    .ZN(_01383_));
 OAI21_X1 _26533_ (.A(_16660_),
    .B1(_01383_),
    .B2(_16460_),
    .ZN(_01384_));
 AND2_X1 _26534_ (.A1(_16527_),
    .A2(_16315_),
    .ZN(_01385_));
 AND2_X1 _26535_ (.A1(_16550_),
    .A2(_16381_),
    .ZN(_01386_));
 NOR4_X1 _26536_ (.A1(_01384_),
    .A2(_01385_),
    .A3(_01386_),
    .A4(_16571_),
    .ZN(_01387_));
 NAND4_X1 _26537_ (.A1(_01370_),
    .A2(_01380_),
    .A3(_01382_),
    .A4(_01387_),
    .ZN(_01388_));
 NOR2_X2 _26538_ (.A1(_01363_),
    .A2(_01388_),
    .ZN(_01389_));
 XOR2_X1 _26539_ (.A(_01020_),
    .B(_01019_),
    .Z(_01390_));
 XNOR2_X1 _26540_ (.A(_01389_),
    .B(_01390_),
    .ZN(_01391_));
 MUX2_X1 _26541_ (.A(_01228_),
    .B(_01391_),
    .S(_16178_),
    .Z(_01077_));
 OAI21_X1 _26542_ (.A(_16381_),
    .B1(_16454_),
    .B2(_16315_),
    .ZN(_01392_));
 AND2_X1 _26543_ (.A1(_16530_),
    .A2(_16426_),
    .ZN(_01393_));
 AOI221_X4 _26544_ (.A(_01393_),
    .B1(_16557_),
    .B2(_16436_),
    .C1(_16522_),
    .C2(_16594_),
    .ZN(_01394_));
 NAND4_X1 _26545_ (.A1(_16334_),
    .A2(_16371_),
    .A3(_11050_),
    .A4(_16379_),
    .ZN(_01395_));
 OAI21_X1 _26546_ (.A(_16381_),
    .B1(_16550_),
    .B2(_16419_),
    .ZN(_01396_));
 AND4_X1 _26547_ (.A1(_01392_),
    .A2(_01394_),
    .A3(_01395_),
    .A4(_01396_),
    .ZN(_01397_));
 AND2_X1 _26548_ (.A1(_16562_),
    .A2(_16445_),
    .ZN(_01398_));
 INV_X1 _26549_ (.A(_01398_),
    .ZN(_01399_));
 OAI21_X1 _26550_ (.A(_16562_),
    .B1(_16397_),
    .B2(_16472_),
    .ZN(_01400_));
 OAI211_X2 _26551_ (.A(_16562_),
    .B(_16435_),
    .C1(_11050_),
    .C2(_11056_),
    .ZN(_01401_));
 NAND4_X1 _26552_ (.A1(_01399_),
    .A2(_16664_),
    .A3(_01400_),
    .A4(_01401_),
    .ZN(_01402_));
 AND2_X1 _26553_ (.A1(_16607_),
    .A2(_16410_),
    .ZN(_01403_));
 NOR4_X1 _26554_ (.A1(_01402_),
    .A2(_16569_),
    .A3(_16668_),
    .A4(_01403_),
    .ZN(_01404_));
 OAI21_X1 _26555_ (.A(_16515_),
    .B1(_16445_),
    .B2(_16383_),
    .ZN(_01405_));
 NAND2_X1 _26556_ (.A1(_16515_),
    .A2(_16655_),
    .ZN(_01406_));
 OAI211_X2 _26557_ (.A(_01405_),
    .B(_01406_),
    .C1(_16629_),
    .C2(_01373_),
    .ZN(_01407_));
 NOR4_X1 _26558_ (.A1(_16508_),
    .A2(_01407_),
    .A3(_16553_),
    .A4(_16675_),
    .ZN(_01408_));
 INV_X1 _26559_ (.A(_01371_),
    .ZN(_01409_));
 OAI211_X2 _26560_ (.A(_16576_),
    .B(_01409_),
    .C1(_16672_),
    .C2(_16529_),
    .ZN(_01410_));
 AOI21_X1 _26561_ (.A(_16579_),
    .B1(_01383_),
    .B2(_16672_),
    .ZN(_01411_));
 AOI21_X1 _26562_ (.A(_16579_),
    .B1(_16554_),
    .B2(_16588_),
    .ZN(_01412_));
 NOR4_X1 _26563_ (.A1(_01410_),
    .A2(_16532_),
    .A3(_01411_),
    .A4(_01412_),
    .ZN(_01413_));
 NAND4_X1 _26564_ (.A1(_01397_),
    .A2(_01404_),
    .A3(_01408_),
    .A4(_01413_),
    .ZN(_01414_));
 INV_X1 _26565_ (.A(_16479_),
    .ZN(_01415_));
 OAI21_X1 _26566_ (.A(_16481_),
    .B1(_16395_),
    .B2(_16328_),
    .ZN(_01416_));
 AND2_X1 _26567_ (.A1(_01415_),
    .A2(_01416_),
    .ZN(_01417_));
 NAND2_X1 _26568_ (.A1(_16445_),
    .A2(_16470_),
    .ZN(_01418_));
 NAND3_X1 _26569_ (.A1(_16383_),
    .A2(_16463_),
    .A3(_16458_),
    .ZN(_01419_));
 AND3_X1 _26570_ (.A1(_16471_),
    .A2(_01418_),
    .A3(_01419_),
    .ZN(_01420_));
 OAI21_X1 _26571_ (.A(_16481_),
    .B1(_16443_),
    .B2(_16340_),
    .ZN(_01421_));
 AND4_X1 _26572_ (.A1(_16625_),
    .A2(_01417_),
    .A3(_01420_),
    .A4(_01421_),
    .ZN(_01422_));
 NAND2_X1 _26573_ (.A1(_16512_),
    .A2(_16617_),
    .ZN(_01423_));
 INV_X1 _26574_ (.A(_16367_),
    .ZN(_01424_));
 NOR3_X1 _26575_ (.A1(_01424_),
    .A2(_16305_),
    .A3(_16302_),
    .ZN(_01425_));
 AND2_X1 _26576_ (.A1(_16366_),
    .A2(_16466_),
    .ZN(_01426_));
 NOR3_X1 _26577_ (.A1(_01425_),
    .A2(_16374_),
    .A3(_01426_),
    .ZN(_01427_));
 OAI211_X2 _26578_ (.A(_16367_),
    .B(_16363_),
    .C1(_16334_),
    .C2(_16357_),
    .ZN(_01428_));
 OAI21_X1 _26579_ (.A(_16617_),
    .B1(_16530_),
    .B2(_16518_),
    .ZN(_01429_));
 AND4_X1 _26580_ (.A1(_01423_),
    .A2(_01427_),
    .A3(_01428_),
    .A4(_01429_),
    .ZN(_01430_));
 AND2_X1 _26581_ (.A1(_16311_),
    .A2(_16530_),
    .ZN(_01431_));
 INV_X1 _26582_ (.A(_01431_),
    .ZN(_01432_));
 NAND2_X1 _26583_ (.A1(_16313_),
    .A2(_16383_),
    .ZN(_01433_));
 OAI21_X1 _26584_ (.A(_16313_),
    .B1(_16390_),
    .B2(_16449_),
    .ZN(_01434_));
 OAI21_X1 _26585_ (.A(_16313_),
    .B1(_16443_),
    .B2(_16598_),
    .ZN(_01435_));
 NAND4_X1 _26586_ (.A1(_01432_),
    .A2(_01433_),
    .A3(_01434_),
    .A4(_01435_),
    .ZN(_01436_));
 INV_X1 _26587_ (.A(_16454_),
    .ZN(_01437_));
 AOI21_X1 _26588_ (.A(_16337_),
    .B1(_01437_),
    .B2(_16336_),
    .ZN(_01438_));
 AND3_X1 _26589_ (.A1(_16610_),
    .A2(_16334_),
    .A3(_16318_),
    .ZN(_01439_));
 INV_X1 _26590_ (.A(_16360_),
    .ZN(_01440_));
 OAI22_X1 _26591_ (.A1(_01440_),
    .A2(_16337_),
    .B1(_16611_),
    .B2(_16305_),
    .ZN(_01441_));
 NOR4_X1 _26592_ (.A1(_01436_),
    .A2(_01438_),
    .A3(_01439_),
    .A4(_01441_),
    .ZN(_01442_));
 OAI21_X1 _26593_ (.A(_16712_),
    .B1(_16530_),
    .B2(_16583_),
    .ZN(_01443_));
 NAND3_X1 _26594_ (.A1(_16712_),
    .A2(_16538_),
    .A3(_16650_),
    .ZN(_01444_));
 OAI211_X2 _26595_ (.A(_16712_),
    .B(_16557_),
    .C1(_16522_),
    .C2(_16388_),
    .ZN(_01445_));
 NAND4_X1 _26596_ (.A1(_16447_),
    .A2(_01443_),
    .A3(_01444_),
    .A4(_01445_),
    .ZN(_01446_));
 AND2_X1 _26597_ (.A1(_16399_),
    .A2(_16496_),
    .ZN(_01447_));
 OR2_X1 _26598_ (.A1(_16718_),
    .A2(_01447_),
    .ZN(_01448_));
 AOI21_X1 _26599_ (.A(_16489_),
    .B1(_16511_),
    .B2(_16386_),
    .ZN(_01449_));
 NOR4_X1 _26600_ (.A1(_01446_),
    .A2(_01448_),
    .A3(_16635_),
    .A4(_01449_),
    .ZN(_01450_));
 NAND4_X1 _26601_ (.A1(_01422_),
    .A2(_01430_),
    .A3(_01442_),
    .A4(_01450_),
    .ZN(_01451_));
 NOR2_X1 _26602_ (.A1(_01414_),
    .A2(_01451_),
    .ZN(_01452_));
 XOR2_X1 _26603_ (.A(_01022_),
    .B(_01021_),
    .Z(_01453_));
 XNOR2_X1 _26604_ (.A(_01452_),
    .B(_01453_),
    .ZN(_01454_));
 MUX2_X1 _26605_ (.A(_01229_),
    .B(_01454_),
    .S(_16178_),
    .Z(_01078_));
 OAI21_X1 _26606_ (.A(_16367_),
    .B1(_01348_),
    .B2(_16435_),
    .ZN(_01455_));
 AOI21_X1 _26607_ (.A(_01438_),
    .B1(_16610_),
    .B2(_16613_),
    .ZN(_01456_));
 AND2_X1 _26608_ (.A1(_16310_),
    .A2(_16360_),
    .ZN(_01457_));
 AOI211_X2 _26609_ (.A(_01457_),
    .B(_16604_),
    .C1(_01381_),
    .C2(_16311_),
    .ZN(_01458_));
 OAI221_X1 _26610_ (.A(_16610_),
    .B1(_16522_),
    .B2(_11056_),
    .C1(_16435_),
    .C2(_16557_),
    .ZN(_01459_));
 OAI21_X1 _26611_ (.A(_16313_),
    .B1(_16748_),
    .B2(_16383_),
    .ZN(_01460_));
 AND4_X1 _26612_ (.A1(_01456_),
    .A2(_01458_),
    .A3(_01459_),
    .A4(_01460_),
    .ZN(_01461_));
 OAI21_X1 _26613_ (.A(_16367_),
    .B1(_16613_),
    .B2(_16685_),
    .ZN(_01462_));
 OAI21_X1 _26614_ (.A(_16353_),
    .B1(_16518_),
    .B2(_16466_),
    .ZN(_01463_));
 NAND2_X1 _26615_ (.A1(_16397_),
    .A2(_16353_),
    .ZN(_01464_));
 NAND2_X1 _26616_ (.A1(_16583_),
    .A2(_16353_),
    .ZN(_01465_));
 AND3_X1 _26617_ (.A1(_01463_),
    .A2(_01464_),
    .A3(_01465_),
    .ZN(_01466_));
 AND4_X2 _26618_ (.A1(_01455_),
    .A2(_01461_),
    .A3(_01462_),
    .A4(_01466_),
    .ZN(_01467_));
 OAI21_X1 _26619_ (.A(_16496_),
    .B1(_16454_),
    .B2(_16328_),
    .ZN(_01468_));
 AND3_X1 _26620_ (.A1(_16445_),
    .A2(_16308_),
    .A3(_16458_),
    .ZN(_01469_));
 AOI211_X4 _26621_ (.A(_01469_),
    .B(_16478_),
    .C1(_16390_),
    .C2(_16477_),
    .ZN(_01470_));
 OAI21_X1 _26622_ (.A(_16470_),
    .B1(_16397_),
    .B2(_16498_),
    .ZN(_01471_));
 OAI21_X1 _26623_ (.A(_16477_),
    .B1(_16360_),
    .B2(_16340_),
    .ZN(_01472_));
 AND4_X1 _26624_ (.A1(_16469_),
    .A2(_01470_),
    .A3(_01471_),
    .A4(_01472_),
    .ZN(_01473_));
 NAND2_X1 _26625_ (.A1(_16442_),
    .A2(_16315_),
    .ZN(_01474_));
 OAI21_X1 _26626_ (.A(_16442_),
    .B1(_16412_),
    .B2(_16419_),
    .ZN(_01475_));
 AND4_X1 _26627_ (.A1(_01474_),
    .A2(_16447_),
    .A3(_16455_),
    .A4(_01475_),
    .ZN(_01476_));
 AND2_X1 _26628_ (.A1(_16583_),
    .A2(_16488_),
    .ZN(_01477_));
 AOI211_X4 _26629_ (.A(_01477_),
    .B(_16718_),
    .C1(_01381_),
    .C2(_16496_),
    .ZN(_01478_));
 AND4_X1 _26630_ (.A1(_01468_),
    .A2(_01473_),
    .A3(_01476_),
    .A4(_01478_),
    .ZN(_01479_));
 NAND2_X1 _26631_ (.A1(_16515_),
    .A2(_16390_),
    .ZN(_01480_));
 NAND2_X1 _26632_ (.A1(_16509_),
    .A2(_16383_),
    .ZN(_01481_));
 NAND4_X1 _26633_ (.A1(_16520_),
    .A2(_16298_),
    .A3(_16301_),
    .A4(_16463_),
    .ZN(_01482_));
 OAI21_X1 _26634_ (.A(_16503_),
    .B1(_16483_),
    .B2(_16370_),
    .ZN(_01483_));
 AND4_X1 _26635_ (.A1(_01481_),
    .A2(_16676_),
    .A3(_01482_),
    .A4(_01483_),
    .ZN(_01484_));
 NAND3_X1 _26636_ (.A1(_16385_),
    .A2(_16640_),
    .A3(_16521_),
    .ZN(_01485_));
 AND4_X1 _26637_ (.A1(_01480_),
    .A2(_01484_),
    .A3(_01374_),
    .A4(_01485_),
    .ZN(_01486_));
 NAND2_X1 _26638_ (.A1(_16526_),
    .A2(_16445_),
    .ZN(_01487_));
 NAND3_X1 _26639_ (.A1(_16397_),
    .A2(_16371_),
    .A3(_16520_),
    .ZN(_01488_));
 AND3_X1 _26640_ (.A1(_16385_),
    .A2(_16371_),
    .A3(_16520_),
    .ZN(_01489_));
 INV_X1 _26641_ (.A(_01489_),
    .ZN(_01490_));
 AND4_X1 _26642_ (.A1(_16576_),
    .A2(_01487_),
    .A3(_01488_),
    .A4(_01490_),
    .ZN(_01491_));
 OAI21_X1 _26643_ (.A(_16527_),
    .B1(_16443_),
    .B2(_16484_),
    .ZN(_01492_));
 AND4_X1 _26644_ (.A1(_16584_),
    .A2(_01491_),
    .A3(_16694_),
    .A4(_01492_),
    .ZN(_01493_));
 OAI21_X1 _26645_ (.A(_16534_),
    .B1(_16449_),
    .B2(_16538_),
    .ZN(_01494_));
 NAND2_X1 _26646_ (.A1(_16534_),
    .A2(_16360_),
    .ZN(_01495_));
 NAND2_X1 _26647_ (.A1(_16534_),
    .A2(_16466_),
    .ZN(_01496_));
 NAND3_X1 _26648_ (.A1(_16340_),
    .A2(_16520_),
    .A3(_16487_),
    .ZN(_01497_));
 AND4_X1 _26649_ (.A1(_16586_),
    .A2(_01495_),
    .A3(_01496_),
    .A4(_01497_),
    .ZN(_01498_));
 AND4_X1 _26650_ (.A1(_01486_),
    .A2(_01493_),
    .A3(_01494_),
    .A4(_01498_),
    .ZN(_01499_));
 AOI211_X4 _26651_ (.A(_16569_),
    .B(_16673_),
    .C1(_16410_),
    .C2(_16324_),
    .ZN(_01500_));
 OAI221_X1 _26652_ (.A(_16661_),
    .B1(_16401_),
    .B2(_16473_),
    .C1(_16659_),
    .C2(_11049_),
    .ZN(_01501_));
 AOI211_X4 _26653_ (.A(_01364_),
    .B(_01501_),
    .C1(_16562_),
    .C2(_16550_),
    .ZN(_01502_));
 OAI21_X1 _26654_ (.A(_16410_),
    .B1(_16492_),
    .B2(_16750_),
    .ZN(_01503_));
 AOI21_X1 _26655_ (.A(_16421_),
    .B1(_16490_),
    .B2(_16403_),
    .ZN(_01504_));
 AND2_X1 _26656_ (.A1(_16380_),
    .A2(_16428_),
    .ZN(_01505_));
 AND2_X1 _26657_ (.A1(_16380_),
    .A2(_16472_),
    .ZN(_01506_));
 OR3_X1 _26658_ (.A1(_01504_),
    .A2(_01505_),
    .A3(_01506_),
    .ZN(_01507_));
 AND2_X1 _26659_ (.A1(_16431_),
    .A2(_16426_),
    .ZN(_01508_));
 OR3_X1 _26660_ (.A1(_01508_),
    .A2(_16594_),
    .A3(_01376_),
    .ZN(_01509_));
 AND3_X1 _26661_ (.A1(_16436_),
    .A2(_16305_),
    .A3(_16301_),
    .ZN(_01510_));
 AND2_X1 _26662_ (.A1(_16436_),
    .A2(_01348_),
    .ZN(_01511_));
 NOR4_X1 _26663_ (.A1(_01507_),
    .A2(_01509_),
    .A3(_01510_),
    .A4(_01511_),
    .ZN(_01512_));
 AND4_X1 _26664_ (.A1(_01500_),
    .A2(_01502_),
    .A3(_01503_),
    .A4(_01512_),
    .ZN(_01513_));
 NAND4_X1 _26665_ (.A1(_01467_),
    .A2(_01479_),
    .A3(_01499_),
    .A4(_01513_),
    .ZN(_01514_));
 NOR2_X2 _26666_ (.A1(_01514_),
    .A2(_16545_),
    .ZN(_01515_));
 XOR2_X1 _26667_ (.A(_01024_),
    .B(_01023_),
    .Z(_01516_));
 XNOR2_X1 _26668_ (.A(_01515_),
    .B(_01516_),
    .ZN(_01517_));
 MUX2_X1 _26669_ (.A(_01230_),
    .B(_01517_),
    .S(_16178_),
    .Z(_01079_));
 AND2_X1 _26670_ (.A1(_16387_),
    .A2(_16503_),
    .ZN(_01518_));
 INV_X1 _26671_ (.A(_16750_),
    .ZN(_01519_));
 OAI211_X2 _26672_ (.A(_16507_),
    .B(_16678_),
    .C1(_16504_),
    .C2(_01519_),
    .ZN(_01520_));
 AOI211_X4 _26673_ (.A(_01518_),
    .B(_01520_),
    .C1(_16509_),
    .C2(_16607_),
    .ZN(_01521_));
 AND4_X1 _26674_ (.A1(_16314_),
    .A2(_16502_),
    .A3(_16323_),
    .A4(_16487_),
    .ZN(_01522_));
 AND2_X1 _26675_ (.A1(_16533_),
    .A2(_16472_),
    .ZN(_01523_));
 AOI211_X2 _26676_ (.A(_01522_),
    .B(_01523_),
    .C1(_16533_),
    .C2(_16324_),
    .ZN(_01524_));
 AND4_X1 _26677_ (.A1(_16697_),
    .A2(_01524_),
    .A3(_01496_),
    .A4(_01497_),
    .ZN(_01525_));
 AND4_X1 _26678_ (.A1(_16680_),
    .A2(_01406_),
    .A3(_16551_),
    .A4(_01485_),
    .ZN(_01526_));
 NOR3_X1 _26679_ (.A1(_01371_),
    .A2(_16525_),
    .A3(_01489_),
    .ZN(_01527_));
 AND4_X1 _26680_ (.A1(_16582_),
    .A2(_01527_),
    .A3(_16584_),
    .A4(_01492_),
    .ZN(_01528_));
 AND4_X1 _26681_ (.A1(_01521_),
    .A2(_01525_),
    .A3(_01526_),
    .A4(_01528_),
    .ZN(_01529_));
 AND2_X1 _26682_ (.A1(_16635_),
    .A2(_16319_),
    .ZN(_01530_));
 AND2_X1 _26683_ (.A1(_16449_),
    .A2(_16496_),
    .ZN(_01531_));
 AND3_X1 _26684_ (.A1(_16488_),
    .A2(_16522_),
    .A3(_16357_),
    .ZN(_01532_));
 OR4_X1 _26685_ (.A1(_01530_),
    .A2(_01447_),
    .A3(_01531_),
    .A4(_01532_),
    .ZN(_01533_));
 AOI21_X1 _26686_ (.A(_16461_),
    .B1(_16712_),
    .B2(_16598_),
    .ZN(_01534_));
 NAND2_X1 _26687_ (.A1(_16712_),
    .A2(_16472_),
    .ZN(_01535_));
 NAND4_X1 _26688_ (.A1(_01534_),
    .A2(_16452_),
    .A3(_16456_),
    .A4(_01535_),
    .ZN(_01536_));
 NAND3_X1 _26689_ (.A1(_16368_),
    .A2(_16363_),
    .A3(_16470_),
    .ZN(_01537_));
 NAND2_X1 _26690_ (.A1(_16492_),
    .A2(_16470_),
    .ZN(_01538_));
 OAI211_X2 _26691_ (.A(_01537_),
    .B(_01538_),
    .C1(_01519_),
    .C2(_16474_),
    .ZN(_01539_));
 NAND4_X1 _26692_ (.A1(_16480_),
    .A2(_16638_),
    .A3(_01355_),
    .A4(_01352_),
    .ZN(_01540_));
 NOR4_X1 _26693_ (.A1(_01533_),
    .A2(_01536_),
    .A3(_01539_),
    .A4(_01540_),
    .ZN(_01541_));
 NAND2_X1 _26694_ (.A1(_16311_),
    .A2(_16484_),
    .ZN(_01542_));
 AND3_X1 _26695_ (.A1(_16603_),
    .A2(_01432_),
    .A3(_01542_),
    .ZN(_01543_));
 OAI211_X2 _26696_ (.A(_01543_),
    .B(_01353_),
    .C1(_16511_),
    .C2(_16317_),
    .ZN(_01544_));
 AND2_X1 _26697_ (.A1(_16353_),
    .A2(_16563_),
    .ZN(_01545_));
 INV_X1 _26698_ (.A(_01545_),
    .ZN(_01546_));
 NAND2_X1 _26699_ (.A1(_16484_),
    .A2(_16617_),
    .ZN(_01547_));
 NAND4_X1 _26700_ (.A1(_01546_),
    .A2(_01547_),
    .A3(_01465_),
    .A4(_01333_),
    .ZN(_01548_));
 OAI21_X1 _26701_ (.A(_16733_),
    .B1(_16337_),
    .B2(_16543_),
    .ZN(_01549_));
 AND2_X1 _26702_ (.A1(_16366_),
    .A2(_16454_),
    .ZN(_01550_));
 AND2_X1 _26703_ (.A1(_16340_),
    .A2(_16366_),
    .ZN(_01551_));
 OR4_X4 _26704_ (.A1(_01550_),
    .A2(_01551_),
    .A3(_16703_),
    .A4(_01426_),
    .ZN(_01552_));
 NOR4_X1 _26705_ (.A1(_01544_),
    .A2(_01548_),
    .A3(_01549_),
    .A4(_01552_),
    .ZN(_01553_));
 OAI21_X1 _26706_ (.A(_16562_),
    .B1(_16492_),
    .B2(_16750_),
    .ZN(_01554_));
 NAND4_X1 _26707_ (.A1(_16538_),
    .A2(_16640_),
    .A3(_16379_),
    .A4(_16650_),
    .ZN(_01555_));
 NAND4_X1 _26708_ (.A1(_16640_),
    .A2(_16334_),
    .A3(_16522_),
    .A4(_16379_),
    .ZN(_01556_));
 AND3_X1 _26709_ (.A1(_01554_),
    .A2(_01555_),
    .A3(_01556_),
    .ZN(_01557_));
 NOR4_X1 _26710_ (.A1(_01375_),
    .A2(_01347_),
    .A3(_16656_),
    .A4(_01506_),
    .ZN(_01558_));
 AOI21_X1 _26711_ (.A(_16433_),
    .B1(_16588_),
    .B2(_01440_),
    .ZN(_01559_));
 AND3_X1 _26712_ (.A1(_16436_),
    .A2(_16321_),
    .A3(_16298_),
    .ZN(_01560_));
 NOR4_X1 _26713_ (.A1(_01559_),
    .A2(_16593_),
    .A3(_01376_),
    .A4(_01560_),
    .ZN(_01561_));
 AND2_X1 _26714_ (.A1(_16406_),
    .A2(_16409_),
    .ZN(_01562_));
 INV_X1 _26715_ (.A(_01562_),
    .ZN(_01563_));
 NAND3_X1 _26716_ (.A1(_16410_),
    .A2(_16305_),
    .A3(_16435_),
    .ZN(_01564_));
 OAI21_X1 _26717_ (.A(_16410_),
    .B1(_16449_),
    .B2(_16454_),
    .ZN(_01565_));
 AND4_X1 _26718_ (.A1(_16415_),
    .A2(_01563_),
    .A3(_01564_),
    .A4(_01565_),
    .ZN(_01566_));
 AND4_X1 _26719_ (.A1(_01557_),
    .A2(_01558_),
    .A3(_01561_),
    .A4(_01566_),
    .ZN(_01567_));
 NAND4_X1 _26720_ (.A1(_01529_),
    .A2(_01541_),
    .A3(_01553_),
    .A4(_01567_),
    .ZN(_01568_));
 NOR2_X2 _26721_ (.A1(_01568_),
    .A2(_16545_),
    .ZN(_01569_));
 XOR2_X1 _26722_ (.A(_01026_),
    .B(_01025_),
    .Z(_01570_));
 XNOR2_X1 _26723_ (.A(_01569_),
    .B(_01570_),
    .ZN(_01571_));
 MUX2_X1 _26724_ (.A(_01231_),
    .B(_01571_),
    .S(_16178_),
    .Z(_01081_));
 AND2_X1 _26725_ (.A1(_16503_),
    .A2(_16394_),
    .ZN(_01572_));
 AOI211_X4 _26726_ (.A(_01572_),
    .B(_01518_),
    .C1(_16550_),
    .C2(_16509_),
    .ZN(_01573_));
 OAI211_X2 _26727_ (.A(_16640_),
    .B(_16521_),
    .C1(_16328_),
    .C2(_16563_),
    .ZN(_01574_));
 OAI211_X2 _26728_ (.A(_16640_),
    .B(_16521_),
    .C1(_16484_),
    .C2(_16598_),
    .ZN(_01575_));
 AND4_X1 _26729_ (.A1(_01374_),
    .A2(_01573_),
    .A3(_01574_),
    .A4(_01575_),
    .ZN(_01576_));
 AND2_X1 _26730_ (.A1(_16516_),
    .A2(_16436_),
    .ZN(_01577_));
 OR4_X1 _26731_ (.A1(_16594_),
    .A2(_01393_),
    .A3(_01577_),
    .A4(_01511_),
    .ZN(_01578_));
 OAI21_X1 _26732_ (.A(_01344_),
    .B1(_16421_),
    .B2(_16473_),
    .ZN(_01579_));
 AOI21_X1 _26733_ (.A(_16421_),
    .B1(_01383_),
    .B2(_16580_),
    .ZN(_01580_));
 OAI21_X1 _26734_ (.A(_16599_),
    .B1(_16302_),
    .B2(_16421_),
    .ZN(_01581_));
 NOR4_X1 _26735_ (.A1(_01578_),
    .A2(_01579_),
    .A3(_01580_),
    .A4(_01581_),
    .ZN(_01582_));
 NAND3_X1 _26736_ (.A1(_16397_),
    .A2(_16640_),
    .A3(_16379_),
    .ZN(_01583_));
 OAI21_X1 _26737_ (.A(_16562_),
    .B1(_16484_),
    .B2(_16466_),
    .ZN(_01584_));
 NAND4_X1 _26738_ (.A1(_01365_),
    .A2(_01399_),
    .A3(_01583_),
    .A4(_01584_),
    .ZN(_01585_));
 AOI211_X4 _26739_ (.A(_16350_),
    .B(_16670_),
    .C1(_16522_),
    .C2(_16388_),
    .ZN(_01586_));
 AOI21_X1 _26740_ (.A(_16670_),
    .B1(_16386_),
    .B2(_16322_),
    .ZN(_01587_));
 NOR4_X1 _26741_ (.A1(_01585_),
    .A2(_01586_),
    .A3(_01562_),
    .A4(_01587_),
    .ZN(_01588_));
 OAI21_X1 _26742_ (.A(_16527_),
    .B1(_16443_),
    .B2(_16466_),
    .ZN(_01589_));
 NAND4_X1 _26743_ (.A1(_01490_),
    .A2(_16582_),
    .A3(_16694_),
    .A4(_01589_),
    .ZN(_01590_));
 NAND2_X1 _26744_ (.A1(_16586_),
    .A2(_01497_),
    .ZN(_01591_));
 NOR4_X1 _26745_ (.A1(_01590_),
    .A2(_01591_),
    .A3(_16535_),
    .A4(_01523_),
    .ZN(_01592_));
 NAND4_X1 _26746_ (.A1(_01576_),
    .A2(_01582_),
    .A3(_01588_),
    .A4(_01592_),
    .ZN(_01593_));
 AND2_X1 _26747_ (.A1(_16477_),
    .A2(_16395_),
    .ZN(_01594_));
 AOI211_X4 _26748_ (.A(_01469_),
    .B(_01594_),
    .C1(_16481_),
    .C2(_16563_),
    .ZN(_01595_));
 OAI21_X1 _26749_ (.A(_16481_),
    .B1(_16555_),
    .B2(_16484_),
    .ZN(_01596_));
 OAI21_X1 _26750_ (.A(_16470_),
    .B1(_16449_),
    .B2(_16454_),
    .ZN(_01597_));
 OAI21_X1 _26751_ (.A(_16470_),
    .B1(_16340_),
    .B2(_16419_),
    .ZN(_01598_));
 AND4_X1 _26752_ (.A1(_01595_),
    .A2(_01596_),
    .A3(_01597_),
    .A4(_01598_),
    .ZN(_01599_));
 OAI21_X1 _26753_ (.A(_16712_),
    .B1(_16530_),
    .B2(_16518_),
    .ZN(_01600_));
 NAND4_X1 _26754_ (.A1(_16451_),
    .A2(_01474_),
    .A3(_01535_),
    .A4(_01600_),
    .ZN(_01601_));
 NAND2_X1 _26755_ (.A1(_16390_),
    .A2(_16496_),
    .ZN(_01602_));
 NAND2_X1 _26756_ (.A1(_16449_),
    .A2(_16496_),
    .ZN(_01603_));
 NAND3_X1 _26757_ (.A1(_01602_),
    .A2(_01603_),
    .A3(_16632_),
    .ZN(_01604_));
 NOR4_X1 _26758_ (.A1(_01601_),
    .A2(_01448_),
    .A3(_01530_),
    .A4(_01604_),
    .ZN(_01605_));
 NAND2_X1 _26759_ (.A1(_16748_),
    .A2(_16313_),
    .ZN(_01606_));
 OAI211_X2 _26760_ (.A(_01606_),
    .B(_16606_),
    .C1(_16672_),
    .C2(_16317_),
    .ZN(_01607_));
 NAND4_X1 _26761_ (.A1(_16605_),
    .A2(_16728_),
    .A3(_16726_),
    .A4(_01542_),
    .ZN(_01608_));
 AND3_X1 _26762_ (.A1(_16747_),
    .A2(_16650_),
    .A3(_16610_),
    .ZN(_01609_));
 AOI211_X4 _26763_ (.A(_16350_),
    .B(_16337_),
    .C1(_11050_),
    .C2(_11056_),
    .ZN(_01610_));
 NOR4_X1 _26764_ (.A1(_01607_),
    .A2(_01608_),
    .A3(_01609_),
    .A4(_01610_),
    .ZN(_01611_));
 OAI21_X1 _26765_ (.A(_16617_),
    .B1(_16340_),
    .B2(_01348_),
    .ZN(_01612_));
 OAI21_X1 _26766_ (.A(_16367_),
    .B1(_16376_),
    .B2(_16492_),
    .ZN(_01613_));
 OAI21_X1 _26767_ (.A(_16367_),
    .B1(_16328_),
    .B2(_16516_),
    .ZN(_01614_));
 OAI211_X2 _26768_ (.A(_16617_),
    .B(_11050_),
    .C1(_16334_),
    .C2(_16357_),
    .ZN(_01615_));
 AND4_X1 _26769_ (.A1(_01612_),
    .A2(_01613_),
    .A3(_01614_),
    .A4(_01615_),
    .ZN(_01616_));
 NAND4_X1 _26770_ (.A1(_01599_),
    .A2(_01605_),
    .A3(_01611_),
    .A4(_01616_),
    .ZN(_01617_));
 NOR2_X1 _26771_ (.A1(_01593_),
    .A2(_01617_),
    .ZN(_01618_));
 XOR2_X1 _26772_ (.A(_01028_),
    .B(_01027_),
    .Z(_01619_));
 XNOR2_X1 _26773_ (.A(_01618_),
    .B(_01619_),
    .ZN(_01620_));
 BUF_X4 _26774_ (.A(_03738_),
    .Z(_01621_));
 MUX2_X1 _26775_ (.A(_01232_),
    .B(_01620_),
    .S(_01621_),
    .Z(_01082_));
 XOR2_X1 _26776_ (.A(_17242_),
    .B(_17077_),
    .Z(_01622_));
 XNOR2_X1 _26777_ (.A(_14014_),
    .B(_12823_),
    .ZN(_01623_));
 XNOR2_X1 _26778_ (.A(_01623_),
    .B(_13275_),
    .ZN(_01624_));
 XNOR2_X1 _26779_ (.A(_01624_),
    .B(_13201_),
    .ZN(_01625_));
 XNOR2_X1 _26780_ (.A(_01625_),
    .B(_17242_),
    .ZN(_01626_));
 MUX2_X1 _26781_ (.A(_01622_),
    .B(_01626_),
    .S(_15306_),
    .Z(_00687_));
 XOR2_X1 _26782_ (.A(_17243_),
    .B(_17078_),
    .Z(_01627_));
 XNOR2_X2 _26783_ (.A(_14014_),
    .B(_12983_),
    .ZN(_01628_));
 XOR2_X1 _26784_ (.A(_13390_),
    .B(_01628_),
    .Z(_01629_));
 XNOR2_X1 _26785_ (.A(_13276_),
    .B(_13621_),
    .ZN(_01630_));
 XNOR2_X1 _26786_ (.A(_01629_),
    .B(_01630_),
    .ZN(_01631_));
 XNOR2_X1 _26787_ (.A(_01631_),
    .B(_17243_),
    .ZN(_01632_));
 MUX2_X1 _26788_ (.A(_01627_),
    .B(_01632_),
    .S(_15306_),
    .Z(_00688_));
 XOR2_X1 _26789_ (.A(_17244_),
    .B(_17079_),
    .Z(_01633_));
 XOR2_X1 _26790_ (.A(_13444_),
    .B(_13903_),
    .Z(_01634_));
 XNOR2_X1 _26791_ (.A(_13622_),
    .B(_01634_),
    .ZN(_01635_));
 XOR2_X1 _26792_ (.A(_01635_),
    .B(_17244_),
    .Z(_01636_));
 MUX2_X1 _26793_ (.A(_01633_),
    .B(_01636_),
    .S(_15306_),
    .Z(_00689_));
 XOR2_X1 _26794_ (.A(_17245_),
    .B(_17080_),
    .Z(_01637_));
 XNOR2_X1 _26795_ (.A(_13685_),
    .B(_13903_),
    .ZN(_01638_));
 XNOR2_X1 _26796_ (.A(_13847_),
    .B(_01638_),
    .ZN(_01639_));
 XNOR2_X1 _26797_ (.A(_01639_),
    .B(_14064_),
    .ZN(_01640_));
 XNOR2_X1 _26798_ (.A(_01640_),
    .B(_17245_),
    .ZN(_01641_));
 MUX2_X1 _26799_ (.A(_01637_),
    .B(_01641_),
    .S(_15306_),
    .Z(_00690_));
 XOR2_X1 _26800_ (.A(_17246_),
    .B(_17081_),
    .Z(_01642_));
 XNOR2_X2 _26801_ (.A(_14064_),
    .B(_13743_),
    .ZN(_01643_));
 XNOR2_X2 _26802_ (.A(_13961_),
    .B(_01643_),
    .ZN(_01644_));
 XNOR2_X1 _26803_ (.A(_01644_),
    .B(_12175_),
    .ZN(_01645_));
 XNOR2_X1 _26804_ (.A(_01645_),
    .B(_17246_),
    .ZN(_01646_));
 MUX2_X1 _26805_ (.A(_01642_),
    .B(_01646_),
    .S(_15306_),
    .Z(_00691_));
 XOR2_X1 _26806_ (.A(_17208_),
    .B(_17176_),
    .Z(_01647_));
 XNOR2_X1 _26807_ (.A(_14296_),
    .B(_01647_),
    .ZN(_01648_));
 MUX2_X1 _26808_ (.A(_01290_),
    .B(_01648_),
    .S(_01621_),
    .Z(_01090_));
 XOR2_X1 _26809_ (.A(_17219_),
    .B(_17187_),
    .Z(_01649_));
 XNOR2_X2 _26810_ (.A(_14400_),
    .B(_01649_),
    .ZN(_01650_));
 MUX2_X1 _26811_ (.A(_01291_),
    .B(_01650_),
    .S(_01621_),
    .Z(_01101_));
 XOR2_X1 _26812_ (.A(_17230_),
    .B(_17198_),
    .Z(_01651_));
 XNOR2_X1 _26813_ (.A(_14484_),
    .B(_01651_),
    .ZN(_01652_));
 MUX2_X1 _26814_ (.A(_01292_),
    .B(_01652_),
    .S(_01621_),
    .Z(_01112_));
 XOR2_X1 _26815_ (.A(_17233_),
    .B(_17201_),
    .Z(_01653_));
 XNOR2_X1 _26816_ (.A(_14560_),
    .B(_01653_),
    .ZN(_01654_));
 MUX2_X1 _26817_ (.A(_01293_),
    .B(_01654_),
    .S(_01621_),
    .Z(_01115_));
 AND2_X1 _26818_ (.A1(_14590_),
    .A2(_14618_),
    .ZN(_01655_));
 XOR2_X1 _26819_ (.A(_17234_),
    .B(_17202_),
    .Z(_01656_));
 XNOR2_X1 _26820_ (.A(_01655_),
    .B(_01656_),
    .ZN(_01657_));
 MUX2_X1 _26821_ (.A(_01294_),
    .B(_01657_),
    .S(_01621_),
    .Z(_01116_));
 XOR2_X1 _26822_ (.A(_17235_),
    .B(_17203_),
    .Z(_01658_));
 XNOR2_X1 _26823_ (.A(_14687_),
    .B(_01658_),
    .ZN(_01659_));
 MUX2_X1 _26824_ (.A(_01295_),
    .B(_01659_),
    .S(_01621_),
    .Z(_01117_));
 XOR2_X1 _26825_ (.A(_17236_),
    .B(_17204_),
    .Z(_01660_));
 XNOR2_X1 _26826_ (.A(_14748_),
    .B(_01660_),
    .ZN(_01661_));
 MUX2_X1 _26827_ (.A(_01297_),
    .B(_01661_),
    .S(_01621_),
    .Z(_01118_));
 XOR2_X1 _26828_ (.A(_17237_),
    .B(_17205_),
    .Z(_01662_));
 XNOR2_X1 _26829_ (.A(_14799_),
    .B(_01662_),
    .ZN(_01663_));
 MUX2_X1 _26830_ (.A(_01298_),
    .B(_01663_),
    .S(_01621_),
    .Z(_01119_));
 XOR2_X1 _26831_ (.A(_17238_),
    .B(_17206_),
    .Z(_01664_));
 XNOR2_X1 _26832_ (.A(_15031_),
    .B(_01664_),
    .ZN(_01665_));
 MUX2_X1 _26833_ (.A(_01299_),
    .B(_01665_),
    .S(_01621_),
    .Z(_01120_));
 NOR2_X1 _26834_ (.A1(_03749_),
    .A2(_01300_),
    .ZN(_01666_));
 XNOR2_X1 _26835_ (.A(_17239_),
    .B(_17207_),
    .ZN(_01667_));
 XNOR2_X1 _26836_ (.A(_15133_),
    .B(_01667_),
    .ZN(_01668_));
 AOI21_X1 _26837_ (.A(_01666_),
    .B1(_01668_),
    .B2(_03749_),
    .ZN(_01121_));
 XOR2_X1 _26838_ (.A(_17209_),
    .B(_17177_),
    .Z(_01669_));
 XNOR2_X1 _26839_ (.A(_15216_),
    .B(_01669_),
    .ZN(_01670_));
 BUF_X4 _26840_ (.A(_03738_),
    .Z(_01671_));
 MUX2_X1 _26841_ (.A(_01301_),
    .B(_01670_),
    .S(_01671_),
    .Z(_01091_));
 XOR2_X1 _26842_ (.A(_17210_),
    .B(_17178_),
    .Z(_01672_));
 XNOR2_X1 _26843_ (.A(_15296_),
    .B(_01672_),
    .ZN(_01673_));
 MUX2_X1 _26844_ (.A(_01302_),
    .B(_01673_),
    .S(_01671_),
    .Z(_01092_));
 XOR2_X1 _26845_ (.A(_17211_),
    .B(_17179_),
    .Z(_01674_));
 XNOR2_X1 _26846_ (.A(_15360_),
    .B(_01674_),
    .ZN(_01675_));
 MUX2_X1 _26847_ (.A(_01303_),
    .B(_01675_),
    .S(_01671_),
    .Z(_01093_));
 XOR2_X1 _26848_ (.A(_17212_),
    .B(_17180_),
    .Z(_01676_));
 XNOR2_X1 _26849_ (.A(_15427_),
    .B(_01676_),
    .ZN(_01677_));
 MUX2_X1 _26850_ (.A(_01304_),
    .B(_01677_),
    .S(_01671_),
    .Z(_01094_));
 XOR2_X1 _26851_ (.A(_17213_),
    .B(_17181_),
    .Z(_01678_));
 XNOR2_X1 _26852_ (.A(_15484_),
    .B(_01678_),
    .ZN(_01679_));
 MUX2_X1 _26853_ (.A(_01305_),
    .B(_01679_),
    .S(_01671_),
    .Z(_01095_));
 XOR2_X1 _26854_ (.A(_17214_),
    .B(_17182_),
    .Z(_01680_));
 XNOR2_X1 _26855_ (.A(_15543_),
    .B(_01680_),
    .ZN(_01681_));
 MUX2_X1 _26856_ (.A(_01306_),
    .B(_01681_),
    .S(_01671_),
    .Z(_01096_));
 XOR2_X1 _26857_ (.A(_17215_),
    .B(_17183_),
    .Z(_01682_));
 XNOR2_X1 _26858_ (.A(_15779_),
    .B(_01682_),
    .ZN(_01683_));
 MUX2_X1 _26859_ (.A(_01308_),
    .B(_01683_),
    .S(_01671_),
    .Z(_01097_));
 NAND2_X1 _26860_ (.A1(_03847_),
    .A2(_01309_),
    .ZN(_01684_));
 XOR2_X1 _26861_ (.A(_17216_),
    .B(_17184_),
    .Z(_01685_));
 XOR2_X1 _26862_ (.A(_15886_),
    .B(_01685_),
    .Z(_01686_));
 OAI21_X1 _26863_ (.A(_01684_),
    .B1(_01686_),
    .B2(_03847_),
    .ZN(_01098_));
 XOR2_X1 _26864_ (.A(_17217_),
    .B(_17185_),
    .Z(_01687_));
 XNOR2_X1 _26865_ (.A(_15969_),
    .B(_01687_),
    .ZN(_01688_));
 MUX2_X1 _26866_ (.A(_01310_),
    .B(_01688_),
    .S(_01671_),
    .Z(_01099_));
 AND2_X1 _26867_ (.A1(_16002_),
    .A2(_16045_),
    .ZN(_01689_));
 XOR2_X1 _26868_ (.A(_17218_),
    .B(_17186_),
    .Z(_01690_));
 XNOR2_X1 _26869_ (.A(_01689_),
    .B(_01690_),
    .ZN(_01691_));
 MUX2_X1 _26870_ (.A(_01311_),
    .B(_01691_),
    .S(_01671_),
    .Z(_01100_));
 XOR2_X1 _26871_ (.A(_17220_),
    .B(_17188_),
    .Z(_01692_));
 XNOR2_X1 _26872_ (.A(_16109_),
    .B(_01692_),
    .ZN(_01693_));
 MUX2_X1 _26873_ (.A(_01312_),
    .B(_01693_),
    .S(_01671_),
    .Z(_01102_));
 NOR2_X1 _26874_ (.A1(_03749_),
    .A2(_01313_),
    .ZN(_01694_));
 XOR2_X1 _26875_ (.A(_17221_),
    .B(_17189_),
    .Z(_01695_));
 XOR2_X1 _26876_ (.A(_16176_),
    .B(_01695_),
    .Z(_01696_));
 AOI21_X1 _26877_ (.A(_01694_),
    .B1(_01696_),
    .B2(_03749_),
    .ZN(_01103_));
 NAND2_X1 _26878_ (.A1(_03847_),
    .A2(_01314_),
    .ZN(_01697_));
 XOR2_X1 _26879_ (.A(_17222_),
    .B(_17190_),
    .Z(_01698_));
 XOR2_X1 _26880_ (.A(_16244_),
    .B(_01698_),
    .Z(_01699_));
 OAI21_X1 _26881_ (.A(_01697_),
    .B1(_01699_),
    .B2(_03847_),
    .ZN(_01104_));
 XOR2_X1 _26882_ (.A(_17223_),
    .B(_17191_),
    .Z(_01700_));
 XNOR2_X1 _26883_ (.A(_16294_),
    .B(_01700_),
    .ZN(_01701_));
 BUF_X4 _26884_ (.A(_03933_),
    .Z(_01702_));
 MUX2_X1 _26885_ (.A(_01315_),
    .B(_01701_),
    .S(_01702_),
    .Z(_01105_));
 XNOR2_X1 _26886_ (.A(_01013_),
    .B(_17192_),
    .ZN(_01703_));
 XNOR2_X1 _26887_ (.A(_01703_),
    .B(_17224_),
    .ZN(_01704_));
 XNOR2_X1 _26888_ (.A(_16547_),
    .B(_01704_),
    .ZN(_01705_));
 MUX2_X1 _26889_ (.A(_01316_),
    .B(_01705_),
    .S(_01702_),
    .Z(_01106_));
 XOR2_X1 _26890_ (.A(_01015_),
    .B(_17193_),
    .Z(_01706_));
 XNOR2_X1 _26891_ (.A(_01706_),
    .B(_17225_),
    .ZN(_01707_));
 XNOR2_X1 _26892_ (.A(_16646_),
    .B(_01707_),
    .ZN(_01708_));
 MUX2_X1 _26893_ (.A(_01317_),
    .B(_01708_),
    .S(_01702_),
    .Z(_01107_));
 XOR2_X1 _26894_ (.A(_01017_),
    .B(_17194_),
    .Z(_01709_));
 XNOR2_X1 _26895_ (.A(_01709_),
    .B(_17226_),
    .ZN(_01710_));
 XNOR2_X1 _26896_ (.A(_16736_),
    .B(_01710_),
    .ZN(_01711_));
 MUX2_X1 _26897_ (.A(_01319_),
    .B(_01711_),
    .S(_01702_),
    .Z(_01108_));
 XNOR2_X1 _26898_ (.A(_01019_),
    .B(_17195_),
    .ZN(_01712_));
 INV_X1 _26899_ (.A(_17227_),
    .ZN(_01713_));
 XNOR2_X1 _26900_ (.A(_01712_),
    .B(_01713_),
    .ZN(_01714_));
 XNOR2_X1 _26901_ (.A(_01389_),
    .B(_01714_),
    .ZN(_01715_));
 MUX2_X1 _26902_ (.A(_01320_),
    .B(_01715_),
    .S(_01702_),
    .Z(_01109_));
 XNOR2_X1 _26903_ (.A(_01021_),
    .B(_17196_),
    .ZN(_01716_));
 INV_X1 _26904_ (.A(_17228_),
    .ZN(_01717_));
 XNOR2_X1 _26905_ (.A(_01716_),
    .B(_01717_),
    .ZN(_01718_));
 XNOR2_X1 _26906_ (.A(_01452_),
    .B(_01718_),
    .ZN(_01719_));
 MUX2_X1 _26907_ (.A(_01321_),
    .B(_01719_),
    .S(_01702_),
    .Z(_01110_));
 XOR2_X1 _26908_ (.A(_01023_),
    .B(_17197_),
    .Z(_01720_));
 XNOR2_X1 _26909_ (.A(_01720_),
    .B(_17229_),
    .ZN(_01721_));
 XNOR2_X1 _26910_ (.A(_01515_),
    .B(_01721_),
    .ZN(_01722_));
 MUX2_X1 _26911_ (.A(_01322_),
    .B(_01722_),
    .S(_01702_),
    .Z(_01111_));
 XOR2_X1 _26912_ (.A(_01025_),
    .B(_17199_),
    .Z(_01723_));
 XNOR2_X1 _26913_ (.A(_01723_),
    .B(_17231_),
    .ZN(_01724_));
 XNOR2_X1 _26914_ (.A(_01569_),
    .B(_01724_),
    .ZN(_01725_));
 MUX2_X1 _26915_ (.A(_01323_),
    .B(_01725_),
    .S(_01702_),
    .Z(_01113_));
 XOR2_X1 _26916_ (.A(_01027_),
    .B(_17200_),
    .Z(_01726_));
 XNOR2_X1 _26917_ (.A(_01726_),
    .B(_17232_),
    .ZN(_01727_));
 XNOR2_X1 _26918_ (.A(_01618_),
    .B(_01727_),
    .ZN(_01728_));
 MUX2_X1 _26919_ (.A(_01324_),
    .B(_01728_),
    .S(_01702_),
    .Z(_01114_));
 XOR2_X1 _26920_ (.A(_17247_),
    .B(_17082_),
    .Z(_01729_));
 XNOR2_X1 _26921_ (.A(_13960_),
    .B(_01029_),
    .ZN(_01730_));
 XOR2_X1 _26922_ (.A(_15300_),
    .B(_01730_),
    .Z(_01731_));
 XOR2_X1 _26923_ (.A(_11857_),
    .B(_12583_),
    .Z(_01732_));
 XNOR2_X1 _26924_ (.A(_01731_),
    .B(_01732_),
    .ZN(_01733_));
 MUX2_X1 _26925_ (.A(_01729_),
    .B(_01733_),
    .S(_15306_),
    .Z(_00652_));
 XOR2_X1 _26926_ (.A(_17248_),
    .B(_17083_),
    .Z(_01734_));
 XNOR2_X1 _26927_ (.A(_12256_),
    .B(_01030_),
    .ZN(_01735_));
 XNOR2_X1 _26928_ (.A(_11387_),
    .B(_13960_),
    .ZN(_01736_));
 XNOR2_X1 _26929_ (.A(_01735_),
    .B(_01736_),
    .ZN(_01737_));
 XNOR2_X1 _26930_ (.A(_15300_),
    .B(_16180_),
    .ZN(_01738_));
 XNOR2_X1 _26931_ (.A(_01737_),
    .B(_01738_),
    .ZN(_01739_));
 MUX2_X1 _26932_ (.A(_01734_),
    .B(_01739_),
    .S(_15306_),
    .Z(_00653_));
 XOR2_X1 _26933_ (.A(_12823_),
    .B(_12661_),
    .Z(_01740_));
 XNOR2_X1 _26934_ (.A(_01740_),
    .B(_13199_),
    .ZN(_01741_));
 XNOR2_X1 _26935_ (.A(_12472_),
    .B(_12357_),
    .ZN(_01742_));
 OAI21_X1 _26936_ (.A(_09098_),
    .B1(_01741_),
    .B2(_01742_),
    .ZN(_01743_));
 AOI21_X1 _26937_ (.A(_01743_),
    .B1(_01741_),
    .B2(_01742_),
    .ZN(_01744_));
 AND2_X1 _26938_ (.A1(_01331_),
    .A2(_17085_),
    .ZN(_01745_));
 NOR2_X1 _26939_ (.A1(_01744_),
    .A2(_01745_),
    .ZN(_01746_));
 XNOR2_X1 _26940_ (.A(_01746_),
    .B(_17249_),
    .ZN(_00654_));
 XOR2_X1 _26941_ (.A(_17250_),
    .B(_17086_),
    .Z(_01747_));
 XNOR2_X1 _26942_ (.A(_13275_),
    .B(_12823_),
    .ZN(_01748_));
 XNOR2_X1 _26943_ (.A(_01748_),
    .B(_01628_),
    .ZN(_01749_));
 XNOR2_X1 _26944_ (.A(_13960_),
    .B(_12736_),
    .ZN(_01750_));
 XOR2_X1 _26945_ (.A(_01750_),
    .B(_13129_),
    .Z(_01751_));
 XNOR2_X1 _26946_ (.A(_01749_),
    .B(_01751_),
    .ZN(_01752_));
 XNOR2_X1 _26947_ (.A(_01752_),
    .B(_17250_),
    .ZN(_01753_));
 MUX2_X1 _26948_ (.A(_01747_),
    .B(_01753_),
    .S(_15306_),
    .Z(_00655_));
 XOR2_X1 _26949_ (.A(_17252_),
    .B(_17087_),
    .Z(_01754_));
 XNOR2_X1 _26950_ (.A(_01628_),
    .B(_13444_),
    .ZN(_01755_));
 XNOR2_X2 _26951_ (.A(_13058_),
    .B(_13960_),
    .ZN(_01756_));
 XOR2_X1 _26952_ (.A(_01756_),
    .B(_13332_),
    .Z(_01757_));
 XNOR2_X1 _26953_ (.A(_01755_),
    .B(_01757_),
    .ZN(_01758_));
 XNOR2_X1 _26954_ (.A(_01758_),
    .B(_13621_),
    .ZN(_01759_));
 INV_X1 _26955_ (.A(_17252_),
    .ZN(_01760_));
 XNOR2_X1 _26956_ (.A(_01759_),
    .B(_01760_),
    .ZN(_01761_));
 BUF_X4 _26957_ (.A(_09099_),
    .Z(_01762_));
 MUX2_X1 _26958_ (.A(_01754_),
    .B(_01761_),
    .S(_01762_),
    .Z(_00656_));
 XOR2_X1 _26959_ (.A(_17253_),
    .B(_17088_),
    .Z(_01763_));
 XNOR2_X1 _26960_ (.A(_01638_),
    .B(_13389_),
    .ZN(_01764_));
 XNOR2_X1 _26961_ (.A(_13444_),
    .B(_01031_),
    .ZN(_01765_));
 XNOR2_X1 _26962_ (.A(_01765_),
    .B(_13508_),
    .ZN(_01766_));
 XNOR2_X1 _26963_ (.A(_01764_),
    .B(_01766_),
    .ZN(_01767_));
 MUX2_X1 _26964_ (.A(_01763_),
    .B(_01767_),
    .S(_01762_),
    .Z(_00657_));
 XOR2_X1 _26965_ (.A(_17254_),
    .B(_17089_),
    .Z(_01768_));
 XNOR2_X1 _26966_ (.A(_13685_),
    .B(_13846_),
    .ZN(_01769_));
 XNOR2_X1 _26967_ (.A(_01769_),
    .B(_14064_),
    .ZN(_01770_));
 XNOR2_X1 _26968_ (.A(_13568_),
    .B(_01032_),
    .ZN(_01771_));
 XOR2_X1 _26969_ (.A(_01771_),
    .B(_13743_),
    .Z(_01772_));
 XNOR2_X1 _26970_ (.A(_01770_),
    .B(_01772_),
    .ZN(_01773_));
 MUX2_X1 _26971_ (.A(_01768_),
    .B(_01773_),
    .S(_01762_),
    .Z(_00658_));
 XOR2_X1 _26972_ (.A(_17255_),
    .B(_17090_),
    .Z(_01774_));
 XOR2_X1 _26973_ (.A(_13743_),
    .B(_11958_),
    .Z(_01775_));
 XNOR2_X1 _26974_ (.A(_14014_),
    .B(_13797_),
    .ZN(_01776_));
 XNOR2_X1 _26975_ (.A(_01775_),
    .B(_01776_),
    .ZN(_01777_));
 XNOR2_X1 _26976_ (.A(_01777_),
    .B(_12175_),
    .ZN(_01778_));
 INV_X1 _26977_ (.A(_17255_),
    .ZN(_01779_));
 XNOR2_X1 _26978_ (.A(_01778_),
    .B(_01779_),
    .ZN(_01780_));
 MUX2_X1 _26979_ (.A(_01774_),
    .B(_01780_),
    .S(_01762_),
    .Z(_00659_));
 XOR2_X1 _26980_ (.A(_01648_),
    .B(_17240_),
    .Z(_01781_));
 MUX2_X1 _26981_ (.A(_01255_),
    .B(_01781_),
    .S(_01702_),
    .Z(_01122_));
 INV_X1 _26982_ (.A(_17251_),
    .ZN(_01782_));
 MUX2_X1 _26983_ (.A(_17251_),
    .B(_01256_),
    .S(_01330_),
    .Z(_01783_));
 NAND2_X1 _26984_ (.A1(_01650_),
    .A2(_03738_),
    .ZN(_01784_));
 MUX2_X1 _26985_ (.A(_01782_),
    .B(_01783_),
    .S(_01784_),
    .Z(_01133_));
 INV_X1 _26986_ (.A(_17262_),
    .ZN(_01785_));
 XNOR2_X1 _26987_ (.A(_01652_),
    .B(_01785_),
    .ZN(_01786_));
 BUF_X4 _26988_ (.A(_03933_),
    .Z(_01787_));
 MUX2_X1 _26989_ (.A(_01257_),
    .B(_01786_),
    .S(_01787_),
    .Z(_01144_));
 BUF_X4 _26990_ (.A(_03933_),
    .Z(_01788_));
 AND3_X1 _26991_ (.A1(_01654_),
    .A2(_01788_),
    .A3(_17265_),
    .ZN(_01789_));
 MUX2_X1 _26992_ (.A(_17265_),
    .B(_01258_),
    .S(_01330_),
    .Z(_01790_));
 AOI21_X1 _26993_ (.A(_01790_),
    .B1(_01654_),
    .B2(_03749_),
    .ZN(_01791_));
 NOR2_X1 _26994_ (.A1(_01789_),
    .A2(_01791_),
    .ZN(_01147_));
 XNOR2_X1 _26995_ (.A(_01656_),
    .B(_17266_),
    .ZN(_01792_));
 XOR2_X1 _26996_ (.A(_01655_),
    .B(_01792_),
    .Z(_01793_));
 MUX2_X1 _26997_ (.A(_01259_),
    .B(_01793_),
    .S(_01787_),
    .Z(_01148_));
 XOR2_X1 _26998_ (.A(_01659_),
    .B(_17267_),
    .Z(_01794_));
 MUX2_X1 _26999_ (.A(_01260_),
    .B(_01794_),
    .S(_01787_),
    .Z(_01149_));
 XOR2_X1 _27000_ (.A(_17268_),
    .B(_17236_),
    .Z(_01795_));
 XOR2_X1 _27001_ (.A(_01795_),
    .B(_17204_),
    .Z(_01796_));
 XNOR2_X1 _27002_ (.A(_14748_),
    .B(_01796_),
    .ZN(_01797_));
 MUX2_X1 _27003_ (.A(_01261_),
    .B(_01797_),
    .S(_01787_),
    .Z(_01150_));
 XNOR2_X1 _27004_ (.A(_01662_),
    .B(_17269_),
    .ZN(_01798_));
 XOR2_X1 _27005_ (.A(_14799_),
    .B(_01798_),
    .Z(_01799_));
 MUX2_X1 _27006_ (.A(_01262_),
    .B(_01799_),
    .S(_01787_),
    .Z(_01151_));
 XNOR2_X1 _27007_ (.A(_01664_),
    .B(_17270_),
    .ZN(_01800_));
 XOR2_X1 _27008_ (.A(_15031_),
    .B(_01800_),
    .Z(_01801_));
 MUX2_X1 _27009_ (.A(_01264_),
    .B(_01801_),
    .S(_01787_),
    .Z(_01152_));
 XNOR2_X1 _27010_ (.A(_01667_),
    .B(_15304_),
    .ZN(_01802_));
 XOR2_X1 _27011_ (.A(_15133_),
    .B(_01802_),
    .Z(_01803_));
 MUX2_X1 _27012_ (.A(_01265_),
    .B(_01803_),
    .S(_01787_),
    .Z(_01153_));
 XOR2_X1 _27013_ (.A(_01670_),
    .B(_17241_),
    .Z(_01804_));
 MUX2_X1 _27014_ (.A(_01266_),
    .B(_01804_),
    .S(_01787_),
    .Z(_01123_));
 XOR2_X1 _27015_ (.A(_01673_),
    .B(_17242_),
    .Z(_01805_));
 MUX2_X1 _27016_ (.A(_01267_),
    .B(_01805_),
    .S(_01787_),
    .Z(_01124_));
 INV_X1 _27017_ (.A(_17243_),
    .ZN(_01806_));
 XNOR2_X1 _27018_ (.A(_01675_),
    .B(_01806_),
    .ZN(_01807_));
 MUX2_X1 _27019_ (.A(_01268_),
    .B(_01807_),
    .S(_01787_),
    .Z(_01125_));
 XOR2_X1 _27020_ (.A(_01677_),
    .B(_17244_),
    .Z(_01808_));
 BUF_X4 _27021_ (.A(_03933_),
    .Z(_01809_));
 MUX2_X1 _27022_ (.A(_01269_),
    .B(_01808_),
    .S(_01809_),
    .Z(_01126_));
 XOR2_X1 _27023_ (.A(_01679_),
    .B(_17245_),
    .Z(_01810_));
 MUX2_X1 _27024_ (.A(_01270_),
    .B(_01810_),
    .S(_01809_),
    .Z(_01127_));
 XOR2_X1 _27025_ (.A(_01681_),
    .B(_17246_),
    .Z(_01811_));
 MUX2_X1 _27026_ (.A(_01271_),
    .B(_01811_),
    .S(_01809_),
    .Z(_01128_));
 XOR2_X1 _27027_ (.A(_17183_),
    .B(_17247_),
    .Z(_01812_));
 XOR2_X1 _27028_ (.A(_01812_),
    .B(_17215_),
    .Z(_01813_));
 XNOR2_X1 _27029_ (.A(_15779_),
    .B(_01813_),
    .ZN(_01814_));
 MUX2_X1 _27030_ (.A(_01272_),
    .B(_01814_),
    .S(_01809_),
    .Z(_01129_));
 XNOR2_X1 _27031_ (.A(_01686_),
    .B(_17248_),
    .ZN(_01815_));
 MUX2_X1 _27032_ (.A(_01273_),
    .B(_01815_),
    .S(_01809_),
    .Z(_01130_));
 XOR2_X1 _27033_ (.A(_17185_),
    .B(_17249_),
    .Z(_01816_));
 XOR2_X1 _27034_ (.A(_01816_),
    .B(_17217_),
    .Z(_01817_));
 XNOR2_X1 _27035_ (.A(_15969_),
    .B(_01817_),
    .ZN(_01818_));
 MUX2_X1 _27036_ (.A(_01275_),
    .B(_01818_),
    .S(_01809_),
    .Z(_01131_));
 XOR2_X1 _27037_ (.A(_17186_),
    .B(_17250_),
    .Z(_01819_));
 INV_X1 _27038_ (.A(_17218_),
    .ZN(_01820_));
 XNOR2_X1 _27039_ (.A(_01819_),
    .B(_01820_),
    .ZN(_01821_));
 XNOR2_X1 _27040_ (.A(_01689_),
    .B(_01821_),
    .ZN(_01822_));
 MUX2_X1 _27041_ (.A(_01276_),
    .B(_01822_),
    .S(_01809_),
    .Z(_01132_));
 MUX2_X1 _27042_ (.A(_17252_),
    .B(_01277_),
    .S(_01330_),
    .Z(_01823_));
 NAND2_X1 _27043_ (.A1(_01693_),
    .A2(_03738_),
    .ZN(_01824_));
 MUX2_X1 _27044_ (.A(_01760_),
    .B(_01823_),
    .S(_01824_),
    .Z(_01134_));
 XNOR2_X1 _27045_ (.A(_01696_),
    .B(_17253_),
    .ZN(_01825_));
 MUX2_X1 _27046_ (.A(_01278_),
    .B(_01825_),
    .S(_01809_),
    .Z(_01135_));
 XNOR2_X1 _27047_ (.A(_01699_),
    .B(_17254_),
    .ZN(_01826_));
 MUX2_X1 _27048_ (.A(_01279_),
    .B(_01826_),
    .S(_01809_),
    .Z(_01136_));
 MUX2_X1 _27049_ (.A(_17255_),
    .B(_01280_),
    .S(_01330_),
    .Z(_01827_));
 NAND2_X1 _27050_ (.A1(_01701_),
    .A2(_03738_),
    .ZN(_01828_));
 MUX2_X1 _27051_ (.A(_01779_),
    .B(_01827_),
    .S(_01828_),
    .Z(_01137_));
 XOR2_X1 _27052_ (.A(_01705_),
    .B(_17256_),
    .Z(_01829_));
 MUX2_X1 _27053_ (.A(_01281_),
    .B(_01829_),
    .S(_01809_),
    .Z(_01138_));
 XOR2_X1 _27054_ (.A(_01708_),
    .B(_17257_),
    .Z(_01830_));
 BUF_X4 _27055_ (.A(_03933_),
    .Z(_01831_));
 MUX2_X1 _27056_ (.A(_01282_),
    .B(_01830_),
    .S(_01831_),
    .Z(_01139_));
 XOR2_X1 _27057_ (.A(_01711_),
    .B(_17258_),
    .Z(_01832_));
 MUX2_X1 _27058_ (.A(_01283_),
    .B(_01832_),
    .S(_01831_),
    .Z(_01140_));
 XOR2_X1 _27059_ (.A(_01715_),
    .B(_17259_),
    .Z(_01833_));
 MUX2_X1 _27060_ (.A(_01284_),
    .B(_01833_),
    .S(_01831_),
    .Z(_01141_));
 XOR2_X1 _27061_ (.A(_01719_),
    .B(_17260_),
    .Z(_01834_));
 MUX2_X1 _27062_ (.A(_01286_),
    .B(_01834_),
    .S(_01831_),
    .Z(_01142_));
 XOR2_X1 _27063_ (.A(_01722_),
    .B(_17261_),
    .Z(_01835_));
 MUX2_X1 _27064_ (.A(_01287_),
    .B(_01835_),
    .S(_01831_),
    .Z(_01143_));
 XOR2_X1 _27065_ (.A(_01725_),
    .B(_17263_),
    .Z(_01836_));
 MUX2_X1 _27066_ (.A(_01288_),
    .B(_01836_),
    .S(_01831_),
    .Z(_01145_));
 XOR2_X1 _27067_ (.A(_01728_),
    .B(_17264_),
    .Z(_01837_));
 MUX2_X1 _27068_ (.A(_01289_),
    .B(_01837_),
    .S(_01831_),
    .Z(_01146_));
 XOR2_X1 _27069_ (.A(_17256_),
    .B(_17091_),
    .Z(_01838_));
 XNOR2_X1 _27070_ (.A(_11625_),
    .B(_13961_),
    .ZN(_01839_));
 XNOR2_X1 _27071_ (.A(_12583_),
    .B(_01033_),
    .ZN(_01840_));
 XNOR2_X1 _27072_ (.A(_01839_),
    .B(_01840_),
    .ZN(_01841_));
 MUX2_X1 _27073_ (.A(_01838_),
    .B(_01841_),
    .S(_01762_),
    .Z(_00620_));
 XOR2_X1 _27074_ (.A(_17257_),
    .B(_17092_),
    .Z(_01842_));
 INV_X1 _27075_ (.A(_01034_),
    .ZN(_01843_));
 XNOR2_X1 _27076_ (.A(_13961_),
    .B(_01843_),
    .ZN(_01844_));
 XNOR2_X1 _27077_ (.A(_01844_),
    .B(_14405_),
    .ZN(_01845_));
 XNOR2_X1 _27078_ (.A(_01742_),
    .B(_12904_),
    .ZN(_01846_));
 XNOR2_X1 _27079_ (.A(_01845_),
    .B(_01846_),
    .ZN(_01847_));
 MUX2_X1 _27080_ (.A(_01842_),
    .B(_01847_),
    .S(_01762_),
    .Z(_00621_));
 XOR2_X1 _27081_ (.A(_17258_),
    .B(_17093_),
    .Z(_01848_));
 XNOR2_X1 _27082_ (.A(_12823_),
    .B(_12736_),
    .ZN(_01849_));
 XNOR2_X1 _27083_ (.A(_12358_),
    .B(_01849_),
    .ZN(_01850_));
 XNOR2_X1 _27084_ (.A(_01850_),
    .B(_13199_),
    .ZN(_01851_));
 XNOR2_X1 _27085_ (.A(_01851_),
    .B(_17258_),
    .ZN(_01852_));
 MUX2_X1 _27086_ (.A(_01848_),
    .B(_01852_),
    .S(_01762_),
    .Z(_00622_));
 XOR2_X1 _27087_ (.A(_17259_),
    .B(_17094_),
    .Z(_01853_));
 XNOR2_X1 _27088_ (.A(_13275_),
    .B(_13058_),
    .ZN(_01854_));
 XNOR2_X1 _27089_ (.A(_01854_),
    .B(_12909_),
    .ZN(_01855_));
 XNOR2_X1 _27090_ (.A(_01750_),
    .B(_12983_),
    .ZN(_01856_));
 XNOR2_X1 _27091_ (.A(_01855_),
    .B(_01856_),
    .ZN(_01857_));
 XNOR2_X1 _27092_ (.A(_01857_),
    .B(_17259_),
    .ZN(_01858_));
 MUX2_X1 _27093_ (.A(_01853_),
    .B(_01858_),
    .S(_01762_),
    .Z(_00623_));
 XOR2_X1 _27094_ (.A(_17260_),
    .B(_17096_),
    .Z(_01859_));
 XNOR2_X2 _27095_ (.A(_13392_),
    .B(_01756_),
    .ZN(_01860_));
 XNOR2_X2 _27096_ (.A(_01860_),
    .B(_13389_),
    .ZN(_01861_));
 XNOR2_X2 _27097_ (.A(_01861_),
    .B(_13444_),
    .ZN(_01862_));
 XNOR2_X2 _27098_ (.A(_01862_),
    .B(_13621_),
    .ZN(_01863_));
 XNOR2_X2 _27099_ (.A(_01863_),
    .B(_17260_),
    .ZN(_01864_));
 MUX2_X2 _27100_ (.A(_01859_),
    .B(_01864_),
    .S(_01762_),
    .Z(_00624_));
 XOR2_X1 _27101_ (.A(_17261_),
    .B(_17097_),
    .Z(_01865_));
 XNOR2_X1 _27102_ (.A(_13685_),
    .B(_13568_),
    .ZN(_01866_));
 INV_X1 _27103_ (.A(_01035_),
    .ZN(_01867_));
 XNOR2_X1 _27104_ (.A(_13903_),
    .B(_01867_),
    .ZN(_01868_));
 XNOR2_X1 _27105_ (.A(_01866_),
    .B(_01868_),
    .ZN(_01869_));
 XOR2_X1 _27106_ (.A(_01869_),
    .B(_13390_),
    .Z(_01870_));
 MUX2_X1 _27107_ (.A(_01865_),
    .B(_01870_),
    .S(_01762_),
    .Z(_00625_));
 XOR2_X1 _27108_ (.A(_17263_),
    .B(_17098_),
    .Z(_01871_));
 XOR2_X1 _27109_ (.A(_14064_),
    .B(_01036_),
    .Z(_01872_));
 XNOR2_X1 _27110_ (.A(_01872_),
    .B(_13569_),
    .ZN(_01873_));
 XOR2_X1 _27111_ (.A(_13797_),
    .B(_13743_),
    .Z(_01874_));
 XNOR2_X1 _27112_ (.A(_01873_),
    .B(_01874_),
    .ZN(_01875_));
 BUF_X4 _27113_ (.A(_09098_),
    .Z(_01876_));
 MUX2_X1 _27114_ (.A(_01871_),
    .B(_01875_),
    .S(_01876_),
    .Z(_00626_));
 XOR2_X1 _27115_ (.A(_17264_),
    .B(_17099_),
    .Z(_01877_));
 XOR2_X1 _27116_ (.A(_14014_),
    .B(_13960_),
    .Z(_01878_));
 XNOR2_X1 _27117_ (.A(_01878_),
    .B(_13847_),
    .ZN(_01879_));
 XNOR2_X1 _27118_ (.A(_01879_),
    .B(_12175_),
    .ZN(_01880_));
 XNOR2_X1 _27119_ (.A(_01880_),
    .B(_17264_),
    .ZN(_01881_));
 MUX2_X1 _27120_ (.A(_01877_),
    .B(_01881_),
    .S(_01876_),
    .Z(_00627_));
 XOR2_X1 _27121_ (.A(_04132_),
    .B(_17240_),
    .Z(_01882_));
 XOR2_X1 _27122_ (.A(_01647_),
    .B(_01882_),
    .Z(_01883_));
 XNOR2_X1 _27123_ (.A(_14296_),
    .B(_01883_),
    .ZN(_01884_));
 MUX2_X1 _27124_ (.A(_01202_),
    .B(_01884_),
    .S(_01831_),
    .Z(_01154_));
 XNOR2_X1 _27125_ (.A(_09101_),
    .B(_17251_),
    .ZN(_01885_));
 XNOR2_X1 _27126_ (.A(_01650_),
    .B(_01885_),
    .ZN(_01886_));
 MUX2_X1 _27127_ (.A(_01241_),
    .B(_01886_),
    .S(_01831_),
    .Z(_01165_));
 XOR2_X1 _27128_ (.A(_17208_),
    .B(_17100_),
    .Z(_01887_));
 AND2_X4 _27129_ (.A1(_16846_),
    .A2(_16847_),
    .ZN(_01888_));
 INV_X1 _27130_ (.A(_01888_),
    .ZN(_01889_));
 NOR2_X4 _27131_ (.A1(_16845_),
    .A2(_16844_),
    .ZN(_01890_));
 BUF_X8 _27132_ (.A(_01890_),
    .Z(_01891_));
 NOR2_X1 _27133_ (.A1(_01889_),
    .A2(_01891_),
    .ZN(_01892_));
 INV_X32 _27134_ (.A(_16851_),
    .ZN(_01893_));
 NOR2_X4 _27135_ (.A1(_01893_),
    .A2(_16850_),
    .ZN(_01894_));
 NOR2_X4 _27136_ (.A1(_16849_),
    .A2(_16848_),
    .ZN(_01895_));
 BUF_X4 _27137_ (.A(_01895_),
    .Z(_01896_));
 AND2_X2 _27138_ (.A1(_01894_),
    .A2(_01896_),
    .ZN(_01897_));
 BUF_X4 _27139_ (.A(_01897_),
    .Z(_01898_));
 AND2_X1 _27140_ (.A1(_01892_),
    .A2(_01898_),
    .ZN(_01899_));
 INV_X1 _27141_ (.A(_01899_),
    .ZN(_01900_));
 INV_X32 _27142_ (.A(_16847_),
    .ZN(_01901_));
 NOR2_X4 _27143_ (.A1(_01901_),
    .A2(_16846_),
    .ZN(_01902_));
 BUF_X4 _27144_ (.A(_01902_),
    .Z(_01903_));
 BUF_X32 _27145_ (.A(_16844_),
    .Z(_01904_));
 AND2_X2 _27146_ (.A1(_01903_),
    .A2(_01904_),
    .ZN(_01905_));
 NOR2_X4 _27147_ (.A1(_16846_),
    .A2(_16847_),
    .ZN(_01906_));
 BUF_X8 _27148_ (.A(_01906_),
    .Z(_01907_));
 BUF_X4 _27149_ (.A(_01907_),
    .Z(_01908_));
 INV_X32 _27150_ (.A(_16844_),
    .ZN(_01909_));
 BUF_X4 _27151_ (.A(_01909_),
    .Z(_01910_));
 AND2_X1 _27152_ (.A1(_01908_),
    .A2(_01910_),
    .ZN(_01911_));
 OAI21_X1 _27153_ (.A(_01898_),
    .B1(_01905_),
    .B2(_01911_),
    .ZN(_01912_));
 AND2_X4 _27154_ (.A1(_16845_),
    .A2(_16844_),
    .ZN(_01913_));
 AND2_X2 _27155_ (.A1(_01888_),
    .A2(_01913_),
    .ZN(_01914_));
 AND2_X4 _27156_ (.A1(_01893_),
    .A2(_16850_),
    .ZN(_01915_));
 BUF_X8 _27157_ (.A(_01915_),
    .Z(_01916_));
 INV_X32 _27158_ (.A(_16849_),
    .ZN(_01917_));
 AND2_X4 _27159_ (.A1(_01917_),
    .A2(_16848_),
    .ZN(_01918_));
 AND3_X1 _27160_ (.A1(_01914_),
    .A2(_01916_),
    .A3(_01918_),
    .ZN(_01919_));
 AND2_X4 _27161_ (.A1(_01918_),
    .A2(_01915_),
    .ZN(_01920_));
 INV_X4 _27162_ (.A(_01891_),
    .ZN(_01921_));
 NAND2_X1 _27163_ (.A1(_01921_),
    .A2(_01907_),
    .ZN(_01922_));
 INV_X1 _27164_ (.A(_01922_),
    .ZN(_01923_));
 AND2_X4 _27165_ (.A1(_16849_),
    .A2(_16848_),
    .ZN(_01924_));
 NOR2_X4 _27166_ (.A1(_16851_),
    .A2(_16850_),
    .ZN(_01925_));
 AND2_X4 _27167_ (.A1(_01924_),
    .A2(_01925_),
    .ZN(_01926_));
 BUF_X8 _27168_ (.A(_01926_),
    .Z(_01927_));
 AOI221_X1 _27169_ (.A(_01919_),
    .B1(_01905_),
    .B2(_01920_),
    .C1(_01923_),
    .C2(_01927_),
    .ZN(_01928_));
 INV_X32 _27170_ (.A(_16846_),
    .ZN(_01929_));
 NOR2_X4 _27171_ (.A1(_01929_),
    .A2(_16847_),
    .ZN(_01930_));
 INV_X1 _27172_ (.A(_01930_),
    .ZN(_01931_));
 INV_X8 _27173_ (.A(_16845_),
    .ZN(_01932_));
 NOR2_X4 _27174_ (.A1(_01932_),
    .A2(_01904_),
    .ZN(_01933_));
 BUF_X4 _27175_ (.A(_01933_),
    .Z(_01934_));
 NOR2_X1 _27176_ (.A1(_01931_),
    .A2(_01934_),
    .ZN(_01935_));
 NAND2_X1 _27177_ (.A1(_01935_),
    .A2(_01898_),
    .ZN(_01936_));
 AND2_X2 _27178_ (.A1(_01915_),
    .A2(_01924_),
    .ZN(_01937_));
 BUF_X4 _27179_ (.A(_01937_),
    .Z(_01938_));
 AND2_X4 _27180_ (.A1(_01902_),
    .A2(_01913_),
    .ZN(_01939_));
 BUF_X4 _27181_ (.A(_01939_),
    .Z(_01940_));
 AND2_X2 _27182_ (.A1(_01933_),
    .A2(_01888_),
    .ZN(_01941_));
 OR2_X1 _27183_ (.A1(_01940_),
    .A2(_01941_),
    .ZN(_01942_));
 NOR2_X4 _27184_ (.A1(_01909_),
    .A2(_16845_),
    .ZN(_01943_));
 BUF_X8 _27185_ (.A(_01943_),
    .Z(_01944_));
 AND2_X4 _27186_ (.A1(_01944_),
    .A2(_01888_),
    .ZN(_01945_));
 OAI21_X1 _27187_ (.A(_01938_),
    .B1(_01942_),
    .B2(_01945_),
    .ZN(_01946_));
 AND4_X1 _27188_ (.A1(_01912_),
    .A2(_01928_),
    .A3(_01936_),
    .A4(_01946_),
    .ZN(_01947_));
 INV_X1 _27189_ (.A(_01939_),
    .ZN(_01948_));
 AND2_X2 _27190_ (.A1(_01902_),
    .A2(_01891_),
    .ZN(_01949_));
 INV_X1 _27191_ (.A(_01949_),
    .ZN(_01950_));
 NAND2_X1 _27192_ (.A1(_01948_),
    .A2(_01950_),
    .ZN(_01951_));
 NOR2_X4 _27193_ (.A1(_01917_),
    .A2(_16848_),
    .ZN(_01952_));
 AND2_X4 _27194_ (.A1(_01915_),
    .A2(_01952_),
    .ZN(_01953_));
 BUF_X4 _27195_ (.A(_01953_),
    .Z(_01954_));
 AND2_X1 _27196_ (.A1(_01951_),
    .A2(_01954_),
    .ZN(_01955_));
 INV_X1 _27197_ (.A(_01955_),
    .ZN(_01956_));
 BUF_X4 _27198_ (.A(_01920_),
    .Z(_01957_));
 INV_X4 _27199_ (.A(_01907_),
    .ZN(_01958_));
 NOR2_X1 _27200_ (.A1(_01958_),
    .A2(_01934_),
    .ZN(_01959_));
 BUF_X4 _27201_ (.A(_01954_),
    .Z(_01960_));
 AND2_X4 _27202_ (.A1(_01944_),
    .A2(_01903_),
    .ZN(_01961_));
 AOI22_X1 _27203_ (.A1(_01957_),
    .A2(_01959_),
    .B1(_01960_),
    .B2(_01961_),
    .ZN(_01962_));
 AND2_X1 _27204_ (.A1(_01956_),
    .A2(_01962_),
    .ZN(_01963_));
 AND2_X4 _27205_ (.A1(_01952_),
    .A2(_01894_),
    .ZN(_01964_));
 BUF_X2 _27206_ (.A(_01964_),
    .Z(_01965_));
 BUF_X4 _27207_ (.A(_01965_),
    .Z(_01966_));
 BUF_X8 _27208_ (.A(_01914_),
    .Z(_01967_));
 AND2_X2 _27209_ (.A1(_01888_),
    .A2(_01932_),
    .ZN(_01968_));
 BUF_X4 _27210_ (.A(_01968_),
    .Z(_01969_));
 OAI21_X1 _27211_ (.A(_01966_),
    .B1(_01967_),
    .B2(_01969_),
    .ZN(_01970_));
 BUF_X4 _27212_ (.A(_01903_),
    .Z(_01971_));
 BUF_X8 _27213_ (.A(_01952_),
    .Z(_01972_));
 BUF_X2 _27214_ (.A(_01894_),
    .Z(_01973_));
 NAND4_X1 _27215_ (.A1(_01944_),
    .A2(_01971_),
    .A3(_01972_),
    .A4(_01973_),
    .ZN(_01974_));
 NAND2_X1 _27216_ (.A1(_01970_),
    .A2(_01974_),
    .ZN(_01975_));
 INV_X1 _27217_ (.A(_01903_),
    .ZN(_01976_));
 NOR2_X1 _27218_ (.A1(_01976_),
    .A2(_01944_),
    .ZN(_01977_));
 AND2_X4 _27219_ (.A1(_16851_),
    .A2(_16850_),
    .ZN(_01978_));
 AND2_X4 _27220_ (.A1(_01972_),
    .A2(_01978_),
    .ZN(_01979_));
 BUF_X8 _27221_ (.A(_01979_),
    .Z(_01980_));
 BUF_X4 _27222_ (.A(_01980_),
    .Z(_01981_));
 AND2_X1 _27223_ (.A1(_01977_),
    .A2(_01981_),
    .ZN(_01982_));
 AND2_X4 _27224_ (.A1(_01894_),
    .A2(_01924_),
    .ZN(_01983_));
 BUF_X8 _27225_ (.A(_01983_),
    .Z(_01984_));
 INV_X4 _27226_ (.A(_01934_),
    .ZN(_01985_));
 BUF_X4 _27227_ (.A(_01930_),
    .Z(_01986_));
 AND3_X1 _27228_ (.A1(_01984_),
    .A2(_01985_),
    .A3(_01986_),
    .ZN(_01987_));
 NOR3_X1 _27229_ (.A1(_01975_),
    .A2(_01982_),
    .A3(_01987_),
    .ZN(_01988_));
 AND4_X1 _27230_ (.A1(_01900_),
    .A2(_01947_),
    .A3(_01963_),
    .A4(_01988_),
    .ZN(_01989_));
 BUF_X8 _27231_ (.A(_01978_),
    .Z(_01990_));
 AND2_X4 _27232_ (.A1(_01918_),
    .A2(_01990_),
    .ZN(_01991_));
 BUF_X4 _27233_ (.A(_01991_),
    .Z(_01992_));
 AND2_X2 _27234_ (.A1(_01943_),
    .A2(_01930_),
    .ZN(_01993_));
 AND2_X2 _27235_ (.A1(_01933_),
    .A2(_01906_),
    .ZN(_01994_));
 BUF_X2 _27236_ (.A(_01994_),
    .Z(_01995_));
 OAI21_X1 _27237_ (.A(_01992_),
    .B1(_01993_),
    .B2(_01995_),
    .ZN(_01996_));
 NAND2_X1 _27238_ (.A1(_01902_),
    .A2(_01932_),
    .ZN(_01997_));
 INV_X1 _27239_ (.A(_01997_),
    .ZN(_01998_));
 BUF_X2 _27240_ (.A(_01998_),
    .Z(_01999_));
 NAND2_X1 _27241_ (.A1(_01992_),
    .A2(_01999_),
    .ZN(_02000_));
 AND2_X2 _27242_ (.A1(_01903_),
    .A2(_01933_),
    .ZN(_02001_));
 NAND2_X1 _27243_ (.A1(_01992_),
    .A2(_02001_),
    .ZN(_02002_));
 NAND2_X1 _27244_ (.A1(_01991_),
    .A2(_01939_),
    .ZN(_02003_));
 AND3_X1 _27245_ (.A1(_02000_),
    .A2(_02002_),
    .A3(_02003_),
    .ZN(_02004_));
 INV_X1 _27246_ (.A(_01913_),
    .ZN(_02005_));
 BUF_X4 _27247_ (.A(_01918_),
    .Z(_02006_));
 NAND4_X1 _27248_ (.A1(_01892_),
    .A2(_02005_),
    .A3(_02006_),
    .A4(_01990_),
    .ZN(_02007_));
 AND2_X4 _27249_ (.A1(_01990_),
    .A2(_01896_),
    .ZN(_02008_));
 BUF_X16 _27250_ (.A(_02008_),
    .Z(_02009_));
 BUF_X16 _27251_ (.A(_02009_),
    .Z(_02010_));
 OAI21_X1 _27252_ (.A(_02010_),
    .B1(_01905_),
    .B2(_01969_),
    .ZN(_02011_));
 AND4_X1 _27253_ (.A1(_01996_),
    .A2(_02004_),
    .A3(_02007_),
    .A4(_02011_),
    .ZN(_02012_));
 AND2_X4 _27254_ (.A1(_01916_),
    .A2(_01896_),
    .ZN(_02013_));
 BUF_X4 _27255_ (.A(_02013_),
    .Z(_02014_));
 BUF_X4 _27256_ (.A(_01941_),
    .Z(_02015_));
 OAI21_X1 _27257_ (.A(_02014_),
    .B1(_02015_),
    .B2(_01969_),
    .ZN(_02016_));
 BUF_X4 _27258_ (.A(_01904_),
    .Z(_02017_));
 NAND4_X1 _27259_ (.A1(_01916_),
    .A2(_01971_),
    .A3(_02017_),
    .A4(_01896_),
    .ZN(_02018_));
 AND2_X1 _27260_ (.A1(_02016_),
    .A2(_02018_),
    .ZN(_02019_));
 AND2_X4 _27261_ (.A1(_01924_),
    .A2(_01978_),
    .ZN(_02020_));
 BUF_X4 _27262_ (.A(_02020_),
    .Z(_02021_));
 BUF_X8 _27263_ (.A(_16845_),
    .Z(_02022_));
 AND2_X2 _27264_ (.A1(_01907_),
    .A2(_02022_),
    .ZN(_02023_));
 AND2_X2 _27265_ (.A1(_02021_),
    .A2(_02023_),
    .ZN(_02024_));
 BUF_X8 _27266_ (.A(_01888_),
    .Z(_02025_));
 AND2_X2 _27267_ (.A1(_02025_),
    .A2(_01904_),
    .ZN(_02026_));
 AOI221_X4 _27268_ (.A(_02024_),
    .B1(_01971_),
    .B2(_02021_),
    .C1(_01981_),
    .C2(_02026_),
    .ZN(_02027_));
 OAI21_X1 _27269_ (.A(_01901_),
    .B1(_01921_),
    .B2(_16846_),
    .ZN(_02028_));
 AND3_X1 _27270_ (.A1(_01896_),
    .A2(_01925_),
    .A3(_01901_),
    .ZN(_02029_));
 AND2_X1 _27271_ (.A1(_02028_),
    .A2(_02029_),
    .ZN(_02030_));
 INV_X1 _27272_ (.A(_02030_),
    .ZN(_02031_));
 NOR2_X4 _27273_ (.A1(_01958_),
    .A2(_01944_),
    .ZN(_02032_));
 AND2_X4 _27274_ (.A1(_02032_),
    .A2(_01985_),
    .ZN(_02033_));
 AND2_X2 _27275_ (.A1(_01930_),
    .A2(_01932_),
    .ZN(_02034_));
 OAI21_X1 _27276_ (.A(_01981_),
    .B1(_02033_),
    .B2(_02034_),
    .ZN(_02035_));
 AND4_X2 _27277_ (.A1(_02019_),
    .A2(_02027_),
    .A3(_02031_),
    .A4(_02035_),
    .ZN(_02036_));
 AND2_X4 _27278_ (.A1(_01972_),
    .A2(_01925_),
    .ZN(_02037_));
 NAND2_X1 _27279_ (.A1(_02037_),
    .A2(_01994_),
    .ZN(_02038_));
 AND2_X1 _27280_ (.A1(_01906_),
    .A2(_01932_),
    .ZN(_02039_));
 NAND3_X1 _27281_ (.A1(_02039_),
    .A2(_01925_),
    .A3(_01972_),
    .ZN(_02040_));
 AND2_X2 _27282_ (.A1(_02038_),
    .A2(_02040_),
    .ZN(_02041_));
 AND2_X2 _27283_ (.A1(_01888_),
    .A2(_01890_),
    .ZN(_02042_));
 NOR2_X1 _27284_ (.A1(_02032_),
    .A2(_02042_),
    .ZN(_02043_));
 INV_X2 _27285_ (.A(_01984_),
    .ZN(_02044_));
 NOR2_X1 _27286_ (.A1(_02043_),
    .A2(_02044_),
    .ZN(_02045_));
 AND2_X2 _27287_ (.A1(_02008_),
    .A2(_02023_),
    .ZN(_02046_));
 AOI221_X1 _27288_ (.A(_02045_),
    .B1(_01910_),
    .B2(_02046_),
    .C1(_02015_),
    .C2(_02009_),
    .ZN(_02047_));
 AND2_X2 _27289_ (.A1(_01921_),
    .A2(_01903_),
    .ZN(_02048_));
 NAND2_X4 _27290_ (.A1(_02048_),
    .A2(_02037_),
    .ZN(_02049_));
 AND2_X4 _27291_ (.A1(_01930_),
    .A2(_01890_),
    .ZN(_02050_));
 AND2_X1 _27292_ (.A1(_02050_),
    .A2(_02020_),
    .ZN(_02051_));
 AND2_X1 _27293_ (.A1(_01943_),
    .A2(_01906_),
    .ZN(_02052_));
 BUF_X2 _27294_ (.A(_02052_),
    .Z(_02053_));
 AND2_X1 _27295_ (.A1(_01888_),
    .A2(_01909_),
    .ZN(_02054_));
 AND2_X1 _27296_ (.A1(_02021_),
    .A2(_02054_),
    .ZN(_02055_));
 AOI221_X4 _27297_ (.A(_02051_),
    .B1(_02053_),
    .B2(_02021_),
    .C1(_02022_),
    .C2(_02055_),
    .ZN(_02056_));
 AND4_X1 _27298_ (.A1(_02041_),
    .A2(_02047_),
    .A3(_02049_),
    .A4(_02056_),
    .ZN(_02057_));
 AND4_X2 _27299_ (.A1(_01989_),
    .A2(_02012_),
    .A3(_02036_),
    .A4(_02057_),
    .ZN(_02058_));
 AND2_X2 _27300_ (.A1(_02013_),
    .A2(_02050_),
    .ZN(_02059_));
 AND2_X2 _27301_ (.A1(_01913_),
    .A2(_01907_),
    .ZN(_02060_));
 BUF_X2 _27302_ (.A(_02060_),
    .Z(_02061_));
 AND2_X1 _27303_ (.A1(_01960_),
    .A2(_02061_),
    .ZN(_02062_));
 AND2_X4 _27304_ (.A1(_01933_),
    .A2(_01930_),
    .ZN(_02063_));
 BUF_X4 _27305_ (.A(_02063_),
    .Z(_02064_));
 AND2_X1 _27306_ (.A1(_01954_),
    .A2(_02064_),
    .ZN(_02065_));
 AND2_X2 _27307_ (.A1(_01954_),
    .A2(_02053_),
    .ZN(_02066_));
 NOR4_X1 _27308_ (.A1(_02059_),
    .A2(_02062_),
    .A3(_02065_),
    .A4(_02066_),
    .ZN(_02067_));
 AND2_X4 _27309_ (.A1(_01918_),
    .A2(_01925_),
    .ZN(_02068_));
 BUF_X4 _27310_ (.A(_02068_),
    .Z(_02069_));
 BUF_X2 _27311_ (.A(_02069_),
    .Z(_02070_));
 NOR3_X4 _27312_ (.A1(_01891_),
    .A2(_01929_),
    .A3(_16847_),
    .ZN(_02071_));
 AND2_X4 _27313_ (.A1(_02071_),
    .A2(_02005_),
    .ZN(_02072_));
 OAI21_X1 _27314_ (.A(_02070_),
    .B1(_01951_),
    .B2(_02072_),
    .ZN(_02073_));
 AND2_X1 _27315_ (.A1(_01918_),
    .A2(_01894_),
    .ZN(_02074_));
 AND4_X1 _27316_ (.A1(_02005_),
    .A2(_02074_),
    .A3(_01921_),
    .A4(_01908_),
    .ZN(_02075_));
 AND2_X2 _27317_ (.A1(_01888_),
    .A2(_16845_),
    .ZN(_02076_));
 BUF_X2 _27318_ (.A(_02076_),
    .Z(_02077_));
 BUF_X2 _27319_ (.A(_02074_),
    .Z(_02078_));
 AOI21_X1 _27320_ (.A(_02075_),
    .B1(_02077_),
    .B2(_02078_),
    .ZN(_02079_));
 BUF_X4 _27321_ (.A(_01938_),
    .Z(_02080_));
 AND2_X2 _27322_ (.A1(_01930_),
    .A2(_01904_),
    .ZN(_02081_));
 AND2_X2 _27323_ (.A1(_01907_),
    .A2(_01904_),
    .ZN(_02082_));
 OAI21_X1 _27324_ (.A(_02080_),
    .B1(_02081_),
    .B2(_02082_),
    .ZN(_02083_));
 BUF_X4 _27325_ (.A(_02037_),
    .Z(_02084_));
 OAI21_X1 _27326_ (.A(_02084_),
    .B1(_02072_),
    .B2(_02077_),
    .ZN(_02085_));
 AND4_X1 _27327_ (.A1(_02073_),
    .A2(_02079_),
    .A3(_02083_),
    .A4(_02085_),
    .ZN(_02086_));
 AND2_X4 _27328_ (.A1(_01960_),
    .A2(_02015_),
    .ZN(_02087_));
 INV_X2 _27329_ (.A(_02087_),
    .ZN(_02088_));
 AND2_X4 _27330_ (.A1(_01930_),
    .A2(_01913_),
    .ZN(_02089_));
 BUF_X4 _27331_ (.A(_02089_),
    .Z(_02090_));
 NAND2_X1 _27332_ (.A1(_01954_),
    .A2(_02090_),
    .ZN(_02091_));
 AND2_X4 _27333_ (.A1(_01891_),
    .A2(_01907_),
    .ZN(_02092_));
 BUF_X8 _27334_ (.A(_02092_),
    .Z(_02093_));
 AOI22_X1 _27335_ (.A1(_02080_),
    .A2(_02093_),
    .B1(_01966_),
    .B2(_02050_),
    .ZN(_02094_));
 NAND3_X1 _27336_ (.A1(_02088_),
    .A2(_02091_),
    .A3(_02094_),
    .ZN(_02095_));
 AND2_X1 _27337_ (.A1(_01895_),
    .A2(_01925_),
    .ZN(_02096_));
 BUF_X4 _27338_ (.A(_02096_),
    .Z(_02097_));
 BUF_X4 _27339_ (.A(_01971_),
    .Z(_02098_));
 BUF_X4 _27340_ (.A(_01986_),
    .Z(_02099_));
 OAI211_X2 _27341_ (.A(_02097_),
    .B(_01944_),
    .C1(_02098_),
    .C2(_02099_),
    .ZN(_02100_));
 INV_X1 _27342_ (.A(_02037_),
    .ZN(_02101_));
 INV_X1 _27343_ (.A(_02042_),
    .ZN(_02102_));
 BUF_X4 _27344_ (.A(_01927_),
    .Z(_02103_));
 INV_X1 _27345_ (.A(_02103_),
    .ZN(_02104_));
 OAI221_X1 _27346_ (.A(_02100_),
    .B1(_02101_),
    .B2(_02102_),
    .C1(_01950_),
    .C2(_02104_),
    .ZN(_02105_));
 BUF_X4 _27347_ (.A(_02023_),
    .Z(_02106_));
 AND2_X1 _27348_ (.A1(_02070_),
    .A2(_02106_),
    .ZN(_02107_));
 INV_X1 _27349_ (.A(_02064_),
    .ZN(_02108_));
 INV_X1 _27350_ (.A(_01914_),
    .ZN(_02109_));
 AOI21_X1 _27351_ (.A(_02104_),
    .B1(_02108_),
    .B2(_02109_),
    .ZN(_02110_));
 NOR4_X1 _27352_ (.A1(_02095_),
    .A2(_02105_),
    .A3(_02107_),
    .A4(_02110_),
    .ZN(_02111_));
 AND2_X2 _27353_ (.A1(_01930_),
    .A2(_02022_),
    .ZN(_02112_));
 BUF_X4 _27354_ (.A(_02039_),
    .Z(_02113_));
 AOI22_X1 _27355_ (.A1(_01957_),
    .A2(_02112_),
    .B1(_02014_),
    .B2(_02113_),
    .ZN(_02114_));
 NAND2_X1 _27356_ (.A1(_01960_),
    .A2(_02034_),
    .ZN(_02115_));
 INV_X1 _27357_ (.A(_01968_),
    .ZN(_02116_));
 OAI211_X2 _27358_ (.A(_02114_),
    .B(_02115_),
    .C1(_02116_),
    .C2(_02104_),
    .ZN(_02117_));
 BUF_X4 _27359_ (.A(_01932_),
    .Z(_02118_));
 INV_X1 _27360_ (.A(_02097_),
    .ZN(_02119_));
 AOI211_X4 _27361_ (.A(_02118_),
    .B(_02119_),
    .C1(_01958_),
    .C2(_01931_),
    .ZN(_02120_));
 AND2_X4 _27362_ (.A1(_01902_),
    .A2(_02022_),
    .ZN(_02121_));
 BUF_X2 _27363_ (.A(_02121_),
    .Z(_02122_));
 BUF_X4 _27364_ (.A(_02097_),
    .Z(_02123_));
 AND2_X1 _27365_ (.A1(_02122_),
    .A2(_02123_),
    .ZN(_02124_));
 AND3_X1 _27366_ (.A1(_01892_),
    .A2(_02005_),
    .A3(_02097_),
    .ZN(_02125_));
 NOR4_X1 _27367_ (.A1(_02117_),
    .A2(_02120_),
    .A3(_02124_),
    .A4(_02125_),
    .ZN(_02126_));
 AND4_X1 _27368_ (.A1(_02067_),
    .A2(_02086_),
    .A3(_02111_),
    .A4(_02126_),
    .ZN(_02127_));
 AND2_X4 _27369_ (.A1(_02058_),
    .A2(_02127_),
    .ZN(_02128_));
 INV_X32 _27370_ (.A(_16809_),
    .ZN(_02129_));
 AND2_X4 _27371_ (.A1(_02129_),
    .A2(_16808_),
    .ZN(_02130_));
 AND2_X4 _27372_ (.A1(_16811_),
    .A2(_16810_),
    .ZN(_02131_));
 BUF_X8 _27373_ (.A(_02131_),
    .Z(_02132_));
 AND2_X2 _27374_ (.A1(_02130_),
    .A2(_02132_),
    .ZN(_02133_));
 BUF_X4 _27375_ (.A(_02133_),
    .Z(_02134_));
 INV_X32 _27376_ (.A(_16806_),
    .ZN(_02135_));
 NOR2_X4 _27377_ (.A1(_02135_),
    .A2(_16807_),
    .ZN(_02136_));
 INV_X32 _27378_ (.A(_16804_),
    .ZN(_02137_));
 NOR2_X4 _27379_ (.A1(_02137_),
    .A2(_16805_),
    .ZN(_02138_));
 BUF_X4 _27380_ (.A(_02138_),
    .Z(_02139_));
 AND2_X1 _27381_ (.A1(_02136_),
    .A2(_02139_),
    .ZN(_02140_));
 BUF_X2 _27382_ (.A(_02140_),
    .Z(_02141_));
 INV_X32 _27383_ (.A(_16805_),
    .ZN(_02142_));
 NOR2_X4 _27384_ (.A1(_02142_),
    .A2(_16804_),
    .ZN(_02143_));
 BUF_X4 _27385_ (.A(_02143_),
    .Z(_02144_));
 NOR2_X4 _27386_ (.A1(_16806_),
    .A2(_16807_),
    .ZN(_02145_));
 BUF_X4 _27387_ (.A(_02145_),
    .Z(_02146_));
 AND2_X2 _27388_ (.A1(_02144_),
    .A2(_02146_),
    .ZN(_02147_));
 NOR2_X1 _27389_ (.A1(_02141_),
    .A2(_02147_),
    .ZN(_02148_));
 INV_X1 _27390_ (.A(_02148_),
    .ZN(_02149_));
 AND2_X4 _27391_ (.A1(_16806_),
    .A2(_16807_),
    .ZN(_02150_));
 BUF_X8 _27392_ (.A(_02150_),
    .Z(_02151_));
 AND2_X4 _27393_ (.A1(_02138_),
    .A2(_02151_),
    .ZN(_02152_));
 BUF_X8 _27394_ (.A(_02152_),
    .Z(_02153_));
 INV_X2 _27395_ (.A(_02153_),
    .ZN(_02154_));
 AND2_X4 _27396_ (.A1(_02143_),
    .A2(_02151_),
    .ZN(_02155_));
 BUF_X8 _27397_ (.A(_02155_),
    .Z(_02156_));
 INV_X1 _27398_ (.A(_02156_),
    .ZN(_02157_));
 INV_X32 _27399_ (.A(_16807_),
    .ZN(_02158_));
 NOR2_X4 _27400_ (.A1(_02158_),
    .A2(_16806_),
    .ZN(_02159_));
 INV_X1 _27401_ (.A(_02159_),
    .ZN(_02160_));
 NAND3_X1 _27402_ (.A1(_02154_),
    .A2(_02157_),
    .A3(_02160_),
    .ZN(_02161_));
 OAI21_X1 _27403_ (.A(_02134_),
    .B1(_02149_),
    .B2(_02161_),
    .ZN(_02162_));
 NOR2_X4 _27404_ (.A1(_16809_),
    .A2(_16808_),
    .ZN(_02163_));
 BUF_X2 _27405_ (.A(_02163_),
    .Z(_02164_));
 AND2_X4 _27406_ (.A1(_02132_),
    .A2(_02164_),
    .ZN(_02165_));
 INV_X2 _27407_ (.A(_02165_),
    .ZN(_02166_));
 INV_X4 _27408_ (.A(_02139_),
    .ZN(_02167_));
 AND2_X4 _27409_ (.A1(_16805_),
    .A2(_16804_),
    .ZN(_02168_));
 BUF_X8 _27410_ (.A(_02168_),
    .Z(_02169_));
 INV_X2 _27411_ (.A(_02169_),
    .ZN(_02170_));
 AOI211_X4 _27412_ (.A(_02160_),
    .B(_02166_),
    .C1(_02167_),
    .C2(_02170_),
    .ZN(_02171_));
 INV_X8 _27413_ (.A(_02151_),
    .ZN(_02172_));
 BUF_X32 _27414_ (.A(_16805_),
    .Z(_02173_));
 BUF_X4 _27415_ (.A(_16804_),
    .Z(_02174_));
 AOI211_X4 _27416_ (.A(_02172_),
    .B(_02166_),
    .C1(_02173_),
    .C2(_02174_),
    .ZN(_02175_));
 BUF_X4 _27417_ (.A(_02165_),
    .Z(_02176_));
 AOI211_X2 _27418_ (.A(_02171_),
    .B(_02175_),
    .C1(_02147_),
    .C2(_02176_),
    .ZN(_02177_));
 NOR2_X1 _27419_ (.A1(_02160_),
    .A2(_02139_),
    .ZN(_02178_));
 NOR2_X4 _27420_ (.A1(_02129_),
    .A2(_16808_),
    .ZN(_02179_));
 AND2_X4 _27421_ (.A1(_02179_),
    .A2(_02132_),
    .ZN(_02180_));
 BUF_X4 _27422_ (.A(_02180_),
    .Z(_02181_));
 BUF_X4 _27423_ (.A(_02181_),
    .Z(_02182_));
 NAND2_X1 _27424_ (.A1(_02178_),
    .A2(_02182_),
    .ZN(_02183_));
 AND2_X1 _27425_ (.A1(_02136_),
    .A2(_02142_),
    .ZN(_02184_));
 BUF_X2 _27426_ (.A(_02184_),
    .Z(_02185_));
 AND2_X1 _27427_ (.A1(_02181_),
    .A2(_02185_),
    .ZN(_02186_));
 INV_X1 _27428_ (.A(_02186_),
    .ZN(_02187_));
 INV_X1 _27429_ (.A(_02145_),
    .ZN(_02188_));
 NOR2_X1 _27430_ (.A1(_02188_),
    .A2(_02144_),
    .ZN(_02189_));
 NAND3_X1 _27431_ (.A1(_02182_),
    .A2(_02189_),
    .A3(_02167_),
    .ZN(_02190_));
 BUF_X4 _27432_ (.A(_02151_),
    .Z(_02191_));
 AND2_X2 _27433_ (.A1(_02191_),
    .A2(_02174_),
    .ZN(_02192_));
 BUF_X4 _27434_ (.A(_02132_),
    .Z(_02193_));
 BUF_X4 _27435_ (.A(_02179_),
    .Z(_02194_));
 NAND3_X1 _27436_ (.A1(_02192_),
    .A2(_02193_),
    .A3(_02194_),
    .ZN(_02195_));
 AND4_X1 _27437_ (.A1(_02183_),
    .A2(_02187_),
    .A3(_02190_),
    .A4(_02195_),
    .ZN(_02196_));
 NOR2_X4 _27438_ (.A1(_16805_),
    .A2(_16804_),
    .ZN(_02197_));
 AND2_X1 _27439_ (.A1(_02136_),
    .A2(_02197_),
    .ZN(_02198_));
 AND2_X4 _27440_ (.A1(_16809_),
    .A2(_16808_),
    .ZN(_02199_));
 AND2_X2 _27441_ (.A1(_02131_),
    .A2(_02199_),
    .ZN(_02200_));
 BUF_X4 _27442_ (.A(_02200_),
    .Z(_02201_));
 BUF_X4 _27443_ (.A(_02201_),
    .Z(_02202_));
 NAND2_X1 _27444_ (.A1(_02198_),
    .A2(_02202_),
    .ZN(_02203_));
 NOR2_X1 _27445_ (.A1(_02158_),
    .A2(_02173_),
    .ZN(_02204_));
 AND2_X2 _27446_ (.A1(_02204_),
    .A2(_02135_),
    .ZN(_02205_));
 BUF_X4 _27447_ (.A(_02205_),
    .Z(_02206_));
 AND2_X2 _27448_ (.A1(_02159_),
    .A2(_16805_),
    .ZN(_02207_));
 BUF_X8 _27449_ (.A(_02207_),
    .Z(_02208_));
 BUF_X4 _27450_ (.A(_02208_),
    .Z(_02209_));
 OAI21_X1 _27451_ (.A(_02202_),
    .B1(_02206_),
    .B2(_02209_),
    .ZN(_02210_));
 BUF_X4 _27452_ (.A(_02146_),
    .Z(_02211_));
 BUF_X4 _27453_ (.A(_02174_),
    .Z(_02212_));
 OAI211_X2 _27454_ (.A(_02202_),
    .B(_02211_),
    .C1(_02173_),
    .C2(_02212_),
    .ZN(_02213_));
 BUF_X4 _27455_ (.A(_02144_),
    .Z(_02214_));
 NAND3_X1 _27456_ (.A1(_02201_),
    .A2(_02214_),
    .A3(_02191_),
    .ZN(_02215_));
 AND4_X1 _27457_ (.A1(_02203_),
    .A2(_02210_),
    .A3(_02213_),
    .A4(_02215_),
    .ZN(_02216_));
 AND4_X1 _27458_ (.A1(_02162_),
    .A2(_02177_),
    .A3(_02196_),
    .A4(_02216_),
    .ZN(_02217_));
 AND2_X2 _27459_ (.A1(_02159_),
    .A2(_02169_),
    .ZN(_02218_));
 BUF_X4 _27460_ (.A(_02159_),
    .Z(_02219_));
 BUF_X4 _27461_ (.A(_02197_),
    .Z(_02220_));
 AND2_X2 _27462_ (.A1(_02219_),
    .A2(_02220_),
    .ZN(_02221_));
 OR2_X1 _27463_ (.A1(_02218_),
    .A2(_02221_),
    .ZN(_02222_));
 NOR2_X4 _27464_ (.A1(_16811_),
    .A2(_16810_),
    .ZN(_02223_));
 AND2_X1 _27465_ (.A1(_02130_),
    .A2(_02223_),
    .ZN(_02224_));
 BUF_X4 _27466_ (.A(_02224_),
    .Z(_02225_));
 BUF_X4 _27467_ (.A(_02225_),
    .Z(_02226_));
 NAND2_X1 _27468_ (.A1(_02222_),
    .A2(_02226_),
    .ZN(_02227_));
 AND2_X1 _27469_ (.A1(_02163_),
    .A2(_02223_),
    .ZN(_02228_));
 AND2_X4 _27470_ (.A1(_02145_),
    .A2(_02173_),
    .ZN(_02229_));
 BUF_X4 _27471_ (.A(_02229_),
    .Z(_02230_));
 AND2_X1 _27472_ (.A1(_02228_),
    .A2(_02230_),
    .ZN(_02231_));
 AND2_X1 _27473_ (.A1(_02136_),
    .A2(_02173_),
    .ZN(_02232_));
 BUF_X2 _27474_ (.A(_02228_),
    .Z(_02233_));
 AND2_X1 _27475_ (.A1(_02232_),
    .A2(_02233_),
    .ZN(_02234_));
 AOI211_X2 _27476_ (.A(_02231_),
    .B(_02234_),
    .C1(_02141_),
    .C2(_02233_),
    .ZN(_02235_));
 INV_X1 _27477_ (.A(_02197_),
    .ZN(_02236_));
 BUF_X4 _27478_ (.A(_02136_),
    .Z(_02237_));
 AND2_X1 _27479_ (.A1(_02236_),
    .A2(_02237_),
    .ZN(_02238_));
 AND2_X1 _27480_ (.A1(_02238_),
    .A2(_02170_),
    .ZN(_02239_));
 OAI21_X1 _27481_ (.A(_02226_),
    .B1(_02239_),
    .B2(_02230_),
    .ZN(_02240_));
 BUF_X4 _27482_ (.A(_02233_),
    .Z(_02241_));
 NOR2_X1 _27483_ (.A1(_02172_),
    .A2(_02169_),
    .ZN(_02242_));
 BUF_X4 _27484_ (.A(_02219_),
    .Z(_02243_));
 OAI221_X1 _27485_ (.A(_02241_),
    .B1(_02173_),
    .B2(_02212_),
    .C1(_02242_),
    .C2(_02243_),
    .ZN(_02244_));
 AND4_X1 _27486_ (.A1(_02227_),
    .A2(_02235_),
    .A3(_02240_),
    .A4(_02244_),
    .ZN(_02245_));
 AND2_X2 _27487_ (.A1(_02179_),
    .A2(_02223_),
    .ZN(_02246_));
 BUF_X4 _27488_ (.A(_02246_),
    .Z(_02247_));
 OAI211_X2 _27489_ (.A(_02170_),
    .B(_02247_),
    .C1(_02238_),
    .C2(_02211_),
    .ZN(_02248_));
 NAND2_X1 _27490_ (.A1(_02247_),
    .A2(_02209_),
    .ZN(_02249_));
 AND2_X4 _27491_ (.A1(_02151_),
    .A2(_02173_),
    .ZN(_02250_));
 BUF_X2 _27492_ (.A(_02250_),
    .Z(_02251_));
 BUF_X2 _27493_ (.A(_02223_),
    .Z(_02252_));
 NAND3_X1 _27494_ (.A1(_02251_),
    .A2(_02194_),
    .A3(_02252_),
    .ZN(_02253_));
 NAND4_X1 _27495_ (.A1(_02139_),
    .A2(_02243_),
    .A3(_02194_),
    .A4(_02252_),
    .ZN(_02254_));
 NAND4_X1 _27496_ (.A1(_02194_),
    .A2(_02220_),
    .A3(_02191_),
    .A4(_02252_),
    .ZN(_02255_));
 AND4_X1 _27497_ (.A1(_02249_),
    .A2(_02253_),
    .A3(_02254_),
    .A4(_02255_),
    .ZN(_02256_));
 AND2_X4 _27498_ (.A1(_02168_),
    .A2(_02151_),
    .ZN(_02257_));
 AND2_X2 _27499_ (.A1(_02199_),
    .A2(_02223_),
    .ZN(_02258_));
 AND2_X4 _27500_ (.A1(_02257_),
    .A2(_02258_),
    .ZN(_02259_));
 AND2_X4 _27501_ (.A1(_02151_),
    .A2(_02142_),
    .ZN(_02260_));
 AND2_X1 _27502_ (.A1(_02260_),
    .A2(_02258_),
    .ZN(_02261_));
 BUF_X4 _27503_ (.A(_02258_),
    .Z(_02262_));
 AOI211_X2 _27504_ (.A(_02259_),
    .B(_02261_),
    .C1(_02262_),
    .C2(_02221_),
    .ZN(_02263_));
 NOR2_X1 _27505_ (.A1(_02188_),
    .A2(_02197_),
    .ZN(_02264_));
 NAND2_X1 _27506_ (.A1(_02264_),
    .A2(_02262_),
    .ZN(_02265_));
 BUF_X4 _27507_ (.A(_02237_),
    .Z(_02266_));
 BUF_X2 _27508_ (.A(_02199_),
    .Z(_02267_));
 BUF_X4 _27509_ (.A(_02267_),
    .Z(_02268_));
 NAND4_X1 _27510_ (.A1(_02214_),
    .A2(_02266_),
    .A3(_02252_),
    .A4(_02268_),
    .ZN(_02269_));
 AND3_X1 _27511_ (.A1(_02263_),
    .A2(_02265_),
    .A3(_02269_),
    .ZN(_02270_));
 AND4_X2 _27512_ (.A1(_02245_),
    .A2(_02248_),
    .A3(_02256_),
    .A4(_02270_),
    .ZN(_02271_));
 INV_X32 _27513_ (.A(_16811_),
    .ZN(_02272_));
 AND2_X4 _27514_ (.A1(_02272_),
    .A2(_16810_),
    .ZN(_02273_));
 AND2_X4 _27515_ (.A1(_02273_),
    .A2(_02163_),
    .ZN(_02274_));
 BUF_X4 _27516_ (.A(_02274_),
    .Z(_02275_));
 BUF_X4 _27517_ (.A(_02260_),
    .Z(_02276_));
 OAI21_X1 _27518_ (.A(_02275_),
    .B1(_02156_),
    .B2(_02276_),
    .ZN(_02277_));
 BUF_X4 _27519_ (.A(_02273_),
    .Z(_02278_));
 BUF_X4 _27520_ (.A(_02278_),
    .Z(_02279_));
 BUF_X2 _27521_ (.A(_02164_),
    .Z(_02280_));
 NAND4_X1 _27522_ (.A1(_02279_),
    .A2(_02212_),
    .A3(_02243_),
    .A4(_02280_),
    .ZN(_02281_));
 AND2_X1 _27523_ (.A1(_02277_),
    .A2(_02281_),
    .ZN(_02282_));
 NAND3_X1 _27524_ (.A1(_02198_),
    .A2(_02164_),
    .A3(_02278_),
    .ZN(_02283_));
 INV_X2 _27525_ (.A(_02274_),
    .ZN(_02284_));
 AND2_X2 _27526_ (.A1(_02145_),
    .A2(_02142_),
    .ZN(_02285_));
 BUF_X4 _27527_ (.A(_02285_),
    .Z(_02286_));
 INV_X1 _27528_ (.A(_02286_),
    .ZN(_02287_));
 OAI211_X2 _27529_ (.A(_02282_),
    .B(_02283_),
    .C1(_02284_),
    .C2(_02287_),
    .ZN(_02288_));
 AND2_X4 _27530_ (.A1(_02273_),
    .A2(_02130_),
    .ZN(_02289_));
 BUF_X8 _27531_ (.A(_02289_),
    .Z(_02290_));
 BUF_X4 _27532_ (.A(_02290_),
    .Z(_02291_));
 AND2_X1 _27533_ (.A1(_02219_),
    .A2(_02174_),
    .ZN(_02292_));
 OAI21_X1 _27534_ (.A(_02291_),
    .B1(_02292_),
    .B2(_02257_),
    .ZN(_02293_));
 BUF_X4 _27535_ (.A(_02232_),
    .Z(_02294_));
 NAND2_X1 _27536_ (.A1(_02291_),
    .A2(_02294_),
    .ZN(_02295_));
 NAND2_X1 _27537_ (.A1(_02291_),
    .A2(_02286_),
    .ZN(_02296_));
 AND2_X2 _27538_ (.A1(_02169_),
    .A2(_02145_),
    .ZN(_02297_));
 NAND2_X2 _27539_ (.A1(_02290_),
    .A2(_02297_),
    .ZN(_02298_));
 NAND4_X1 _27540_ (.A1(_02293_),
    .A2(_02295_),
    .A3(_02296_),
    .A4(_02298_),
    .ZN(_02299_));
 AND2_X4 _27541_ (.A1(_02273_),
    .A2(_02179_),
    .ZN(_02300_));
 BUF_X4 _27542_ (.A(_02300_),
    .Z(_02301_));
 BUF_X4 _27543_ (.A(_02301_),
    .Z(_02302_));
 OAI21_X1 _27544_ (.A(_02302_),
    .B1(_02294_),
    .B2(_02185_),
    .ZN(_02303_));
 AND2_X1 _27545_ (.A1(_02138_),
    .A2(_02145_),
    .ZN(_02304_));
 BUF_X4 _27546_ (.A(_02304_),
    .Z(_02305_));
 BUF_X4 _27547_ (.A(_02297_),
    .Z(_02306_));
 OAI21_X1 _27548_ (.A(_02302_),
    .B1(_02305_),
    .B2(_02306_),
    .ZN(_02307_));
 NAND2_X1 _27549_ (.A1(_02301_),
    .A2(_02155_),
    .ZN(_02308_));
 NOR2_X1 _27550_ (.A1(_02160_),
    .A2(_02144_),
    .ZN(_02309_));
 NAND2_X1 _27551_ (.A1(_02309_),
    .A2(_02301_),
    .ZN(_02310_));
 NAND4_X1 _27552_ (.A1(_02303_),
    .A2(_02307_),
    .A3(_02308_),
    .A4(_02310_),
    .ZN(_02311_));
 AND2_X4 _27553_ (.A1(_02273_),
    .A2(_02199_),
    .ZN(_02312_));
 BUF_X2 _27554_ (.A(_02312_),
    .Z(_02313_));
 NOR2_X4 _27555_ (.A1(_02172_),
    .A2(_02220_),
    .ZN(_02314_));
 NAND3_X1 _27556_ (.A1(_02313_),
    .A2(_02170_),
    .A3(_02314_),
    .ZN(_02315_));
 OAI211_X2 _27557_ (.A(_02279_),
    .B(_02268_),
    .C1(_02306_),
    .C2(_02286_),
    .ZN(_02316_));
 NOR2_X1 _27558_ (.A1(_02137_),
    .A2(_16807_),
    .ZN(_02317_));
 AND2_X2 _27559_ (.A1(_02317_),
    .A2(_16806_),
    .ZN(_02318_));
 NAND3_X1 _27560_ (.A1(_02318_),
    .A2(_02279_),
    .A3(_02268_),
    .ZN(_02319_));
 BUF_X4 _27561_ (.A(_02218_),
    .Z(_02320_));
 NAND3_X1 _27562_ (.A1(_02320_),
    .A2(_02279_),
    .A3(_02268_),
    .ZN(_02321_));
 NAND4_X1 _27563_ (.A1(_02315_),
    .A2(_02316_),
    .A3(_02319_),
    .A4(_02321_),
    .ZN(_02322_));
 NOR4_X1 _27564_ (.A1(_02288_),
    .A2(_02299_),
    .A3(_02311_),
    .A4(_02322_),
    .ZN(_02323_));
 BUF_X2 _27565_ (.A(_02130_),
    .Z(_02324_));
 NOR2_X4 _27566_ (.A1(_02272_),
    .A2(_16810_),
    .ZN(_02325_));
 BUF_X8 _27567_ (.A(_02325_),
    .Z(_02326_));
 AND2_X2 _27568_ (.A1(_02324_),
    .A2(_02326_),
    .ZN(_02327_));
 BUF_X2 _27569_ (.A(_02327_),
    .Z(_02328_));
 AND3_X1 _27570_ (.A1(_02328_),
    .A2(_02170_),
    .A3(_02264_),
    .ZN(_02329_));
 AOI21_X1 _27571_ (.A(_02329_),
    .B1(_02328_),
    .B2(_02251_),
    .ZN(_02330_));
 AND2_X2 _27572_ (.A1(_02179_),
    .A2(_02325_),
    .ZN(_02331_));
 AND2_X1 _27573_ (.A1(_02331_),
    .A2(_02257_),
    .ZN(_02332_));
 INV_X1 _27574_ (.A(_02332_),
    .ZN(_02333_));
 BUF_X4 _27575_ (.A(_02331_),
    .Z(_02334_));
 AND2_X2 _27576_ (.A1(_02138_),
    .A2(_02159_),
    .ZN(_02335_));
 OAI21_X1 _27577_ (.A(_02334_),
    .B1(_02335_),
    .B2(_02276_),
    .ZN(_02336_));
 INV_X1 _27578_ (.A(_02334_),
    .ZN(_02337_));
 INV_X1 _27579_ (.A(_02198_),
    .ZN(_02338_));
 OAI211_X2 _27580_ (.A(_02333_),
    .B(_02336_),
    .C1(_02337_),
    .C2(_02338_),
    .ZN(_02339_));
 INV_X1 _27581_ (.A(_02136_),
    .ZN(_02340_));
 NOR2_X1 _27582_ (.A1(_02340_),
    .A2(_02144_),
    .ZN(_02341_));
 AND2_X4 _27583_ (.A1(_02326_),
    .A2(_02199_),
    .ZN(_02342_));
 AND2_X1 _27584_ (.A1(_02341_),
    .A2(_02342_),
    .ZN(_02343_));
 NOR2_X1 _27585_ (.A1(_02188_),
    .A2(_02139_),
    .ZN(_02344_));
 AND2_X1 _27586_ (.A1(_02342_),
    .A2(_02344_),
    .ZN(_02345_));
 AND2_X4 _27587_ (.A1(_02151_),
    .A2(_02197_),
    .ZN(_02346_));
 BUF_X2 _27588_ (.A(_02326_),
    .Z(_02347_));
 AND3_X1 _27589_ (.A1(_02346_),
    .A2(_02347_),
    .A3(_02268_),
    .ZN(_02348_));
 NOR4_X1 _27590_ (.A1(_02339_),
    .A2(_02343_),
    .A3(_02345_),
    .A4(_02348_),
    .ZN(_02349_));
 BUF_X4 _27591_ (.A(_02137_),
    .Z(_02350_));
 AND4_X1 _27592_ (.A1(_02350_),
    .A2(_02347_),
    .A3(_02211_),
    .A4(_02280_),
    .ZN(_02351_));
 AND2_X2 _27593_ (.A1(_02326_),
    .A2(_02164_),
    .ZN(_02352_));
 BUF_X4 _27594_ (.A(_02352_),
    .Z(_02353_));
 AOI21_X1 _27595_ (.A(_02351_),
    .B1(_02353_),
    .B2(_02341_),
    .ZN(_02354_));
 OAI21_X1 _27596_ (.A(_02353_),
    .B1(_02314_),
    .B2(_02292_),
    .ZN(_02355_));
 AND4_X1 _27597_ (.A1(_02330_),
    .A2(_02349_),
    .A3(_02354_),
    .A4(_02355_),
    .ZN(_02356_));
 NAND4_X1 _27598_ (.A1(_02217_),
    .A2(_02271_),
    .A3(_02323_),
    .A4(_02356_),
    .ZN(_02357_));
 AND2_X1 _27599_ (.A1(_02145_),
    .A2(_02197_),
    .ZN(_02358_));
 BUF_X2 _27600_ (.A(_02358_),
    .Z(_02359_));
 AND2_X1 _27601_ (.A1(_02241_),
    .A2(_02359_),
    .ZN(_02360_));
 OR2_X2 _27602_ (.A1(_02357_),
    .A2(_02360_),
    .ZN(_02361_));
 XOR2_X2 _27603_ (.A(_02128_),
    .B(_02361_),
    .Z(_02362_));
 BUF_X32 _27604_ (.A(_16764_),
    .Z(_02363_));
 NOR2_X4 _27605_ (.A1(_16765_),
    .A2(_02363_),
    .ZN(_02364_));
 INV_X2 _27606_ (.A(_02364_),
    .ZN(_02365_));
 INV_X16 _27607_ (.A(_16767_),
    .ZN(_02366_));
 NOR2_X4 _27608_ (.A1(_02366_),
    .A2(_16766_),
    .ZN(_02367_));
 AND2_X4 _27609_ (.A1(_02365_),
    .A2(_02367_),
    .ZN(_02368_));
 AND2_X4 _27610_ (.A1(_16765_),
    .A2(_16764_),
    .ZN(_02369_));
 INV_X1 _27611_ (.A(_02369_),
    .ZN(_02370_));
 BUF_X4 _27612_ (.A(_02370_),
    .Z(_02371_));
 AND2_X4 _27613_ (.A1(_02368_),
    .A2(_02371_),
    .ZN(_02372_));
 INV_X32 _27614_ (.A(_16769_),
    .ZN(_02373_));
 AND2_X4 _27615_ (.A1(_02373_),
    .A2(_16768_),
    .ZN(_02374_));
 BUF_X8 _27616_ (.A(_02374_),
    .Z(_02375_));
 INV_X32 _27617_ (.A(_16771_),
    .ZN(_02376_));
 NOR2_X4 _27618_ (.A1(_02376_),
    .A2(_16770_),
    .ZN(_02377_));
 BUF_X8 _27619_ (.A(_02377_),
    .Z(_02378_));
 AND2_X4 _27620_ (.A1(_02375_),
    .A2(_02378_),
    .ZN(_02379_));
 BUF_X4 _27621_ (.A(_02379_),
    .Z(_02380_));
 AND2_X1 _27622_ (.A1(_02372_),
    .A2(_02380_),
    .ZN(_02381_));
 NOR2_X4 _27623_ (.A1(_16766_),
    .A2(_16767_),
    .ZN(_02382_));
 BUF_X4 _27624_ (.A(_02382_),
    .Z(_02383_));
 NAND4_X1 _27625_ (.A1(_02375_),
    .A2(_02378_),
    .A3(_02363_),
    .A4(_02383_),
    .ZN(_02384_));
 INV_X1 _27626_ (.A(_02379_),
    .ZN(_02385_));
 INV_X32 _27627_ (.A(_16766_),
    .ZN(_02386_));
 NOR2_X4 _27628_ (.A1(_02386_),
    .A2(_16767_),
    .ZN(_02387_));
 BUF_X32 _27629_ (.A(_16765_),
    .Z(_02388_));
 AND2_X4 _27630_ (.A1(_02387_),
    .A2(_02388_),
    .ZN(_02389_));
 BUF_X4 _27631_ (.A(_02389_),
    .Z(_02390_));
 INV_X1 _27632_ (.A(_02390_),
    .ZN(_02391_));
 OAI21_X1 _27633_ (.A(_02384_),
    .B1(_02385_),
    .B2(_02391_),
    .ZN(_02392_));
 AND2_X4 _27634_ (.A1(_16766_),
    .A2(_16767_),
    .ZN(_02393_));
 BUF_X4 _27635_ (.A(_02393_),
    .Z(_02394_));
 INV_X1 _27636_ (.A(_02394_),
    .ZN(_02395_));
 INV_X32 _27637_ (.A(_16765_),
    .ZN(_02396_));
 NOR2_X4 _27638_ (.A1(_02396_),
    .A2(_02363_),
    .ZN(_02397_));
 BUF_X4 _27639_ (.A(_02397_),
    .Z(_02398_));
 NOR2_X1 _27640_ (.A1(_02395_),
    .A2(_02398_),
    .ZN(_02399_));
 INV_X16 _27641_ (.A(_02363_),
    .ZN(_02400_));
 NOR2_X4 _27642_ (.A1(_02400_),
    .A2(_02388_),
    .ZN(_02401_));
 BUF_X8 _27643_ (.A(_02401_),
    .Z(_02402_));
 INV_X1 _27644_ (.A(_02402_),
    .ZN(_02403_));
 AND3_X1 _27645_ (.A1(_02380_),
    .A2(_02399_),
    .A3(_02403_),
    .ZN(_02404_));
 OR3_X1 _27646_ (.A1(_02381_),
    .A2(_02392_),
    .A3(_02404_),
    .ZN(_02405_));
 AND2_X4 _27647_ (.A1(_16771_),
    .A2(_16770_),
    .ZN(_02406_));
 AND2_X2 _27648_ (.A1(_02374_),
    .A2(_02406_),
    .ZN(_02407_));
 NOR3_X1 _27649_ (.A1(_02396_),
    .A2(_02363_),
    .A3(_16767_),
    .ZN(_02408_));
 AND2_X1 _27650_ (.A1(_02407_),
    .A2(_02408_),
    .ZN(_02409_));
 AND2_X4 _27651_ (.A1(_02393_),
    .A2(_02388_),
    .ZN(_02410_));
 NOR2_X4 _27652_ (.A1(_16769_),
    .A2(_16768_),
    .ZN(_02411_));
 AND2_X4 _27653_ (.A1(_02406_),
    .A2(_02411_),
    .ZN(_02412_));
 BUF_X8 _27654_ (.A(_02412_),
    .Z(_02413_));
 AND2_X2 _27655_ (.A1(_02378_),
    .A2(_02411_),
    .ZN(_02414_));
 AND2_X2 _27656_ (.A1(_02369_),
    .A2(_02382_),
    .ZN(_02415_));
 BUF_X8 _27657_ (.A(_02415_),
    .Z(_02416_));
 INV_X4 _27658_ (.A(_02416_),
    .ZN(_02417_));
 AND2_X2 _27659_ (.A1(_02364_),
    .A2(_02382_),
    .ZN(_02418_));
 BUF_X8 _27660_ (.A(_02418_),
    .Z(_02419_));
 INV_X4 _27661_ (.A(_02419_),
    .ZN(_02420_));
 NAND2_X4 _27662_ (.A1(_02417_),
    .A2(_02420_),
    .ZN(_02421_));
 AOI221_X1 _27663_ (.A(_02409_),
    .B1(_02410_),
    .B2(_02413_),
    .C1(_02414_),
    .C2(_02421_),
    .ZN(_02422_));
 AND2_X2 _27664_ (.A1(_02393_),
    .A2(_02369_),
    .ZN(_02423_));
 INV_X2 _27665_ (.A(_02423_),
    .ZN(_02424_));
 AND2_X4 _27666_ (.A1(_02393_),
    .A2(_02364_),
    .ZN(_02425_));
 INV_X1 _27667_ (.A(_02425_),
    .ZN(_02426_));
 NAND2_X1 _27668_ (.A1(_02424_),
    .A2(_02426_),
    .ZN(_02427_));
 NOR2_X4 _27669_ (.A1(_02373_),
    .A2(_16768_),
    .ZN(_02428_));
 BUF_X4 _27670_ (.A(_02428_),
    .Z(_02429_));
 AND2_X2 _27671_ (.A1(_02429_),
    .A2(_02406_),
    .ZN(_02430_));
 BUF_X4 _27672_ (.A(_02430_),
    .Z(_02431_));
 NAND2_X1 _27673_ (.A1(_02427_),
    .A2(_02431_),
    .ZN(_02432_));
 AND2_X2 _27674_ (.A1(_02367_),
    .A2(_02396_),
    .ZN(_02433_));
 BUF_X2 _27675_ (.A(_02433_),
    .Z(_02434_));
 BUF_X4 _27676_ (.A(_02413_),
    .Z(_02435_));
 OAI21_X1 _27677_ (.A(_02434_),
    .B1(_02414_),
    .B2(_02435_),
    .ZN(_02436_));
 BUF_X8 _27678_ (.A(_02387_),
    .Z(_02437_));
 AND2_X4 _27679_ (.A1(_02437_),
    .A2(_02363_),
    .ZN(_02438_));
 BUF_X4 _27680_ (.A(_02438_),
    .Z(_02439_));
 AND2_X1 _27681_ (.A1(_02382_),
    .A2(_02396_),
    .ZN(_02440_));
 BUF_X4 _27682_ (.A(_02440_),
    .Z(_02441_));
 OAI21_X1 _27683_ (.A(_02431_),
    .B1(_02439_),
    .B2(_02441_),
    .ZN(_02442_));
 NAND4_X1 _27684_ (.A1(_02422_),
    .A2(_02432_),
    .A3(_02436_),
    .A4(_02442_),
    .ZN(_02443_));
 AND2_X1 _27685_ (.A1(_02393_),
    .A2(_02396_),
    .ZN(_02444_));
 BUF_X2 _27686_ (.A(_02444_),
    .Z(_02445_));
 NOR2_X4 _27687_ (.A1(_16771_),
    .A2(_16770_),
    .ZN(_02446_));
 AND2_X1 _27688_ (.A1(_02446_),
    .A2(_02411_),
    .ZN(_02447_));
 BUF_X2 _27689_ (.A(_02447_),
    .Z(_02448_));
 BUF_X4 _27690_ (.A(_02448_),
    .Z(_02449_));
 AND2_X1 _27691_ (.A1(_02445_),
    .A2(_02449_),
    .ZN(_02450_));
 AND2_X4 _27692_ (.A1(_02374_),
    .A2(_02446_),
    .ZN(_02451_));
 AND2_X1 _27693_ (.A1(_02451_),
    .A2(_02444_),
    .ZN(_02452_));
 INV_X4 _27694_ (.A(_02451_),
    .ZN(_02453_));
 AND2_X2 _27695_ (.A1(_02397_),
    .A2(_02382_),
    .ZN(_02454_));
 INV_X2 _27696_ (.A(_02454_),
    .ZN(_02455_));
 AOI21_X2 _27697_ (.A(_02453_),
    .B1(_02424_),
    .B2(_02455_),
    .ZN(_02456_));
 AND2_X1 _27698_ (.A1(_02367_),
    .A2(_02388_),
    .ZN(_02457_));
 AOI211_X2 _27699_ (.A(_02452_),
    .B(_02456_),
    .C1(_02457_),
    .C2(_02451_),
    .ZN(_02458_));
 AND2_X4 _27700_ (.A1(_02376_),
    .A2(_16770_),
    .ZN(_02459_));
 AND2_X4 _27701_ (.A1(_16769_),
    .A2(_16768_),
    .ZN(_02460_));
 AND2_X4 _27702_ (.A1(_02459_),
    .A2(_02460_),
    .ZN(_02461_));
 BUF_X4 _27703_ (.A(_02461_),
    .Z(_02462_));
 AND2_X2 _27704_ (.A1(_02437_),
    .A2(_02396_),
    .ZN(_02463_));
 AND2_X2 _27705_ (.A1(_02459_),
    .A2(_02428_),
    .ZN(_02464_));
 CLKBUF_X3 _27706_ (.A(_02464_),
    .Z(_02465_));
 BUF_X4 _27707_ (.A(_02410_),
    .Z(_02466_));
 AOI22_X1 _27708_ (.A1(_02462_),
    .A2(_02463_),
    .B1(_02465_),
    .B2(_02466_),
    .ZN(_02467_));
 INV_X1 _27709_ (.A(_02382_),
    .ZN(_02468_));
 INV_X2 _27710_ (.A(_02464_),
    .ZN(_02469_));
 OAI211_X2 _27711_ (.A(_02458_),
    .B(_02467_),
    .C1(_02468_),
    .C2(_02469_),
    .ZN(_02470_));
 OR4_X4 _27712_ (.A1(_02405_),
    .A2(_02443_),
    .A3(_02450_),
    .A4(_02470_),
    .ZN(_02471_));
 BUF_X2 _27713_ (.A(_02406_),
    .Z(_02472_));
 AND3_X1 _27714_ (.A1(_02399_),
    .A2(_02375_),
    .A3(_02472_),
    .ZN(_02473_));
 AND2_X2 _27715_ (.A1(_02378_),
    .A2(_02460_),
    .ZN(_02474_));
 NAND2_X1 _27716_ (.A1(_02457_),
    .A2(_02474_),
    .ZN(_02475_));
 AND2_X2 _27717_ (.A1(_02397_),
    .A2(_02393_),
    .ZN(_02476_));
 BUF_X4 _27718_ (.A(_02476_),
    .Z(_02477_));
 NAND2_X1 _27719_ (.A1(_02477_),
    .A2(_02474_),
    .ZN(_02478_));
 NAND2_X1 _27720_ (.A1(_02475_),
    .A2(_02478_),
    .ZN(_02479_));
 AND2_X1 _27721_ (.A1(_02474_),
    .A2(_02463_),
    .ZN(_02480_));
 AND2_X2 _27722_ (.A1(_02437_),
    .A2(_02369_),
    .ZN(_02481_));
 AND2_X1 _27723_ (.A1(_02481_),
    .A2(_02474_),
    .ZN(_02482_));
 OR4_X4 _27724_ (.A1(_02473_),
    .A2(_02479_),
    .A3(_02480_),
    .A4(_02482_),
    .ZN(_02483_));
 INV_X1 _27725_ (.A(_02481_),
    .ZN(_02484_));
 AND2_X2 _27726_ (.A1(_02387_),
    .A2(_02364_),
    .ZN(_02485_));
 INV_X1 _27727_ (.A(_02485_),
    .ZN(_02486_));
 NAND2_X1 _27728_ (.A1(_02484_),
    .A2(_02486_),
    .ZN(_02487_));
 OAI21_X1 _27729_ (.A(_02449_),
    .B1(_02487_),
    .B2(_02477_),
    .ZN(_02488_));
 INV_X2 _27730_ (.A(_02462_),
    .ZN(_02489_));
 BUF_X2 _27731_ (.A(_02394_),
    .Z(_02490_));
 NAND2_X1 _27732_ (.A1(_02365_),
    .A2(_02490_),
    .ZN(_02491_));
 OAI21_X1 _27733_ (.A(_02488_),
    .B1(_02489_),
    .B2(_02491_),
    .ZN(_02492_));
 INV_X1 _27734_ (.A(_02433_),
    .ZN(_02493_));
 AND2_X2 _27735_ (.A1(_02428_),
    .A2(_02446_),
    .ZN(_02494_));
 INV_X1 _27736_ (.A(_02494_),
    .ZN(_02495_));
 NOR2_X1 _27737_ (.A1(_02468_),
    .A2(_02369_),
    .ZN(_02496_));
 INV_X1 _27738_ (.A(_02496_),
    .ZN(_02497_));
 OAI22_X1 _27739_ (.A1(_02489_),
    .A2(_02493_),
    .B1(_02495_),
    .B2(_02497_),
    .ZN(_02498_));
 BUF_X4 _27740_ (.A(_02367_),
    .Z(_02499_));
 AND2_X4 _27741_ (.A1(_02499_),
    .A2(_02398_),
    .ZN(_02500_));
 AND2_X1 _27742_ (.A1(_02462_),
    .A2(_02500_),
    .ZN(_02501_));
 OR2_X1 _27743_ (.A1(_02498_),
    .A2(_02501_),
    .ZN(_02502_));
 AND2_X1 _27744_ (.A1(_02460_),
    .A2(_02446_),
    .ZN(_02503_));
 BUF_X4 _27745_ (.A(_02503_),
    .Z(_02504_));
 BUF_X2 _27746_ (.A(_02457_),
    .Z(_02505_));
 BUF_X4 _27747_ (.A(_02400_),
    .Z(_02506_));
 AND2_X1 _27748_ (.A1(_02394_),
    .A2(_02506_),
    .ZN(_02507_));
 OAI21_X1 _27749_ (.A(_02504_),
    .B1(_02505_),
    .B2(_02507_),
    .ZN(_02508_));
 NOR3_X2 _27750_ (.A1(_02364_),
    .A2(_02386_),
    .A3(_16767_),
    .ZN(_02509_));
 OAI21_X1 _27751_ (.A(_02413_),
    .B1(_02509_),
    .B2(_02419_),
    .ZN(_02510_));
 NAND2_X1 _27752_ (.A1(_02368_),
    .A2(_02494_),
    .ZN(_02511_));
 NOR3_X1 _27753_ (.A1(_02402_),
    .A2(_16766_),
    .A3(_02366_),
    .ZN(_02512_));
 NAND2_X1 _27754_ (.A1(_02512_),
    .A2(_02431_),
    .ZN(_02513_));
 NAND4_X1 _27755_ (.A1(_02508_),
    .A2(_02510_),
    .A3(_02511_),
    .A4(_02513_),
    .ZN(_02514_));
 NOR4_X4 _27756_ (.A1(_02483_),
    .A2(_02492_),
    .A3(_02502_),
    .A4(_02514_),
    .ZN(_02515_));
 BUF_X4 _27757_ (.A(_02451_),
    .Z(_02516_));
 AND2_X1 _27758_ (.A1(_02487_),
    .A2(_02516_),
    .ZN(_02517_));
 INV_X1 _27759_ (.A(_02517_),
    .ZN(_02518_));
 AND2_X1 _27760_ (.A1(_02389_),
    .A2(_02494_),
    .ZN(_02519_));
 AND2_X2 _27761_ (.A1(_02451_),
    .A2(_02440_),
    .ZN(_02520_));
 AOI211_X4 _27762_ (.A(_02519_),
    .B(_02520_),
    .C1(_02451_),
    .C2(_02433_),
    .ZN(_02521_));
 BUF_X4 _27763_ (.A(_02504_),
    .Z(_02522_));
 AND2_X4 _27764_ (.A1(_02460_),
    .A2(_02406_),
    .ZN(_02523_));
 BUF_X8 _27765_ (.A(_02523_),
    .Z(_02524_));
 BUF_X4 _27766_ (.A(_02524_),
    .Z(_02525_));
 AOI22_X1 _27767_ (.A1(_02522_),
    .A2(_02439_),
    .B1(_02525_),
    .B2(_02507_),
    .ZN(_02526_));
 BUF_X4 _27768_ (.A(_02463_),
    .Z(_02527_));
 AND2_X2 _27769_ (.A1(_02382_),
    .A2(_02363_),
    .ZN(_02528_));
 AOI22_X1 _27770_ (.A1(_02527_),
    .A2(_02525_),
    .B1(_02522_),
    .B2(_02528_),
    .ZN(_02529_));
 AND4_X2 _27771_ (.A1(_02518_),
    .A2(_02521_),
    .A3(_02526_),
    .A4(_02529_),
    .ZN(_02530_));
 AND2_X2 _27772_ (.A1(_02459_),
    .A2(_02374_),
    .ZN(_02531_));
 BUF_X2 _27773_ (.A(_02531_),
    .Z(_02532_));
 OAI21_X1 _27774_ (.A(_02532_),
    .B1(_02372_),
    .B2(_02423_),
    .ZN(_02533_));
 BUF_X4 _27775_ (.A(_02459_),
    .Z(_02534_));
 BUF_X4 _27776_ (.A(_02363_),
    .Z(_02535_));
 NAND4_X1 _27777_ (.A1(_02534_),
    .A2(_02375_),
    .A3(_02535_),
    .A4(_02383_),
    .ZN(_02536_));
 AND2_X4 _27778_ (.A1(_02401_),
    .A2(_02387_),
    .ZN(_02537_));
 BUF_X8 _27779_ (.A(_02537_),
    .Z(_02538_));
 AND2_X2 _27780_ (.A1(_02398_),
    .A2(_02437_),
    .ZN(_02539_));
 OAI21_X1 _27781_ (.A(_02531_),
    .B1(_02538_),
    .B2(_02539_),
    .ZN(_02540_));
 AND3_X1 _27782_ (.A1(_02533_),
    .A2(_02536_),
    .A3(_02540_),
    .ZN(_02541_));
 AND2_X1 _27783_ (.A1(_02459_),
    .A2(_02411_),
    .ZN(_02542_));
 INV_X1 _27784_ (.A(_02542_),
    .ZN(_02543_));
 INV_X1 _27785_ (.A(_02457_),
    .ZN(_02544_));
 AND2_X2 _27786_ (.A1(_02393_),
    .A2(_02363_),
    .ZN(_02545_));
 INV_X1 _27787_ (.A(_02545_),
    .ZN(_02546_));
 AOI21_X1 _27788_ (.A(_02543_),
    .B1(_02544_),
    .B2(_02546_),
    .ZN(_02547_));
 BUF_X4 _27789_ (.A(_02542_),
    .Z(_02548_));
 AND2_X4 _27790_ (.A1(_02402_),
    .A2(_02382_),
    .ZN(_02549_));
 INV_X1 _27791_ (.A(_02549_),
    .ZN(_02550_));
 NAND2_X1 _27792_ (.A1(_02484_),
    .A2(_02550_),
    .ZN(_02551_));
 AOI21_X1 _27793_ (.A(_02547_),
    .B1(_02548_),
    .B2(_02551_),
    .ZN(_02552_));
 BUF_X4 _27794_ (.A(_02378_),
    .Z(_02553_));
 NAND3_X1 _27795_ (.A1(_02445_),
    .A2(_02553_),
    .A3(_02429_),
    .ZN(_02554_));
 AND2_X2 _27796_ (.A1(_02377_),
    .A2(_02428_),
    .ZN(_02555_));
 BUF_X2 _27797_ (.A(_02555_),
    .Z(_02556_));
 BUF_X4 _27798_ (.A(_02474_),
    .Z(_02557_));
 AOI22_X1 _27799_ (.A1(_02434_),
    .A2(_02556_),
    .B1(_02557_),
    .B2(_02441_),
    .ZN(_02558_));
 AND4_X1 _27800_ (.A1(_02541_),
    .A2(_02552_),
    .A3(_02554_),
    .A4(_02558_),
    .ZN(_02559_));
 AND2_X4 _27801_ (.A1(_02367_),
    .A2(_02402_),
    .ZN(_02560_));
 AND2_X1 _27802_ (.A1(_02560_),
    .A2(_02524_),
    .ZN(_02561_));
 AOI221_X1 _27803_ (.A(_02561_),
    .B1(_02481_),
    .B2(_02464_),
    .C1(_02524_),
    .C2(_02496_),
    .ZN(_02562_));
 AND2_X1 _27804_ (.A1(_02555_),
    .A2(_02476_),
    .ZN(_02563_));
 AND2_X4 _27805_ (.A1(_02402_),
    .A2(_02394_),
    .ZN(_02564_));
 AOI221_X4 _27806_ (.A(_02563_),
    .B1(_02564_),
    .B2(_02413_),
    .C1(_02555_),
    .C2(_02419_),
    .ZN(_02565_));
 NAND2_X1 _27807_ (.A1(_02464_),
    .A2(_02560_),
    .ZN(_02566_));
 NAND2_X1 _27808_ (.A1(_02462_),
    .A2(_02528_),
    .ZN(_02567_));
 NAND2_X1 _27809_ (.A1(_02462_),
    .A2(_02481_),
    .ZN(_02568_));
 NAND2_X1 _27810_ (.A1(_02494_),
    .A2(_02564_),
    .ZN(_02569_));
 AND4_X1 _27811_ (.A1(_02566_),
    .A2(_02567_),
    .A3(_02568_),
    .A4(_02569_),
    .ZN(_02570_));
 AND2_X4 _27812_ (.A1(_02367_),
    .A2(_02369_),
    .ZN(_02571_));
 BUF_X4 _27813_ (.A(_02571_),
    .Z(_02572_));
 AND2_X1 _27814_ (.A1(_02407_),
    .A2(_02572_),
    .ZN(_02573_));
 AND2_X1 _27815_ (.A1(_02500_),
    .A2(_02555_),
    .ZN(_02574_));
 AND2_X1 _27816_ (.A1(_02538_),
    .A2(_02414_),
    .ZN(_02575_));
 AND3_X1 _27817_ (.A1(_02408_),
    .A2(_02429_),
    .A3(_02472_),
    .ZN(_02576_));
 NOR4_X1 _27818_ (.A1(_02573_),
    .A2(_02574_),
    .A3(_02575_),
    .A4(_02576_),
    .ZN(_02577_));
 AND4_X2 _27819_ (.A1(_02562_),
    .A2(_02565_),
    .A3(_02570_),
    .A4(_02577_),
    .ZN(_02578_));
 NAND4_X4 _27820_ (.A1(_02515_),
    .A2(_02530_),
    .A3(_02559_),
    .A4(_02578_),
    .ZN(_02579_));
 NOR2_X4 _27821_ (.A1(_02471_),
    .A2(_02579_),
    .ZN(_02580_));
 BUF_X4 _27822_ (.A(_02437_),
    .Z(_02581_));
 OAI21_X1 _27823_ (.A(_02465_),
    .B1(_02528_),
    .B2(_02581_),
    .ZN(_02582_));
 NAND2_X1 _27824_ (.A1(_02531_),
    .A2(_02416_),
    .ZN(_02583_));
 NAND3_X1 _27825_ (.A1(_02440_),
    .A2(_02459_),
    .A3(_02375_),
    .ZN(_02584_));
 NAND2_X1 _27826_ (.A1(_02583_),
    .A2(_02584_),
    .ZN(_02585_));
 AND2_X1 _27827_ (.A1(_02367_),
    .A2(_02363_),
    .ZN(_02586_));
 OAI21_X2 _27828_ (.A(_02531_),
    .B1(_02586_),
    .B2(_02423_),
    .ZN(_02587_));
 NAND3_X1 _27829_ (.A1(_02485_),
    .A2(_02459_),
    .A3(_02411_),
    .ZN(_02588_));
 INV_X1 _27830_ (.A(_02440_),
    .ZN(_02589_));
 OAI211_X2 _27831_ (.A(_02587_),
    .B(_02588_),
    .C1(_02589_),
    .C2(_02543_),
    .ZN(_02590_));
 NOR3_X1 _27832_ (.A1(_02398_),
    .A2(_16766_),
    .A3(_02366_),
    .ZN(_02591_));
 AOI211_X2 _27833_ (.A(_02585_),
    .B(_02590_),
    .C1(_02465_),
    .C2(_02591_),
    .ZN(_02592_));
 BUF_X2 _27834_ (.A(_02460_),
    .Z(_02593_));
 NAND3_X1 _27835_ (.A1(_02439_),
    .A2(_02534_),
    .A3(_02593_),
    .ZN(_02594_));
 NAND2_X1 _27836_ (.A1(_02462_),
    .A2(_02416_),
    .ZN(_02595_));
 AND2_X1 _27837_ (.A1(_02594_),
    .A2(_02595_),
    .ZN(_02596_));
 INV_X1 _27838_ (.A(_02437_),
    .ZN(_02597_));
 BUF_X4 _27839_ (.A(_02398_),
    .Z(_02598_));
 NOR2_X1 _27840_ (.A1(_02597_),
    .A2(_02598_),
    .ZN(_02599_));
 NAND2_X1 _27841_ (.A1(_02599_),
    .A2(_02414_),
    .ZN(_02600_));
 AND4_X1 _27842_ (.A1(_02582_),
    .A2(_02592_),
    .A3(_02596_),
    .A4(_02600_),
    .ZN(_02601_));
 NOR2_X2 _27843_ (.A1(_02468_),
    .A2(_02402_),
    .ZN(_02602_));
 AND2_X1 _27844_ (.A1(_02474_),
    .A2(_02602_),
    .ZN(_02603_));
 OAI21_X2 _27845_ (.A(_02462_),
    .B1(_02477_),
    .B2(_02564_),
    .ZN(_02604_));
 NAND3_X1 _27846_ (.A1(_02571_),
    .A2(_02534_),
    .A3(_02593_),
    .ZN(_02605_));
 INV_X1 _27847_ (.A(_02555_),
    .ZN(_02606_));
 INV_X1 _27848_ (.A(_02397_),
    .ZN(_02607_));
 AOI22_X1 _27849_ (.A1(_02607_),
    .A2(_02394_),
    .B1(_02499_),
    .B2(_02402_),
    .ZN(_02608_));
 OAI211_X2 _27850_ (.A(_02604_),
    .B(_02605_),
    .C1(_02606_),
    .C2(_02608_),
    .ZN(_02609_));
 BUF_X4 _27851_ (.A(_02414_),
    .Z(_02610_));
 AND2_X1 _27852_ (.A1(_02382_),
    .A2(_02400_),
    .ZN(_02611_));
 OR4_X1 _27853_ (.A1(_02410_),
    .A2(_02586_),
    .A3(_02545_),
    .A4(_02611_),
    .ZN(_02612_));
 AOI211_X2 _27854_ (.A(_02603_),
    .B(_02609_),
    .C1(_02610_),
    .C2(_02612_),
    .ZN(_02613_));
 CLKBUF_X3 _27855_ (.A(_02494_),
    .Z(_02614_));
 AND2_X1 _27856_ (.A1(_02509_),
    .A2(_02371_),
    .ZN(_02615_));
 OAI21_X1 _27857_ (.A(_02614_),
    .B1(_02615_),
    .B2(_02507_),
    .ZN(_02616_));
 OAI21_X1 _27858_ (.A(_02431_),
    .B1(_02421_),
    .B2(_02463_),
    .ZN(_02617_));
 AND2_X1 _27859_ (.A1(_02382_),
    .A2(_02388_),
    .ZN(_02618_));
 BUF_X4 _27860_ (.A(_02618_),
    .Z(_02619_));
 AOI22_X1 _27861_ (.A1(_02516_),
    .A2(_02619_),
    .B1(_02390_),
    .B2(_02448_),
    .ZN(_02620_));
 BUF_X4 _27862_ (.A(_02364_),
    .Z(_02621_));
 NOR3_X1 _27863_ (.A1(_02468_),
    .A2(_02369_),
    .A3(_02621_),
    .ZN(_02622_));
 OAI21_X1 _27864_ (.A(_02380_),
    .B1(_02622_),
    .B2(_02466_),
    .ZN(_02623_));
 AND4_X1 _27865_ (.A1(_02616_),
    .A2(_02617_),
    .A3(_02620_),
    .A4(_02623_),
    .ZN(_02624_));
 AOI22_X1 _27866_ (.A1(_02556_),
    .A2(_02485_),
    .B1(_02474_),
    .B2(_02425_),
    .ZN(_02625_));
 NAND2_X1 _27867_ (.A1(_02448_),
    .A2(_02619_),
    .ZN(_02626_));
 NAND2_X1 _27868_ (.A1(_02423_),
    .A2(_02504_),
    .ZN(_02627_));
 NAND3_X1 _27869_ (.A1(_02625_),
    .A2(_02626_),
    .A3(_02627_),
    .ZN(_02628_));
 NAND2_X1 _27870_ (.A1(_02494_),
    .A2(_02423_),
    .ZN(_02629_));
 NAND2_X1 _27871_ (.A1(_02560_),
    .A2(_02413_),
    .ZN(_02630_));
 INV_X1 _27872_ (.A(_02476_),
    .ZN(_02631_));
 OAI211_X2 _27873_ (.A(_02629_),
    .B(_02630_),
    .C1(_02469_),
    .C2(_02631_),
    .ZN(_02632_));
 NOR4_X1 _27874_ (.A1(_02628_),
    .A2(_02632_),
    .A3(_02480_),
    .A4(_02482_),
    .ZN(_02633_));
 AND4_X1 _27875_ (.A1(_02601_),
    .A2(_02613_),
    .A3(_02624_),
    .A4(_02633_),
    .ZN(_02634_));
 NOR2_X4 _27876_ (.A1(_02477_),
    .A2(_02564_),
    .ZN(_02635_));
 AND2_X1 _27877_ (.A1(_02635_),
    .A2(_02544_),
    .ZN(_02636_));
 INV_X1 _27878_ (.A(_02636_),
    .ZN(_02637_));
 INV_X1 _27879_ (.A(_02499_),
    .ZN(_02638_));
 AOI21_X1 _27880_ (.A(_02403_),
    .B1(_02638_),
    .B2(_02597_),
    .ZN(_02639_));
 OAI21_X1 _27881_ (.A(_02449_),
    .B1(_02637_),
    .B2(_02639_),
    .ZN(_02640_));
 AND2_X1 _27882_ (.A1(_02494_),
    .A2(_02496_),
    .ZN(_02641_));
 INV_X1 _27883_ (.A(_02524_),
    .ZN(_02642_));
 AOI21_X1 _27884_ (.A(_02642_),
    .B1(_02631_),
    .B2(_02486_),
    .ZN(_02643_));
 AND2_X2 _27885_ (.A1(_02571_),
    .A2(_02413_),
    .ZN(_02644_));
 AND2_X4 _27886_ (.A1(_02549_),
    .A2(_02524_),
    .ZN(_02645_));
 OR4_X2 _27887_ (.A1(_02641_),
    .A2(_02643_),
    .A3(_02644_),
    .A4(_02645_),
    .ZN(_02646_));
 AND2_X1 _27888_ (.A1(_02512_),
    .A2(_02607_),
    .ZN(_02647_));
 OAI21_X1 _27889_ (.A(_02516_),
    .B1(_02647_),
    .B2(_02615_),
    .ZN(_02648_));
 NAND2_X1 _27890_ (.A1(_02504_),
    .A2(_02445_),
    .ZN(_02649_));
 AND2_X1 _27891_ (.A1(_02499_),
    .A2(_02621_),
    .ZN(_02650_));
 OAI21_X1 _27892_ (.A(_02504_),
    .B1(_02539_),
    .B2(_02650_),
    .ZN(_02651_));
 NAND3_X1 _27893_ (.A1(_02648_),
    .A2(_02649_),
    .A3(_02651_),
    .ZN(_02652_));
 AND3_X1 _27894_ (.A1(_02370_),
    .A2(_02472_),
    .A3(_02411_),
    .ZN(_02653_));
 OAI21_X1 _27895_ (.A(_02653_),
    .B1(_02490_),
    .B2(_02619_),
    .ZN(_02654_));
 NAND2_X1 _27896_ (.A1(_02531_),
    .A2(_02390_),
    .ZN(_02655_));
 OAI211_X2 _27897_ (.A(_02654_),
    .B(_02655_),
    .C1(_02489_),
    .C2(_02589_),
    .ZN(_02656_));
 INV_X1 _27898_ (.A(_02504_),
    .ZN(_02657_));
 NOR2_X1 _27899_ (.A1(_02468_),
    .A2(_02621_),
    .ZN(_02658_));
 INV_X1 _27900_ (.A(_02658_),
    .ZN(_02659_));
 OAI211_X2 _27901_ (.A(_02511_),
    .B(_02513_),
    .C1(_02657_),
    .C2(_02659_),
    .ZN(_02660_));
 NOR4_X2 _27902_ (.A1(_02646_),
    .A2(_02652_),
    .A3(_02656_),
    .A4(_02660_),
    .ZN(_02661_));
 BUF_X4 _27903_ (.A(_02407_),
    .Z(_02662_));
 OAI21_X1 _27904_ (.A(_02662_),
    .B1(_02538_),
    .B2(_02454_),
    .ZN(_02663_));
 BUF_X4 _27905_ (.A(_02396_),
    .Z(_02664_));
 AOI21_X1 _27906_ (.A(_16766_),
    .B1(_02664_),
    .B2(_02366_),
    .ZN(_02665_));
 AOI22_X1 _27907_ (.A1(_02431_),
    .A2(_02545_),
    .B1(_02525_),
    .B2(_02665_),
    .ZN(_02666_));
 OAI21_X1 _27908_ (.A(_02407_),
    .B1(_02505_),
    .B2(_02433_),
    .ZN(_02667_));
 OAI21_X1 _27909_ (.A(_02407_),
    .B1(_02477_),
    .B2(_02564_),
    .ZN(_02668_));
 AND4_X1 _27910_ (.A1(_02663_),
    .A2(_02666_),
    .A3(_02667_),
    .A4(_02668_),
    .ZN(_02669_));
 AND2_X4 _27911_ (.A1(_02419_),
    .A2(_02448_),
    .ZN(_02670_));
 INV_X1 _27912_ (.A(_02670_),
    .ZN(_02671_));
 BUF_X4 _27913_ (.A(_02534_),
    .Z(_02672_));
 NAND4_X1 _27914_ (.A1(_02672_),
    .A2(_02499_),
    .A3(_02535_),
    .A4(_02411_),
    .ZN(_02673_));
 OAI21_X1 _27915_ (.A(_02548_),
    .B1(_02477_),
    .B2(_02445_),
    .ZN(_02674_));
 AND3_X1 _27916_ (.A1(_02671_),
    .A2(_02673_),
    .A3(_02674_),
    .ZN(_02675_));
 AND4_X2 _27917_ (.A1(_02640_),
    .A2(_02661_),
    .A3(_02669_),
    .A4(_02675_),
    .ZN(_02676_));
 AND2_X4 _27918_ (.A1(_02634_),
    .A2(_02676_),
    .ZN(_02677_));
 XNOR2_X2 _27919_ (.A(_02580_),
    .B(_02677_),
    .ZN(_02678_));
 XNOR2_X1 _27920_ (.A(_02362_),
    .B(_02678_),
    .ZN(_02679_));
 INV_X32 _27921_ (.A(_16859_),
    .ZN(_02680_));
 AND2_X4 _27922_ (.A1(_02680_),
    .A2(_16858_),
    .ZN(_02681_));
 AND2_X4 _27923_ (.A1(_16857_),
    .A2(_16856_),
    .ZN(_02682_));
 BUF_X8 _27924_ (.A(_02682_),
    .Z(_02683_));
 AND2_X4 _27925_ (.A1(_02681_),
    .A2(_02683_),
    .ZN(_02684_));
 INV_X32 _27926_ (.A(_16853_),
    .ZN(_02685_));
 BUF_X32 _27927_ (.A(_16852_),
    .Z(_02686_));
 NOR2_X4 _27928_ (.A1(_02685_),
    .A2(_02686_),
    .ZN(_02687_));
 INV_X32 _27929_ (.A(_16855_),
    .ZN(_02688_));
 NOR2_X4 _27930_ (.A1(_02688_),
    .A2(_16854_),
    .ZN(_02689_));
 BUF_X4 _27931_ (.A(_02689_),
    .Z(_02690_));
 AND2_X1 _27932_ (.A1(_02687_),
    .A2(_02690_),
    .ZN(_02691_));
 AND2_X1 _27933_ (.A1(_02684_),
    .A2(_02691_),
    .ZN(_02692_));
 INV_X1 _27934_ (.A(_02692_),
    .ZN(_02693_));
 AND2_X1 _27935_ (.A1(_02689_),
    .A2(_02685_),
    .ZN(_02694_));
 AND2_X1 _27936_ (.A1(_02684_),
    .A2(_02694_),
    .ZN(_02695_));
 INV_X1 _27937_ (.A(_02695_),
    .ZN(_02696_));
 BUF_X4 _27938_ (.A(_02684_),
    .Z(_02697_));
 INV_X32 _27939_ (.A(_16852_),
    .ZN(_02698_));
 NOR2_X4 _27940_ (.A1(_02698_),
    .A2(_16853_),
    .ZN(_02699_));
 AND2_X4 _27941_ (.A1(_16854_),
    .A2(_16855_),
    .ZN(_02700_));
 AND2_X1 _27942_ (.A1(_02699_),
    .A2(_02700_),
    .ZN(_02701_));
 BUF_X2 _27943_ (.A(_02701_),
    .Z(_02702_));
 AND2_X2 _27944_ (.A1(_02700_),
    .A2(_16853_),
    .ZN(_02703_));
 BUF_X4 _27945_ (.A(_02703_),
    .Z(_02704_));
 OAI21_X1 _27946_ (.A(_02697_),
    .B1(_02702_),
    .B2(_02704_),
    .ZN(_02705_));
 AND3_X1 _27947_ (.A1(_02693_),
    .A2(_02696_),
    .A3(_02705_),
    .ZN(_02706_));
 INV_X4 _27948_ (.A(_16854_),
    .ZN(_02707_));
 NOR2_X4 _27949_ (.A1(_02707_),
    .A2(_16855_),
    .ZN(_02708_));
 AND2_X4 _27950_ (.A1(_02686_),
    .A2(_16853_),
    .ZN(_02709_));
 AND2_X4 _27951_ (.A1(_02708_),
    .A2(_02709_),
    .ZN(_02710_));
 NAND2_X1 _27952_ (.A1(_02697_),
    .A2(_02710_),
    .ZN(_02711_));
 BUF_X4 _27953_ (.A(_02699_),
    .Z(_02712_));
 NOR2_X4 _27954_ (.A1(_16854_),
    .A2(_16855_),
    .ZN(_02713_));
 BUF_X4 _27955_ (.A(_02713_),
    .Z(_02714_));
 AND2_X2 _27956_ (.A1(_02712_),
    .A2(_02714_),
    .ZN(_02715_));
 NAND2_X1 _27957_ (.A1(_02697_),
    .A2(_02715_),
    .ZN(_02716_));
 AND2_X4 _27958_ (.A1(_02709_),
    .A2(_02713_),
    .ZN(_02717_));
 NAND2_X1 _27959_ (.A1(_02684_),
    .A2(_02717_),
    .ZN(_02718_));
 AND2_X2 _27960_ (.A1(_02708_),
    .A2(_02685_),
    .ZN(_02719_));
 NAND2_X1 _27961_ (.A1(_02684_),
    .A2(_02719_),
    .ZN(_02720_));
 AND4_X1 _27962_ (.A1(_02711_),
    .A2(_02716_),
    .A3(_02718_),
    .A4(_02720_),
    .ZN(_02721_));
 INV_X32 _27963_ (.A(_16857_),
    .ZN(_02722_));
 NOR2_X1 _27964_ (.A1(_02722_),
    .A2(_16856_),
    .ZN(_02723_));
 BUF_X2 _27965_ (.A(_02723_),
    .Z(_02724_));
 AND2_X1 _27966_ (.A1(_02681_),
    .A2(_02724_),
    .ZN(_02725_));
 BUF_X4 _27967_ (.A(_02725_),
    .Z(_02726_));
 BUF_X4 _27968_ (.A(_02726_),
    .Z(_02727_));
 BUF_X4 _27969_ (.A(_02714_),
    .Z(_02728_));
 OAI21_X1 _27970_ (.A(_02727_),
    .B1(_02710_),
    .B2(_02728_),
    .ZN(_02729_));
 AND2_X1 _27971_ (.A1(_02699_),
    .A2(_02690_),
    .ZN(_02730_));
 BUF_X2 _27972_ (.A(_02730_),
    .Z(_02731_));
 BUF_X4 _27973_ (.A(_02704_),
    .Z(_02732_));
 OAI21_X1 _27974_ (.A(_02727_),
    .B1(_02731_),
    .B2(_02732_),
    .ZN(_02733_));
 AND4_X1 _27975_ (.A1(_02706_),
    .A2(_02721_),
    .A3(_02729_),
    .A4(_02733_),
    .ZN(_02734_));
 NOR2_X4 _27976_ (.A1(_02686_),
    .A2(_16853_),
    .ZN(_02735_));
 AND2_X2 _27977_ (.A1(_02708_),
    .A2(_02735_),
    .ZN(_02736_));
 INV_X1 _27978_ (.A(_02736_),
    .ZN(_02737_));
 INV_X4 _27979_ (.A(_02710_),
    .ZN(_02738_));
 NAND2_X1 _27980_ (.A1(_02737_),
    .A2(_02738_),
    .ZN(_02739_));
 INV_X32 _27981_ (.A(_16856_),
    .ZN(_02740_));
 NOR2_X2 _27982_ (.A1(_02740_),
    .A2(_16857_),
    .ZN(_02741_));
 NOR2_X4 _27983_ (.A1(_16859_),
    .A2(_16858_),
    .ZN(_02742_));
 BUF_X4 _27984_ (.A(_02742_),
    .Z(_02743_));
 AND2_X2 _27985_ (.A1(_02741_),
    .A2(_02743_),
    .ZN(_02744_));
 AND2_X1 _27986_ (.A1(_02739_),
    .A2(_02744_),
    .ZN(_02745_));
 AND2_X1 _27987_ (.A1(_02713_),
    .A2(_02685_),
    .ZN(_02746_));
 BUF_X4 _27988_ (.A(_02746_),
    .Z(_02747_));
 AND2_X1 _27989_ (.A1(_02744_),
    .A2(_02747_),
    .ZN(_02748_));
 AND2_X2 _27990_ (.A1(_02687_),
    .A2(_02713_),
    .ZN(_02749_));
 AND2_X1 _27991_ (.A1(_02749_),
    .A2(_02744_),
    .ZN(_02750_));
 OR3_X4 _27992_ (.A1(_02745_),
    .A2(_02748_),
    .A3(_02750_),
    .ZN(_02751_));
 BUF_X4 _27993_ (.A(_02744_),
    .Z(_02752_));
 BUF_X4 _27994_ (.A(_02690_),
    .Z(_02753_));
 AND2_X1 _27995_ (.A1(_02752_),
    .A2(_02753_),
    .ZN(_02754_));
 BUF_X8 _27996_ (.A(_02700_),
    .Z(_02755_));
 AND2_X4 _27997_ (.A1(_02755_),
    .A2(_02685_),
    .ZN(_02756_));
 NOR2_X4 _27998_ (.A1(_16857_),
    .A2(_16856_),
    .ZN(_02757_));
 AND2_X1 _27999_ (.A1(_02757_),
    .A2(_02743_),
    .ZN(_02758_));
 BUF_X4 _28000_ (.A(_02758_),
    .Z(_02759_));
 NAND2_X1 _28001_ (.A1(_02756_),
    .A2(_02759_),
    .ZN(_02760_));
 AND2_X2 _28002_ (.A1(_02687_),
    .A2(_02755_),
    .ZN(_02761_));
 AND2_X1 _28003_ (.A1(_02761_),
    .A2(_02759_),
    .ZN(_02762_));
 INV_X2 _28004_ (.A(_02762_),
    .ZN(_02763_));
 INV_X1 _28005_ (.A(_02739_),
    .ZN(_02764_));
 INV_X1 _28006_ (.A(_02759_),
    .ZN(_02765_));
 OAI211_X2 _28007_ (.A(_02760_),
    .B(_02763_),
    .C1(_02764_),
    .C2(_02765_),
    .ZN(_02766_));
 AND2_X2 _28008_ (.A1(_02755_),
    .A2(_02709_),
    .ZN(_02767_));
 NAND2_X2 _28009_ (.A1(_02744_),
    .A2(_02767_),
    .ZN(_02768_));
 INV_X4 _28010_ (.A(_02744_),
    .ZN(_02769_));
 INV_X1 _28011_ (.A(_02756_),
    .ZN(_02770_));
 OAI21_X1 _28012_ (.A(_02768_),
    .B1(_02769_),
    .B2(_02770_),
    .ZN(_02771_));
 NOR4_X2 _28013_ (.A1(_02751_),
    .A2(_02754_),
    .A3(_02766_),
    .A4(_02771_),
    .ZN(_02772_));
 BUF_X4 _28014_ (.A(_02681_),
    .Z(_02773_));
 AND2_X4 _28015_ (.A1(_02773_),
    .A2(_02741_),
    .ZN(_02774_));
 AND2_X2 _28016_ (.A1(_02712_),
    .A2(_02708_),
    .ZN(_02775_));
 NAND2_X1 _28017_ (.A1(_02774_),
    .A2(_02775_),
    .ZN(_02776_));
 INV_X1 _28018_ (.A(_02774_),
    .ZN(_02777_));
 AND2_X2 _28019_ (.A1(_02687_),
    .A2(_02708_),
    .ZN(_02778_));
 INV_X2 _28020_ (.A(_02778_),
    .ZN(_02779_));
 OAI21_X1 _28021_ (.A(_02776_),
    .B1(_02777_),
    .B2(_02779_),
    .ZN(_02780_));
 AND2_X2 _28022_ (.A1(_02714_),
    .A2(_02686_),
    .ZN(_02781_));
 AOI21_X1 _28023_ (.A(_02780_),
    .B1(_02781_),
    .B2(_02774_),
    .ZN(_02782_));
 NOR2_X1 _28024_ (.A1(_02691_),
    .A2(_02730_),
    .ZN(_02783_));
 INV_X1 _28025_ (.A(_02783_),
    .ZN(_02784_));
 OAI21_X1 _28026_ (.A(_02774_),
    .B1(_02784_),
    .B2(_02767_),
    .ZN(_02785_));
 AND2_X2 _28027_ (.A1(_02681_),
    .A2(_02757_),
    .ZN(_02786_));
 BUF_X4 _28028_ (.A(_02786_),
    .Z(_02787_));
 OAI21_X1 _28029_ (.A(_02787_),
    .B1(_02710_),
    .B2(_02715_),
    .ZN(_02788_));
 AND2_X1 _28030_ (.A1(_02690_),
    .A2(_16853_),
    .ZN(_02789_));
 BUF_X2 _28031_ (.A(_02789_),
    .Z(_02790_));
 AND2_X2 _28032_ (.A1(_02755_),
    .A2(_02686_),
    .ZN(_02791_));
 OAI21_X1 _28033_ (.A(_02787_),
    .B1(_02790_),
    .B2(_02791_),
    .ZN(_02792_));
 AND4_X1 _28034_ (.A1(_02782_),
    .A2(_02785_),
    .A3(_02788_),
    .A4(_02792_),
    .ZN(_02793_));
 AND2_X4 _28035_ (.A1(_02683_),
    .A2(_02742_),
    .ZN(_02794_));
 BUF_X8 _28036_ (.A(_02794_),
    .Z(_02795_));
 BUF_X4 _28037_ (.A(_02795_),
    .Z(_02796_));
 AND2_X1 _28038_ (.A1(_02755_),
    .A2(_02698_),
    .ZN(_02797_));
 OAI21_X1 _28039_ (.A(_02796_),
    .B1(_02790_),
    .B2(_02797_),
    .ZN(_02798_));
 AND2_X2 _28040_ (.A1(_02723_),
    .A2(_02743_),
    .ZN(_02799_));
 BUF_X4 _28041_ (.A(_16853_),
    .Z(_02800_));
 AND2_X2 _28042_ (.A1(_02708_),
    .A2(_02800_),
    .ZN(_02801_));
 NAND2_X1 _28043_ (.A1(_02799_),
    .A2(_02801_),
    .ZN(_02802_));
 NAND2_X1 _28044_ (.A1(_02749_),
    .A2(_02799_),
    .ZN(_02803_));
 NAND3_X1 _28045_ (.A1(_02747_),
    .A2(_02724_),
    .A3(_02743_),
    .ZN(_02804_));
 AND3_X1 _28046_ (.A1(_02802_),
    .A2(_02803_),
    .A3(_02804_),
    .ZN(_02805_));
 BUF_X2 _28047_ (.A(_02799_),
    .Z(_02806_));
 INV_X1 _28048_ (.A(_02735_),
    .ZN(_02807_));
 NAND2_X1 _28049_ (.A1(_02807_),
    .A2(_02753_),
    .ZN(_02808_));
 INV_X1 _28050_ (.A(_02808_),
    .ZN(_02809_));
 OAI21_X1 _28051_ (.A(_02806_),
    .B1(_02809_),
    .B2(_02702_),
    .ZN(_02810_));
 BUF_X4 _28052_ (.A(_02686_),
    .Z(_02811_));
 BUF_X4 _28053_ (.A(_02708_),
    .Z(_02812_));
 OAI211_X2 _28054_ (.A(_02795_),
    .B(_02811_),
    .C1(_02728_),
    .C2(_02812_),
    .ZN(_02813_));
 AND4_X1 _28055_ (.A1(_02798_),
    .A2(_02805_),
    .A3(_02810_),
    .A4(_02813_),
    .ZN(_02814_));
 AND4_X1 _28056_ (.A1(_02734_),
    .A2(_02772_),
    .A3(_02793_),
    .A4(_02814_),
    .ZN(_02815_));
 AND2_X4 _28057_ (.A1(_16859_),
    .A2(_16858_),
    .ZN(_02816_));
 BUF_X8 _28058_ (.A(_02816_),
    .Z(_02817_));
 AND2_X4 _28059_ (.A1(_02817_),
    .A2(_02682_),
    .ZN(_02818_));
 AND2_X1 _28060_ (.A1(_02731_),
    .A2(_02818_),
    .ZN(_02819_));
 INV_X1 _28061_ (.A(_02819_),
    .ZN(_02820_));
 AND2_X1 _28062_ (.A1(_02719_),
    .A2(_02818_),
    .ZN(_02821_));
 INV_X1 _28063_ (.A(_02821_),
    .ZN(_02822_));
 BUF_X8 _28064_ (.A(_02818_),
    .Z(_02823_));
 NAND2_X1 _28065_ (.A1(_02823_),
    .A2(_02797_),
    .ZN(_02824_));
 INV_X1 _28066_ (.A(_02709_),
    .ZN(_02825_));
 NAND3_X1 _28067_ (.A1(_02823_),
    .A2(_02825_),
    .A3(_02728_),
    .ZN(_02826_));
 NAND4_X1 _28068_ (.A1(_02820_),
    .A2(_02822_),
    .A3(_02824_),
    .A4(_02826_),
    .ZN(_02827_));
 AND2_X1 _28069_ (.A1(_02723_),
    .A2(_02816_),
    .ZN(_02828_));
 BUF_X4 _28070_ (.A(_02828_),
    .Z(_02829_));
 AND2_X4 _28071_ (.A1(_02700_),
    .A2(_02735_),
    .ZN(_02830_));
 BUF_X8 _28072_ (.A(_02830_),
    .Z(_02831_));
 AND2_X4 _28073_ (.A1(_02829_),
    .A2(_02831_),
    .ZN(_02832_));
 AND3_X1 _28074_ (.A1(_02767_),
    .A2(_02724_),
    .A3(_02817_),
    .ZN(_02833_));
 OR2_X1 _28075_ (.A1(_02832_),
    .A2(_02833_),
    .ZN(_02834_));
 BUF_X4 _28076_ (.A(_02829_),
    .Z(_02835_));
 OAI211_X2 _28077_ (.A(_02835_),
    .B(_02812_),
    .C1(_02811_),
    .C2(_02800_),
    .ZN(_02836_));
 NAND2_X1 _28078_ (.A1(_02829_),
    .A2(_02747_),
    .ZN(_02837_));
 INV_X1 _28079_ (.A(_02829_),
    .ZN(_02838_));
 INV_X1 _28080_ (.A(_02749_),
    .ZN(_02839_));
 OAI211_X2 _28081_ (.A(_02836_),
    .B(_02837_),
    .C1(_02838_),
    .C2(_02839_),
    .ZN(_02840_));
 INV_X4 _28082_ (.A(_02712_),
    .ZN(_02841_));
 NAND2_X1 _28083_ (.A1(_02841_),
    .A2(_02753_),
    .ZN(_02842_));
 NOR2_X1 _28084_ (.A1(_02838_),
    .A2(_02842_),
    .ZN(_02843_));
 NOR4_X1 _28085_ (.A1(_02827_),
    .A2(_02834_),
    .A3(_02840_),
    .A4(_02843_),
    .ZN(_02844_));
 NOR2_X4 _28086_ (.A1(_02680_),
    .A2(_16858_),
    .ZN(_02845_));
 AND2_X2 _28087_ (.A1(_02724_),
    .A2(_02845_),
    .ZN(_02846_));
 BUF_X2 _28088_ (.A(_02846_),
    .Z(_02847_));
 AND2_X2 _28089_ (.A1(_02735_),
    .A2(_02714_),
    .ZN(_02848_));
 NAND2_X1 _28090_ (.A1(_02847_),
    .A2(_02848_),
    .ZN(_02849_));
 AND2_X2 _28091_ (.A1(_02845_),
    .A2(_02682_),
    .ZN(_02850_));
 BUF_X4 _28092_ (.A(_02850_),
    .Z(_02851_));
 AND2_X1 _28093_ (.A1(_02851_),
    .A2(_02761_),
    .ZN(_02852_));
 INV_X1 _28094_ (.A(_02852_),
    .ZN(_02853_));
 NAND2_X1 _28095_ (.A1(_02790_),
    .A2(_02851_),
    .ZN(_02854_));
 AND2_X1 _28096_ (.A1(_02853_),
    .A2(_02854_),
    .ZN(_02855_));
 BUF_X4 _28097_ (.A(_02698_),
    .Z(_02856_));
 BUF_X4 _28098_ (.A(_02685_),
    .Z(_02857_));
 BUF_X4 _28099_ (.A(_02755_),
    .Z(_02858_));
 BUF_X4 _28100_ (.A(_02690_),
    .Z(_02859_));
 OAI221_X1 _28101_ (.A(_02847_),
    .B1(_02856_),
    .B2(_02857_),
    .C1(_02858_),
    .C2(_02859_),
    .ZN(_02860_));
 BUF_X4 _28102_ (.A(_02851_),
    .Z(_02861_));
 BUF_X4 _28103_ (.A(_02687_),
    .Z(_02862_));
 INV_X1 _28104_ (.A(_02862_),
    .ZN(_02863_));
 AND2_X4 _28105_ (.A1(_02863_),
    .A2(_02812_),
    .ZN(_02864_));
 OAI21_X1 _28106_ (.A(_02861_),
    .B1(_02864_),
    .B2(_02747_),
    .ZN(_02865_));
 AND4_X1 _28107_ (.A1(_02849_),
    .A2(_02855_),
    .A3(_02860_),
    .A4(_02865_),
    .ZN(_02866_));
 AND2_X2 _28108_ (.A1(_02741_),
    .A2(_02817_),
    .ZN(_02867_));
 BUF_X4 _28109_ (.A(_02867_),
    .Z(_02868_));
 AND2_X4 _28110_ (.A1(_02689_),
    .A2(_02709_),
    .ZN(_02869_));
 BUF_X4 _28111_ (.A(_02869_),
    .Z(_02870_));
 AND2_X1 _28112_ (.A1(_02868_),
    .A2(_02870_),
    .ZN(_02871_));
 INV_X1 _28113_ (.A(_02871_),
    .ZN(_02872_));
 NAND2_X1 _28114_ (.A1(_02749_),
    .A2(_02868_),
    .ZN(_02873_));
 NAND2_X1 _28115_ (.A1(_02778_),
    .A2(_02868_),
    .ZN(_02874_));
 OAI211_X2 _28116_ (.A(_02868_),
    .B(_02858_),
    .C1(_02811_),
    .C2(_02857_),
    .ZN(_02875_));
 NAND4_X1 _28117_ (.A1(_02872_),
    .A2(_02873_),
    .A3(_02874_),
    .A4(_02875_),
    .ZN(_02876_));
 AND2_X4 _28118_ (.A1(_02817_),
    .A2(_02757_),
    .ZN(_02877_));
 AND2_X1 _28119_ (.A1(_02702_),
    .A2(_02877_),
    .ZN(_02878_));
 AND2_X1 _28120_ (.A1(_02704_),
    .A2(_02877_),
    .ZN(_02879_));
 OR2_X1 _28121_ (.A1(_02878_),
    .A2(_02879_),
    .ZN(_02880_));
 BUF_X2 _28122_ (.A(_02694_),
    .Z(_02881_));
 AND2_X1 _28123_ (.A1(_02881_),
    .A2(_02877_),
    .ZN(_02882_));
 BUF_X4 _28124_ (.A(_02877_),
    .Z(_02883_));
 NAND2_X1 _28125_ (.A1(_02883_),
    .A2(_02848_),
    .ZN(_02884_));
 NAND4_X1 _28126_ (.A1(_02712_),
    .A2(_02812_),
    .A3(_02817_),
    .A4(_02757_),
    .ZN(_02885_));
 INV_X1 _28127_ (.A(_02801_),
    .ZN(_02886_));
 INV_X1 _28128_ (.A(_02877_),
    .ZN(_02887_));
 OAI211_X2 _28129_ (.A(_02884_),
    .B(_02885_),
    .C1(_02886_),
    .C2(_02887_),
    .ZN(_02888_));
 NOR4_X1 _28130_ (.A1(_02876_),
    .A2(_02880_),
    .A3(_02882_),
    .A4(_02888_),
    .ZN(_02889_));
 AND2_X2 _28131_ (.A1(_02845_),
    .A2(_02741_),
    .ZN(_02890_));
 BUF_X4 _28132_ (.A(_02890_),
    .Z(_02891_));
 OAI21_X1 _28133_ (.A(_02891_),
    .B1(_02801_),
    .B2(_02781_),
    .ZN(_02892_));
 INV_X1 _28134_ (.A(_02767_),
    .ZN(_02893_));
 INV_X1 _28135_ (.A(_02831_),
    .ZN(_02894_));
 NAND2_X1 _28136_ (.A1(_02893_),
    .A2(_02894_),
    .ZN(_02895_));
 OAI21_X1 _28137_ (.A(_02891_),
    .B1(_02784_),
    .B2(_02895_),
    .ZN(_02896_));
 AND2_X2 _28138_ (.A1(_02845_),
    .A2(_02757_),
    .ZN(_02897_));
 BUF_X4 _28139_ (.A(_02897_),
    .Z(_02898_));
 NAND2_X1 _28140_ (.A1(_02898_),
    .A2(_02881_),
    .ZN(_02899_));
 INV_X1 _28141_ (.A(_02717_),
    .ZN(_02900_));
 INV_X2 _28142_ (.A(_02848_),
    .ZN(_02901_));
 NAND2_X1 _28143_ (.A1(_02900_),
    .A2(_02901_),
    .ZN(_02902_));
 BUF_X4 _28144_ (.A(_02775_),
    .Z(_02903_));
 OAI21_X1 _28145_ (.A(_02897_),
    .B1(_02902_),
    .B2(_02903_),
    .ZN(_02904_));
 AND4_X1 _28146_ (.A1(_02892_),
    .A2(_02896_),
    .A3(_02899_),
    .A4(_02904_),
    .ZN(_02905_));
 AND4_X1 _28147_ (.A1(_02844_),
    .A2(_02866_),
    .A3(_02889_),
    .A4(_02905_),
    .ZN(_02906_));
 NAND2_X4 _28148_ (.A1(_02815_),
    .A2(_02906_),
    .ZN(_02907_));
 XNOR2_X1 _28149_ (.A(_02679_),
    .B(_02907_),
    .ZN(_02908_));
 INV_X1 _28150_ (.A(_17208_),
    .ZN(_02909_));
 XNOR2_X1 _28151_ (.A(_02908_),
    .B(_02909_),
    .ZN(_02910_));
 MUX2_X1 _28152_ (.A(_01887_),
    .B(_02910_),
    .S(_01876_),
    .Z(_00708_));
 XOR2_X1 _28153_ (.A(_17166_),
    .B(_17262_),
    .Z(_02911_));
 XOR2_X1 _28154_ (.A(_01651_),
    .B(_02911_),
    .Z(_02912_));
 XNOR2_X1 _28155_ (.A(_14484_),
    .B(_02912_),
    .ZN(_02913_));
 MUX2_X1 _28156_ (.A(_01252_),
    .B(_02913_),
    .S(_01831_),
    .Z(_01176_));
 XNOR2_X1 _28157_ (.A(_17169_),
    .B(_17265_),
    .ZN(_02914_));
 XNOR2_X1 _28158_ (.A(_01654_),
    .B(_02914_),
    .ZN(_02915_));
 BUF_X4 _28159_ (.A(_03933_),
    .Z(_02916_));
 MUX2_X1 _28160_ (.A(_01263_),
    .B(_02915_),
    .S(_02916_),
    .Z(_01179_));
 XNOR2_X1 _28161_ (.A(_17170_),
    .B(_17266_),
    .ZN(_02917_));
 XNOR2_X1 _28162_ (.A(_01657_),
    .B(_02917_),
    .ZN(_02918_));
 MUX2_X1 _28163_ (.A(_01274_),
    .B(_02918_),
    .S(_02916_),
    .Z(_01180_));
 XOR2_X1 _28164_ (.A(_17171_),
    .B(_17267_),
    .Z(_02919_));
 XOR2_X1 _28165_ (.A(_01658_),
    .B(_02919_),
    .Z(_02920_));
 XNOR2_X1 _28166_ (.A(_14687_),
    .B(_02920_),
    .ZN(_02921_));
 MUX2_X1 _28167_ (.A(_01285_),
    .B(_02921_),
    .S(_02916_),
    .Z(_01181_));
 XNOR2_X1 _28168_ (.A(_17172_),
    .B(_17268_),
    .ZN(_02922_));
 NOR2_X1 _28169_ (.A1(_03933_),
    .A2(_01296_),
    .ZN(_02923_));
 AOI21_X1 _28170_ (.A(_02923_),
    .B1(_02922_),
    .B2(_01788_),
    .ZN(_02924_));
 NAND2_X1 _28171_ (.A1(_01661_),
    .A2(_03738_),
    .ZN(_02925_));
 MUX2_X1 _28172_ (.A(_02922_),
    .B(_02924_),
    .S(_02925_),
    .Z(_01182_));
 XNOR2_X1 _28173_ (.A(_17173_),
    .B(_17269_),
    .ZN(_02926_));
 XNOR2_X1 _28174_ (.A(_01663_),
    .B(_02926_),
    .ZN(_02927_));
 MUX2_X1 _28175_ (.A(_01307_),
    .B(_02927_),
    .S(_02916_),
    .Z(_01183_));
 XNOR2_X1 _28176_ (.A(_10997_),
    .B(_17270_),
    .ZN(_02928_));
 XNOR2_X1 _28177_ (.A(_01665_),
    .B(_02928_),
    .ZN(_02929_));
 MUX2_X1 _28178_ (.A(_01318_),
    .B(_02929_),
    .S(_02916_),
    .Z(_01184_));
 XOR2_X1 _28179_ (.A(_11004_),
    .B(_17271_),
    .Z(_02930_));
 XNOR2_X1 _28180_ (.A(_01668_),
    .B(_02930_),
    .ZN(_02931_));
 MUX2_X1 _28181_ (.A(_01329_),
    .B(_02931_),
    .S(_02916_),
    .Z(_01185_));
 XOR2_X1 _28182_ (.A(_17145_),
    .B(_17241_),
    .Z(_02932_));
 XOR2_X1 _28183_ (.A(_01669_),
    .B(_02932_),
    .Z(_02933_));
 XNOR2_X1 _28184_ (.A(_15216_),
    .B(_02933_),
    .ZN(_02934_));
 MUX2_X1 _28185_ (.A(_01213_),
    .B(_02934_),
    .S(_02916_),
    .Z(_01155_));
 XOR2_X1 _28186_ (.A(_17146_),
    .B(_17242_),
    .Z(_02935_));
 XOR2_X1 _28187_ (.A(_01672_),
    .B(_02935_),
    .Z(_02936_));
 XNOR2_X1 _28188_ (.A(_15296_),
    .B(_02936_),
    .ZN(_02937_));
 MUX2_X1 _28189_ (.A(_01224_),
    .B(_02937_),
    .S(_02916_),
    .Z(_01156_));
 XOR2_X1 _28190_ (.A(_17219_),
    .B(_17101_),
    .Z(_02938_));
 AND2_X1 _28191_ (.A1(_02380_),
    .A2(_02463_),
    .ZN(_02939_));
 AND2_X1 _28192_ (.A1(_02379_),
    .A2(_02394_),
    .ZN(_02940_));
 AND2_X2 _28193_ (.A1(_02379_),
    .A2(_02433_),
    .ZN(_02941_));
 AND4_X1 _28194_ (.A1(_02375_),
    .A2(_02398_),
    .A3(_02378_),
    .A4(_02383_),
    .ZN(_02942_));
 NOR4_X1 _28195_ (.A1(_02939_),
    .A2(_02940_),
    .A3(_02941_),
    .A4(_02942_),
    .ZN(_02943_));
 BUF_X2 _28196_ (.A(_02411_),
    .Z(_02944_));
 NAND4_X1 _28197_ (.A1(_02598_),
    .A2(_02553_),
    .A3(_02383_),
    .A4(_02944_),
    .ZN(_02945_));
 OAI21_X1 _28198_ (.A(_02610_),
    .B1(_02372_),
    .B2(_02423_),
    .ZN(_02946_));
 NAND4_X1 _28199_ (.A1(_02943_),
    .A2(_02600_),
    .A3(_02945_),
    .A4(_02946_),
    .ZN(_02947_));
 AND2_X1 _28200_ (.A1(_02555_),
    .A2(_02618_),
    .ZN(_02948_));
 AND2_X1 _28201_ (.A1(_02537_),
    .A2(_02555_),
    .ZN(_02949_));
 AOI211_X2 _28202_ (.A(_02948_),
    .B(_02949_),
    .C1(_02549_),
    .C2(_02555_),
    .ZN(_02950_));
 AND2_X1 _28203_ (.A1(_02591_),
    .A2(_02555_),
    .ZN(_02951_));
 INV_X1 _28204_ (.A(_02951_),
    .ZN(_02952_));
 INV_X2 _28205_ (.A(_02635_),
    .ZN(_02953_));
 OAI21_X1 _28206_ (.A(_02557_),
    .B1(_02953_),
    .B2(_02586_),
    .ZN(_02954_));
 OAI21_X1 _28207_ (.A(_02557_),
    .B1(_02539_),
    .B2(_02611_),
    .ZN(_02955_));
 NAND4_X1 _28208_ (.A1(_02950_),
    .A2(_02952_),
    .A3(_02954_),
    .A4(_02955_),
    .ZN(_02956_));
 AND2_X4 _28209_ (.A1(_02425_),
    .A2(_02413_),
    .ZN(_02957_));
 AOI211_X2 _28210_ (.A(_02957_),
    .B(_02644_),
    .C1(_02466_),
    .C2(_02413_),
    .ZN(_02958_));
 INV_X1 _28211_ (.A(_02407_),
    .ZN(_02959_));
 AOI21_X1 _28212_ (.A(_02959_),
    .B1(_02424_),
    .B2(_02426_),
    .ZN(_02960_));
 AOI21_X1 _28213_ (.A(_02960_),
    .B1(_02500_),
    .B2(_02407_),
    .ZN(_02961_));
 NAND3_X1 _28214_ (.A1(_02390_),
    .A2(_02375_),
    .A3(_02472_),
    .ZN(_02962_));
 INV_X4 _28215_ (.A(_02538_),
    .ZN(_02963_));
 OAI21_X1 _28216_ (.A(_02962_),
    .B1(_02959_),
    .B2(_02963_),
    .ZN(_02964_));
 AOI21_X1 _28217_ (.A(_02964_),
    .B1(_02528_),
    .B2(_02407_),
    .ZN(_02965_));
 OAI21_X1 _28218_ (.A(_02435_),
    .B1(_02421_),
    .B2(_02439_),
    .ZN(_02966_));
 NAND4_X1 _28219_ (.A1(_02958_),
    .A2(_02961_),
    .A3(_02965_),
    .A4(_02966_),
    .ZN(_02967_));
 OAI21_X1 _28220_ (.A(_02524_),
    .B1(_02572_),
    .B2(_02466_),
    .ZN(_02968_));
 NAND2_X1 _28221_ (.A1(_02463_),
    .A2(_02524_),
    .ZN(_02969_));
 NAND4_X1 _28222_ (.A1(_02398_),
    .A2(_02437_),
    .A3(_02593_),
    .A4(_02472_),
    .ZN(_02970_));
 AND3_X1 _28223_ (.A1(_02968_),
    .A2(_02969_),
    .A3(_02970_),
    .ZN(_02971_));
 NAND2_X1 _28224_ (.A1(_02539_),
    .A2(_02431_),
    .ZN(_02972_));
 OAI211_X2 _28225_ (.A(_02431_),
    .B(_02499_),
    .C1(_02664_),
    .C2(_02506_),
    .ZN(_02973_));
 NAND4_X1 _28226_ (.A1(_02971_),
    .A2(_02432_),
    .A3(_02972_),
    .A4(_02973_),
    .ZN(_02974_));
 NOR4_X2 _28227_ (.A1(_02947_),
    .A2(_02956_),
    .A3(_02967_),
    .A4(_02974_),
    .ZN(_02975_));
 AND2_X1 _28228_ (.A1(_02371_),
    .A2(_02437_),
    .ZN(_02976_));
 NAND2_X1 _28229_ (.A1(_02976_),
    .A2(_02448_),
    .ZN(_02977_));
 NAND2_X1 _28230_ (.A1(_02505_),
    .A2(_02448_),
    .ZN(_02978_));
 NAND2_X1 _28231_ (.A1(_02448_),
    .A2(_02490_),
    .ZN(_02979_));
 AND4_X1 _28232_ (.A1(_02626_),
    .A2(_02977_),
    .A3(_02978_),
    .A4(_02979_),
    .ZN(_02980_));
 AND2_X1 _28233_ (.A1(_02438_),
    .A2(_02504_),
    .ZN(_02981_));
 OAI211_X2 _28234_ (.A(_02504_),
    .B(_02394_),
    .C1(_02396_),
    .C2(_02400_),
    .ZN(_02982_));
 NAND2_X1 _28235_ (.A1(_02571_),
    .A2(_02503_),
    .ZN(_02983_));
 OAI211_X2 _28236_ (.A(_02982_),
    .B(_02983_),
    .C1(_02657_),
    .C2(_02493_),
    .ZN(_02984_));
 AOI211_X2 _28237_ (.A(_02981_),
    .B(_02984_),
    .C1(_02504_),
    .C2(_02658_),
    .ZN(_02985_));
 AOI21_X1 _28238_ (.A(_02453_),
    .B1(_02544_),
    .B2(_02631_),
    .ZN(_02986_));
 AND2_X1 _28239_ (.A1(_02437_),
    .A2(_02506_),
    .ZN(_02987_));
 AOI211_X4 _28240_ (.A(_02520_),
    .B(_02986_),
    .C1(_02451_),
    .C2(_02987_),
    .ZN(_02988_));
 OAI21_X1 _28241_ (.A(_02614_),
    .B1(_02976_),
    .B2(_02602_),
    .ZN(_02989_));
 AND4_X4 _28242_ (.A1(_02980_),
    .A2(_02985_),
    .A3(_02988_),
    .A4(_02989_),
    .ZN(_02990_));
 BUF_X4 _28243_ (.A(_02499_),
    .Z(_02991_));
 NAND3_X1 _28244_ (.A1(_02672_),
    .A2(_02991_),
    .A3(_02944_),
    .ZN(_02992_));
 NAND2_X1 _28245_ (.A1(_02532_),
    .A2(_02500_),
    .ZN(_02993_));
 OAI211_X2 _28246_ (.A(_02534_),
    .B(_02375_),
    .C1(_02481_),
    .C2(_02419_),
    .ZN(_02994_));
 NAND2_X1 _28247_ (.A1(_02531_),
    .A2(_02433_),
    .ZN(_02995_));
 NAND4_X1 _28248_ (.A1(_02399_),
    .A2(_02534_),
    .A3(_02375_),
    .A4(_02403_),
    .ZN(_02996_));
 AND4_X1 _28249_ (.A1(_02993_),
    .A2(_02994_),
    .A3(_02995_),
    .A4(_02996_),
    .ZN(_02997_));
 OAI21_X1 _28250_ (.A(_02548_),
    .B1(_02976_),
    .B2(_02528_),
    .ZN(_02998_));
 BUF_X4 _28251_ (.A(_02564_),
    .Z(_02999_));
 OAI21_X1 _28252_ (.A(_02548_),
    .B1(_02477_),
    .B2(_02999_),
    .ZN(_03000_));
 AND4_X1 _28253_ (.A1(_02992_),
    .A2(_02997_),
    .A3(_02998_),
    .A4(_03000_),
    .ZN(_03001_));
 NAND3_X1 _28254_ (.A1(_02462_),
    .A2(_02368_),
    .A3(_02371_),
    .ZN(_03002_));
 BUF_X4 _28255_ (.A(_02462_),
    .Z(_03003_));
 NAND2_X1 _28256_ (.A1(_03003_),
    .A2(_02999_),
    .ZN(_03004_));
 INV_X1 _28257_ (.A(_02466_),
    .ZN(_03005_));
 OAI211_X2 _28258_ (.A(_03002_),
    .B(_03004_),
    .C1(_02489_),
    .C2(_03005_),
    .ZN(_03006_));
 NAND2_X1 _28259_ (.A1(_02465_),
    .A2(_02549_),
    .ZN(_03007_));
 NAND3_X1 _28260_ (.A1(_02619_),
    .A2(_02534_),
    .A3(_02429_),
    .ZN(_03008_));
 INV_X1 _28261_ (.A(_02987_),
    .ZN(_03009_));
 OAI211_X2 _28262_ (.A(_03007_),
    .B(_03008_),
    .C1(_02469_),
    .C2(_03009_),
    .ZN(_03010_));
 AOI21_X1 _28263_ (.A(_02469_),
    .B1(_02544_),
    .B2(_02631_),
    .ZN(_03011_));
 OAI21_X1 _28264_ (.A(_02567_),
    .B1(_02489_),
    .B2(_02486_),
    .ZN(_03012_));
 NOR4_X1 _28265_ (.A1(_03006_),
    .A2(_03010_),
    .A3(_03011_),
    .A4(_03012_),
    .ZN(_03013_));
 NAND4_X2 _28266_ (.A1(_02975_),
    .A2(_02990_),
    .A3(_03001_),
    .A4(_03013_),
    .ZN(_03014_));
 NOR2_X4 _28267_ (.A1(_03014_),
    .A2(_02670_),
    .ZN(_03015_));
 AND3_X1 _28268_ (.A1(_02232_),
    .A2(_02324_),
    .A3(_02132_),
    .ZN(_03016_));
 AND3_X1 _28269_ (.A1(_02140_),
    .A2(_02324_),
    .A3(_02132_),
    .ZN(_03017_));
 AND2_X1 _28270_ (.A1(_02146_),
    .A2(_02174_),
    .ZN(_03018_));
 AOI211_X4 _28271_ (.A(_03016_),
    .B(_03017_),
    .C1(_02134_),
    .C2(_03018_),
    .ZN(_03019_));
 AND2_X4 _28272_ (.A1(_02184_),
    .A2(_02201_),
    .ZN(_03020_));
 INV_X1 _28273_ (.A(_03020_),
    .ZN(_03021_));
 AND2_X2 _28274_ (.A1(_02205_),
    .A2(_02181_),
    .ZN(_03022_));
 NOR2_X4 _28275_ (.A1(_02172_),
    .A2(_02143_),
    .ZN(_03023_));
 AND3_X1 _28276_ (.A1(_03023_),
    .A2(_02180_),
    .A3(_02167_),
    .ZN(_03024_));
 AND2_X1 _28277_ (.A1(_02143_),
    .A2(_02136_),
    .ZN(_03025_));
 AND2_X1 _28278_ (.A1(_03025_),
    .A2(_02180_),
    .ZN(_03026_));
 AND4_X1 _28279_ (.A1(_02132_),
    .A2(_02144_),
    .A3(_02159_),
    .A4(_02179_),
    .ZN(_03027_));
 NOR4_X1 _28280_ (.A1(_03022_),
    .A2(_03024_),
    .A3(_03026_),
    .A4(_03027_),
    .ZN(_03028_));
 NAND4_X1 _28281_ (.A1(_02214_),
    .A2(_02237_),
    .A3(_02193_),
    .A4(_02267_),
    .ZN(_03029_));
 OAI21_X1 _28282_ (.A(_02201_),
    .B1(_02320_),
    .B2(_02250_),
    .ZN(_03030_));
 AND4_X1 _28283_ (.A1(_03021_),
    .A2(_03028_),
    .A3(_03029_),
    .A4(_03030_),
    .ZN(_03031_));
 BUF_X4 _28284_ (.A(_02324_),
    .Z(_03032_));
 NAND3_X1 _28285_ (.A1(_02346_),
    .A2(_03032_),
    .A3(_02193_),
    .ZN(_03033_));
 INV_X1 _28286_ (.A(_02133_),
    .ZN(_03034_));
 INV_X1 _28287_ (.A(_02257_),
    .ZN(_03035_));
 OAI21_X1 _28288_ (.A(_03033_),
    .B1(_03034_),
    .B2(_03035_),
    .ZN(_03036_));
 AND2_X2 _28289_ (.A1(_02144_),
    .A2(_02159_),
    .ZN(_03037_));
 AOI21_X1 _28290_ (.A(_03036_),
    .B1(_02134_),
    .B2(_03037_),
    .ZN(_03038_));
 INV_X4 _28291_ (.A(_02359_),
    .ZN(_03039_));
 INV_X1 _28292_ (.A(_02297_),
    .ZN(_03040_));
 AOI21_X1 _28293_ (.A(_02166_),
    .B1(_03039_),
    .B2(_03040_),
    .ZN(_03041_));
 NAND2_X1 _28294_ (.A1(_02346_),
    .A2(_02176_),
    .ZN(_03042_));
 NAND2_X1 _28295_ (.A1(_02165_),
    .A2(_02250_),
    .ZN(_03043_));
 NAND2_X1 _28296_ (.A1(_03042_),
    .A2(_03043_),
    .ZN(_03044_));
 AND2_X1 _28297_ (.A1(_02218_),
    .A2(_02176_),
    .ZN(_03045_));
 AND4_X1 _28298_ (.A1(_02174_),
    .A2(_02237_),
    .A3(_02132_),
    .A4(_02164_),
    .ZN(_03046_));
 NOR4_X1 _28299_ (.A1(_03041_),
    .A2(_03044_),
    .A3(_03045_),
    .A4(_03046_),
    .ZN(_03047_));
 AND4_X2 _28300_ (.A1(_03019_),
    .A2(_03031_),
    .A3(_03038_),
    .A4(_03047_),
    .ZN(_03048_));
 OAI21_X1 _28301_ (.A(_02225_),
    .B1(_02156_),
    .B2(_02208_),
    .ZN(_03049_));
 AND2_X1 _28302_ (.A1(_02136_),
    .A2(_02350_),
    .ZN(_03050_));
 OAI21_X1 _28303_ (.A(_02225_),
    .B1(_03050_),
    .B2(_02285_),
    .ZN(_03051_));
 AND2_X1 _28304_ (.A1(_03049_),
    .A2(_03051_),
    .ZN(_03052_));
 AND2_X1 _28305_ (.A1(_02318_),
    .A2(_02258_),
    .ZN(_03053_));
 INV_X1 _28306_ (.A(_03053_),
    .ZN(_03054_));
 BUF_X4 _28307_ (.A(_02142_),
    .Z(_03055_));
 OAI211_X2 _28308_ (.A(_02262_),
    .B(_02219_),
    .C1(_03055_),
    .C2(_02174_),
    .ZN(_03056_));
 OAI211_X2 _28309_ (.A(_02258_),
    .B(_02191_),
    .C1(_03055_),
    .C2(_02350_),
    .ZN(_03057_));
 AND4_X1 _28310_ (.A1(_02265_),
    .A2(_03054_),
    .A3(_03056_),
    .A4(_03057_),
    .ZN(_03058_));
 AND2_X1 _28311_ (.A1(_02170_),
    .A2(_02136_),
    .ZN(_03059_));
 OAI21_X1 _28312_ (.A(_02247_),
    .B1(_03059_),
    .B2(_02344_),
    .ZN(_03060_));
 AND2_X1 _28313_ (.A1(_03059_),
    .A2(_02233_),
    .ZN(_03061_));
 AND2_X1 _28314_ (.A1(_02260_),
    .A2(_02233_),
    .ZN(_03062_));
 AND2_X1 _28315_ (.A1(_02173_),
    .A2(_16807_),
    .ZN(_03063_));
 AND2_X1 _28316_ (.A1(_02233_),
    .A2(_03063_),
    .ZN(_03064_));
 NOR4_X1 _28317_ (.A1(_03061_),
    .A2(_02231_),
    .A3(_03062_),
    .A4(_03064_),
    .ZN(_03065_));
 AND4_X1 _28318_ (.A1(_03052_),
    .A2(_03058_),
    .A3(_03060_),
    .A4(_03065_),
    .ZN(_03066_));
 AND2_X1 _28319_ (.A1(_03059_),
    .A2(_02275_),
    .ZN(_03067_));
 OAI21_X1 _28320_ (.A(_02275_),
    .B1(_02205_),
    .B2(_02207_),
    .ZN(_03068_));
 NAND3_X1 _28321_ (.A1(_02156_),
    .A2(_02164_),
    .A3(_02273_),
    .ZN(_03069_));
 OAI211_X2 _28322_ (.A(_03068_),
    .B(_03069_),
    .C1(_02154_),
    .C2(_02284_),
    .ZN(_03070_));
 AOI211_X2 _28323_ (.A(_03067_),
    .B(_03070_),
    .C1(_02275_),
    .C2(_03018_),
    .ZN(_03071_));
 AND2_X1 _28324_ (.A1(_02313_),
    .A2(_02314_),
    .ZN(_03072_));
 NAND2_X2 _28325_ (.A1(_02312_),
    .A2(_02297_),
    .ZN(_03073_));
 NAND3_X1 _28326_ (.A1(_02304_),
    .A2(_02273_),
    .A3(_02267_),
    .ZN(_03074_));
 INV_X2 _28327_ (.A(_02313_),
    .ZN(_03075_));
 OAI211_X2 _28328_ (.A(_03073_),
    .B(_03074_),
    .C1(_03075_),
    .C2(_02338_),
    .ZN(_03076_));
 AND2_X1 _28329_ (.A1(_02236_),
    .A2(_02159_),
    .ZN(_03077_));
 AND2_X4 _28330_ (.A1(_03077_),
    .A2(_02170_),
    .ZN(_03078_));
 AOI211_X2 _28331_ (.A(_03072_),
    .B(_03076_),
    .C1(_02313_),
    .C2(_03078_),
    .ZN(_03079_));
 NAND2_X1 _28332_ (.A1(_02290_),
    .A2(_03037_),
    .ZN(_03080_));
 AND2_X4 _28333_ (.A1(_02136_),
    .A2(_02169_),
    .ZN(_03081_));
 OAI211_X2 _28334_ (.A(_03032_),
    .B(_02278_),
    .C1(_03081_),
    .C2(_02359_),
    .ZN(_03082_));
 BUF_X4 _28335_ (.A(_03023_),
    .Z(_03083_));
 NAND4_X1 _28336_ (.A1(_03083_),
    .A2(_03032_),
    .A3(_02167_),
    .A4(_02278_),
    .ZN(_03084_));
 NAND2_X1 _28337_ (.A1(_02290_),
    .A2(_02205_),
    .ZN(_03085_));
 AND4_X1 _28338_ (.A1(_03080_),
    .A2(_03082_),
    .A3(_03084_),
    .A4(_03085_),
    .ZN(_03086_));
 AND2_X1 _28339_ (.A1(_02301_),
    .A2(_02264_),
    .ZN(_03087_));
 INV_X1 _28340_ (.A(_02301_),
    .ZN(_03088_));
 INV_X4 _28341_ (.A(_02208_),
    .ZN(_03089_));
 OAI21_X1 _28342_ (.A(_02308_),
    .B1(_03088_),
    .B2(_03089_),
    .ZN(_03090_));
 AOI211_X2 _28343_ (.A(_03087_),
    .B(_03090_),
    .C1(_02301_),
    .C2(_03050_),
    .ZN(_03091_));
 AND4_X4 _28344_ (.A1(_03071_),
    .A2(_03079_),
    .A3(_03086_),
    .A4(_03091_),
    .ZN(_03092_));
 NAND2_X1 _28345_ (.A1(_02153_),
    .A2(_02342_),
    .ZN(_03093_));
 INV_X1 _28346_ (.A(_02342_),
    .ZN(_03094_));
 OAI21_X1 _28347_ (.A(_03093_),
    .B1(_02157_),
    .B2(_03094_),
    .ZN(_03095_));
 BUF_X2 _28348_ (.A(_03025_),
    .Z(_03096_));
 BUF_X4 _28349_ (.A(_02342_),
    .Z(_03097_));
 NAND2_X1 _28350_ (.A1(_03096_),
    .A2(_03097_),
    .ZN(_03098_));
 NAND4_X1 _28351_ (.A1(_02326_),
    .A2(_02350_),
    .A3(_02267_),
    .A4(_02146_),
    .ZN(_03099_));
 NAND2_X1 _28352_ (.A1(_03098_),
    .A2(_03099_),
    .ZN(_03100_));
 AND4_X1 _28353_ (.A1(_02174_),
    .A2(_02219_),
    .A3(_02326_),
    .A4(_02267_),
    .ZN(_03101_));
 NOR3_X1 _28354_ (.A1(_03095_),
    .A2(_03100_),
    .A3(_03101_),
    .ZN(_03102_));
 NAND2_X1 _28355_ (.A1(_02341_),
    .A2(_02352_),
    .ZN(_03103_));
 NAND4_X1 _28356_ (.A1(_02144_),
    .A2(_02326_),
    .A3(_02146_),
    .A4(_02164_),
    .ZN(_03104_));
 AND2_X1 _28357_ (.A1(_03103_),
    .A2(_03104_),
    .ZN(_03105_));
 OAI21_X1 _28358_ (.A(_02352_),
    .B1(_03078_),
    .B2(_02257_),
    .ZN(_03106_));
 OAI21_X1 _28359_ (.A(_02327_),
    .B1(_02147_),
    .B2(_02184_),
    .ZN(_03107_));
 OAI21_X1 _28360_ (.A(_02327_),
    .B1(_02205_),
    .B2(_02191_),
    .ZN(_03108_));
 AND4_X1 _28361_ (.A1(_03105_),
    .A2(_03106_),
    .A3(_03107_),
    .A4(_03108_),
    .ZN(_03109_));
 NAND2_X1 _28362_ (.A1(_02309_),
    .A2(_02334_),
    .ZN(_03110_));
 AND2_X1 _28363_ (.A1(_02331_),
    .A2(_02229_),
    .ZN(_03111_));
 AND2_X1 _28364_ (.A1(_02331_),
    .A2(_02305_),
    .ZN(_03112_));
 AOI211_X4 _28365_ (.A(_03111_),
    .B(_03112_),
    .C1(_02141_),
    .C2(_02331_),
    .ZN(_03113_));
 AND4_X4 _28366_ (.A1(_03102_),
    .A2(_03109_),
    .A3(_03110_),
    .A4(_03113_),
    .ZN(_03114_));
 NAND4_X4 _28367_ (.A1(_03048_),
    .A2(_03066_),
    .A3(_03092_),
    .A4(_03114_),
    .ZN(_03115_));
 NOR2_X2 _28368_ (.A1(_03115_),
    .A2(_02360_),
    .ZN(_03116_));
 XNOR2_X2 _28369_ (.A(_03015_),
    .B(_03116_),
    .ZN(_03117_));
 XOR2_X1 _28370_ (.A(_02678_),
    .B(_03117_),
    .Z(_03118_));
 MUX2_X1 _28371_ (.A(_02099_),
    .B(_01908_),
    .S(_01934_),
    .Z(_03119_));
 NAND2_X1 _28372_ (.A1(_03119_),
    .A2(_01898_),
    .ZN(_03120_));
 AND2_X1 _28373_ (.A1(_01998_),
    .A2(_01965_),
    .ZN(_03121_));
 AND2_X1 _28374_ (.A1(_01965_),
    .A2(_01940_),
    .ZN(_03122_));
 NOR2_X1 _28375_ (.A1(_03121_),
    .A2(_03122_),
    .ZN(_03123_));
 AND2_X4 _28376_ (.A1(_01941_),
    .A2(_01984_),
    .ZN(_03124_));
 AND2_X1 _28377_ (.A1(_01945_),
    .A2(_01983_),
    .ZN(_03125_));
 AOI211_X2 _28378_ (.A(_03124_),
    .B(_03125_),
    .C1(_01905_),
    .C2(_01984_),
    .ZN(_03126_));
 AND2_X1 _28379_ (.A1(_01965_),
    .A2(_02052_),
    .ZN(_03127_));
 AND2_X1 _28380_ (.A1(_01993_),
    .A2(_01965_),
    .ZN(_03128_));
 AOI211_X2 _28381_ (.A(_03127_),
    .B(_03128_),
    .C1(_02106_),
    .C2(_01966_),
    .ZN(_03129_));
 BUF_X4 _28382_ (.A(_01984_),
    .Z(_03130_));
 OAI21_X1 _28383_ (.A(_03130_),
    .B1(_02064_),
    .B2(_01911_),
    .ZN(_03131_));
 AND4_X4 _28384_ (.A1(_03123_),
    .A2(_03126_),
    .A3(_03129_),
    .A4(_03131_),
    .ZN(_03132_));
 NOR3_X1 _28385_ (.A1(_01913_),
    .A2(_16846_),
    .A3(_01901_),
    .ZN(_03133_));
 AND2_X2 _28386_ (.A1(_03133_),
    .A2(_01921_),
    .ZN(_03134_));
 OAI21_X1 _28387_ (.A(_01898_),
    .B1(_03134_),
    .B2(_01967_),
    .ZN(_03135_));
 AND2_X1 _28388_ (.A1(_02074_),
    .A2(_02025_),
    .ZN(_03136_));
 AND2_X1 _28389_ (.A1(_02078_),
    .A2(_02034_),
    .ZN(_03137_));
 AND2_X1 _28390_ (.A1(_02074_),
    .A2(_01998_),
    .ZN(_03138_));
 AND3_X1 _28391_ (.A1(_01995_),
    .A2(_02006_),
    .A3(_01973_),
    .ZN(_03139_));
 NOR4_X1 _28392_ (.A1(_03136_),
    .A2(_03137_),
    .A3(_03138_),
    .A4(_03139_),
    .ZN(_03140_));
 AND4_X4 _28393_ (.A1(_03120_),
    .A2(_03132_),
    .A3(_03135_),
    .A4(_03140_),
    .ZN(_03141_));
 AND2_X1 _28394_ (.A1(_01957_),
    .A2(_01999_),
    .ZN(_03142_));
 INV_X1 _28395_ (.A(_01920_),
    .ZN(_03143_));
 INV_X1 _28396_ (.A(_02093_),
    .ZN(_03144_));
 INV_X1 _28397_ (.A(_02090_),
    .ZN(_03145_));
 AOI21_X1 _28398_ (.A(_03143_),
    .B1(_03144_),
    .B2(_03145_),
    .ZN(_03146_));
 AOI21_X1 _28399_ (.A(_03143_),
    .B1(_02102_),
    .B2(_02109_),
    .ZN(_03147_));
 AND2_X1 _28400_ (.A1(_01957_),
    .A2(_02001_),
    .ZN(_03148_));
 OR4_X2 _28401_ (.A1(_03142_),
    .A2(_03146_),
    .A3(_03147_),
    .A4(_03148_),
    .ZN(_03149_));
 AND2_X4 _28402_ (.A1(_02072_),
    .A2(_02013_),
    .ZN(_03150_));
 NOR2_X2 _28403_ (.A1(_03150_),
    .A2(_02059_),
    .ZN(_03151_));
 NAND4_X1 _28404_ (.A1(_01916_),
    .A2(_02017_),
    .A3(_01896_),
    .A4(_01908_),
    .ZN(_03152_));
 OAI21_X1 _28405_ (.A(_02014_),
    .B1(_01999_),
    .B2(_02122_),
    .ZN(_03153_));
 BUF_X4 _28406_ (.A(_01945_),
    .Z(_03154_));
 OAI21_X1 _28407_ (.A(_02014_),
    .B1(_03154_),
    .B2(_02015_),
    .ZN(_03155_));
 NAND4_X1 _28408_ (.A1(_03151_),
    .A2(_03152_),
    .A3(_03153_),
    .A4(_03155_),
    .ZN(_03156_));
 AND2_X1 _28409_ (.A1(_01954_),
    .A2(_02023_),
    .ZN(_03157_));
 NOR2_X1 _28410_ (.A1(_02066_),
    .A2(_03157_),
    .ZN(_03158_));
 BUF_X4 _28411_ (.A(_01910_),
    .Z(_03159_));
 NAND4_X1 _28412_ (.A1(_01916_),
    .A2(_01972_),
    .A3(_02099_),
    .A4(_03159_),
    .ZN(_03160_));
 BUF_X4 _28413_ (.A(_02022_),
    .Z(_03161_));
 NAND4_X1 _28414_ (.A1(_01916_),
    .A2(_02098_),
    .A3(_01972_),
    .A4(_03161_),
    .ZN(_03162_));
 NAND4_X1 _28415_ (.A1(_03158_),
    .A2(_02088_),
    .A3(_03160_),
    .A4(_03162_),
    .ZN(_03163_));
 OAI21_X1 _28416_ (.A(_02080_),
    .B1(_02050_),
    .B2(_02082_),
    .ZN(_03164_));
 OAI21_X1 _28417_ (.A(_01937_),
    .B1(_01945_),
    .B2(_02076_),
    .ZN(_03165_));
 INV_X1 _28418_ (.A(_03134_),
    .ZN(_03166_));
 INV_X1 _28419_ (.A(_02080_),
    .ZN(_03167_));
 OAI211_X2 _28420_ (.A(_03164_),
    .B(_03165_),
    .C1(_03166_),
    .C2(_03167_),
    .ZN(_03168_));
 NOR4_X1 _28421_ (.A1(_03149_),
    .A2(_03156_),
    .A3(_03163_),
    .A4(_03168_),
    .ZN(_03169_));
 AND3_X1 _28422_ (.A1(_02097_),
    .A2(_01934_),
    .A3(_01986_),
    .ZN(_03170_));
 NAND3_X1 _28423_ (.A1(_02097_),
    .A2(_01891_),
    .A3(_01986_),
    .ZN(_03171_));
 INV_X1 _28424_ (.A(_01993_),
    .ZN(_03172_));
 OAI21_X1 _28425_ (.A(_03171_),
    .B1(_03172_),
    .B2(_02119_),
    .ZN(_03173_));
 AOI211_X4 _28426_ (.A(_03170_),
    .B(_03173_),
    .C1(_02106_),
    .C2(_02123_),
    .ZN(_03174_));
 OAI211_X2 _28427_ (.A(_02123_),
    .B(_16847_),
    .C1(_03161_),
    .C2(_16846_),
    .ZN(_03175_));
 AND2_X1 _28428_ (.A1(_01986_),
    .A2(_03159_),
    .ZN(_03176_));
 AND2_X1 _28429_ (.A1(_02070_),
    .A2(_03176_),
    .ZN(_03177_));
 AND2_X1 _28430_ (.A1(_02068_),
    .A2(_02121_),
    .ZN(_03178_));
 AND2_X1 _28431_ (.A1(_02068_),
    .A2(_01941_),
    .ZN(_03179_));
 AND2_X1 _28432_ (.A1(_02068_),
    .A2(_02039_),
    .ZN(_03180_));
 NOR4_X1 _28433_ (.A1(_03177_),
    .A2(_03178_),
    .A3(_03179_),
    .A4(_03180_),
    .ZN(_03181_));
 NAND2_X1 _28434_ (.A1(_02005_),
    .A2(_01986_),
    .ZN(_03182_));
 INV_X1 _28435_ (.A(_03182_),
    .ZN(_03183_));
 OAI21_X1 _28436_ (.A(_02084_),
    .B1(_03183_),
    .B2(_02032_),
    .ZN(_03184_));
 OAI21_X1 _28437_ (.A(_02103_),
    .B1(_01923_),
    .B2(_02081_),
    .ZN(_03185_));
 OAI211_X2 _28438_ (.A(_02103_),
    .B(_02098_),
    .C1(_02118_),
    .C2(_02017_),
    .ZN(_03186_));
 OAI211_X2 _28439_ (.A(_02103_),
    .B(_02025_),
    .C1(_02118_),
    .C2(_03159_),
    .ZN(_03187_));
 AND4_X1 _28440_ (.A1(_03184_),
    .A2(_03185_),
    .A3(_03186_),
    .A4(_03187_),
    .ZN(_03188_));
 AND4_X1 _28441_ (.A1(_03174_),
    .A2(_03175_),
    .A3(_03181_),
    .A4(_03188_),
    .ZN(_03189_));
 OAI21_X1 _28442_ (.A(_02010_),
    .B1(_02033_),
    .B2(_02081_),
    .ZN(_03190_));
 AND2_X1 _28443_ (.A1(_01940_),
    .A2(_02010_),
    .ZN(_03191_));
 INV_X1 _28444_ (.A(_03191_),
    .ZN(_03192_));
 OAI211_X2 _28445_ (.A(_02010_),
    .B(_02025_),
    .C1(_03161_),
    .C2(_03159_),
    .ZN(_03193_));
 AND3_X1 _28446_ (.A1(_03190_),
    .A2(_03192_),
    .A3(_03193_),
    .ZN(_03194_));
 BUF_X4 _28447_ (.A(_02021_),
    .Z(_03195_));
 AND2_X1 _28448_ (.A1(_01940_),
    .A2(_03195_),
    .ZN(_03196_));
 AND2_X1 _28449_ (.A1(_02064_),
    .A2(_03195_),
    .ZN(_03197_));
 AND2_X1 _28450_ (.A1(_02034_),
    .A2(_02020_),
    .ZN(_03198_));
 AND2_X1 _28451_ (.A1(_03195_),
    .A2(_02077_),
    .ZN(_03199_));
 NOR4_X1 _28452_ (.A1(_03196_),
    .A2(_03197_),
    .A3(_03198_),
    .A4(_03199_),
    .ZN(_03200_));
 OAI21_X1 _28453_ (.A(_01992_),
    .B1(_02082_),
    .B2(_02071_),
    .ZN(_03201_));
 BUF_X4 _28454_ (.A(_02042_),
    .Z(_03202_));
 OAI21_X1 _28455_ (.A(_01992_),
    .B1(_03202_),
    .B2(_01967_),
    .ZN(_03203_));
 AND3_X1 _28456_ (.A1(_03201_),
    .A2(_03203_),
    .A3(_02002_),
    .ZN(_03204_));
 OAI21_X1 _28457_ (.A(_01981_),
    .B1(_01999_),
    .B2(_02001_),
    .ZN(_03205_));
 NAND2_X1 _28458_ (.A1(_02063_),
    .A2(_01980_),
    .ZN(_03206_));
 NAND3_X1 _28459_ (.A1(_01967_),
    .A2(_01972_),
    .A3(_01990_),
    .ZN(_03207_));
 NAND3_X1 _28460_ (.A1(_01981_),
    .A2(_03159_),
    .A3(_01969_),
    .ZN(_03208_));
 AND4_X1 _28461_ (.A1(_03205_),
    .A2(_03206_),
    .A3(_03207_),
    .A4(_03208_),
    .ZN(_03209_));
 AND4_X1 _28462_ (.A1(_03194_),
    .A2(_03200_),
    .A3(_03204_),
    .A4(_03209_),
    .ZN(_03210_));
 NAND4_X1 _28463_ (.A1(_03141_),
    .A2(_03169_),
    .A3(_03189_),
    .A4(_03210_),
    .ZN(_03211_));
 NOR2_X2 _28464_ (.A1(_03211_),
    .A2(_02030_),
    .ZN(_03212_));
 XNOR2_X1 _28465_ (.A(_03118_),
    .B(_03212_),
    .ZN(_03213_));
 INV_X4 _28466_ (.A(_02851_),
    .ZN(_03214_));
 OAI22_X1 _28467_ (.A1(_02894_),
    .A2(_03214_),
    .B1(_02839_),
    .B2(_02887_),
    .ZN(_03215_));
 NAND2_X1 _28468_ (.A1(_02684_),
    .A2(_02848_),
    .ZN(_03216_));
 INV_X1 _28469_ (.A(_02846_),
    .ZN(_03217_));
 OAI21_X1 _28470_ (.A(_03216_),
    .B1(_03217_),
    .B2(_02737_),
    .ZN(_03218_));
 AOI211_X2 _28471_ (.A(_03215_),
    .B(_03218_),
    .C1(_02806_),
    .C2(_02809_),
    .ZN(_03219_));
 AND2_X1 _28472_ (.A1(_02806_),
    .A2(_02831_),
    .ZN(_03220_));
 INV_X1 _28473_ (.A(_03220_),
    .ZN(_03221_));
 BUF_X2 _28474_ (.A(_02759_),
    .Z(_03222_));
 OAI21_X1 _28475_ (.A(_03222_),
    .B1(_02731_),
    .B2(_02903_),
    .ZN(_03223_));
 AND2_X1 _28476_ (.A1(_03221_),
    .A2(_03223_),
    .ZN(_03224_));
 AND2_X1 _28477_ (.A1(_02697_),
    .A2(_02781_),
    .ZN(_03225_));
 INV_X1 _28478_ (.A(_03225_),
    .ZN(_03226_));
 NAND2_X1 _28479_ (.A1(_02736_),
    .A2(_02823_),
    .ZN(_03227_));
 OAI211_X2 _28480_ (.A(_02759_),
    .B(_02800_),
    .C1(_02728_),
    .C2(_02812_),
    .ZN(_03228_));
 AND4_X1 _28481_ (.A1(_02873_),
    .A2(_03226_),
    .A3(_03227_),
    .A4(_03228_),
    .ZN(_03229_));
 AND2_X1 _28482_ (.A1(_02689_),
    .A2(_02735_),
    .ZN(_03230_));
 NAND2_X1 _28483_ (.A1(_03230_),
    .A2(_02796_),
    .ZN(_03231_));
 AOI22_X1 _28484_ (.A1(_02787_),
    .A2(_02736_),
    .B1(_02767_),
    .B2(_02795_),
    .ZN(_03232_));
 BUF_X2 _28485_ (.A(_02812_),
    .Z(_03233_));
 NAND3_X1 _28486_ (.A1(_02795_),
    .A2(_02862_),
    .A3(_03233_),
    .ZN(_03234_));
 NAND3_X1 _28487_ (.A1(_02726_),
    .A2(_02856_),
    .A3(_02704_),
    .ZN(_03235_));
 AND4_X1 _28488_ (.A1(_03231_),
    .A2(_03232_),
    .A3(_03234_),
    .A4(_03235_),
    .ZN(_03236_));
 NAND4_X1 _28489_ (.A1(_03219_),
    .A2(_03224_),
    .A3(_03229_),
    .A4(_03236_),
    .ZN(_03237_));
 AND2_X1 _28490_ (.A1(_02715_),
    .A2(_02818_),
    .ZN(_03238_));
 AND2_X1 _28491_ (.A1(_02803_),
    .A2(_02804_),
    .ZN(_03239_));
 INV_X1 _28492_ (.A(_03239_),
    .ZN(_03240_));
 AND3_X1 _28493_ (.A1(_02883_),
    .A2(_02858_),
    .A3(_02862_),
    .ZN(_03241_));
 AND3_X1 _28494_ (.A1(_02823_),
    .A2(_02704_),
    .A3(_02856_),
    .ZN(_03242_));
 OR4_X4 _28495_ (.A1(_03238_),
    .A2(_03240_),
    .A3(_03241_),
    .A4(_03242_),
    .ZN(_03243_));
 AND2_X1 _28496_ (.A1(_02756_),
    .A2(_02794_),
    .ZN(_03244_));
 AOI221_X1 _28497_ (.A(_03244_),
    .B1(_02747_),
    .B2(_02786_),
    .C1(_02801_),
    .C2(_02774_),
    .ZN(_03245_));
 XNOR2_X1 _28498_ (.A(_02686_),
    .B(_16853_),
    .ZN(_03246_));
 INV_X1 _28499_ (.A(_02755_),
    .ZN(_03247_));
 NOR2_X1 _28500_ (.A1(_03246_),
    .A2(_03247_),
    .ZN(_03248_));
 OAI21_X1 _28501_ (.A(_03222_),
    .B1(_03248_),
    .B2(_02790_),
    .ZN(_03249_));
 AND2_X1 _28502_ (.A1(_02754_),
    .A2(_03246_),
    .ZN(_03250_));
 INV_X1 _28503_ (.A(_03250_),
    .ZN(_03251_));
 NOR2_X1 _28504_ (.A1(_02778_),
    .A2(_02775_),
    .ZN(_03252_));
 INV_X1 _28505_ (.A(_03252_),
    .ZN(_03253_));
 AND2_X2 _28506_ (.A1(_02714_),
    .A2(_02800_),
    .ZN(_03254_));
 OAI21_X1 _28507_ (.A(_02752_),
    .B1(_03253_),
    .B2(_03254_),
    .ZN(_03255_));
 NAND4_X1 _28508_ (.A1(_03245_),
    .A2(_03249_),
    .A3(_03251_),
    .A4(_03255_),
    .ZN(_03256_));
 OAI21_X1 _28509_ (.A(_02806_),
    .B1(_03253_),
    .B2(_02732_),
    .ZN(_03257_));
 NAND2_X1 _28510_ (.A1(_02807_),
    .A2(_02714_),
    .ZN(_03258_));
 INV_X1 _28511_ (.A(_03258_),
    .ZN(_03259_));
 NAND2_X1 _28512_ (.A1(_03259_),
    .A2(_02796_),
    .ZN(_03260_));
 INV_X1 _28513_ (.A(_02842_),
    .ZN(_03261_));
 AOI22_X1 _28514_ (.A1(_03261_),
    .A2(_02835_),
    .B1(_02864_),
    .B2(_02861_),
    .ZN(_03262_));
 NAND3_X1 _28515_ (.A1(_03257_),
    .A2(_03260_),
    .A3(_03262_),
    .ZN(_03263_));
 NOR4_X4 _28516_ (.A1(_03237_),
    .A2(_03243_),
    .A3(_03256_),
    .A4(_03263_),
    .ZN(_03264_));
 AOI21_X1 _28517_ (.A(_16855_),
    .B1(_02735_),
    .B2(_02707_),
    .ZN(_03265_));
 NAND3_X1 _28518_ (.A1(_02757_),
    .A2(_02743_),
    .A3(_02688_),
    .ZN(_03266_));
 NOR2_X2 _28519_ (.A1(_03265_),
    .A2(_03266_),
    .ZN(_03267_));
 INV_X1 _28520_ (.A(_02890_),
    .ZN(_03268_));
 NAND3_X2 _28521_ (.A1(_02825_),
    .A2(_02807_),
    .A3(_02714_),
    .ZN(_03269_));
 NOR2_X1 _28522_ (.A1(_03268_),
    .A2(_03269_),
    .ZN(_03270_));
 AND2_X2 _28523_ (.A1(_02690_),
    .A2(_02686_),
    .ZN(_03271_));
 AOI211_X2 _28524_ (.A(_03267_),
    .B(_03270_),
    .C1(_03271_),
    .C2(_02883_),
    .ZN(_03272_));
 AND2_X2 _28525_ (.A1(_02708_),
    .A2(_02686_),
    .ZN(_03273_));
 NAND2_X1 _28526_ (.A1(_02697_),
    .A2(_03273_),
    .ZN(_03274_));
 AND2_X1 _28527_ (.A1(_02829_),
    .A2(_02719_),
    .ZN(_03275_));
 AND2_X1 _28528_ (.A1(_02756_),
    .A2(_02877_),
    .ZN(_03276_));
 NOR2_X1 _28529_ (.A1(_03275_),
    .A2(_03276_),
    .ZN(_03277_));
 NAND3_X1 _28530_ (.A1(_02732_),
    .A2(_02845_),
    .A3(_02741_),
    .ZN(_03278_));
 BUF_X8 _28531_ (.A(_02868_),
    .Z(_03279_));
 OAI21_X1 _28532_ (.A(_03279_),
    .B1(_02790_),
    .B2(_02881_),
    .ZN(_03280_));
 AND4_X2 _28533_ (.A1(_03274_),
    .A2(_03277_),
    .A3(_03278_),
    .A4(_03280_),
    .ZN(_03281_));
 OAI21_X1 _28534_ (.A(_02835_),
    .B1(_02902_),
    .B2(_02791_),
    .ZN(_03282_));
 OAI21_X1 _28535_ (.A(_02787_),
    .B1(_02761_),
    .B2(_02756_),
    .ZN(_03283_));
 NAND4_X1 _28536_ (.A1(_02773_),
    .A2(_02686_),
    .A3(_02753_),
    .A4(_02757_),
    .ZN(_03284_));
 NAND2_X1 _28537_ (.A1(_03283_),
    .A2(_03284_),
    .ZN(_03285_));
 AND2_X1 _28538_ (.A1(_02789_),
    .A2(_02818_),
    .ZN(_03286_));
 NOR2_X1 _28539_ (.A1(_03285_),
    .A2(_03286_),
    .ZN(_03287_));
 NAND4_X1 _28540_ (.A1(_03272_),
    .A2(_03281_),
    .A3(_03282_),
    .A4(_03287_),
    .ZN(_03288_));
 OAI21_X1 _28541_ (.A(_02847_),
    .B1(_02767_),
    .B2(_02756_),
    .ZN(_03289_));
 NAND2_X1 _28542_ (.A1(_02731_),
    .A2(_02847_),
    .ZN(_03290_));
 AND2_X1 _28543_ (.A1(_03289_),
    .A2(_03290_),
    .ZN(_03291_));
 OAI21_X1 _28544_ (.A(_03279_),
    .B1(_03248_),
    .B2(_02903_),
    .ZN(_03292_));
 OAI21_X1 _28545_ (.A(_02823_),
    .B1(_02881_),
    .B2(_03254_),
    .ZN(_03293_));
 NAND2_X2 _28546_ (.A1(_02841_),
    .A2(_02714_),
    .ZN(_03294_));
 INV_X1 _28547_ (.A(_03294_),
    .ZN(_03295_));
 NAND2_X1 _28548_ (.A1(_03295_),
    .A2(_02851_),
    .ZN(_03296_));
 NAND4_X1 _28549_ (.A1(_03291_),
    .A2(_03292_),
    .A3(_03293_),
    .A4(_03296_),
    .ZN(_03297_));
 NAND2_X1 _28550_ (.A1(_03248_),
    .A2(_02697_),
    .ZN(_03298_));
 NAND3_X1 _28551_ (.A1(_02870_),
    .A2(_02683_),
    .A3(_02773_),
    .ZN(_03299_));
 AND2_X1 _28552_ (.A1(_03298_),
    .A2(_03299_),
    .ZN(_03300_));
 AND2_X1 _28553_ (.A1(_02714_),
    .A2(_02698_),
    .ZN(_03301_));
 OAI21_X1 _28554_ (.A(_02898_),
    .B1(_03271_),
    .B2(_03301_),
    .ZN(_03302_));
 NAND2_X1 _28555_ (.A1(_02807_),
    .A2(_02858_),
    .ZN(_03303_));
 INV_X1 _28556_ (.A(_03303_),
    .ZN(_03304_));
 AND2_X1 _28557_ (.A1(_03304_),
    .A2(_02897_),
    .ZN(_03305_));
 INV_X1 _28558_ (.A(_03305_),
    .ZN(_03306_));
 NAND2_X1 _28559_ (.A1(_02864_),
    .A2(_02898_),
    .ZN(_03307_));
 NAND4_X1 _28560_ (.A1(_03300_),
    .A2(_03302_),
    .A3(_03306_),
    .A4(_03307_),
    .ZN(_03308_));
 BUF_X4 _28561_ (.A(_02774_),
    .Z(_03309_));
 OAI21_X1 _28562_ (.A(_03309_),
    .B1(_03271_),
    .B2(_02767_),
    .ZN(_03310_));
 OAI21_X1 _28563_ (.A(_02727_),
    .B1(_02781_),
    .B2(_03233_),
    .ZN(_03311_));
 NAND3_X1 _28564_ (.A1(_03309_),
    .A2(_02728_),
    .A3(_02863_),
    .ZN(_03312_));
 NAND3_X1 _28565_ (.A1(_02726_),
    .A2(_02863_),
    .A3(_02859_),
    .ZN(_03313_));
 NAND4_X1 _28566_ (.A1(_03310_),
    .A2(_03311_),
    .A3(_03312_),
    .A4(_03313_),
    .ZN(_03314_));
 NOR4_X2 _28567_ (.A1(_03288_),
    .A2(_03297_),
    .A3(_03308_),
    .A4(_03314_),
    .ZN(_03315_));
 NAND2_X2 _28568_ (.A1(_03264_),
    .A2(_03315_),
    .ZN(_03316_));
 XOR2_X2 _28569_ (.A(_02907_),
    .B(_03316_),
    .Z(_03317_));
 XNOR2_X1 _28570_ (.A(_03213_),
    .B(_03317_),
    .ZN(_03318_));
 XNOR2_X1 _28571_ (.A(_03318_),
    .B(_17219_),
    .ZN(_03319_));
 MUX2_X1 _28572_ (.A(_02938_),
    .B(_03319_),
    .S(_01876_),
    .Z(_00709_));
 XOR2_X1 _28573_ (.A(_17147_),
    .B(_17243_),
    .Z(_03320_));
 XOR2_X1 _28574_ (.A(_01674_),
    .B(_03320_),
    .Z(_03321_));
 XNOR2_X1 _28575_ (.A(_15360_),
    .B(_03321_),
    .ZN(_03322_));
 MUX2_X1 _28576_ (.A(_01233_),
    .B(_03322_),
    .S(_02916_),
    .Z(_01157_));
 XOR2_X1 _28577_ (.A(_17148_),
    .B(_17244_),
    .Z(_03323_));
 XOR2_X1 _28578_ (.A(_01676_),
    .B(_03323_),
    .Z(_03324_));
 XNOR2_X1 _28579_ (.A(_15427_),
    .B(_03324_),
    .ZN(_03325_));
 MUX2_X1 _28580_ (.A(_01234_),
    .B(_03325_),
    .S(_02916_),
    .Z(_01158_));
 XOR2_X1 _28581_ (.A(_17149_),
    .B(_17245_),
    .Z(_03326_));
 XOR2_X1 _28582_ (.A(_01678_),
    .B(_03326_),
    .Z(_03327_));
 XNOR2_X1 _28583_ (.A(_15484_),
    .B(_03327_),
    .ZN(_03328_));
 BUF_X4 _28584_ (.A(_03933_),
    .Z(_03329_));
 MUX2_X1 _28585_ (.A(_01235_),
    .B(_03328_),
    .S(_03329_),
    .Z(_01159_));
 XOR2_X1 _28586_ (.A(_17150_),
    .B(_17246_),
    .Z(_03330_));
 XOR2_X1 _28587_ (.A(_01680_),
    .B(_03330_),
    .Z(_03331_));
 XNOR2_X1 _28588_ (.A(_15543_),
    .B(_03331_),
    .ZN(_03332_));
 MUX2_X1 _28589_ (.A(_01236_),
    .B(_03332_),
    .S(_03329_),
    .Z(_01160_));
 XOR2_X1 _28590_ (.A(_11050_),
    .B(_17215_),
    .Z(_03333_));
 XNOR2_X1 _28591_ (.A(_01812_),
    .B(_03333_),
    .ZN(_03334_));
 XOR2_X1 _28592_ (.A(_15779_),
    .B(_03334_),
    .Z(_03335_));
 MUX2_X1 _28593_ (.A(_01237_),
    .B(_03335_),
    .S(_03329_),
    .Z(_01161_));
 XNOR2_X1 _28594_ (.A(_17184_),
    .B(_17248_),
    .ZN(_03336_));
 XNOR2_X1 _28595_ (.A(_11056_),
    .B(_17216_),
    .ZN(_03337_));
 XOR2_X1 _28596_ (.A(_03336_),
    .B(_03337_),
    .Z(_03338_));
 XNOR2_X1 _28597_ (.A(_15886_),
    .B(_03338_),
    .ZN(_03339_));
 MUX2_X1 _28598_ (.A(_01238_),
    .B(_03339_),
    .S(_03329_),
    .Z(_01162_));
 XOR2_X1 _28599_ (.A(_17153_),
    .B(_17217_),
    .Z(_03340_));
 XNOR2_X1 _28600_ (.A(_01816_),
    .B(_03340_),
    .ZN(_03341_));
 XOR2_X1 _28601_ (.A(_15969_),
    .B(_03341_),
    .Z(_03342_));
 MUX2_X1 _28602_ (.A(_01239_),
    .B(_03342_),
    .S(_03329_),
    .Z(_01163_));
 XOR2_X1 _28603_ (.A(_17154_),
    .B(_17218_),
    .Z(_03343_));
 XOR2_X1 _28604_ (.A(_01819_),
    .B(_03343_),
    .Z(_03344_));
 XNOR2_X1 _28605_ (.A(_01689_),
    .B(_03344_),
    .ZN(_03345_));
 MUX2_X1 _28606_ (.A(_01240_),
    .B(_03345_),
    .S(_03329_),
    .Z(_01164_));
 XOR2_X1 _28607_ (.A(_17188_),
    .B(_17252_),
    .Z(_03346_));
 XOR2_X1 _28608_ (.A(_17156_),
    .B(_17220_),
    .Z(_03347_));
 XNOR2_X1 _28609_ (.A(_03346_),
    .B(_03347_),
    .ZN(_03348_));
 XOR2_X1 _28610_ (.A(_16109_),
    .B(_03348_),
    .Z(_03349_));
 MUX2_X1 _28611_ (.A(_01242_),
    .B(_03349_),
    .S(_03329_),
    .Z(_01166_));
 XOR2_X1 _28612_ (.A(_17189_),
    .B(_17253_),
    .Z(_03350_));
 XOR2_X1 _28613_ (.A(_17157_),
    .B(_17221_),
    .Z(_03351_));
 XNOR2_X1 _28614_ (.A(_03350_),
    .B(_03351_),
    .ZN(_03352_));
 XOR2_X1 _28615_ (.A(_16176_),
    .B(_03352_),
    .Z(_03353_));
 MUX2_X1 _28616_ (.A(_01243_),
    .B(_03353_),
    .S(_03329_),
    .Z(_01167_));
 XOR2_X1 _28617_ (.A(_17230_),
    .B(_17102_),
    .Z(_03354_));
 AND2_X1 _28618_ (.A1(_02133_),
    .A2(_02250_),
    .ZN(_03355_));
 INV_X1 _28619_ (.A(_03355_),
    .ZN(_03356_));
 INV_X1 _28620_ (.A(_03078_),
    .ZN(_03357_));
 OAI211_X2 _28621_ (.A(_03356_),
    .B(_03033_),
    .C1(_03357_),
    .C2(_03034_),
    .ZN(_03358_));
 NAND3_X1 _28622_ (.A1(_02305_),
    .A2(_03032_),
    .A3(_02193_),
    .ZN(_03359_));
 INV_X1 _28623_ (.A(_02230_),
    .ZN(_03360_));
 OAI21_X1 _28624_ (.A(_03359_),
    .B1(_03034_),
    .B2(_03360_),
    .ZN(_03361_));
 OR3_X1 _28625_ (.A1(_03358_),
    .A2(_03016_),
    .A3(_03361_),
    .ZN(_03362_));
 AOI21_X1 _28626_ (.A(_02166_),
    .B1(_02340_),
    .B2(_03360_),
    .ZN(_03363_));
 OAI211_X2 _28627_ (.A(_02176_),
    .B(_02243_),
    .C1(_02173_),
    .C2(_02212_),
    .ZN(_03364_));
 NAND2_X1 _28628_ (.A1(_02153_),
    .A2(_02165_),
    .ZN(_03365_));
 NAND2_X1 _28629_ (.A1(_03364_),
    .A2(_03365_),
    .ZN(_03366_));
 NOR3_X1 _28630_ (.A1(_03362_),
    .A2(_03363_),
    .A3(_03366_),
    .ZN(_03367_));
 NAND2_X1 _28631_ (.A1(_02294_),
    .A2(_02182_),
    .ZN(_03368_));
 OAI21_X1 _28632_ (.A(_02182_),
    .B1(_03078_),
    .B2(_03083_),
    .ZN(_03369_));
 OAI21_X1 _28633_ (.A(_02202_),
    .B1(_02209_),
    .B2(_02192_),
    .ZN(_03370_));
 NAND2_X1 _28634_ (.A1(_03040_),
    .A2(_03039_),
    .ZN(_03371_));
 OAI21_X1 _28635_ (.A(_02202_),
    .B1(_03371_),
    .B2(_02185_),
    .ZN(_03372_));
 AND4_X1 _28636_ (.A1(_03368_),
    .A2(_03369_),
    .A3(_03370_),
    .A4(_03372_),
    .ZN(_03373_));
 OAI21_X1 _28637_ (.A(_02353_),
    .B1(_02294_),
    .B2(_02185_),
    .ZN(_03374_));
 OAI21_X1 _28638_ (.A(_02328_),
    .B1(_02206_),
    .B2(_02320_),
    .ZN(_03375_));
 NAND3_X1 _28639_ (.A1(_02276_),
    .A2(_03032_),
    .A3(_02347_),
    .ZN(_03376_));
 NAND2_X1 _28640_ (.A1(_02327_),
    .A2(_02230_),
    .ZN(_03377_));
 AND3_X1 _28641_ (.A1(_03375_),
    .A2(_03376_),
    .A3(_03377_),
    .ZN(_03378_));
 OAI21_X1 _28642_ (.A(_02353_),
    .B1(_02297_),
    .B2(_02285_),
    .ZN(_03379_));
 OAI211_X2 _28643_ (.A(_02353_),
    .B(_16807_),
    .C1(_03055_),
    .C2(_02135_),
    .ZN(_03380_));
 AND4_X1 _28644_ (.A1(_03374_),
    .A2(_03378_),
    .A3(_03379_),
    .A4(_03380_),
    .ZN(_03381_));
 OAI21_X1 _28645_ (.A(_02334_),
    .B1(_02141_),
    .B2(_02294_),
    .ZN(_03382_));
 AND2_X1 _28646_ (.A1(_03096_),
    .A2(_03097_),
    .ZN(_03383_));
 AOI211_X2 _28647_ (.A(_02345_),
    .B(_03383_),
    .C1(_02185_),
    .C2(_03097_),
    .ZN(_03384_));
 AND2_X1 _28648_ (.A1(_02242_),
    .A2(_02236_),
    .ZN(_03385_));
 OAI21_X1 _28649_ (.A(_02334_),
    .B1(_03385_),
    .B2(_03037_),
    .ZN(_03386_));
 NAND2_X1 _28650_ (.A1(_02206_),
    .A2(_03097_),
    .ZN(_03387_));
 NAND4_X1 _28651_ (.A1(_02214_),
    .A2(_02243_),
    .A3(_02347_),
    .A4(_02268_),
    .ZN(_03388_));
 NAND4_X1 _28652_ (.A1(_02347_),
    .A2(_02191_),
    .A3(_02268_),
    .A4(_02350_),
    .ZN(_03389_));
 AND3_X1 _28653_ (.A1(_03387_),
    .A2(_03388_),
    .A3(_03389_),
    .ZN(_03390_));
 AND4_X1 _28654_ (.A1(_03382_),
    .A2(_03384_),
    .A3(_03386_),
    .A4(_03390_),
    .ZN(_03391_));
 NAND4_X1 _28655_ (.A1(_03367_),
    .A2(_03373_),
    .A3(_03381_),
    .A4(_03391_),
    .ZN(_03392_));
 OAI21_X1 _28656_ (.A(_02262_),
    .B1(_02239_),
    .B2(_02286_),
    .ZN(_03393_));
 INV_X1 _28657_ (.A(_02247_),
    .ZN(_03394_));
 INV_X1 _28658_ (.A(_03037_),
    .ZN(_03395_));
 INV_X1 _28659_ (.A(_02206_),
    .ZN(_03396_));
 AOI21_X1 _28660_ (.A(_03394_),
    .B1(_03395_),
    .B2(_03396_),
    .ZN(_03397_));
 AOI21_X1 _28661_ (.A(_03397_),
    .B1(_02257_),
    .B2(_02247_),
    .ZN(_03398_));
 OAI21_X1 _28662_ (.A(_02262_),
    .B1(_02221_),
    .B2(_02192_),
    .ZN(_03399_));
 OAI21_X1 _28663_ (.A(_02247_),
    .B1(_02189_),
    .B2(_02266_),
    .ZN(_03400_));
 AND4_X1 _28664_ (.A1(_03393_),
    .A2(_03398_),
    .A3(_03399_),
    .A4(_03400_),
    .ZN(_03401_));
 OAI21_X1 _28665_ (.A(_02302_),
    .B1(_02320_),
    .B2(_02221_),
    .ZN(_03402_));
 NAND3_X1 _28666_ (.A1(_02153_),
    .A2(_02194_),
    .A3(_02279_),
    .ZN(_03403_));
 NAND3_X1 _28667_ (.A1(_03402_),
    .A2(_02308_),
    .A3(_03403_),
    .ZN(_03404_));
 NAND2_X1 _28668_ (.A1(_02302_),
    .A2(_02305_),
    .ZN(_03405_));
 NAND2_X1 _28669_ (.A1(_02301_),
    .A2(_03081_),
    .ZN(_03406_));
 INV_X1 _28670_ (.A(_02141_),
    .ZN(_03407_));
 OAI211_X2 _28671_ (.A(_03405_),
    .B(_03406_),
    .C1(_03088_),
    .C2(_03407_),
    .ZN(_03408_));
 AOI21_X1 _28672_ (.A(_03075_),
    .B1(_02154_),
    .B2(_03396_),
    .ZN(_03409_));
 NAND2_X1 _28673_ (.A1(_03073_),
    .A2(_02319_),
    .ZN(_03410_));
 NOR4_X1 _28674_ (.A1(_03404_),
    .A2(_03408_),
    .A3(_03409_),
    .A4(_03410_),
    .ZN(_03411_));
 OAI21_X1 _28675_ (.A(_02275_),
    .B1(_02141_),
    .B2(_02147_),
    .ZN(_03412_));
 OAI21_X1 _28676_ (.A(_02291_),
    .B1(_02141_),
    .B2(_02306_),
    .ZN(_03413_));
 OAI21_X1 _28677_ (.A(_02291_),
    .B1(_03037_),
    .B2(_02192_),
    .ZN(_03414_));
 OAI21_X1 _28678_ (.A(_02275_),
    .B1(_03037_),
    .B2(_02251_),
    .ZN(_03415_));
 AND4_X1 _28679_ (.A1(_03412_),
    .A2(_03413_),
    .A3(_03414_),
    .A4(_03415_),
    .ZN(_03416_));
 AND2_X1 _28680_ (.A1(_03083_),
    .A2(_02241_),
    .ZN(_03417_));
 AND4_X1 _28681_ (.A1(_02214_),
    .A2(_02219_),
    .A3(_02164_),
    .A4(_02252_),
    .ZN(_03418_));
 OR2_X1 _28682_ (.A1(_03417_),
    .A2(_03418_),
    .ZN(_03419_));
 OAI21_X1 _28683_ (.A(_02226_),
    .B1(_02206_),
    .B2(_02320_),
    .ZN(_03420_));
 OAI21_X1 _28684_ (.A(_02226_),
    .B1(_03096_),
    .B2(_02306_),
    .ZN(_03421_));
 NAND3_X1 _28685_ (.A1(_02276_),
    .A2(_03032_),
    .A3(_02252_),
    .ZN(_03422_));
 NAND3_X1 _28686_ (.A1(_03420_),
    .A2(_03421_),
    .A3(_03422_),
    .ZN(_03423_));
 AND3_X1 _28687_ (.A1(_02264_),
    .A2(_02170_),
    .A3(_02241_),
    .ZN(_03424_));
 NOR4_X1 _28688_ (.A1(_03419_),
    .A2(_03423_),
    .A3(_02234_),
    .A4(_03424_),
    .ZN(_03425_));
 NAND4_X1 _28689_ (.A1(_03401_),
    .A2(_03411_),
    .A3(_03416_),
    .A4(_03425_),
    .ZN(_03426_));
 NOR2_X2 _28690_ (.A1(_03392_),
    .A2(_03426_),
    .ZN(_03427_));
 OAI21_X1 _28691_ (.A(_02610_),
    .B1(_02390_),
    .B2(_02527_),
    .ZN(_03428_));
 AND2_X1 _28692_ (.A1(_02380_),
    .A2(_02445_),
    .ZN(_03429_));
 AND2_X2 _28693_ (.A1(_02380_),
    .A2(_02619_),
    .ZN(_03430_));
 BUF_X4 _28694_ (.A(_02375_),
    .Z(_03431_));
 AND3_X1 _28695_ (.A1(_02572_),
    .A2(_03431_),
    .A3(_02378_),
    .ZN(_03432_));
 NOR4_X1 _28696_ (.A1(_03429_),
    .A2(_02941_),
    .A3(_03430_),
    .A4(_03432_),
    .ZN(_03433_));
 OAI21_X1 _28697_ (.A(_02610_),
    .B1(_02416_),
    .B2(_02441_),
    .ZN(_03434_));
 OAI211_X2 _28698_ (.A(_02610_),
    .B(_16767_),
    .C1(_02664_),
    .C2(_02386_),
    .ZN(_03435_));
 AND4_X1 _28699_ (.A1(_03428_),
    .A2(_03433_),
    .A3(_03434_),
    .A4(_03435_),
    .ZN(_03436_));
 BUF_X4 _28700_ (.A(_02466_),
    .Z(_03437_));
 OAI21_X1 _28701_ (.A(_02662_),
    .B1(_02425_),
    .B2(_03437_),
    .ZN(_03438_));
 INV_X1 _28702_ (.A(_02372_),
    .ZN(_03439_));
 OAI21_X1 _28703_ (.A(_03438_),
    .B1(_03439_),
    .B2(_02959_),
    .ZN(_03440_));
 INV_X1 _28704_ (.A(_02413_),
    .ZN(_03441_));
 AOI211_X4 _28705_ (.A(_16767_),
    .B(_03441_),
    .C1(_02664_),
    .C2(_02386_),
    .ZN(_03442_));
 OAI211_X2 _28706_ (.A(_02435_),
    .B(_02991_),
    .C1(_02388_),
    .C2(_02535_),
    .ZN(_03443_));
 NAND2_X1 _28707_ (.A1(_02999_),
    .A2(_02435_),
    .ZN(_03444_));
 NAND2_X1 _28708_ (.A1(_03443_),
    .A2(_03444_),
    .ZN(_03445_));
 NAND3_X1 _28709_ (.A1(_02549_),
    .A2(_03431_),
    .A3(_02472_),
    .ZN(_03446_));
 NAND3_X1 _28710_ (.A1(_02619_),
    .A2(_03431_),
    .A3(_02472_),
    .ZN(_03447_));
 NAND3_X1 _28711_ (.A1(_03446_),
    .A2(_02962_),
    .A3(_03447_),
    .ZN(_03448_));
 NOR4_X1 _28712_ (.A1(_03440_),
    .A2(_03442_),
    .A3(_03445_),
    .A4(_03448_),
    .ZN(_03449_));
 BUF_X4 _28713_ (.A(_02431_),
    .Z(_03450_));
 NAND2_X1 _28714_ (.A1(_02399_),
    .A2(_03450_),
    .ZN(_03451_));
 OAI21_X1 _28715_ (.A(_03450_),
    .B1(_02372_),
    .B2(_02390_),
    .ZN(_03452_));
 OAI21_X1 _28716_ (.A(_02525_),
    .B1(_02505_),
    .B2(_02545_),
    .ZN(_03453_));
 NAND3_X1 _28717_ (.A1(_02602_),
    .A2(_02525_),
    .A3(_02607_),
    .ZN(_03454_));
 AND2_X1 _28718_ (.A1(_03454_),
    .A2(_02969_),
    .ZN(_03455_));
 AND4_X1 _28719_ (.A1(_03451_),
    .A2(_03452_),
    .A3(_03453_),
    .A4(_03455_),
    .ZN(_03456_));
 AND2_X1 _28720_ (.A1(_02539_),
    .A2(_02557_),
    .ZN(_03457_));
 OR3_X1 _28721_ (.A1(_02480_),
    .A2(_03457_),
    .A3(_02603_),
    .ZN(_03458_));
 AOI21_X1 _28722_ (.A(_02606_),
    .B1(_02963_),
    .B2(_02391_),
    .ZN(_03459_));
 INV_X1 _28723_ (.A(_02500_),
    .ZN(_03460_));
 AOI21_X1 _28724_ (.A(_02606_),
    .B1(_02635_),
    .B2(_03460_),
    .ZN(_03461_));
 NAND2_X1 _28725_ (.A1(_02433_),
    .A2(_02474_),
    .ZN(_03462_));
 NAND4_X1 _28726_ (.A1(_02991_),
    .A2(_02598_),
    .A3(_02553_),
    .A4(_02593_),
    .ZN(_03463_));
 INV_X1 _28727_ (.A(_02507_),
    .ZN(_03464_));
 INV_X2 _28728_ (.A(_02474_),
    .ZN(_03465_));
 OAI211_X2 _28729_ (.A(_03462_),
    .B(_03463_),
    .C1(_03464_),
    .C2(_03465_),
    .ZN(_03466_));
 NOR4_X1 _28730_ (.A1(_03458_),
    .A2(_03459_),
    .A3(_03461_),
    .A4(_03466_),
    .ZN(_03467_));
 NAND4_X1 _28731_ (.A1(_03436_),
    .A2(_03449_),
    .A3(_03456_),
    .A4(_03467_),
    .ZN(_03468_));
 OAI21_X1 _28732_ (.A(_02465_),
    .B1(_02953_),
    .B2(_02647_),
    .ZN(_03469_));
 OAI21_X1 _28733_ (.A(_03003_),
    .B1(_02999_),
    .B2(_02434_),
    .ZN(_03470_));
 OAI21_X1 _28734_ (.A(_02465_),
    .B1(_02538_),
    .B2(_02481_),
    .ZN(_03471_));
 AND2_X1 _28735_ (.A1(_03471_),
    .A2(_03007_),
    .ZN(_03472_));
 AND4_X1 _28736_ (.A1(_02596_),
    .A2(_03469_),
    .A3(_03470_),
    .A4(_03472_),
    .ZN(_03473_));
 MUX2_X1 _28737_ (.A(_02490_),
    .B(_02991_),
    .S(_02598_),
    .Z(_03474_));
 AND2_X1 _28738_ (.A1(_03474_),
    .A2(_02449_),
    .ZN(_03475_));
 NAND2_X1 _28739_ (.A1(_02516_),
    .A2(_02434_),
    .ZN(_03476_));
 NAND3_X1 _28740_ (.A1(_02572_),
    .A2(_03431_),
    .A3(_02446_),
    .ZN(_03477_));
 INV_X1 _28741_ (.A(_02445_),
    .ZN(_03478_));
 OAI211_X2 _28742_ (.A(_03476_),
    .B(_03477_),
    .C1(_02453_),
    .C2(_03478_),
    .ZN(_03479_));
 INV_X1 _28743_ (.A(_02539_),
    .ZN(_03480_));
 AOI21_X1 _28744_ (.A(_02453_),
    .B1(_03480_),
    .B2(_02417_),
    .ZN(_03481_));
 NAND2_X1 _28745_ (.A1(_02658_),
    .A2(_02449_),
    .ZN(_03482_));
 INV_X1 _28746_ (.A(_02449_),
    .ZN(_03483_));
 OAI22_X1 _28747_ (.A1(_03482_),
    .A2(_02369_),
    .B1(_02391_),
    .B2(_03483_),
    .ZN(_03484_));
 NOR4_X1 _28748_ (.A1(_03475_),
    .A2(_03479_),
    .A3(_03481_),
    .A4(_03484_),
    .ZN(_03485_));
 OAI21_X1 _28749_ (.A(_02548_),
    .B1(_02538_),
    .B2(_02454_),
    .ZN(_03486_));
 OAI21_X1 _28750_ (.A(_02532_),
    .B1(_02538_),
    .B2(_02416_),
    .ZN(_03487_));
 OAI21_X1 _28751_ (.A(_02532_),
    .B1(_02500_),
    .B2(_02545_),
    .ZN(_03488_));
 OAI21_X1 _28752_ (.A(_02548_),
    .B1(_02500_),
    .B2(_03437_),
    .ZN(_03489_));
 AND4_X1 _28753_ (.A1(_03486_),
    .A2(_03487_),
    .A3(_03488_),
    .A4(_03489_),
    .ZN(_03490_));
 OAI21_X1 _28754_ (.A(_02522_),
    .B1(_02650_),
    .B2(_02545_),
    .ZN(_03491_));
 NAND4_X1 _28755_ (.A1(_02593_),
    .A2(_02383_),
    .A3(_02446_),
    .A4(_02664_),
    .ZN(_03492_));
 NAND3_X1 _28756_ (.A1(_02522_),
    .A2(_02509_),
    .A3(_02371_),
    .ZN(_03493_));
 NAND3_X1 _28757_ (.A1(_03491_),
    .A2(_03492_),
    .A3(_03493_),
    .ZN(_03494_));
 NAND2_X1 _28758_ (.A1(_02614_),
    .A2(_02434_),
    .ZN(_03495_));
 OAI211_X2 _28759_ (.A(_03495_),
    .B(_02629_),
    .C1(_03460_),
    .C2(_02495_),
    .ZN(_03496_));
 INV_X1 _28760_ (.A(_02527_),
    .ZN(_03497_));
 AOI21_X1 _28761_ (.A(_02495_),
    .B1(_02391_),
    .B2(_03497_),
    .ZN(_03498_));
 NOR2_X1 _28762_ (.A1(_02468_),
    .A2(_02598_),
    .ZN(_03499_));
 AND2_X1 _28763_ (.A1(_02614_),
    .A2(_03499_),
    .ZN(_03500_));
 NOR4_X1 _28764_ (.A1(_03494_),
    .A2(_03496_),
    .A3(_03498_),
    .A4(_03500_),
    .ZN(_03501_));
 NAND4_X1 _28765_ (.A1(_03473_),
    .A2(_03485_),
    .A3(_03490_),
    .A4(_03501_),
    .ZN(_03502_));
 NOR2_X2 _28766_ (.A1(_03468_),
    .A2(_03502_),
    .ZN(_03503_));
 XNOR2_X1 _28767_ (.A(_03427_),
    .B(_03503_),
    .ZN(_03504_));
 AND2_X1 _28768_ (.A1(_02001_),
    .A2(_01965_),
    .ZN(_03505_));
 INV_X1 _28769_ (.A(_01965_),
    .ZN(_03506_));
 AOI211_X4 _28770_ (.A(_01931_),
    .B(_03506_),
    .C1(_02118_),
    .C2(_01910_),
    .ZN(_03507_));
 AND2_X1 _28771_ (.A1(_01892_),
    .A2(_02005_),
    .ZN(_03508_));
 AOI211_X4 _28772_ (.A(_03505_),
    .B(_03507_),
    .C1(_03508_),
    .C2(_01966_),
    .ZN(_03509_));
 AND4_X1 _28773_ (.A1(_01924_),
    .A2(_01973_),
    .A3(_01891_),
    .A4(_01908_),
    .ZN(_03510_));
 AOI211_X4 _28774_ (.A(_01931_),
    .B(_02044_),
    .C1(_02022_),
    .C2(_01904_),
    .ZN(_03511_));
 AOI211_X4 _28775_ (.A(_03510_),
    .B(_03511_),
    .C1(_02106_),
    .C2(_03130_),
    .ZN(_03512_));
 OAI211_X2 _28776_ (.A(_03130_),
    .B(_02098_),
    .C1(_02118_),
    .C2(_03159_),
    .ZN(_03513_));
 OAI21_X1 _28777_ (.A(_03130_),
    .B1(_02015_),
    .B2(_03202_),
    .ZN(_03514_));
 NAND4_X1 _28778_ (.A1(_03509_),
    .A2(_03512_),
    .A3(_03513_),
    .A4(_03514_),
    .ZN(_03515_));
 OAI21_X1 _28779_ (.A(_03195_),
    .B1(_02033_),
    .B2(_02034_),
    .ZN(_03516_));
 NOR2_X1 _28780_ (.A1(_01889_),
    .A2(_01934_),
    .ZN(_03517_));
 OAI21_X1 _28781_ (.A(_01981_),
    .B1(_03134_),
    .B2(_03517_),
    .ZN(_03518_));
 AND2_X1 _28782_ (.A1(_02112_),
    .A2(_01979_),
    .ZN(_03519_));
 INV_X1 _28783_ (.A(_03519_),
    .ZN(_03520_));
 OAI21_X1 _28784_ (.A(_03195_),
    .B1(_02122_),
    .B2(_02026_),
    .ZN(_03521_));
 NAND4_X1 _28785_ (.A1(_03516_),
    .A2(_03518_),
    .A3(_03520_),
    .A4(_03521_),
    .ZN(_03522_));
 NAND2_X1 _28786_ (.A1(_03134_),
    .A2(_01992_),
    .ZN(_03523_));
 NAND3_X1 _28787_ (.A1(_02112_),
    .A2(_02006_),
    .A3(_01990_),
    .ZN(_03524_));
 OAI21_X1 _28788_ (.A(_01992_),
    .B1(_02053_),
    .B2(_02106_),
    .ZN(_03525_));
 OAI21_X1 _28789_ (.A(_01991_),
    .B1(_03202_),
    .B2(_02077_),
    .ZN(_03526_));
 NAND4_X1 _28790_ (.A1(_03523_),
    .A2(_03524_),
    .A3(_03525_),
    .A4(_03526_),
    .ZN(_03527_));
 NAND2_X1 _28791_ (.A1(_03154_),
    .A2(_02010_),
    .ZN(_03528_));
 NAND3_X1 _28792_ (.A1(_02010_),
    .A2(_01971_),
    .A3(_01921_),
    .ZN(_03529_));
 NAND2_X1 _28793_ (.A1(_03528_),
    .A2(_03529_),
    .ZN(_03530_));
 NAND2_X1 _28794_ (.A1(_02050_),
    .A2(_02008_),
    .ZN(_03531_));
 NAND3_X1 _28795_ (.A1(_02010_),
    .A2(_01944_),
    .A3(_02099_),
    .ZN(_03532_));
 NAND3_X1 _28796_ (.A1(_02009_),
    .A2(_03161_),
    .A3(_02099_),
    .ZN(_03533_));
 NAND3_X1 _28797_ (.A1(_03531_),
    .A2(_03532_),
    .A3(_03533_),
    .ZN(_03534_));
 OR4_X2 _28798_ (.A1(_02046_),
    .A2(_03527_),
    .A3(_03530_),
    .A4(_03534_),
    .ZN(_03535_));
 AND3_X4 _28799_ (.A1(_01940_),
    .A2(_02006_),
    .A3(_01973_),
    .ZN(_03536_));
 AOI211_X4 _28800_ (.A(_03536_),
    .B(_03138_),
    .C1(_01969_),
    .C2(_02078_),
    .ZN(_03537_));
 NAND2_X1 _28801_ (.A1(_02074_),
    .A2(_02023_),
    .ZN(_03538_));
 OAI21_X1 _28802_ (.A(_01898_),
    .B1(_01959_),
    .B2(_02099_),
    .ZN(_03539_));
 OAI211_X2 _28803_ (.A(_01898_),
    .B(_16847_),
    .C1(_02118_),
    .C2(_01929_),
    .ZN(_03540_));
 NAND4_X1 _28804_ (.A1(_03537_),
    .A2(_03538_),
    .A3(_03539_),
    .A4(_03540_),
    .ZN(_03541_));
 NOR4_X4 _28805_ (.A1(_03515_),
    .A2(_03522_),
    .A3(_03535_),
    .A4(_03541_),
    .ZN(_03542_));
 INV_X1 _28806_ (.A(_02066_),
    .ZN(_03543_));
 INV_X1 _28807_ (.A(_01960_),
    .ZN(_03544_));
 OAI211_X2 _28808_ (.A(_03543_),
    .B(_02091_),
    .C1(_03172_),
    .C2(_03544_),
    .ZN(_03545_));
 AND2_X1 _28809_ (.A1(_01953_),
    .A2(_01945_),
    .ZN(_03546_));
 OR2_X1 _28810_ (.A1(_02087_),
    .A2(_03546_),
    .ZN(_03547_));
 OAI21_X1 _28811_ (.A(_02080_),
    .B1(_02081_),
    .B2(_02061_),
    .ZN(_03548_));
 NAND2_X1 _28812_ (.A1(_02080_),
    .A2(_03154_),
    .ZN(_03549_));
 OAI211_X2 _28813_ (.A(_03548_),
    .B(_03549_),
    .C1(_03167_),
    .C2(_01997_),
    .ZN(_03550_));
 NOR4_X1 _28814_ (.A1(_03545_),
    .A2(_03547_),
    .A3(_01955_),
    .A4(_03550_),
    .ZN(_03551_));
 OAI211_X2 _28815_ (.A(_02070_),
    .B(_02098_),
    .C1(_02118_),
    .C2(_02017_),
    .ZN(_03552_));
 OAI21_X1 _28816_ (.A(_02070_),
    .B1(_02064_),
    .B2(_02061_),
    .ZN(_03553_));
 NAND3_X1 _28817_ (.A1(_01969_),
    .A2(_01925_),
    .A3(_02006_),
    .ZN(_03554_));
 NAND3_X1 _28818_ (.A1(_03552_),
    .A2(_03553_),
    .A3(_03554_),
    .ZN(_03555_));
 AND2_X1 _28819_ (.A1(_02112_),
    .A2(_02123_),
    .ZN(_03556_));
 NAND2_X1 _28820_ (.A1(_03517_),
    .A2(_02123_),
    .ZN(_03557_));
 NAND3_X1 _28821_ (.A1(_02123_),
    .A2(_02098_),
    .A3(_01934_),
    .ZN(_03558_));
 NAND2_X1 _28822_ (.A1(_03557_),
    .A2(_03558_),
    .ZN(_03559_));
 NOR2_X1 _28823_ (.A1(_01995_),
    .A2(_02053_),
    .ZN(_03560_));
 NOR2_X1 _28824_ (.A1(_03560_),
    .A2(_02119_),
    .ZN(_03561_));
 NOR4_X1 _28825_ (.A1(_03555_),
    .A2(_03556_),
    .A3(_03559_),
    .A4(_03561_),
    .ZN(_03562_));
 OAI21_X1 _28826_ (.A(_02014_),
    .B1(_01993_),
    .B2(_01995_),
    .ZN(_03563_));
 OAI21_X1 _28827_ (.A(_01957_),
    .B1(_01993_),
    .B2(_02061_),
    .ZN(_03564_));
 OAI21_X1 _28828_ (.A(_01957_),
    .B1(_02001_),
    .B2(_02026_),
    .ZN(_03565_));
 OAI21_X1 _28829_ (.A(_02014_),
    .B1(_02001_),
    .B2(_02077_),
    .ZN(_03566_));
 AND4_X1 _28830_ (.A1(_03563_),
    .A2(_03564_),
    .A3(_03565_),
    .A4(_03566_),
    .ZN(_03567_));
 OAI21_X1 _28831_ (.A(_02084_),
    .B1(_03133_),
    .B2(_01967_),
    .ZN(_03568_));
 NAND2_X1 _28832_ (.A1(_02084_),
    .A2(_02034_),
    .ZN(_03569_));
 NAND2_X1 _28833_ (.A1(_02037_),
    .A2(_02112_),
    .ZN(_03570_));
 NAND2_X1 _28834_ (.A1(_02037_),
    .A2(_01959_),
    .ZN(_03571_));
 AND3_X1 _28835_ (.A1(_03569_),
    .A2(_03570_),
    .A3(_03571_),
    .ZN(_03572_));
 OAI21_X1 _28836_ (.A(_02103_),
    .B1(_02072_),
    .B2(_02113_),
    .ZN(_03573_));
 OAI21_X1 _28837_ (.A(_02103_),
    .B1(_01949_),
    .B2(_02026_),
    .ZN(_03574_));
 AND4_X1 _28838_ (.A1(_03568_),
    .A2(_03572_),
    .A3(_03573_),
    .A4(_03574_),
    .ZN(_03575_));
 AND4_X1 _28839_ (.A1(_03551_),
    .A2(_03562_),
    .A3(_03567_),
    .A4(_03575_),
    .ZN(_03576_));
 NAND2_X4 _28840_ (.A1(_03542_),
    .A2(_03576_),
    .ZN(_03577_));
 XNOR2_X1 _28841_ (.A(_03504_),
    .B(_03577_),
    .ZN(_03578_));
 NAND3_X1 _28842_ (.A1(_03222_),
    .A2(_02712_),
    .A3(_03233_),
    .ZN(_03579_));
 NAND3_X1 _28843_ (.A1(_03222_),
    .A2(_02735_),
    .A3(_03233_),
    .ZN(_03580_));
 NAND3_X1 _28844_ (.A1(_03222_),
    .A2(_02862_),
    .A3(_03233_),
    .ZN(_03581_));
 NAND3_X1 _28845_ (.A1(_03579_),
    .A2(_03580_),
    .A3(_03581_),
    .ZN(_03582_));
 AND2_X1 _28846_ (.A1(_02790_),
    .A2(_03222_),
    .ZN(_03583_));
 AND2_X1 _28847_ (.A1(_02758_),
    .A2(_02755_),
    .ZN(_03584_));
 AND2_X1 _28848_ (.A1(_03222_),
    .A2(_03254_),
    .ZN(_03585_));
 NOR4_X1 _28849_ (.A1(_03582_),
    .A2(_03583_),
    .A3(_03584_),
    .A4(_03585_),
    .ZN(_03586_));
 NAND2_X1 _28850_ (.A1(_02761_),
    .A2(_02744_),
    .ZN(_03587_));
 INV_X1 _28851_ (.A(_02789_),
    .ZN(_03588_));
 OAI21_X1 _28852_ (.A(_03587_),
    .B1(_03588_),
    .B2(_02769_),
    .ZN(_03589_));
 AND2_X1 _28853_ (.A1(_02812_),
    .A2(_02698_),
    .ZN(_03590_));
 AOI211_X4 _28854_ (.A(_02748_),
    .B(_03589_),
    .C1(_02752_),
    .C2(_03590_),
    .ZN(_03591_));
 INV_X1 _28855_ (.A(_02799_),
    .ZN(_03592_));
 NAND2_X1 _28856_ (.A1(_02825_),
    .A2(_02812_),
    .ZN(_03593_));
 NOR2_X1 _28857_ (.A1(_03592_),
    .A2(_03593_),
    .ZN(_03594_));
 BUF_X4 _28858_ (.A(_02717_),
    .Z(_03595_));
 NAND2_X1 _28859_ (.A1(_02799_),
    .A2(_03595_),
    .ZN(_03596_));
 NAND2_X1 _28860_ (.A1(_02803_),
    .A2(_03596_),
    .ZN(_03597_));
 AOI211_X4 _28861_ (.A(_03594_),
    .B(_03597_),
    .C1(_02848_),
    .C2(_02806_),
    .ZN(_03598_));
 OAI21_X1 _28862_ (.A(_02796_),
    .B1(_03259_),
    .B2(_03273_),
    .ZN(_03599_));
 OAI211_X2 _28863_ (.A(_02796_),
    .B(_02859_),
    .C1(_02735_),
    .C2(_02712_),
    .ZN(_03600_));
 NAND2_X1 _28864_ (.A1(_02869_),
    .A2(_02794_),
    .ZN(_03601_));
 OAI211_X2 _28865_ (.A(_02796_),
    .B(_02858_),
    .C1(_02856_),
    .C2(_02857_),
    .ZN(_03602_));
 AND4_X1 _28866_ (.A1(_03599_),
    .A2(_03600_),
    .A3(_03601_),
    .A4(_03602_),
    .ZN(_03603_));
 AND4_X1 _28867_ (.A1(_03586_),
    .A2(_03591_),
    .A3(_03598_),
    .A4(_03603_),
    .ZN(_03604_));
 AND3_X1 _28868_ (.A1(_02702_),
    .A2(_02757_),
    .A3(_02773_),
    .ZN(_03605_));
 AND2_X1 _28869_ (.A1(_02786_),
    .A2(_02753_),
    .ZN(_03606_));
 AOI211_X4 _28870_ (.A(_03605_),
    .B(_03606_),
    .C1(_02761_),
    .C2(_02787_),
    .ZN(_03607_));
 INV_X1 _28871_ (.A(_03593_),
    .ZN(_03608_));
 NAND2_X1 _28872_ (.A1(_03608_),
    .A2(_02786_),
    .ZN(_03609_));
 INV_X1 _28873_ (.A(_02781_),
    .ZN(_03610_));
 INV_X1 _28874_ (.A(_02787_),
    .ZN(_03611_));
 OAI211_X2 _28875_ (.A(_03607_),
    .B(_03609_),
    .C1(_03610_),
    .C2(_03611_),
    .ZN(_03612_));
 AND2_X1 _28876_ (.A1(_02774_),
    .A2(_02881_),
    .ZN(_03613_));
 AOI21_X1 _28877_ (.A(_02777_),
    .B1(_02901_),
    .B2(_02738_),
    .ZN(_03614_));
 AOI21_X1 _28878_ (.A(_02777_),
    .B1(_02893_),
    .B2(_02894_),
    .ZN(_03615_));
 BUF_X4 _28879_ (.A(_02691_),
    .Z(_03616_));
 AND2_X1 _28880_ (.A1(_02774_),
    .A2(_03616_),
    .ZN(_03617_));
 OR4_X2 _28881_ (.A1(_03613_),
    .A2(_03614_),
    .A3(_03615_),
    .A4(_03617_),
    .ZN(_03618_));
 AND2_X1 _28882_ (.A1(_03259_),
    .A2(_02726_),
    .ZN(_03619_));
 INV_X1 _28883_ (.A(_03619_),
    .ZN(_03620_));
 OAI21_X1 _28884_ (.A(_02727_),
    .B1(_02761_),
    .B2(_02790_),
    .ZN(_03621_));
 INV_X1 _28885_ (.A(_02726_),
    .ZN(_03622_));
 INV_X1 _28886_ (.A(_03590_),
    .ZN(_03623_));
 OAI211_X2 _28887_ (.A(_03620_),
    .B(_03621_),
    .C1(_03622_),
    .C2(_03623_),
    .ZN(_03624_));
 NAND4_X1 _28888_ (.A1(_02773_),
    .A2(_02735_),
    .A3(_03233_),
    .A4(_02683_),
    .ZN(_03625_));
 OAI21_X1 _28889_ (.A(_02697_),
    .B1(_03616_),
    .B2(_02731_),
    .ZN(_03626_));
 NAND4_X1 _28890_ (.A1(_03226_),
    .A2(_02705_),
    .A3(_03625_),
    .A4(_03626_),
    .ZN(_03627_));
 NOR4_X2 _28891_ (.A1(_03612_),
    .A2(_03618_),
    .A3(_03624_),
    .A4(_03627_),
    .ZN(_03628_));
 NAND2_X1 _28892_ (.A1(_02903_),
    .A2(_03279_),
    .ZN(_03629_));
 NAND2_X1 _28893_ (.A1(_03279_),
    .A2(_02801_),
    .ZN(_03630_));
 NAND4_X1 _28894_ (.A1(_02741_),
    .A2(_02811_),
    .A3(_02817_),
    .A4(_02728_),
    .ZN(_03631_));
 AND3_X1 _28895_ (.A1(_03629_),
    .A2(_03630_),
    .A3(_03631_),
    .ZN(_03632_));
 OAI21_X1 _28896_ (.A(_02823_),
    .B1(_02870_),
    .B2(_02732_),
    .ZN(_03633_));
 INV_X2 _28897_ (.A(_02818_),
    .ZN(_03634_));
 OAI211_X2 _28898_ (.A(_02822_),
    .B(_03633_),
    .C1(_02779_),
    .C2(_03634_),
    .ZN(_03635_));
 INV_X1 _28899_ (.A(_02690_),
    .ZN(_03636_));
 AOI211_X4 _28900_ (.A(_03636_),
    .B(_02838_),
    .C1(_02811_),
    .C2(_02800_),
    .ZN(_03637_));
 AND2_X1 _28901_ (.A1(_02778_),
    .A2(_02829_),
    .ZN(_03638_));
 NOR4_X1 _28902_ (.A1(_03635_),
    .A2(_03637_),
    .A3(_02834_),
    .A4(_03638_),
    .ZN(_03639_));
 INV_X1 _28903_ (.A(_02879_),
    .ZN(_03640_));
 OAI21_X1 _28904_ (.A(_02883_),
    .B1(_02902_),
    .B2(_03273_),
    .ZN(_03641_));
 NAND2_X1 _28905_ (.A1(_02831_),
    .A2(_02883_),
    .ZN(_03642_));
 AND2_X2 _28906_ (.A1(_02870_),
    .A2(_02877_),
    .ZN(_03643_));
 INV_X1 _28907_ (.A(_03643_),
    .ZN(_03644_));
 AND4_X1 _28908_ (.A1(_03640_),
    .A2(_03641_),
    .A3(_03642_),
    .A4(_03644_),
    .ZN(_03645_));
 OAI21_X1 _28909_ (.A(_03279_),
    .B1(_02895_),
    .B2(_03616_),
    .ZN(_03646_));
 AND4_X1 _28910_ (.A1(_03632_),
    .A2(_03639_),
    .A3(_03645_),
    .A4(_03646_),
    .ZN(_03647_));
 AND2_X1 _28911_ (.A1(_02846_),
    .A2(_02775_),
    .ZN(_03648_));
 AND2_X1 _28912_ (.A1(_02847_),
    .A2(_03254_),
    .ZN(_03649_));
 AND2_X1 _28913_ (.A1(_02847_),
    .A2(_02715_),
    .ZN(_03650_));
 NOR3_X1 _28914_ (.A1(_03648_),
    .A2(_03649_),
    .A3(_03650_),
    .ZN(_03651_));
 AND2_X2 _28915_ (.A1(_02846_),
    .A2(_02870_),
    .ZN(_03652_));
 INV_X2 _28916_ (.A(_03652_),
    .ZN(_03653_));
 NAND2_X1 _28917_ (.A1(_02846_),
    .A2(_02881_),
    .ZN(_03654_));
 AND2_X2 _28918_ (.A1(_03653_),
    .A2(_03654_),
    .ZN(_03655_));
 OAI21_X1 _28919_ (.A(_02861_),
    .B1(_03248_),
    .B2(_03271_),
    .ZN(_03656_));
 OAI21_X1 _28920_ (.A(_02861_),
    .B1(_02778_),
    .B2(_03301_),
    .ZN(_03657_));
 NAND4_X1 _28921_ (.A1(_03651_),
    .A2(_03655_),
    .A3(_03656_),
    .A4(_03657_),
    .ZN(_03658_));
 AND2_X1 _28922_ (.A1(_02891_),
    .A2(_02719_),
    .ZN(_03659_));
 AND2_X1 _28923_ (.A1(_02891_),
    .A2(_02749_),
    .ZN(_03660_));
 AND2_X1 _28924_ (.A1(_02891_),
    .A2(_02858_),
    .ZN(_03661_));
 AND2_X4 _28925_ (.A1(_02891_),
    .A2(_02694_),
    .ZN(_03662_));
 OR4_X1 _28926_ (.A1(_03659_),
    .A2(_03660_),
    .A3(_03661_),
    .A4(_03662_),
    .ZN(_03663_));
 INV_X1 _28927_ (.A(_02897_),
    .ZN(_03664_));
 AOI21_X1 _28928_ (.A(_03664_),
    .B1(_02783_),
    .B2(_02893_),
    .ZN(_03665_));
 NAND4_X1 _28929_ (.A1(_02845_),
    .A2(_02862_),
    .A3(_02757_),
    .A4(_02728_),
    .ZN(_03666_));
 NAND2_X1 _28930_ (.A1(_03307_),
    .A2(_03666_),
    .ZN(_03667_));
 NOR4_X1 _28931_ (.A1(_03658_),
    .A2(_03663_),
    .A3(_03665_),
    .A4(_03667_),
    .ZN(_03668_));
 AND4_X1 _28932_ (.A1(_03604_),
    .A2(_03628_),
    .A3(_03647_),
    .A4(_03668_),
    .ZN(_03669_));
 INV_X1 _28933_ (.A(_03267_),
    .ZN(_03670_));
 NAND2_X2 _28934_ (.A1(_03669_),
    .A2(_03670_),
    .ZN(_03671_));
 XNOR2_X1 _28935_ (.A(_03671_),
    .B(_03015_),
    .ZN(_03672_));
 XNOR2_X1 _28936_ (.A(_03578_),
    .B(_03672_),
    .ZN(_03673_));
 XNOR2_X1 _28937_ (.A(_03673_),
    .B(_17230_),
    .ZN(_03674_));
 MUX2_X1 _28938_ (.A(_03354_),
    .B(_03674_),
    .S(_01876_),
    .Z(_00710_));
 XOR2_X1 _28939_ (.A(_17190_),
    .B(_17254_),
    .Z(_03675_));
 XOR2_X1 _28940_ (.A(_17158_),
    .B(_17222_),
    .Z(_03676_));
 XNOR2_X1 _28941_ (.A(_03675_),
    .B(_03676_),
    .ZN(_03677_));
 XOR2_X1 _28942_ (.A(_16244_),
    .B(_03677_),
    .Z(_03678_));
 MUX2_X1 _28943_ (.A(_01244_),
    .B(_03678_),
    .S(_03329_),
    .Z(_01168_));
 XOR2_X1 _28944_ (.A(_17191_),
    .B(_17255_),
    .Z(_03679_));
 XOR2_X1 _28945_ (.A(_17159_),
    .B(_17223_),
    .Z(_03680_));
 XNOR2_X1 _28946_ (.A(_03679_),
    .B(_03680_),
    .ZN(_03681_));
 XOR2_X1 _28947_ (.A(_16294_),
    .B(_03681_),
    .Z(_03682_));
 MUX2_X1 _28948_ (.A(_01245_),
    .B(_03682_),
    .S(_03329_),
    .Z(_01169_));
 XNOR2_X1 _28949_ (.A(_11105_),
    .B(_01013_),
    .ZN(_03683_));
 XNOR2_X1 _28950_ (.A(_03683_),
    .B(_17192_),
    .ZN(_03684_));
 XOR2_X1 _28951_ (.A(_17224_),
    .B(_17256_),
    .Z(_03685_));
 XOR2_X1 _28952_ (.A(_03684_),
    .B(_03685_),
    .Z(_03686_));
 XNOR2_X1 _28953_ (.A(_16547_),
    .B(_03686_),
    .ZN(_03687_));
 MUX2_X1 _28954_ (.A(_01246_),
    .B(_03687_),
    .S(_01788_),
    .Z(_01170_));
 XNOR2_X1 _28955_ (.A(_11111_),
    .B(_01015_),
    .ZN(_03688_));
 XNOR2_X1 _28956_ (.A(_03688_),
    .B(_17193_),
    .ZN(_03689_));
 XNOR2_X1 _28957_ (.A(_17225_),
    .B(_17257_),
    .ZN(_03690_));
 XOR2_X1 _28958_ (.A(_03689_),
    .B(_03690_),
    .Z(_03691_));
 XNOR2_X1 _28959_ (.A(_16646_),
    .B(_03691_),
    .ZN(_03692_));
 MUX2_X1 _28960_ (.A(_01247_),
    .B(_03692_),
    .S(_01788_),
    .Z(_01171_));
 XNOR2_X1 _28961_ (.A(_17162_),
    .B(_01017_),
    .ZN(_03693_));
 INV_X1 _28962_ (.A(_17194_),
    .ZN(_03694_));
 XNOR2_X1 _28963_ (.A(_03693_),
    .B(_03694_),
    .ZN(_03695_));
 XOR2_X1 _28964_ (.A(_17226_),
    .B(_17258_),
    .Z(_03696_));
 XOR2_X1 _28965_ (.A(_03695_),
    .B(_03696_),
    .Z(_03697_));
 XNOR2_X1 _28966_ (.A(_16736_),
    .B(_03697_),
    .ZN(_03698_));
 MUX2_X1 _28967_ (.A(_01248_),
    .B(_03698_),
    .S(_01788_),
    .Z(_01172_));
 XNOR2_X1 _28968_ (.A(_17163_),
    .B(_01019_),
    .ZN(_03699_));
 XNOR2_X1 _28969_ (.A(_03699_),
    .B(_17195_),
    .ZN(_03700_));
 XOR2_X1 _28970_ (.A(_17227_),
    .B(_17259_),
    .Z(_03701_));
 XNOR2_X1 _28971_ (.A(_03700_),
    .B(_03701_),
    .ZN(_03702_));
 XNOR2_X1 _28972_ (.A(_01389_),
    .B(_03702_),
    .ZN(_03703_));
 MUX2_X1 _28973_ (.A(_01249_),
    .B(_03703_),
    .S(_01788_),
    .Z(_01173_));
 XNOR2_X1 _28974_ (.A(_17164_),
    .B(_01021_),
    .ZN(_03704_));
 XNOR2_X1 _28975_ (.A(_03704_),
    .B(_17196_),
    .ZN(_03705_));
 XNOR2_X1 _28976_ (.A(_17228_),
    .B(_17260_),
    .ZN(_03706_));
 XOR2_X1 _28977_ (.A(_03705_),
    .B(_03706_),
    .Z(_03707_));
 XNOR2_X1 _28978_ (.A(_01452_),
    .B(_03707_),
    .ZN(_03708_));
 MUX2_X1 _28979_ (.A(_01250_),
    .B(_03708_),
    .S(_01788_),
    .Z(_01174_));
 XOR2_X1 _28980_ (.A(_17165_),
    .B(_01023_),
    .Z(_03709_));
 XNOR2_X1 _28981_ (.A(_03709_),
    .B(_17197_),
    .ZN(_03710_));
 XOR2_X1 _28982_ (.A(_17229_),
    .B(_17261_),
    .Z(_03711_));
 XOR2_X1 _28983_ (.A(_03710_),
    .B(_03711_),
    .Z(_03712_));
 XNOR2_X1 _28984_ (.A(_01515_),
    .B(_03712_),
    .ZN(_03713_));
 MUX2_X1 _28985_ (.A(_01251_),
    .B(_03713_),
    .S(_01788_),
    .Z(_01175_));
 XNOR2_X1 _28986_ (.A(_17167_),
    .B(_01025_),
    .ZN(_03714_));
 XNOR2_X1 _28987_ (.A(_03714_),
    .B(_17199_),
    .ZN(_03715_));
 XOR2_X1 _28988_ (.A(_17231_),
    .B(_17263_),
    .Z(_03716_));
 XNOR2_X1 _28989_ (.A(_03715_),
    .B(_03716_),
    .ZN(_03717_));
 XNOR2_X1 _28990_ (.A(_01569_),
    .B(_03717_),
    .ZN(_03718_));
 MUX2_X1 _28991_ (.A(_01253_),
    .B(_03718_),
    .S(_01788_),
    .Z(_01177_));
 XOR2_X1 _28992_ (.A(_17168_),
    .B(_01027_),
    .Z(_03719_));
 XNOR2_X1 _28993_ (.A(_03719_),
    .B(_17200_),
    .ZN(_03720_));
 XOR2_X1 _28994_ (.A(_17232_),
    .B(_17264_),
    .Z(_03721_));
 XOR2_X1 _28995_ (.A(_03720_),
    .B(_03721_),
    .Z(_03722_));
 XNOR2_X1 _28996_ (.A(_01618_),
    .B(_03722_),
    .ZN(_03723_));
 MUX2_X1 _28997_ (.A(_01254_),
    .B(_03723_),
    .S(_01788_),
    .Z(_01178_));
 XOR2_X1 _28998_ (.A(_17233_),
    .B(_17103_),
    .Z(_03724_));
 XOR2_X2 _28999_ (.A(_02580_),
    .B(_03503_),
    .Z(_03725_));
 NAND4_X1 _29000_ (.A1(_01973_),
    .A2(_02017_),
    .A3(_01924_),
    .A4(_01908_),
    .ZN(_03726_));
 NAND2_X1 _29001_ (.A1(_01965_),
    .A2(_01914_),
    .ZN(_03728_));
 AND2_X1 _29002_ (.A1(_01965_),
    .A2(_02050_),
    .ZN(_03729_));
 AND2_X4 _29003_ (.A1(_01964_),
    .A2(_02090_),
    .ZN(_03730_));
 NOR2_X4 _29004_ (.A1(_03729_),
    .A2(_03730_),
    .ZN(_03731_));
 NAND2_X1 _29005_ (.A1(_01965_),
    .A2(_02106_),
    .ZN(_03732_));
 INV_X1 _29006_ (.A(_03505_),
    .ZN(_03733_));
 AND4_X2 _29007_ (.A1(_03728_),
    .A2(_03731_),
    .A3(_03732_),
    .A4(_03733_),
    .ZN(_03734_));
 OAI211_X2 _29008_ (.A(_03130_),
    .B(_02099_),
    .C1(_03161_),
    .C2(_03159_),
    .ZN(_03735_));
 AND4_X1 _29009_ (.A1(_02022_),
    .A2(_01894_),
    .A3(_01924_),
    .A4(_01888_),
    .ZN(_03736_));
 AOI211_X2 _29010_ (.A(_03736_),
    .B(_03125_),
    .C1(_01951_),
    .C2(_01984_),
    .ZN(_03737_));
 AND4_X4 _29011_ (.A1(_03726_),
    .A2(_03734_),
    .A3(_03735_),
    .A4(_03737_),
    .ZN(_03739_));
 NAND2_X1 _29012_ (.A1(_02015_),
    .A2(_02021_),
    .ZN(_03740_));
 OAI211_X2 _29013_ (.A(_02021_),
    .B(_01903_),
    .C1(_02022_),
    .C2(_01904_),
    .ZN(_03741_));
 OAI211_X2 _29014_ (.A(_02021_),
    .B(_01986_),
    .C1(_01913_),
    .C2(_01891_),
    .ZN(_03742_));
 OAI21_X1 _29015_ (.A(_02021_),
    .B1(_02093_),
    .B2(_02023_),
    .ZN(_03743_));
 AND4_X1 _29016_ (.A1(_03740_),
    .A2(_03741_),
    .A3(_03742_),
    .A4(_03743_),
    .ZN(_03744_));
 NAND2_X1 _29017_ (.A1(_02050_),
    .A2(_01980_),
    .ZN(_03745_));
 OAI211_X2 _29018_ (.A(_01980_),
    .B(_01907_),
    .C1(_01944_),
    .C2(_01934_),
    .ZN(_03746_));
 NAND2_X1 _29019_ (.A1(_01993_),
    .A2(_01980_),
    .ZN(_03747_));
 AND4_X1 _29020_ (.A1(_03745_),
    .A2(_03746_),
    .A3(_03747_),
    .A4(_03206_),
    .ZN(_03748_));
 OAI211_X2 _29021_ (.A(_01981_),
    .B(_01971_),
    .C1(_02118_),
    .C2(_02017_),
    .ZN(_03750_));
 OAI21_X1 _29022_ (.A(_01981_),
    .B1(_03202_),
    .B2(_02077_),
    .ZN(_03751_));
 AND4_X1 _29023_ (.A1(_03744_),
    .A2(_03748_),
    .A3(_03750_),
    .A4(_03751_),
    .ZN(_03752_));
 OAI21_X1 _29024_ (.A(_02008_),
    .B1(_01968_),
    .B2(_02076_),
    .ZN(_03753_));
 OAI211_X2 _29025_ (.A(_02008_),
    .B(_01903_),
    .C1(_01932_),
    .C2(_01904_),
    .ZN(_03754_));
 OAI21_X1 _29026_ (.A(_02008_),
    .B1(_02060_),
    .B2(_02039_),
    .ZN(_03755_));
 AND4_X1 _29027_ (.A1(_03531_),
    .A2(_03753_),
    .A3(_03754_),
    .A4(_03755_),
    .ZN(_03756_));
 NAND2_X1 _29028_ (.A1(_01991_),
    .A2(_02077_),
    .ZN(_03757_));
 OR2_X4 _29029_ (.A1(_02089_),
    .A2(_02050_),
    .ZN(_03758_));
 OAI21_X1 _29030_ (.A(_01991_),
    .B1(_03758_),
    .B2(_02053_),
    .ZN(_03759_));
 AND4_X1 _29031_ (.A1(_02003_),
    .A2(_03756_),
    .A3(_03757_),
    .A4(_03759_),
    .ZN(_03761_));
 OAI21_X1 _29032_ (.A(_01897_),
    .B1(_02050_),
    .B2(_01959_),
    .ZN(_03762_));
 OAI21_X1 _29033_ (.A(_01897_),
    .B1(_03508_),
    .B2(_02122_),
    .ZN(_03763_));
 OAI21_X1 _29034_ (.A(_02078_),
    .B1(_02081_),
    .B2(_02106_),
    .ZN(_03764_));
 OAI21_X1 _29035_ (.A(_02074_),
    .B1(_03134_),
    .B2(_02025_),
    .ZN(_03765_));
 AND4_X1 _29036_ (.A1(_03762_),
    .A2(_03763_),
    .A3(_03764_),
    .A4(_03765_),
    .ZN(_03766_));
 NAND4_X4 _29037_ (.A1(_03739_),
    .A2(_03752_),
    .A3(_03761_),
    .A4(_03766_),
    .ZN(_03767_));
 AND2_X1 _29038_ (.A1(_01903_),
    .A2(_01909_),
    .ZN(_03768_));
 OAI21_X1 _29039_ (.A(_01938_),
    .B1(_03154_),
    .B2(_03768_),
    .ZN(_03769_));
 AND2_X1 _29040_ (.A1(_01953_),
    .A2(_02076_),
    .ZN(_03770_));
 AOI211_X2 _29041_ (.A(_03770_),
    .B(_03546_),
    .C1(_01905_),
    .C2(_01954_),
    .ZN(_03772_));
 OAI21_X1 _29042_ (.A(_01938_),
    .B1(_02072_),
    .B2(_02061_),
    .ZN(_03773_));
 AND2_X1 _29043_ (.A1(_01954_),
    .A2(_01993_),
    .ZN(_03774_));
 NOR3_X1 _29044_ (.A1(_03157_),
    .A2(_03774_),
    .A3(_02066_),
    .ZN(_03775_));
 AND4_X1 _29045_ (.A1(_03769_),
    .A2(_03772_),
    .A3(_03773_),
    .A4(_03775_),
    .ZN(_03776_));
 OAI211_X2 _29046_ (.A(_02013_),
    .B(_01908_),
    .C1(_02022_),
    .C2(_01910_),
    .ZN(_03777_));
 OAI21_X1 _29047_ (.A(_02014_),
    .B1(_01961_),
    .B2(_02054_),
    .ZN(_03778_));
 NAND3_X1 _29048_ (.A1(_03151_),
    .A2(_03777_),
    .A3(_03778_),
    .ZN(_03779_));
 OAI21_X1 _29049_ (.A(_01920_),
    .B1(_02015_),
    .B2(_01967_),
    .ZN(_03780_));
 OAI21_X1 _29050_ (.A(_03780_),
    .B1(_02116_),
    .B2(_03143_),
    .ZN(_03781_));
 INV_X1 _29051_ (.A(_02121_),
    .ZN(_03783_));
 AOI21_X1 _29052_ (.A(_03143_),
    .B1(_03783_),
    .B2(_01997_),
    .ZN(_03784_));
 AND2_X1 _29053_ (.A1(_01920_),
    .A2(_02060_),
    .ZN(_03785_));
 AND2_X1 _29054_ (.A1(_01920_),
    .A2(_02081_),
    .ZN(_03786_));
 OR2_X2 _29055_ (.A1(_03785_),
    .A2(_03786_),
    .ZN(_03787_));
 NOR4_X4 _29056_ (.A1(_03779_),
    .A2(_03781_),
    .A3(_03784_),
    .A4(_03787_),
    .ZN(_03788_));
 NAND2_X1 _29057_ (.A1(_01940_),
    .A2(_02097_),
    .ZN(_03789_));
 OAI21_X1 _29058_ (.A(_02069_),
    .B1(_01939_),
    .B2(_01949_),
    .ZN(_03790_));
 NAND2_X2 _29059_ (.A1(_02069_),
    .A2(_03202_),
    .ZN(_03791_));
 NAND2_X1 _29060_ (.A1(_02069_),
    .A2(_02034_),
    .ZN(_03792_));
 NAND2_X1 _29061_ (.A1(_02069_),
    .A2(_02032_),
    .ZN(_03793_));
 AND4_X2 _29062_ (.A1(_03790_),
    .A2(_03791_),
    .A3(_03792_),
    .A4(_03793_),
    .ZN(_03794_));
 OAI21_X1 _29063_ (.A(_02097_),
    .B1(_02072_),
    .B2(_02082_),
    .ZN(_03795_));
 OAI211_X2 _29064_ (.A(_02097_),
    .B(_02025_),
    .C1(_01934_),
    .C2(_01891_),
    .ZN(_03796_));
 AND4_X1 _29065_ (.A1(_03789_),
    .A2(_03794_),
    .A3(_03795_),
    .A4(_03796_),
    .ZN(_03797_));
 NAND2_X1 _29066_ (.A1(_03202_),
    .A2(_02103_),
    .ZN(_03798_));
 OAI21_X1 _29067_ (.A(_02103_),
    .B1(_02090_),
    .B2(_02050_),
    .ZN(_03799_));
 OAI21_X1 _29068_ (.A(_02037_),
    .B1(_02053_),
    .B2(_02081_),
    .ZN(_03800_));
 NAND2_X1 _29069_ (.A1(_02037_),
    .A2(_01945_),
    .ZN(_03801_));
 AND4_X1 _29070_ (.A1(_03798_),
    .A2(_03799_),
    .A3(_03800_),
    .A4(_03801_),
    .ZN(_03802_));
 NAND4_X4 _29071_ (.A1(_03776_),
    .A2(_03788_),
    .A3(_03797_),
    .A4(_03802_),
    .ZN(_03804_));
 NOR2_X4 _29072_ (.A1(_03767_),
    .A2(_03804_),
    .ZN(_03805_));
 XNOR2_X1 _29073_ (.A(_03725_),
    .B(_03805_),
    .ZN(_03806_));
 INV_X2 _29074_ (.A(_02327_),
    .ZN(_03807_));
 INV_X1 _29075_ (.A(_02318_),
    .ZN(_03808_));
 OAI21_X1 _29076_ (.A(_03377_),
    .B1(_03807_),
    .B2(_03808_),
    .ZN(_03809_));
 AND2_X1 _29077_ (.A1(_03078_),
    .A2(_02327_),
    .ZN(_03810_));
 AOI211_X2 _29078_ (.A(_03809_),
    .B(_03810_),
    .C1(_02191_),
    .C2(_02328_),
    .ZN(_03811_));
 OAI21_X1 _29079_ (.A(_02353_),
    .B1(_03385_),
    .B2(_02208_),
    .ZN(_03812_));
 NAND4_X1 _29080_ (.A1(_02237_),
    .A2(_02347_),
    .A3(_02220_),
    .A4(_02280_),
    .ZN(_03813_));
 AND3_X1 _29081_ (.A1(_03812_),
    .A2(_03379_),
    .A3(_03813_),
    .ZN(_03815_));
 AOI211_X2 _29082_ (.A(_02340_),
    .B(_03094_),
    .C1(_03055_),
    .C2(_02174_),
    .ZN(_03816_));
 AND4_X1 _29083_ (.A1(_02212_),
    .A2(_02347_),
    .A3(_02146_),
    .A4(_02267_),
    .ZN(_03817_));
 OAI211_X2 _29084_ (.A(_03097_),
    .B(_02219_),
    .C1(_02220_),
    .C2(_02169_),
    .ZN(_03818_));
 INV_X1 _29085_ (.A(_02251_),
    .ZN(_03819_));
 OAI211_X2 _29086_ (.A(_03818_),
    .B(_03093_),
    .C1(_03819_),
    .C2(_03094_),
    .ZN(_03820_));
 NOR3_X1 _29087_ (.A1(_03816_),
    .A2(_03817_),
    .A3(_03820_),
    .ZN(_03821_));
 AND2_X1 _29088_ (.A1(_02331_),
    .A2(_02198_),
    .ZN(_03822_));
 AND2_X4 _29089_ (.A1(_02331_),
    .A2(_03081_),
    .ZN(_03823_));
 NOR2_X1 _29090_ (.A1(_03822_),
    .A2(_03823_),
    .ZN(_03824_));
 INV_X1 _29091_ (.A(_03824_),
    .ZN(_03826_));
 AND2_X1 _29092_ (.A1(_03037_),
    .A2(_02331_),
    .ZN(_03827_));
 NOR4_X4 _29093_ (.A1(_03826_),
    .A2(_02332_),
    .A3(_03111_),
    .A4(_03827_),
    .ZN(_03828_));
 NAND4_X2 _29094_ (.A1(_03811_),
    .A2(_03815_),
    .A3(_03821_),
    .A4(_03828_),
    .ZN(_03829_));
 OAI211_X2 _29095_ (.A(_02181_),
    .B(_02146_),
    .C1(_02214_),
    .C2(_02139_),
    .ZN(_03830_));
 OAI211_X2 _29096_ (.A(_02181_),
    .B(_02237_),
    .C1(_03055_),
    .C2(_02350_),
    .ZN(_03831_));
 OAI211_X2 _29097_ (.A(_02181_),
    .B(_02243_),
    .C1(_03055_),
    .C2(_02212_),
    .ZN(_03832_));
 OAI21_X1 _29098_ (.A(_02181_),
    .B1(_02346_),
    .B2(_02250_),
    .ZN(_03833_));
 AND4_X1 _29099_ (.A1(_03830_),
    .A2(_03831_),
    .A3(_03832_),
    .A4(_03833_),
    .ZN(_03834_));
 NAND2_X1 _29100_ (.A1(_02335_),
    .A2(_02201_),
    .ZN(_03835_));
 NAND2_X1 _29101_ (.A1(_02208_),
    .A2(_02202_),
    .ZN(_03837_));
 AND3_X1 _29102_ (.A1(_03835_),
    .A2(_03837_),
    .A3(_02215_),
    .ZN(_03838_));
 OAI21_X1 _29103_ (.A(_02202_),
    .B1(_02359_),
    .B2(_02230_),
    .ZN(_03839_));
 OAI211_X2 _29104_ (.A(_02202_),
    .B(_02266_),
    .C1(_02220_),
    .C2(_02169_),
    .ZN(_03840_));
 NAND4_X1 _29105_ (.A1(_03834_),
    .A2(_03838_),
    .A3(_03839_),
    .A4(_03840_),
    .ZN(_03841_));
 OAI21_X1 _29106_ (.A(_02176_),
    .B1(_02276_),
    .B2(_02251_),
    .ZN(_03842_));
 OAI211_X2 _29107_ (.A(_02176_),
    .B(_02243_),
    .C1(_03055_),
    .C2(_02212_),
    .ZN(_03843_));
 OAI21_X1 _29108_ (.A(_02176_),
    .B1(_02306_),
    .B2(_02286_),
    .ZN(_03844_));
 NAND4_X1 _29109_ (.A1(_02266_),
    .A2(_02193_),
    .A3(_02220_),
    .A4(_02280_),
    .ZN(_03845_));
 NAND4_X1 _29110_ (.A1(_03842_),
    .A2(_03843_),
    .A3(_03844_),
    .A4(_03845_),
    .ZN(_03846_));
 AND3_X1 _29111_ (.A1(_02305_),
    .A2(_03032_),
    .A3(_02193_),
    .ZN(_03848_));
 AND3_X2 _29112_ (.A1(_02341_),
    .A2(_02134_),
    .A3(_02167_),
    .ZN(_03849_));
 AND2_X1 _29113_ (.A1(_02133_),
    .A2(_02218_),
    .ZN(_03850_));
 OR4_X4 _29114_ (.A1(_03848_),
    .A2(_03849_),
    .A3(_03355_),
    .A4(_03850_),
    .ZN(_03851_));
 NOR4_X4 _29115_ (.A1(_03829_),
    .A2(_03841_),
    .A3(_03846_),
    .A4(_03851_),
    .ZN(_03852_));
 NAND2_X1 _29116_ (.A1(_02226_),
    .A2(_02185_),
    .ZN(_03853_));
 OAI21_X1 _29117_ (.A(_02225_),
    .B1(_02359_),
    .B2(_02230_),
    .ZN(_03854_));
 AND3_X1 _29118_ (.A1(_02346_),
    .A2(_02324_),
    .A3(_02223_),
    .ZN(_03855_));
 INV_X1 _29119_ (.A(_03855_),
    .ZN(_03856_));
 AND4_X1 _29120_ (.A1(_02227_),
    .A2(_03853_),
    .A3(_03854_),
    .A4(_03856_),
    .ZN(_03857_));
 NAND4_X1 _29121_ (.A1(_02211_),
    .A2(_02280_),
    .A3(_02252_),
    .A4(_02212_),
    .ZN(_03858_));
 OAI211_X2 _29122_ (.A(_02241_),
    .B(_02266_),
    .C1(_02214_),
    .C2(_02139_),
    .ZN(_03859_));
 AND2_X1 _29123_ (.A1(_02346_),
    .A2(_02233_),
    .ZN(_03860_));
 AND3_X1 _29124_ (.A1(_02233_),
    .A2(_02144_),
    .A3(_02151_),
    .ZN(_03861_));
 AOI211_X2 _29125_ (.A(_03860_),
    .B(_03861_),
    .C1(_02320_),
    .C2(_02233_),
    .ZN(_03862_));
 NAND4_X1 _29126_ (.A1(_03857_),
    .A2(_03858_),
    .A3(_03859_),
    .A4(_03862_),
    .ZN(_03863_));
 OAI21_X1 _29127_ (.A(_02290_),
    .B1(_02205_),
    .B2(_02208_),
    .ZN(_03864_));
 NAND2_X1 _29128_ (.A1(_02290_),
    .A2(_02318_),
    .ZN(_03865_));
 NAND2_X1 _29129_ (.A1(_02290_),
    .A2(_02191_),
    .ZN(_03866_));
 NAND4_X1 _29130_ (.A1(_03864_),
    .A2(_02298_),
    .A3(_03865_),
    .A4(_03866_),
    .ZN(_03867_));
 AOI21_X1 _29131_ (.A(_02284_),
    .B1(_03039_),
    .B2(_03360_),
    .ZN(_03869_));
 NAND4_X1 _29132_ (.A1(_02273_),
    .A2(_02139_),
    .A3(_02219_),
    .A4(_02164_),
    .ZN(_03870_));
 AND2_X4 _29133_ (.A1(_02151_),
    .A2(_02137_),
    .ZN(_03871_));
 INV_X1 _29134_ (.A(_03871_),
    .ZN(_03872_));
 OAI21_X1 _29135_ (.A(_03870_),
    .B1(_02284_),
    .B2(_03872_),
    .ZN(_03873_));
 OR4_X1 _29136_ (.A1(_03067_),
    .A2(_03867_),
    .A3(_03869_),
    .A4(_03873_),
    .ZN(_03874_));
 OAI21_X1 _29137_ (.A(_02313_),
    .B1(_02239_),
    .B2(_02306_),
    .ZN(_03875_));
 OAI21_X1 _29138_ (.A(_02301_),
    .B1(_02314_),
    .B2(_02292_),
    .ZN(_03876_));
 AND2_X1 _29139_ (.A1(_02219_),
    .A2(_02137_),
    .ZN(_03877_));
 OAI21_X1 _29140_ (.A(_02313_),
    .B1(_02153_),
    .B2(_03877_),
    .ZN(_03878_));
 OAI21_X1 _29141_ (.A(_02301_),
    .B1(_02141_),
    .B2(_02264_),
    .ZN(_03880_));
 NAND4_X1 _29142_ (.A1(_03875_),
    .A2(_03876_),
    .A3(_03878_),
    .A4(_03880_),
    .ZN(_03881_));
 AND2_X4 _29143_ (.A1(_02346_),
    .A2(_02258_),
    .ZN(_03882_));
 INV_X1 _29144_ (.A(_03081_),
    .ZN(_03883_));
 NAND2_X1 _29145_ (.A1(_02338_),
    .A2(_03883_),
    .ZN(_03884_));
 AOI21_X1 _29146_ (.A(_03882_),
    .B1(_03884_),
    .B2(_02262_),
    .ZN(_03885_));
 NAND2_X1 _29147_ (.A1(_02247_),
    .A2(_02318_),
    .ZN(_03886_));
 NAND2_X1 _29148_ (.A1(_02305_),
    .A2(_02246_),
    .ZN(_03887_));
 NAND2_X1 _29149_ (.A1(_02247_),
    .A2(_02153_),
    .ZN(_03888_));
 NAND4_X1 _29150_ (.A1(_03885_),
    .A2(_03886_),
    .A3(_03887_),
    .A4(_03888_),
    .ZN(_03889_));
 NOR4_X1 _29151_ (.A1(_03863_),
    .A2(_03874_),
    .A3(_03881_),
    .A4(_03889_),
    .ZN(_03891_));
 NAND2_X1 _29152_ (.A1(_03852_),
    .A2(_03891_),
    .ZN(_03892_));
 AND2_X1 _29153_ (.A1(_02499_),
    .A2(_02506_),
    .ZN(_03893_));
 OAI21_X1 _29154_ (.A(_03003_),
    .B1(_02999_),
    .B2(_03893_),
    .ZN(_03894_));
 AND2_X1 _29155_ (.A1(_02464_),
    .A2(_02564_),
    .ZN(_03895_));
 INV_X1 _29156_ (.A(_02571_),
    .ZN(_03896_));
 OAI21_X1 _29157_ (.A(_02566_),
    .B1(_02469_),
    .B2(_03896_),
    .ZN(_03897_));
 AOI211_X2 _29158_ (.A(_03895_),
    .B(_03897_),
    .C1(_02466_),
    .C2(_02465_),
    .ZN(_03898_));
 OAI21_X1 _29159_ (.A(_03003_),
    .B1(_02615_),
    .B2(_02416_),
    .ZN(_03899_));
 NAND3_X1 _29160_ (.A1(_02538_),
    .A2(_02672_),
    .A3(_02429_),
    .ZN(_03900_));
 AND3_X1 _29161_ (.A1(_03007_),
    .A2(_03900_),
    .A3(_03008_),
    .ZN(_03901_));
 AND4_X1 _29162_ (.A1(_03894_),
    .A2(_03898_),
    .A3(_03899_),
    .A4(_03901_),
    .ZN(_03902_));
 AOI21_X1 _29163_ (.A(_03483_),
    .B1(_02963_),
    .B2(_03480_),
    .ZN(_03903_));
 AOI21_X1 _29164_ (.A(_03903_),
    .B1(_02528_),
    .B2(_02449_),
    .ZN(_03904_));
 OAI21_X1 _29165_ (.A(_02516_),
    .B1(_02647_),
    .B2(_02425_),
    .ZN(_03905_));
 AND2_X1 _29166_ (.A1(_02451_),
    .A2(_02463_),
    .ZN(_03906_));
 INV_X1 _29167_ (.A(_03906_),
    .ZN(_03907_));
 OAI21_X1 _29168_ (.A(_02516_),
    .B1(_02419_),
    .B2(_02619_),
    .ZN(_03908_));
 AND3_X1 _29169_ (.A1(_03905_),
    .A2(_03907_),
    .A3(_03908_),
    .ZN(_03909_));
 AND2_X1 _29170_ (.A1(_02425_),
    .A2(_02448_),
    .ZN(_03910_));
 AND3_X1 _29171_ (.A1(_02447_),
    .A2(_02394_),
    .A3(_02398_),
    .ZN(_03912_));
 AOI211_X2 _29172_ (.A(_03910_),
    .B(_03912_),
    .C1(_02572_),
    .C2(_02448_),
    .ZN(_03913_));
 NAND2_X1 _29173_ (.A1(_02425_),
    .A2(_02522_),
    .ZN(_03914_));
 OAI21_X1 _29174_ (.A(_02614_),
    .B1(_02549_),
    .B2(_02439_),
    .ZN(_03915_));
 NAND3_X1 _29175_ (.A1(_02599_),
    .A2(_02403_),
    .A3(_02504_),
    .ZN(_03916_));
 AND4_X1 _29176_ (.A1(_03914_),
    .A2(_03915_),
    .A3(_03916_),
    .A4(_02569_),
    .ZN(_03917_));
 AND4_X1 _29177_ (.A1(_03904_),
    .A2(_03909_),
    .A3(_03913_),
    .A4(_03917_),
    .ZN(_03918_));
 AOI211_X4 _29178_ (.A(_02468_),
    .B(_02543_),
    .C1(_02664_),
    .C2(_02535_),
    .ZN(_03919_));
 AND2_X1 _29179_ (.A1(_02976_),
    .A2(_02548_),
    .ZN(_03920_));
 AND4_X1 _29180_ (.A1(_02506_),
    .A2(_02672_),
    .A3(_02490_),
    .A4(_02944_),
    .ZN(_03921_));
 AND4_X1 _29181_ (.A1(_02672_),
    .A2(_02991_),
    .A3(_02402_),
    .A4(_02944_),
    .ZN(_03923_));
 NOR4_X1 _29182_ (.A1(_03919_),
    .A2(_03920_),
    .A3(_03921_),
    .A4(_03923_),
    .ZN(_03924_));
 OAI21_X1 _29183_ (.A(_02532_),
    .B1(_02466_),
    .B2(_02445_),
    .ZN(_03925_));
 OAI211_X2 _29184_ (.A(_02672_),
    .B(_03431_),
    .C1(_02439_),
    .C2(_02416_),
    .ZN(_03926_));
 NAND2_X1 _29185_ (.A1(_02532_),
    .A2(_02505_),
    .ZN(_03927_));
 AND4_X1 _29186_ (.A1(_02995_),
    .A2(_03925_),
    .A3(_03926_),
    .A4(_03927_),
    .ZN(_03928_));
 AND4_X2 _29187_ (.A1(_03902_),
    .A2(_03918_),
    .A3(_03924_),
    .A4(_03928_),
    .ZN(_03929_));
 AND2_X1 _29188_ (.A1(_02485_),
    .A2(_02525_),
    .ZN(_03930_));
 AND2_X1 _29189_ (.A1(_02457_),
    .A2(_02524_),
    .ZN(_03931_));
 AND3_X1 _29190_ (.A1(_02524_),
    .A2(_02394_),
    .A3(_02398_),
    .ZN(_03932_));
 OR3_X2 _29191_ (.A1(_02561_),
    .A2(_03931_),
    .A3(_03932_),
    .ZN(_03934_));
 AND2_X1 _29192_ (.A1(_02481_),
    .A2(_02525_),
    .ZN(_03935_));
 AOI211_X4 _29193_ (.A(_02468_),
    .B(_02642_),
    .C1(_02664_),
    .C2(_02535_),
    .ZN(_03936_));
 OR4_X4 _29194_ (.A1(_03930_),
    .A2(_03934_),
    .A3(_03935_),
    .A4(_03936_),
    .ZN(_03937_));
 AND2_X1 _29195_ (.A1(_02487_),
    .A2(_02556_),
    .ZN(_03938_));
 AND2_X1 _29196_ (.A1(_02556_),
    .A2(_02423_),
    .ZN(_03939_));
 NOR4_X1 _29197_ (.A1(_03938_),
    .A2(_02574_),
    .A3(_03939_),
    .A4(_02948_),
    .ZN(_03940_));
 AND2_X1 _29198_ (.A1(_02505_),
    .A2(_02414_),
    .ZN(_03941_));
 AOI21_X1 _29199_ (.A(_03941_),
    .B1(_02953_),
    .B2(_02610_),
    .ZN(_03942_));
 NAND4_X1 _29200_ (.A1(_02581_),
    .A2(_02553_),
    .A3(_02621_),
    .A4(_02944_),
    .ZN(_03943_));
 AND3_X1 _29201_ (.A1(_03942_),
    .A2(_03434_),
    .A3(_03943_),
    .ZN(_03945_));
 AND3_X1 _29202_ (.A1(_02439_),
    .A2(_03431_),
    .A3(_02378_),
    .ZN(_03946_));
 NOR4_X1 _29203_ (.A1(_02381_),
    .A2(_02940_),
    .A3(_03430_),
    .A4(_03946_),
    .ZN(_03947_));
 NAND4_X1 _29204_ (.A1(_02553_),
    .A2(_02535_),
    .A3(_02593_),
    .A4(_02383_),
    .ZN(_03948_));
 NAND4_X1 _29205_ (.A1(_02581_),
    .A2(_02553_),
    .A3(_02621_),
    .A4(_02593_),
    .ZN(_03949_));
 OAI211_X2 _29206_ (.A(_03948_),
    .B(_03949_),
    .C1(_02391_),
    .C2(_03465_),
    .ZN(_03950_));
 NAND2_X1 _29207_ (.A1(_02999_),
    .A2(_02557_),
    .ZN(_03951_));
 OAI21_X1 _29208_ (.A(_03951_),
    .B1(_03465_),
    .B2(_03005_),
    .ZN(_03952_));
 AND3_X1 _29209_ (.A1(_02591_),
    .A2(_02557_),
    .A3(_02403_),
    .ZN(_03953_));
 NOR3_X1 _29210_ (.A1(_03950_),
    .A2(_03952_),
    .A3(_03953_),
    .ZN(_03954_));
 NAND4_X1 _29211_ (.A1(_03940_),
    .A2(_03945_),
    .A3(_03947_),
    .A4(_03954_),
    .ZN(_03956_));
 OAI211_X2 _29212_ (.A(_03450_),
    .B(_02383_),
    .C1(_02598_),
    .C2(_02402_),
    .ZN(_03957_));
 OAI211_X2 _29213_ (.A(_03450_),
    .B(_02581_),
    .C1(_02664_),
    .C2(_02506_),
    .ZN(_03958_));
 OAI211_X2 _29214_ (.A(_03450_),
    .B(_02991_),
    .C1(_02664_),
    .C2(_02535_),
    .ZN(_03959_));
 OAI21_X1 _29215_ (.A(_03450_),
    .B1(_02425_),
    .B2(_03437_),
    .ZN(_03960_));
 NAND4_X1 _29216_ (.A1(_03957_),
    .A2(_03958_),
    .A3(_03959_),
    .A4(_03960_),
    .ZN(_03961_));
 AOI21_X1 _29217_ (.A(_03441_),
    .B1(_03005_),
    .B2(_03478_),
    .ZN(_03962_));
 AND2_X1 _29218_ (.A1(_02434_),
    .A2(_02435_),
    .ZN(_03963_));
 NOR3_X1 _29219_ (.A1(_03962_),
    .A2(_03963_),
    .A3(_02644_),
    .ZN(_03964_));
 OAI21_X1 _29220_ (.A(_02435_),
    .B1(_02485_),
    .B2(_03499_),
    .ZN(_03965_));
 OAI21_X1 _29221_ (.A(_02662_),
    .B1(_02487_),
    .B2(_02549_),
    .ZN(_03967_));
 OAI21_X1 _29222_ (.A(_02662_),
    .B1(_02572_),
    .B2(_03437_),
    .ZN(_03968_));
 NAND4_X1 _29223_ (.A1(_03964_),
    .A2(_03965_),
    .A3(_03967_),
    .A4(_03968_),
    .ZN(_03969_));
 NOR4_X4 _29224_ (.A1(_03937_),
    .A2(_03956_),
    .A3(_03961_),
    .A4(_03969_),
    .ZN(_03970_));
 NAND2_X4 _29225_ (.A1(_03929_),
    .A2(_03970_),
    .ZN(_03971_));
 XOR2_X1 _29226_ (.A(_03892_),
    .B(_03971_),
    .Z(_03972_));
 AND2_X1 _29227_ (.A1(_02829_),
    .A2(_02791_),
    .ZN(_03973_));
 NOR2_X1 _29228_ (.A1(_03973_),
    .A2(_02832_),
    .ZN(_03974_));
 OAI21_X1 _29229_ (.A(_02835_),
    .B1(_03616_),
    .B2(_02731_),
    .ZN(_03975_));
 OAI211_X2 _29230_ (.A(_03974_),
    .B(_03975_),
    .C1(_02838_),
    .C2(_02886_),
    .ZN(_03976_));
 NAND4_X1 _29231_ (.A1(_02858_),
    .A2(_02817_),
    .A3(_02683_),
    .A4(_02811_),
    .ZN(_03978_));
 OAI21_X1 _29232_ (.A(_03978_),
    .B1(_03588_),
    .B2(_03634_),
    .ZN(_03979_));
 AND4_X1 _29233_ (.A1(_02841_),
    .A2(_02823_),
    .A3(_02728_),
    .A4(_02863_),
    .ZN(_03980_));
 NOR4_X1 _29234_ (.A1(_03976_),
    .A2(_02821_),
    .A3(_03979_),
    .A4(_03980_),
    .ZN(_03981_));
 NAND2_X1 _29235_ (.A1(_02863_),
    .A2(_02714_),
    .ZN(_03982_));
 OR2_X1 _29236_ (.A1(_03664_),
    .A2(_03982_),
    .ZN(_03983_));
 AND2_X1 _29237_ (.A1(_02891_),
    .A2(_02870_),
    .ZN(_03984_));
 AND2_X1 _29238_ (.A1(_02891_),
    .A2(_02756_),
    .ZN(_03985_));
 AND2_X1 _29239_ (.A1(_02891_),
    .A2(_03254_),
    .ZN(_03986_));
 NOR4_X1 _29240_ (.A1(_03984_),
    .A2(_03985_),
    .A3(_03986_),
    .A4(_03662_),
    .ZN(_03987_));
 NAND2_X1 _29241_ (.A1(_02898_),
    .A2(_03233_),
    .ZN(_03988_));
 OAI211_X2 _29242_ (.A(_02898_),
    .B(_16855_),
    .C1(_02857_),
    .C2(_02707_),
    .ZN(_03989_));
 AND4_X1 _29243_ (.A1(_03983_),
    .A2(_03987_),
    .A3(_03988_),
    .A4(_03989_),
    .ZN(_03990_));
 INV_X1 _29244_ (.A(_02878_),
    .ZN(_03991_));
 OAI211_X2 _29245_ (.A(_02883_),
    .B(_02859_),
    .C1(_02811_),
    .C2(_02800_),
    .ZN(_03992_));
 NAND2_X1 _29246_ (.A1(_03991_),
    .A2(_03992_),
    .ZN(_03993_));
 OAI211_X2 _29247_ (.A(_03279_),
    .B(_02859_),
    .C1(_02712_),
    .C2(_02862_),
    .ZN(_03994_));
 OAI21_X1 _29248_ (.A(_02868_),
    .B1(_02715_),
    .B2(_03254_),
    .ZN(_03995_));
 OAI21_X1 _29249_ (.A(_02868_),
    .B1(_02831_),
    .B2(_02704_),
    .ZN(_03996_));
 NAND4_X1 _29250_ (.A1(_03994_),
    .A2(_03995_),
    .A3(_03996_),
    .A4(_03630_),
    .ZN(_03997_));
 AND3_X1 _29251_ (.A1(_03233_),
    .A2(_02817_),
    .A3(_02757_),
    .ZN(_03999_));
 AOI21_X1 _29252_ (.A(_02887_),
    .B1(_02839_),
    .B2(_02900_),
    .ZN(_04000_));
 NOR4_X1 _29253_ (.A1(_03993_),
    .A2(_03997_),
    .A3(_03999_),
    .A4(_04000_),
    .ZN(_04001_));
 INV_X1 _29254_ (.A(_03648_),
    .ZN(_04002_));
 OAI21_X1 _29255_ (.A(_02847_),
    .B1(_03248_),
    .B2(_03616_),
    .ZN(_04003_));
 OAI211_X2 _29256_ (.A(_04002_),
    .B(_04003_),
    .C1(_02886_),
    .C2(_03217_),
    .ZN(_04004_));
 AOI211_X4 _29257_ (.A(_03636_),
    .B(_03214_),
    .C1(_02811_),
    .C2(_02800_),
    .ZN(_04005_));
 NAND2_X1 _29258_ (.A1(_02851_),
    .A2(_02719_),
    .ZN(_04006_));
 OAI211_X2 _29259_ (.A(_03296_),
    .B(_04006_),
    .C1(_02779_),
    .C2(_03214_),
    .ZN(_04007_));
 INV_X1 _29260_ (.A(_02761_),
    .ZN(_04008_));
 AOI21_X1 _29261_ (.A(_03214_),
    .B1(_02894_),
    .B2(_04008_),
    .ZN(_04009_));
 NOR4_X1 _29262_ (.A1(_04004_),
    .A2(_04005_),
    .A3(_04007_),
    .A4(_04009_),
    .ZN(_04010_));
 AND4_X1 _29263_ (.A1(_03981_),
    .A2(_03990_),
    .A3(_04001_),
    .A4(_04010_),
    .ZN(_04011_));
 NAND3_X1 _29264_ (.A1(_02702_),
    .A2(_02683_),
    .A3(_02773_),
    .ZN(_04012_));
 NAND4_X1 _29265_ (.A1(_02696_),
    .A2(_03274_),
    .A3(_02718_),
    .A4(_04012_),
    .ZN(_04013_));
 AND4_X1 _29266_ (.A1(_02724_),
    .A2(_03246_),
    .A3(_02859_),
    .A4(_02773_),
    .ZN(_04014_));
 INV_X1 _29267_ (.A(_02701_),
    .ZN(_04015_));
 AOI21_X1 _29268_ (.A(_03622_),
    .B1(_04015_),
    .B2(_04008_),
    .ZN(_04016_));
 NAND2_X1 _29269_ (.A1(_02726_),
    .A2(_02715_),
    .ZN(_04017_));
 NAND2_X1 _29270_ (.A1(_02726_),
    .A2(_02903_),
    .ZN(_04018_));
 OAI211_X2 _29271_ (.A(_04017_),
    .B(_04018_),
    .C1(_03622_),
    .C2(_02738_),
    .ZN(_04020_));
 NOR4_X1 _29272_ (.A1(_04013_),
    .A2(_04014_),
    .A3(_04016_),
    .A4(_04020_),
    .ZN(_04021_));
 OAI21_X1 _29273_ (.A(_02796_),
    .B1(_03253_),
    .B2(_02747_),
    .ZN(_04022_));
 AND4_X1 _29274_ (.A1(_02755_),
    .A2(_02724_),
    .A3(_02709_),
    .A4(_02743_),
    .ZN(_04023_));
 AND4_X1 _29275_ (.A1(_02724_),
    .A2(_02687_),
    .A3(_02690_),
    .A4(_02743_),
    .ZN(_04024_));
 AOI211_X4 _29276_ (.A(_04023_),
    .B(_04024_),
    .C1(_02881_),
    .C2(_02806_),
    .ZN(_04025_));
 OAI21_X1 _29277_ (.A(_02796_),
    .B1(_03230_),
    .B2(_02791_),
    .ZN(_04026_));
 NAND2_X1 _29278_ (.A1(_02806_),
    .A2(_02719_),
    .ZN(_04027_));
 AND4_X1 _29279_ (.A1(_02802_),
    .A2(_04027_),
    .A3(_03596_),
    .A4(_02804_),
    .ZN(_04028_));
 AND4_X1 _29280_ (.A1(_04022_),
    .A2(_04025_),
    .A3(_04026_),
    .A4(_04028_),
    .ZN(_04029_));
 OAI21_X1 _29281_ (.A(_02787_),
    .B1(_02903_),
    .B2(_02749_),
    .ZN(_04030_));
 OAI21_X1 _29282_ (.A(_02787_),
    .B1(_03616_),
    .B2(_02732_),
    .ZN(_04031_));
 OAI21_X1 _29283_ (.A(_03309_),
    .B1(_02903_),
    .B2(_03595_),
    .ZN(_04032_));
 OAI21_X1 _29284_ (.A(_03309_),
    .B1(_03616_),
    .B2(_02791_),
    .ZN(_04033_));
 AND4_X1 _29285_ (.A1(_04030_),
    .A2(_04031_),
    .A3(_04032_),
    .A4(_04033_),
    .ZN(_04034_));
 NAND2_X1 _29286_ (.A1(_03584_),
    .A2(_02863_),
    .ZN(_04035_));
 NAND3_X1 _29287_ (.A1(_02759_),
    .A2(_02862_),
    .A3(_02859_),
    .ZN(_04036_));
 NAND2_X1 _29288_ (.A1(_04035_),
    .A2(_04036_),
    .ZN(_04037_));
 OAI211_X2 _29289_ (.A(_02752_),
    .B(_02753_),
    .C1(_02811_),
    .C2(_02857_),
    .ZN(_04038_));
 OAI21_X1 _29290_ (.A(_04038_),
    .B1(_02770_),
    .B2(_02769_),
    .ZN(_04039_));
 AOI21_X1 _29291_ (.A(_02765_),
    .B1(_02886_),
    .B2(_03269_),
    .ZN(_04041_));
 AOI21_X1 _29292_ (.A(_02769_),
    .B1(_02900_),
    .B2(_02779_),
    .ZN(_04042_));
 NOR4_X1 _29293_ (.A1(_04037_),
    .A2(_04039_),
    .A3(_04041_),
    .A4(_04042_),
    .ZN(_04043_));
 AND4_X1 _29294_ (.A1(_04021_),
    .A2(_04029_),
    .A3(_04034_),
    .A4(_04043_),
    .ZN(_04044_));
 NAND2_X1 _29295_ (.A1(_04011_),
    .A2(_04044_),
    .ZN(_04045_));
 XOR2_X1 _29296_ (.A(_02907_),
    .B(_04045_),
    .Z(_04046_));
 XNOR2_X2 _29297_ (.A(_03972_),
    .B(_04046_),
    .ZN(_04047_));
 XOR2_X1 _29298_ (.A(_03806_),
    .B(_04047_),
    .Z(_04048_));
 XNOR2_X1 _29299_ (.A(_04048_),
    .B(_17233_),
    .ZN(_04049_));
 MUX2_X1 _29300_ (.A(_03724_),
    .B(_04049_),
    .S(_01876_),
    .Z(_00711_));
 XOR2_X1 _29301_ (.A(_17234_),
    .B(_17104_),
    .Z(_04050_));
 XOR2_X2 _29302_ (.A(_02580_),
    .B(_03971_),
    .Z(_04051_));
 AND2_X1 _29303_ (.A1(_01957_),
    .A2(_02113_),
    .ZN(_04052_));
 AND2_X2 _29304_ (.A1(_01920_),
    .A2(_01993_),
    .ZN(_04053_));
 AOI211_X4 _29305_ (.A(_04052_),
    .B(_04053_),
    .C1(_02112_),
    .C2(_01957_),
    .ZN(_04054_));
 AND3_X1 _29306_ (.A1(_02064_),
    .A2(_01916_),
    .A3(_01896_),
    .ZN(_04055_));
 AOI211_X4 _29307_ (.A(_04055_),
    .B(_02059_),
    .C1(_02014_),
    .C2(_02061_),
    .ZN(_04056_));
 OAI21_X1 _29308_ (.A(_01957_),
    .B1(_02015_),
    .B2(_02122_),
    .ZN(_04057_));
 AND4_X4 _29309_ (.A1(_03153_),
    .A2(_04054_),
    .A3(_04056_),
    .A4(_04057_),
    .ZN(_04058_));
 OAI21_X1 _29310_ (.A(_02080_),
    .B1(_01969_),
    .B2(_02077_),
    .ZN(_04059_));
 NAND2_X1 _29311_ (.A1(_01960_),
    .A2(_01905_),
    .ZN(_04060_));
 OAI21_X1 _29312_ (.A(_01960_),
    .B1(_02033_),
    .B2(_02064_),
    .ZN(_04061_));
 OAI21_X1 _29313_ (.A(_01960_),
    .B1(_03154_),
    .B2(_03202_),
    .ZN(_04062_));
 AND4_X2 _29314_ (.A1(_04060_),
    .A2(_04061_),
    .A3(_02088_),
    .A4(_04062_),
    .ZN(_04063_));
 NAND2_X1 _29315_ (.A1(_01938_),
    .A2(_03133_),
    .ZN(_04064_));
 OAI211_X2 _29316_ (.A(_01916_),
    .B(_01924_),
    .C1(_02093_),
    .C2(_02099_),
    .ZN(_04065_));
 AND4_X1 _29317_ (.A1(_04059_),
    .A2(_04063_),
    .A3(_04064_),
    .A4(_04065_),
    .ZN(_04066_));
 INV_X1 _29318_ (.A(_03179_),
    .ZN(_04067_));
 NAND2_X2 _29319_ (.A1(_02069_),
    .A2(_01961_),
    .ZN(_04068_));
 NAND3_X1 _29320_ (.A1(_04067_),
    .A2(_04068_),
    .A3(_03791_),
    .ZN(_04069_));
 AND2_X1 _29321_ (.A1(_02070_),
    .A2(_02061_),
    .ZN(_04070_));
 AND2_X1 _29322_ (.A1(_01935_),
    .A2(_02070_),
    .ZN(_04071_));
 NAND2_X1 _29323_ (.A1(_01923_),
    .A2(_02123_),
    .ZN(_04072_));
 NAND3_X1 _29324_ (.A1(_02123_),
    .A2(_02098_),
    .A3(_01891_),
    .ZN(_04073_));
 NAND4_X1 _29325_ (.A1(_04072_),
    .A2(_03171_),
    .A3(_03557_),
    .A4(_04073_),
    .ZN(_04074_));
 NOR4_X1 _29326_ (.A1(_04069_),
    .A2(_04070_),
    .A3(_04071_),
    .A4(_04074_),
    .ZN(_04075_));
 NAND3_X1 _29327_ (.A1(_01977_),
    .A2(_01985_),
    .A3(_02084_),
    .ZN(_04076_));
 AND2_X1 _29328_ (.A1(_02076_),
    .A2(_01927_),
    .ZN(_04077_));
 AND3_X1 _29329_ (.A1(_01927_),
    .A2(_01944_),
    .A3(_01903_),
    .ZN(_04078_));
 AOI211_X2 _29330_ (.A(_04077_),
    .B(_04078_),
    .C1(_02103_),
    .C2(_01935_),
    .ZN(_04079_));
 OAI211_X2 _29331_ (.A(_02084_),
    .B(_02005_),
    .C1(_01908_),
    .C2(_02099_),
    .ZN(_04081_));
 OAI21_X1 _29332_ (.A(_02084_),
    .B1(_01969_),
    .B2(_02077_),
    .ZN(_04082_));
 AND4_X1 _29333_ (.A1(_04076_),
    .A2(_04079_),
    .A3(_04081_),
    .A4(_04082_),
    .ZN(_04083_));
 NAND4_X1 _29334_ (.A1(_04058_),
    .A2(_04066_),
    .A3(_04075_),
    .A4(_04083_),
    .ZN(_04084_));
 INV_X1 _29335_ (.A(_01975_),
    .ZN(_04085_));
 AOI211_X2 _29336_ (.A(_03127_),
    .B(_03730_),
    .C1(_01995_),
    .C2(_01966_),
    .ZN(_04086_));
 OAI21_X1 _29337_ (.A(_03130_),
    .B1(_01993_),
    .B2(_01995_),
    .ZN(_04087_));
 OAI21_X1 _29338_ (.A(_03130_),
    .B1(_03134_),
    .B2(_03154_),
    .ZN(_04088_));
 AND4_X1 _29339_ (.A1(_04085_),
    .A2(_04086_),
    .A3(_04087_),
    .A4(_04088_),
    .ZN(_04089_));
 INV_X1 _29340_ (.A(_02051_),
    .ZN(_04090_));
 OAI21_X1 _29341_ (.A(_01981_),
    .B1(_01923_),
    .B2(_02081_),
    .ZN(_04091_));
 OAI211_X2 _29342_ (.A(_03195_),
    .B(_16847_),
    .C1(_16846_),
    .C2(_01944_),
    .ZN(_04092_));
 OAI21_X1 _29343_ (.A(_01981_),
    .B1(_01999_),
    .B2(_02026_),
    .ZN(_04093_));
 AND4_X1 _29344_ (.A1(_04090_),
    .A2(_04091_),
    .A3(_04092_),
    .A4(_04093_),
    .ZN(_04094_));
 AND2_X2 _29345_ (.A1(_01991_),
    .A2(_02063_),
    .ZN(_04095_));
 INV_X2 _29346_ (.A(_04095_),
    .ZN(_04096_));
 OAI21_X1 _29347_ (.A(_01992_),
    .B1(_01995_),
    .B2(_02113_),
    .ZN(_04097_));
 OAI211_X2 _29348_ (.A(_01992_),
    .B(_02098_),
    .C1(_03161_),
    .C2(_02017_),
    .ZN(_04098_));
 NAND4_X1 _29349_ (.A1(_04096_),
    .A2(_03757_),
    .A3(_04097_),
    .A4(_04098_),
    .ZN(_04099_));
 AND2_X1 _29350_ (.A1(_02009_),
    .A2(_02113_),
    .ZN(_04100_));
 AND2_X1 _29351_ (.A1(_03176_),
    .A2(_02010_),
    .ZN(_04101_));
 NOR4_X1 _29352_ (.A1(_04099_),
    .A2(_04100_),
    .A3(_04101_),
    .A4(_03530_),
    .ZN(_04102_));
 AOI22_X1 _29353_ (.A1(_03136_),
    .A2(_01985_),
    .B1(_02122_),
    .B2(_02078_),
    .ZN(_04103_));
 OAI21_X1 _29354_ (.A(_02078_),
    .B1(_02064_),
    .B2(_02061_),
    .ZN(_04104_));
 OAI21_X1 _29355_ (.A(_01898_),
    .B1(_01892_),
    .B2(_02122_),
    .ZN(_04105_));
 AND4_X1 _29356_ (.A1(_03120_),
    .A2(_04103_),
    .A3(_04104_),
    .A4(_04105_),
    .ZN(_04106_));
 NAND4_X1 _29357_ (.A1(_04089_),
    .A2(_04094_),
    .A3(_04102_),
    .A4(_04106_),
    .ZN(_04107_));
 NOR2_X4 _29358_ (.A1(_04084_),
    .A2(_04107_),
    .ZN(_04108_));
 XNOR2_X1 _29359_ (.A(_04051_),
    .B(_04108_),
    .ZN(_04109_));
 NAND2_X1 _29360_ (.A1(_02264_),
    .A2(_02241_),
    .ZN(_04110_));
 AND3_X1 _29361_ (.A1(_02335_),
    .A2(_02324_),
    .A3(_02223_),
    .ZN(_04111_));
 AOI211_X2 _29362_ (.A(_03855_),
    .B(_04111_),
    .C1(_02156_),
    .C2(_02225_),
    .ZN(_04112_));
 NAND2_X1 _29363_ (.A1(_02226_),
    .A2(_02297_),
    .ZN(_04113_));
 NAND4_X1 _29364_ (.A1(_03032_),
    .A2(_02237_),
    .A3(_02169_),
    .A4(_02252_),
    .ZN(_04114_));
 AND4_X1 _29365_ (.A1(_03853_),
    .A2(_04112_),
    .A3(_04113_),
    .A4(_04114_),
    .ZN(_04115_));
 NAND3_X1 _29366_ (.A1(_02241_),
    .A2(_02266_),
    .A3(_02220_),
    .ZN(_04116_));
 OAI21_X1 _29367_ (.A(_02241_),
    .B1(_03083_),
    .B2(_02221_),
    .ZN(_04117_));
 AND4_X1 _29368_ (.A1(_04110_),
    .A2(_04115_),
    .A3(_04116_),
    .A4(_04117_),
    .ZN(_04118_));
 NAND2_X1 _29369_ (.A1(_03371_),
    .A2(_02302_),
    .ZN(_04119_));
 NAND2_X1 _29370_ (.A1(_02302_),
    .A2(_02292_),
    .ZN(_04120_));
 NAND2_X1 _29371_ (.A1(_02302_),
    .A2(_03096_),
    .ZN(_04122_));
 OAI21_X1 _29372_ (.A(_02302_),
    .B1(_02156_),
    .B2(_02276_),
    .ZN(_04123_));
 NAND4_X1 _29373_ (.A1(_04119_),
    .A2(_04120_),
    .A3(_04122_),
    .A4(_04123_),
    .ZN(_04124_));
 AND2_X1 _29374_ (.A1(_02313_),
    .A2(_02205_),
    .ZN(_04125_));
 AND2_X1 _29375_ (.A1(_02313_),
    .A2(_03037_),
    .ZN(_04126_));
 OR2_X1 _29376_ (.A1(_04125_),
    .A2(_04126_),
    .ZN(_04127_));
 NAND4_X1 _29377_ (.A1(_02279_),
    .A2(_03055_),
    .A3(_02191_),
    .A4(_02268_),
    .ZN(_04128_));
 OAI21_X1 _29378_ (.A(_04128_),
    .B1(_03075_),
    .B2(_03819_),
    .ZN(_04129_));
 NAND2_X1 _29379_ (.A1(_02313_),
    .A2(_02294_),
    .ZN(_04130_));
 NAND4_X1 _29380_ (.A1(_02279_),
    .A2(_02211_),
    .A3(_02220_),
    .A4(_02268_),
    .ZN(_04131_));
 INV_X1 _29381_ (.A(_02185_),
    .ZN(_04133_));
 OAI211_X2 _29382_ (.A(_04130_),
    .B(_04131_),
    .C1(_03075_),
    .C2(_04133_),
    .ZN(_04134_));
 NOR4_X1 _29383_ (.A1(_04124_),
    .A2(_04127_),
    .A3(_04129_),
    .A4(_04134_),
    .ZN(_04135_));
 AND2_X1 _29384_ (.A1(_02291_),
    .A2(_02141_),
    .ZN(_04136_));
 INV_X1 _29385_ (.A(_04136_),
    .ZN(_04137_));
 AND3_X1 _29386_ (.A1(_04137_),
    .A2(_02295_),
    .A3(_02296_),
    .ZN(_04138_));
 INV_X1 _29387_ (.A(_03096_),
    .ZN(_04139_));
 OAI21_X1 _29388_ (.A(_02283_),
    .B1(_02284_),
    .B2(_04139_),
    .ZN(_04140_));
 AOI21_X1 _29389_ (.A(_04140_),
    .B1(_02275_),
    .B2(_02306_),
    .ZN(_04141_));
 OAI21_X1 _29390_ (.A(_02291_),
    .B1(_02156_),
    .B2(_02209_),
    .ZN(_04142_));
 AND4_X1 _29391_ (.A1(_03068_),
    .A2(_04138_),
    .A3(_04141_),
    .A4(_04142_),
    .ZN(_04144_));
 OAI211_X2 _29392_ (.A(_02262_),
    .B(_02266_),
    .C1(_03055_),
    .C2(_02212_),
    .ZN(_04145_));
 AND3_X1 _29393_ (.A1(_02250_),
    .A2(_02179_),
    .A3(_02252_),
    .ZN(_04146_));
 AND3_X1 _29394_ (.A1(_02309_),
    .A2(_02167_),
    .A3(_02246_),
    .ZN(_04147_));
 AOI211_X4 _29395_ (.A(_04146_),
    .B(_04147_),
    .C1(_02276_),
    .C2(_02246_),
    .ZN(_04148_));
 OAI21_X1 _29396_ (.A(_02262_),
    .B1(_02335_),
    .B2(_02251_),
    .ZN(_04149_));
 OAI211_X2 _29397_ (.A(_02247_),
    .B(_02170_),
    .C1(_02211_),
    .C2(_02266_),
    .ZN(_04150_));
 AND4_X1 _29398_ (.A1(_04145_),
    .A2(_04148_),
    .A3(_04149_),
    .A4(_04150_),
    .ZN(_04151_));
 NAND4_X2 _29399_ (.A1(_04118_),
    .A2(_04135_),
    .A3(_04144_),
    .A4(_04151_),
    .ZN(_04152_));
 AOI21_X1 _29400_ (.A(_03094_),
    .B1(_03357_),
    .B2(_02154_),
    .ZN(_04153_));
 AOI21_X1 _29401_ (.A(_04153_),
    .B1(_02149_),
    .B2(_03097_),
    .ZN(_04155_));
 AOI221_X1 _29402_ (.A(_03823_),
    .B1(_02334_),
    .B2(_02305_),
    .C1(_02350_),
    .C2(_03111_),
    .ZN(_04156_));
 AND4_X1 _29403_ (.A1(_02333_),
    .A2(_04155_),
    .A3(_02336_),
    .A4(_04156_),
    .ZN(_04157_));
 OAI21_X1 _29404_ (.A(_02202_),
    .B1(_02276_),
    .B2(_02251_),
    .ZN(_04158_));
 AND3_X1 _29405_ (.A1(_04158_),
    .A2(_02203_),
    .A3(_03835_),
    .ZN(_04159_));
 NAND2_X1 _29406_ (.A1(_02206_),
    .A2(_02182_),
    .ZN(_04160_));
 OAI21_X1 _29407_ (.A(_02182_),
    .B1(_02317_),
    .B2(_02230_),
    .ZN(_04161_));
 AND4_X1 _29408_ (.A1(_02195_),
    .A2(_04159_),
    .A3(_04160_),
    .A4(_04161_),
    .ZN(_04162_));
 NAND4_X1 _29409_ (.A1(_03032_),
    .A2(_02139_),
    .A3(_02243_),
    .A4(_02193_),
    .ZN(_04163_));
 OAI211_X2 _29410_ (.A(_03356_),
    .B(_04163_),
    .C1(_03034_),
    .C2(_03089_),
    .ZN(_04164_));
 NAND4_X1 _29411_ (.A1(_02266_),
    .A2(_02350_),
    .A3(_02193_),
    .A4(_02280_),
    .ZN(_04166_));
 OAI21_X1 _29412_ (.A(_04166_),
    .B1(_02166_),
    .B2(_02287_),
    .ZN(_04167_));
 NAND3_X1 _29413_ (.A1(_03096_),
    .A2(_02324_),
    .A3(_02132_),
    .ZN(_04168_));
 NAND3_X1 _29414_ (.A1(_02147_),
    .A2(_02324_),
    .A3(_02132_),
    .ZN(_04169_));
 OAI211_X2 _29415_ (.A(_04168_),
    .B(_04169_),
    .C1(_03034_),
    .C2(_02287_),
    .ZN(_04170_));
 NOR4_X1 _29416_ (.A1(_04164_),
    .A2(_03366_),
    .A3(_04167_),
    .A4(_04170_),
    .ZN(_04171_));
 OAI21_X1 _29417_ (.A(_02328_),
    .B1(_03096_),
    .B2(_02306_),
    .ZN(_04172_));
 OAI21_X1 _29418_ (.A(_02353_),
    .B1(_02314_),
    .B2(_02209_),
    .ZN(_04173_));
 OAI21_X1 _29419_ (.A(_02328_),
    .B1(_03083_),
    .B2(_02209_),
    .ZN(_04174_));
 AND4_X1 _29420_ (.A1(_03105_),
    .A2(_04172_),
    .A3(_04173_),
    .A4(_04174_),
    .ZN(_04175_));
 NAND4_X2 _29421_ (.A1(_04157_),
    .A2(_04162_),
    .A3(_04171_),
    .A4(_04175_),
    .ZN(_04177_));
 NOR2_X4 _29422_ (.A1(_04152_),
    .A2(_04177_),
    .ZN(_04178_));
 AND2_X1 _29423_ (.A1(_02556_),
    .A2(_02549_),
    .ZN(_04179_));
 AND2_X1 _29424_ (.A1(_02555_),
    .A2(_02454_),
    .ZN(_04180_));
 AOI211_X2 _29425_ (.A(_04179_),
    .B(_04180_),
    .C1(_02481_),
    .C2(_02556_),
    .ZN(_04181_));
 OAI21_X1 _29426_ (.A(_02557_),
    .B1(_02538_),
    .B2(_02454_),
    .ZN(_04182_));
 NAND3_X1 _29427_ (.A1(_02368_),
    .A2(_02557_),
    .A3(_02371_),
    .ZN(_04183_));
 AND3_X1 _29428_ (.A1(_04182_),
    .A2(_03951_),
    .A3(_04183_),
    .ZN(_04184_));
 OAI211_X2 _29429_ (.A(_04181_),
    .B(_04184_),
    .C1(_02606_),
    .C2(_02608_),
    .ZN(_04185_));
 NAND2_X1 _29430_ (.A1(_02435_),
    .A2(_02441_),
    .ZN(_04186_));
 NAND3_X1 _29431_ (.A1(_02435_),
    .A2(_02506_),
    .A3(_02581_),
    .ZN(_04188_));
 AND4_X1 _29432_ (.A1(_03444_),
    .A2(_03443_),
    .A3(_04186_),
    .A4(_04188_),
    .ZN(_04189_));
 NAND2_X1 _29433_ (.A1(_02662_),
    .A2(_02539_),
    .ZN(_04190_));
 OAI21_X1 _29434_ (.A(_02662_),
    .B1(_02368_),
    .B2(_03437_),
    .ZN(_04191_));
 OAI21_X1 _29435_ (.A(_02662_),
    .B1(_02454_),
    .B2(_02441_),
    .ZN(_04192_));
 NAND4_X1 _29436_ (.A1(_04189_),
    .A2(_04190_),
    .A3(_04191_),
    .A4(_04192_),
    .ZN(_04193_));
 OAI21_X1 _29437_ (.A(_02525_),
    .B1(_02560_),
    .B2(_02490_),
    .ZN(_04194_));
 OAI21_X1 _29438_ (.A(_03450_),
    .B1(_02439_),
    .B2(_02658_),
    .ZN(_04195_));
 OAI21_X1 _29439_ (.A(_03450_),
    .B1(_02434_),
    .B2(_02545_),
    .ZN(_04196_));
 NAND2_X1 _29440_ (.A1(_02485_),
    .A2(_02525_),
    .ZN(_04197_));
 NAND4_X1 _29441_ (.A1(_04194_),
    .A2(_04195_),
    .A3(_04196_),
    .A4(_04197_),
    .ZN(_04199_));
 AND4_X1 _29442_ (.A1(_02388_),
    .A2(_02553_),
    .A3(_02490_),
    .A4(_02944_),
    .ZN(_04200_));
 AND4_X1 _29443_ (.A1(_02490_),
    .A2(_02402_),
    .A3(_02553_),
    .A4(_02944_),
    .ZN(_04201_));
 NOR3_X1 _29444_ (.A1(_03941_),
    .A2(_04200_),
    .A3(_04201_),
    .ZN(_04202_));
 OAI21_X1 _29445_ (.A(_02417_),
    .B1(_02607_),
    .B2(_02597_),
    .ZN(_04203_));
 OAI21_X1 _29446_ (.A(_02380_),
    .B1(_04203_),
    .B2(_02505_),
    .ZN(_04204_));
 AND2_X1 _29447_ (.A1(_02600_),
    .A2(_02945_),
    .ZN(_04205_));
 NAND2_X1 _29448_ (.A1(_02380_),
    .A2(_02399_),
    .ZN(_04206_));
 NAND4_X1 _29449_ (.A1(_04202_),
    .A2(_04204_),
    .A3(_04205_),
    .A4(_04206_),
    .ZN(_04207_));
 NOR4_X1 _29450_ (.A1(_04185_),
    .A2(_04193_),
    .A3(_04199_),
    .A4(_04207_),
    .ZN(_04208_));
 AOI21_X1 _29451_ (.A(_02469_),
    .B1(_02631_),
    .B2(_03478_),
    .ZN(_04210_));
 AND2_X1 _29452_ (.A1(_02465_),
    .A2(_02539_),
    .ZN(_04211_));
 AND4_X1 _29453_ (.A1(_02672_),
    .A2(_02602_),
    .A3(_02607_),
    .A4(_02429_),
    .ZN(_04212_));
 NOR4_X4 _29454_ (.A1(_04210_),
    .A2(_03897_),
    .A3(_04211_),
    .A4(_04212_),
    .ZN(_04213_));
 AND4_X1 _29455_ (.A1(_02534_),
    .A2(_02621_),
    .A3(_02383_),
    .A4(_02593_),
    .ZN(_04214_));
 AND2_X4 _29456_ (.A1(_02462_),
    .A2(_02390_),
    .ZN(_04215_));
 AOI211_X4 _29457_ (.A(_04214_),
    .B(_04215_),
    .C1(_03003_),
    .C2(_02527_),
    .ZN(_04216_));
 OAI21_X1 _29458_ (.A(_03003_),
    .B1(_02500_),
    .B2(_02434_),
    .ZN(_04217_));
 OAI21_X1 _29459_ (.A(_03003_),
    .B1(_03437_),
    .B2(_02445_),
    .ZN(_04218_));
 NAND4_X2 _29460_ (.A1(_04213_),
    .A2(_04216_),
    .A3(_04217_),
    .A4(_04218_),
    .ZN(_04219_));
 AND2_X4 _29461_ (.A1(_02451_),
    .A2(_02416_),
    .ZN(_04221_));
 AOI211_X2 _29462_ (.A(_04221_),
    .B(_03906_),
    .C1(_02481_),
    .C2(_02516_),
    .ZN(_04222_));
 AND2_X1 _29463_ (.A1(_02650_),
    .A2(_02448_),
    .ZN(_04223_));
 INV_X1 _29464_ (.A(_04223_),
    .ZN(_04224_));
 OR2_X1 _29465_ (.A1(_02979_),
    .A2(_02598_),
    .ZN(_04225_));
 NAND3_X1 _29466_ (.A1(_02449_),
    .A2(_02621_),
    .A3(_02581_),
    .ZN(_04226_));
 AND4_X2 _29467_ (.A1(_03482_),
    .A2(_04224_),
    .A3(_04225_),
    .A4(_04226_),
    .ZN(_04227_));
 OAI21_X1 _29468_ (.A(_02516_),
    .B1(_02477_),
    .B2(_02425_),
    .ZN(_04228_));
 NAND3_X1 _29469_ (.A1(_02560_),
    .A2(_03431_),
    .A3(_02446_),
    .ZN(_04229_));
 NAND4_X1 _29470_ (.A1(_04222_),
    .A2(_04227_),
    .A3(_04228_),
    .A4(_04229_),
    .ZN(_04230_));
 AND2_X1 _29471_ (.A1(_02532_),
    .A2(_02538_),
    .ZN(_04232_));
 INV_X1 _29472_ (.A(_04232_),
    .ZN(_04233_));
 AND3_X1 _29473_ (.A1(_04233_),
    .A2(_02655_),
    .A3(_02584_),
    .ZN(_04234_));
 OAI21_X1 _29474_ (.A(_02548_),
    .B1(_02987_),
    .B2(_02416_),
    .ZN(_04235_));
 OAI21_X1 _29475_ (.A(_02532_),
    .B1(_02505_),
    .B2(_02477_),
    .ZN(_04236_));
 NAND4_X1 _29476_ (.A1(_04234_),
    .A2(_02992_),
    .A3(_04235_),
    .A4(_04236_),
    .ZN(_04237_));
 OAI21_X1 _29477_ (.A(_02614_),
    .B1(_02647_),
    .B2(_02490_),
    .ZN(_04238_));
 OAI21_X1 _29478_ (.A(_02522_),
    .B1(_02560_),
    .B2(_02466_),
    .ZN(_04239_));
 OAI211_X2 _29479_ (.A(_02522_),
    .B(_02581_),
    .C1(_02664_),
    .C2(_02535_),
    .ZN(_04240_));
 AND2_X1 _29480_ (.A1(_04239_),
    .A2(_04240_),
    .ZN(_04241_));
 OAI211_X2 _29481_ (.A(_02614_),
    .B(_02371_),
    .C1(_02383_),
    .C2(_02581_),
    .ZN(_04243_));
 NAND3_X1 _29482_ (.A1(_04238_),
    .A2(_04241_),
    .A3(_04243_),
    .ZN(_04244_));
 NOR4_X2 _29483_ (.A1(_04219_),
    .A2(_04230_),
    .A3(_04237_),
    .A4(_04244_),
    .ZN(_04245_));
 NAND2_X1 _29484_ (.A1(_04208_),
    .A2(_04245_),
    .ZN(_04246_));
 XNOR2_X1 _29485_ (.A(_04178_),
    .B(_04246_),
    .ZN(_04247_));
 AOI21_X1 _29486_ (.A(_03634_),
    .B1(_02764_),
    .B2(_03294_),
    .ZN(_04248_));
 AND3_X1 _29487_ (.A1(_02818_),
    .A2(_02858_),
    .A3(_02862_),
    .ZN(_04249_));
 NOR4_X1 _29488_ (.A1(_04248_),
    .A2(_02819_),
    .A3(_03286_),
    .A4(_04249_),
    .ZN(_04250_));
 INV_X1 _29489_ (.A(_03638_),
    .ZN(_04251_));
 OAI21_X1 _29490_ (.A(_02829_),
    .B1(_02775_),
    .B2(_02736_),
    .ZN(_04252_));
 OAI211_X2 _29491_ (.A(_02829_),
    .B(_02728_),
    .C1(_02712_),
    .C2(_02862_),
    .ZN(_04254_));
 AND3_X1 _29492_ (.A1(_04251_),
    .A2(_04252_),
    .A3(_04254_),
    .ZN(_04255_));
 OAI211_X2 _29493_ (.A(_02835_),
    .B(_02859_),
    .C1(_02811_),
    .C2(_02857_),
    .ZN(_04256_));
 OAI21_X1 _29494_ (.A(_02835_),
    .B1(_02831_),
    .B2(_02732_),
    .ZN(_04257_));
 AND4_X1 _29495_ (.A1(_04250_),
    .A2(_04255_),
    .A3(_04256_),
    .A4(_04257_),
    .ZN(_04258_));
 OAI21_X1 _29496_ (.A(_03279_),
    .B1(_02870_),
    .B2(_02704_),
    .ZN(_04259_));
 AND2_X1 _29497_ (.A1(_02867_),
    .A2(_02746_),
    .ZN(_04260_));
 INV_X1 _29498_ (.A(_04260_),
    .ZN(_04261_));
 INV_X1 _29499_ (.A(_03279_),
    .ZN(_04262_));
 OAI221_X1 _29500_ (.A(_04259_),
    .B1(_04261_),
    .B2(_02856_),
    .C1(_02764_),
    .C2(_04262_),
    .ZN(_04263_));
 OR4_X4 _29501_ (.A1(_02882_),
    .A2(_03643_),
    .A3(_02879_),
    .A4(_03276_),
    .ZN(_04265_));
 AND2_X1 _29502_ (.A1(_02736_),
    .A2(_02883_),
    .ZN(_04266_));
 NAND2_X1 _29503_ (.A1(_02883_),
    .A2(_02747_),
    .ZN(_04267_));
 OAI21_X1 _29504_ (.A(_04267_),
    .B1(_02900_),
    .B2(_02887_),
    .ZN(_04268_));
 NOR4_X4 _29505_ (.A1(_04263_),
    .A2(_04265_),
    .A3(_04266_),
    .A4(_04268_),
    .ZN(_04269_));
 NOR2_X1 _29506_ (.A1(_02783_),
    .A2(_03268_),
    .ZN(_04270_));
 AND2_X1 _29507_ (.A1(_02891_),
    .A2(_03273_),
    .ZN(_04271_));
 NOR4_X1 _29508_ (.A1(_04270_),
    .A2(_03986_),
    .A3(_03661_),
    .A4(_04271_),
    .ZN(_04272_));
 NAND2_X1 _29509_ (.A1(_02898_),
    .A2(_02736_),
    .ZN(_04273_));
 OAI21_X1 _29510_ (.A(_02898_),
    .B1(_03248_),
    .B2(_02790_),
    .ZN(_04274_));
 AND4_X1 _29511_ (.A1(_03983_),
    .A2(_04272_),
    .A3(_04273_),
    .A4(_04274_),
    .ZN(_04276_));
 AND2_X1 _29512_ (.A1(_02846_),
    .A2(_02736_),
    .ZN(_04277_));
 AND2_X1 _29513_ (.A1(_02846_),
    .A2(_02710_),
    .ZN(_04278_));
 NOR2_X4 _29514_ (.A1(_04277_),
    .A2(_04278_),
    .ZN(_04279_));
 OAI21_X1 _29515_ (.A(_02847_),
    .B1(_03616_),
    .B2(_02767_),
    .ZN(_04280_));
 INV_X1 _29516_ (.A(_03254_),
    .ZN(_04281_));
 OAI211_X2 _29517_ (.A(_04279_),
    .B(_04280_),
    .C1(_04281_),
    .C2(_03217_),
    .ZN(_04282_));
 OAI211_X2 _29518_ (.A(_02851_),
    .B(_02812_),
    .C1(_02856_),
    .C2(_02800_),
    .ZN(_04283_));
 OAI21_X1 _29519_ (.A(_04283_),
    .B1(_03610_),
    .B2(_03214_),
    .ZN(_04284_));
 AOI211_X4 _29520_ (.A(_03247_),
    .B(_03214_),
    .C1(_02856_),
    .C2(_02857_),
    .ZN(_04285_));
 AND4_X1 _29521_ (.A1(_02845_),
    .A2(_03246_),
    .A3(_02753_),
    .A4(_02683_),
    .ZN(_04287_));
 NOR4_X1 _29522_ (.A1(_04282_),
    .A2(_04284_),
    .A3(_04285_),
    .A4(_04287_),
    .ZN(_04288_));
 NAND4_X2 _29523_ (.A1(_04258_),
    .A2(_04269_),
    .A3(_04276_),
    .A4(_04288_),
    .ZN(_04289_));
 OAI21_X1 _29524_ (.A(_02752_),
    .B1(_03295_),
    .B2(_02719_),
    .ZN(_04290_));
 AND2_X1 _29525_ (.A1(_02830_),
    .A2(_02758_),
    .ZN(_04291_));
 AOI221_X1 _29526_ (.A(_04291_),
    .B1(_02870_),
    .B2(_02759_),
    .C1(_02862_),
    .C2(_03584_),
    .ZN(_04292_));
 OAI21_X1 _29527_ (.A(_03222_),
    .B1(_03253_),
    .B2(_02781_),
    .ZN(_04293_));
 AOI22_X1 _29528_ (.A1(_02754_),
    .A2(_03246_),
    .B1(_02831_),
    .B2(_02752_),
    .ZN(_04294_));
 AND4_X1 _29529_ (.A1(_04290_),
    .A2(_04292_),
    .A3(_04293_),
    .A4(_04294_),
    .ZN(_04295_));
 NAND2_X1 _29530_ (.A1(_02727_),
    .A2(_03271_),
    .ZN(_04296_));
 OAI21_X1 _29531_ (.A(_02697_),
    .B1(_02778_),
    .B2(_02775_),
    .ZN(_04298_));
 NAND4_X1 _29532_ (.A1(_02773_),
    .A2(_02698_),
    .A3(_02690_),
    .A4(_02683_),
    .ZN(_04299_));
 AND4_X2 _29533_ (.A1(_02718_),
    .A2(_04298_),
    .A3(_04012_),
    .A4(_04299_),
    .ZN(_04300_));
 OAI21_X1 _29534_ (.A(_02727_),
    .B1(_03259_),
    .B2(_02903_),
    .ZN(_04301_));
 OAI21_X1 _29535_ (.A(_02727_),
    .B1(_02702_),
    .B2(_02732_),
    .ZN(_04302_));
 AND4_X1 _29536_ (.A1(_04296_),
    .A2(_04300_),
    .A3(_04301_),
    .A4(_04302_),
    .ZN(_04303_));
 NAND2_X1 _29537_ (.A1(_03309_),
    .A2(_02858_),
    .ZN(_04304_));
 OAI211_X2 _29538_ (.A(_02786_),
    .B(_02728_),
    .C1(_02698_),
    .C2(_02800_),
    .ZN(_04305_));
 OAI21_X1 _29539_ (.A(_02786_),
    .B1(_02731_),
    .B2(_02797_),
    .ZN(_04306_));
 AND3_X1 _29540_ (.A1(_04305_),
    .A2(_03609_),
    .A3(_04306_),
    .ZN(_04307_));
 OAI21_X1 _29541_ (.A(_03309_),
    .B1(_02790_),
    .B2(_02881_),
    .ZN(_04309_));
 OAI21_X1 _29542_ (.A(_03309_),
    .B1(_03273_),
    .B2(_03595_),
    .ZN(_04310_));
 AND4_X1 _29543_ (.A1(_04304_),
    .A2(_04307_),
    .A3(_04309_),
    .A4(_04310_),
    .ZN(_04311_));
 NAND2_X4 _29544_ (.A1(_02831_),
    .A2(_02795_),
    .ZN(_04312_));
 OAI21_X1 _29545_ (.A(_02806_),
    .B1(_02715_),
    .B2(_03273_),
    .ZN(_04313_));
 OAI21_X1 _29546_ (.A(_02795_),
    .B1(_02736_),
    .B2(_02710_),
    .ZN(_04314_));
 NAND2_X1 _29547_ (.A1(_02702_),
    .A2(_02806_),
    .ZN(_04315_));
 AND4_X1 _29548_ (.A1(_04312_),
    .A2(_04313_),
    .A3(_04314_),
    .A4(_04315_),
    .ZN(_04316_));
 NAND4_X1 _29549_ (.A1(_04295_),
    .A2(_04303_),
    .A3(_04311_),
    .A4(_04316_),
    .ZN(_04317_));
 NOR2_X4 _29550_ (.A1(_04289_),
    .A2(_04317_),
    .ZN(_04318_));
 XOR2_X2 _29551_ (.A(_04318_),
    .B(_02907_),
    .Z(_04320_));
 XNOR2_X2 _29552_ (.A(_04247_),
    .B(_04320_),
    .ZN(_04321_));
 XNOR2_X1 _29553_ (.A(_04109_),
    .B(_04321_),
    .ZN(_04322_));
 XOR2_X1 _29554_ (.A(_04322_),
    .B(_17234_),
    .Z(_04323_));
 MUX2_X1 _29555_ (.A(_04050_),
    .B(_04323_),
    .S(_01876_),
    .Z(_00712_));
 XOR2_X1 _29556_ (.A(_17235_),
    .B(_17105_),
    .Z(_04324_));
 NAND2_X1 _29557_ (.A1(_02372_),
    .A2(_02380_),
    .ZN(_04325_));
 OAI21_X1 _29558_ (.A(_02610_),
    .B1(_02427_),
    .B2(_02368_),
    .ZN(_04326_));
 NAND2_X1 _29559_ (.A1(_02610_),
    .A2(_02416_),
    .ZN(_04327_));
 OAI21_X1 _29560_ (.A(_02380_),
    .B1(_02527_),
    .B2(_02419_),
    .ZN(_04328_));
 AND4_X1 _29561_ (.A1(_04325_),
    .A2(_04326_),
    .A3(_04327_),
    .A4(_04328_),
    .ZN(_04330_));
 AND4_X1 _29562_ (.A1(_02398_),
    .A2(_02437_),
    .A3(_02378_),
    .A4(_02429_),
    .ZN(_04331_));
 AOI211_X4 _29563_ (.A(_04331_),
    .B(_04180_),
    .C1(_02556_),
    .C2(_02441_),
    .ZN(_04332_));
 OAI21_X1 _29564_ (.A(_02556_),
    .B1(_02505_),
    .B2(_03437_),
    .ZN(_04333_));
 NAND2_X1 _29565_ (.A1(_04332_),
    .A2(_04333_),
    .ZN(_04334_));
 OAI211_X2 _29566_ (.A(_02557_),
    .B(_02499_),
    .C1(_02388_),
    .C2(_02506_),
    .ZN(_04335_));
 OAI211_X2 _29567_ (.A(_04335_),
    .B(_02478_),
    .C1(_03478_),
    .C2(_03465_),
    .ZN(_04336_));
 NOR4_X1 _29568_ (.A1(_04334_),
    .A2(_02482_),
    .A3(_02603_),
    .A4(_04336_),
    .ZN(_04337_));
 OAI21_X1 _29569_ (.A(_02435_),
    .B1(_02999_),
    .B2(_03893_),
    .ZN(_04338_));
 OAI21_X1 _29570_ (.A(_02413_),
    .B1(_02441_),
    .B2(_02619_),
    .ZN(_04339_));
 NAND3_X1 _29571_ (.A1(_02435_),
    .A2(_02509_),
    .A3(_02371_),
    .ZN(_04341_));
 AND3_X1 _29572_ (.A1(_04338_),
    .A2(_04339_),
    .A3(_04341_),
    .ZN(_04342_));
 OAI211_X2 _29573_ (.A(_03431_),
    .B(_02472_),
    .C1(_02441_),
    .C2(_02619_),
    .ZN(_04343_));
 OAI21_X1 _29574_ (.A(_02662_),
    .B1(_02572_),
    .B2(_02434_),
    .ZN(_04344_));
 AND4_X1 _29575_ (.A1(_04190_),
    .A2(_04342_),
    .A3(_04343_),
    .A4(_04344_),
    .ZN(_04345_));
 OAI21_X1 _29576_ (.A(_03450_),
    .B1(_02572_),
    .B2(_02477_),
    .ZN(_04346_));
 NAND2_X1 _29577_ (.A1(_03450_),
    .A2(_02441_),
    .ZN(_04347_));
 NAND4_X1 _29578_ (.A1(_02581_),
    .A2(_02429_),
    .A3(_02621_),
    .A4(_02472_),
    .ZN(_04348_));
 NAND3_X1 _29579_ (.A1(_04346_),
    .A2(_04347_),
    .A3(_04348_),
    .ZN(_04349_));
 OAI21_X1 _29580_ (.A(_02969_),
    .B1(_02484_),
    .B2(_02642_),
    .ZN(_04350_));
 AOI21_X1 _29581_ (.A(_02642_),
    .B1(_03460_),
    .B2(_03464_),
    .ZN(_04352_));
 NOR4_X1 _29582_ (.A1(_04349_),
    .A2(_04350_),
    .A3(_04352_),
    .A4(_02645_),
    .ZN(_04353_));
 AND4_X1 _29583_ (.A1(_04330_),
    .A2(_04337_),
    .A3(_04345_),
    .A4(_04353_),
    .ZN(_04354_));
 OAI22_X1 _29584_ (.A1(_03476_),
    .A2(_02535_),
    .B1(_02453_),
    .B2(_02544_),
    .ZN(_04355_));
 NOR2_X1 _29585_ (.A1(_02635_),
    .A2(_02453_),
    .ZN(_04356_));
 NOR4_X1 _29586_ (.A1(_02517_),
    .A2(_04355_),
    .A3(_04356_),
    .A4(_04221_),
    .ZN(_04357_));
 OAI221_X1 _29587_ (.A(_02449_),
    .B1(_02388_),
    .B2(_02506_),
    .C1(_02490_),
    .C2(_02991_),
    .ZN(_04358_));
 AND4_X1 _29588_ (.A1(_03482_),
    .A2(_04357_),
    .A3(_02977_),
    .A4(_04358_),
    .ZN(_04359_));
 NAND3_X1 _29589_ (.A1(_02522_),
    .A2(_02598_),
    .A3(_02383_),
    .ZN(_04360_));
 NAND2_X1 _29590_ (.A1(_02522_),
    .A2(_03437_),
    .ZN(_04361_));
 NAND4_X1 _29591_ (.A1(_02983_),
    .A2(_04360_),
    .A3(_02649_),
    .A4(_04361_),
    .ZN(_04363_));
 AOI21_X1 _29592_ (.A(_02495_),
    .B1(_03464_),
    .B2(_02638_),
    .ZN(_04364_));
 AND2_X1 _29593_ (.A1(_02976_),
    .A2(_02614_),
    .ZN(_04365_));
 NOR4_X1 _29594_ (.A1(_04363_),
    .A2(_04364_),
    .A3(_04365_),
    .A4(_03500_),
    .ZN(_04366_));
 OAI21_X1 _29595_ (.A(_02548_),
    .B1(_02454_),
    .B2(_02439_),
    .ZN(_04367_));
 AND3_X1 _29596_ (.A1(_04367_),
    .A2(_02674_),
    .A3(_02673_),
    .ZN(_04368_));
 OAI211_X2 _29597_ (.A(_03007_),
    .B(_03008_),
    .C1(_02469_),
    .C2(_03480_),
    .ZN(_04369_));
 AOI211_X2 _29598_ (.A(_03897_),
    .B(_04369_),
    .C1(_02545_),
    .C2(_02465_),
    .ZN(_04370_));
 OAI21_X1 _29599_ (.A(_02532_),
    .B1(_02539_),
    .B2(_02527_),
    .ZN(_04371_));
 NAND4_X1 _29600_ (.A1(_02672_),
    .A2(_03431_),
    .A3(_02991_),
    .A4(_02621_),
    .ZN(_04372_));
 AND4_X1 _29601_ (.A1(_02583_),
    .A2(_04371_),
    .A3(_03927_),
    .A4(_04372_),
    .ZN(_04374_));
 NAND2_X1 _29602_ (.A1(_03003_),
    .A2(_02434_),
    .ZN(_04375_));
 OAI21_X1 _29603_ (.A(_03003_),
    .B1(_02549_),
    .B2(_02390_),
    .ZN(_04376_));
 AND4_X1 _29604_ (.A1(_04375_),
    .A2(_02604_),
    .A3(_04376_),
    .A4(_02605_),
    .ZN(_04377_));
 AND4_X1 _29605_ (.A1(_04368_),
    .A2(_04370_),
    .A3(_04374_),
    .A4(_04377_),
    .ZN(_04378_));
 NAND4_X1 _29606_ (.A1(_04354_),
    .A2(_04359_),
    .A3(_04366_),
    .A4(_04378_),
    .ZN(_04379_));
 NOR2_X4 _29607_ (.A1(_04379_),
    .A2(_02670_),
    .ZN(_04380_));
 NAND4_X1 _29608_ (.A1(_02278_),
    .A2(_02211_),
    .A3(_02214_),
    .A4(_02280_),
    .ZN(_04381_));
 OAI21_X1 _29609_ (.A(_04381_),
    .B1(_02284_),
    .B2(_03808_),
    .ZN(_04382_));
 AND2_X1 _29610_ (.A1(_02218_),
    .A2(_02258_),
    .ZN(_04383_));
 AND2_X1 _29611_ (.A1(_02258_),
    .A2(_02250_),
    .ZN(_04385_));
 OR3_X4 _29612_ (.A1(_04383_),
    .A2(_02261_),
    .A3(_04385_),
    .ZN(_04386_));
 AND4_X1 _29613_ (.A1(_02211_),
    .A2(_02214_),
    .A3(_02252_),
    .A4(_02267_),
    .ZN(_04387_));
 NAND2_X1 _29614_ (.A1(_02156_),
    .A2(_02342_),
    .ZN(_04388_));
 NAND2_X1 _29615_ (.A1(_02208_),
    .A2(_02342_),
    .ZN(_04389_));
 NAND2_X1 _29616_ (.A1(_04388_),
    .A2(_04389_),
    .ZN(_04390_));
 OR4_X4 _29617_ (.A1(_04382_),
    .A2(_04386_),
    .A3(_04387_),
    .A4(_04390_),
    .ZN(_04391_));
 AND2_X1 _29618_ (.A1(_03059_),
    .A2(_02246_),
    .ZN(_04392_));
 AND2_X1 _29619_ (.A1(_02246_),
    .A2(_02189_),
    .ZN(_04393_));
 OR4_X1 _29620_ (.A1(_03061_),
    .A2(_04392_),
    .A3(_03087_),
    .A4(_04393_),
    .ZN(_04394_));
 AOI21_X1 _29621_ (.A(_03394_),
    .B1(_03872_),
    .B2(_02160_),
    .ZN(_04396_));
 NOR4_X2 _29622_ (.A1(_04391_),
    .A2(_04394_),
    .A3(_02360_),
    .A4(_04396_),
    .ZN(_04397_));
 AND4_X1 _29623_ (.A1(_02144_),
    .A2(_02237_),
    .A3(_02194_),
    .A4(_02326_),
    .ZN(_04398_));
 AOI221_X4 _29624_ (.A(_04398_),
    .B1(_02334_),
    .B2(_02286_),
    .C1(_03111_),
    .C2(_02350_),
    .ZN(_04399_));
 OAI21_X1 _29625_ (.A(_02334_),
    .B1(_02209_),
    .B2(_02251_),
    .ZN(_04400_));
 OAI21_X1 _29626_ (.A(_02353_),
    .B1(_02257_),
    .B2(_02346_),
    .ZN(_04401_));
 NAND2_X1 _29627_ (.A1(_02353_),
    .A2(_02209_),
    .ZN(_04402_));
 NAND4_X1 _29628_ (.A1(_02139_),
    .A2(_02243_),
    .A3(_02347_),
    .A4(_02280_),
    .ZN(_04403_));
 NAND3_X1 _29629_ (.A1(_04401_),
    .A2(_04402_),
    .A3(_04403_),
    .ZN(_04404_));
 AND3_X1 _29630_ (.A1(_02306_),
    .A2(_02347_),
    .A3(_02280_),
    .ZN(_04405_));
 NOR2_X1 _29631_ (.A1(_04404_),
    .A2(_04405_),
    .ZN(_04407_));
 OAI21_X1 _29632_ (.A(_02291_),
    .B1(_03096_),
    .B2(_02185_),
    .ZN(_04408_));
 OAI21_X1 _29633_ (.A(_02291_),
    .B1(_02221_),
    .B2(_02209_),
    .ZN(_04409_));
 AND3_X1 _29634_ (.A1(_04408_),
    .A2(_04409_),
    .A3(_02298_),
    .ZN(_04410_));
 AND4_X1 _29635_ (.A1(_04399_),
    .A2(_04400_),
    .A3(_04407_),
    .A4(_04410_),
    .ZN(_04411_));
 AOI22_X1 _29636_ (.A1(_03078_),
    .A2(_02328_),
    .B1(_02134_),
    .B2(_02286_),
    .ZN(_04412_));
 NAND2_X1 _29637_ (.A1(_02201_),
    .A2(_03871_),
    .ZN(_04413_));
 NAND3_X1 _29638_ (.A1(_02192_),
    .A2(_02194_),
    .A3(_02279_),
    .ZN(_04414_));
 NAND2_X1 _29639_ (.A1(_03097_),
    .A2(_02276_),
    .ZN(_04415_));
 AND4_X1 _29640_ (.A1(_04130_),
    .A2(_04413_),
    .A3(_04414_),
    .A4(_04415_),
    .ZN(_04416_));
 OAI21_X1 _29641_ (.A(_02226_),
    .B1(_03385_),
    .B2(_02178_),
    .ZN(_04418_));
 AND4_X1 _29642_ (.A1(_02282_),
    .A2(_04412_),
    .A3(_04416_),
    .A4(_04418_),
    .ZN(_04419_));
 OAI211_X2 _29643_ (.A(_04113_),
    .B(_04110_),
    .C1(_03807_),
    .C2(_03039_),
    .ZN(_04420_));
 NAND2_X1 _29644_ (.A1(_02315_),
    .A2(_02321_),
    .ZN(_04421_));
 NOR4_X1 _29645_ (.A1(_04420_),
    .A2(_04421_),
    .A3(_02345_),
    .A4(_03860_),
    .ZN(_04422_));
 NAND4_X2 _29646_ (.A1(_04397_),
    .A2(_04411_),
    .A3(_04419_),
    .A4(_04422_),
    .ZN(_04423_));
 AOI22_X1 _29647_ (.A1(_02302_),
    .A2(_03096_),
    .B1(_02134_),
    .B2(_02320_),
    .ZN(_04424_));
 OAI211_X2 _29648_ (.A(_04424_),
    .B(_03365_),
    .C1(_03883_),
    .C2(_03094_),
    .ZN(_04425_));
 OAI211_X2 _29649_ (.A(_02305_),
    .B(_02268_),
    .C1(_02193_),
    .C2(_02279_),
    .ZN(_04426_));
 OAI21_X1 _29650_ (.A(_02221_),
    .B1(_03097_),
    .B2(_02241_),
    .ZN(_04427_));
 OAI211_X2 _29651_ (.A(_04426_),
    .B(_04427_),
    .C1(_03807_),
    .C2(_04133_),
    .ZN(_04429_));
 NOR4_X1 _29652_ (.A1(_04425_),
    .A2(_04429_),
    .A3(_03064_),
    .A4(_04125_),
    .ZN(_04430_));
 OR2_X1 _29653_ (.A1(_02239_),
    .A2(_03877_),
    .ZN(_04431_));
 OAI21_X1 _29654_ (.A(_02176_),
    .B1(_04431_),
    .B2(_02211_),
    .ZN(_04432_));
 AOI22_X1 _29655_ (.A1(_03884_),
    .A2(_02226_),
    .B1(_02292_),
    .B2(_02302_),
    .ZN(_04433_));
 OAI21_X1 _29656_ (.A(_02202_),
    .B1(_02341_),
    .B2(_03037_),
    .ZN(_04434_));
 NAND2_X1 _29657_ (.A1(_04139_),
    .A2(_03396_),
    .ZN(_04435_));
 OAI21_X1 _29658_ (.A(_02134_),
    .B1(_04435_),
    .B2(_02230_),
    .ZN(_04436_));
 OAI21_X1 _29659_ (.A(_02182_),
    .B1(_02198_),
    .B2(_02286_),
    .ZN(_04437_));
 OAI21_X1 _29660_ (.A(_02182_),
    .B1(_02156_),
    .B2(_02320_),
    .ZN(_04438_));
 AND4_X1 _29661_ (.A1(_04434_),
    .A2(_04436_),
    .A3(_04437_),
    .A4(_04438_),
    .ZN(_04440_));
 NAND4_X1 _29662_ (.A1(_04430_),
    .A2(_04432_),
    .A3(_04433_),
    .A4(_04440_),
    .ZN(_04441_));
 NOR2_X4 _29663_ (.A1(_04423_),
    .A2(_04441_),
    .ZN(_04442_));
 XNOR2_X2 _29664_ (.A(_04380_),
    .B(_04442_),
    .ZN(_04443_));
 AND2_X1 _29665_ (.A1(_03134_),
    .A2(_02078_),
    .ZN(_04444_));
 INV_X1 _29666_ (.A(_04444_),
    .ZN(_04445_));
 NAND3_X1 _29667_ (.A1(_02061_),
    .A2(_01896_),
    .A3(_01973_),
    .ZN(_04446_));
 NAND2_X1 _29668_ (.A1(_02109_),
    .A2(_02102_),
    .ZN(_04447_));
 OAI21_X1 _29669_ (.A(_01898_),
    .B1(_04447_),
    .B2(_02048_),
    .ZN(_04448_));
 OAI21_X1 _29670_ (.A(_02078_),
    .B1(_02034_),
    .B2(_02093_),
    .ZN(_04449_));
 NAND4_X1 _29671_ (.A1(_04445_),
    .A2(_04446_),
    .A3(_04448_),
    .A4(_04449_),
    .ZN(_04451_));
 OAI221_X1 _29672_ (.A(_01966_),
    .B1(_02025_),
    .B2(_01971_),
    .C1(_01913_),
    .C2(_01934_),
    .ZN(_04452_));
 NAND2_X1 _29673_ (.A1(_02064_),
    .A2(_01966_),
    .ZN(_04453_));
 OAI211_X2 _29674_ (.A(_01966_),
    .B(_01908_),
    .C1(_02118_),
    .C2(_03159_),
    .ZN(_04454_));
 NAND3_X1 _29675_ (.A1(_04452_),
    .A2(_04453_),
    .A3(_04454_),
    .ZN(_04455_));
 INV_X1 _29676_ (.A(_01945_),
    .ZN(_04456_));
 AOI21_X1 _29677_ (.A(_02044_),
    .B1(_04456_),
    .B2(_02102_),
    .ZN(_04457_));
 AND2_X1 _29678_ (.A1(_01949_),
    .A2(_01984_),
    .ZN(_04458_));
 AND2_X4 _29679_ (.A1(_02121_),
    .A2(_01984_),
    .ZN(_04459_));
 OR4_X4 _29680_ (.A1(_03124_),
    .A2(_04457_),
    .A3(_04458_),
    .A4(_04459_),
    .ZN(_04460_));
 OAI21_X1 _29681_ (.A(_03130_),
    .B1(_02093_),
    .B2(_02106_),
    .ZN(_04462_));
 OAI21_X1 _29682_ (.A(_04462_),
    .B1(_03145_),
    .B2(_02044_),
    .ZN(_04463_));
 OR4_X4 _29683_ (.A1(_04451_),
    .A2(_04455_),
    .A3(_04460_),
    .A4(_04463_),
    .ZN(_04464_));
 NAND2_X1 _29684_ (.A1(_02001_),
    .A2(_03195_),
    .ZN(_04465_));
 AND2_X1 _29685_ (.A1(_02052_),
    .A2(_02020_),
    .ZN(_04466_));
 AOI211_X4 _29686_ (.A(_04466_),
    .B(_03198_),
    .C1(_02090_),
    .C2(_02021_),
    .ZN(_04467_));
 INV_X1 _29687_ (.A(_02055_),
    .ZN(_04468_));
 OAI21_X1 _29688_ (.A(_01980_),
    .B1(_01940_),
    .B2(_02015_),
    .ZN(_04469_));
 NAND2_X1 _29689_ (.A1(_01980_),
    .A2(_02113_),
    .ZN(_04470_));
 AND3_X1 _29690_ (.A1(_04469_),
    .A2(_03745_),
    .A3(_04470_),
    .ZN(_04471_));
 AND4_X2 _29691_ (.A1(_04465_),
    .A2(_04467_),
    .A3(_04468_),
    .A4(_04471_),
    .ZN(_04473_));
 AOI211_X4 _29692_ (.A(_02046_),
    .B(_04100_),
    .C1(_02072_),
    .C2(_02010_),
    .ZN(_04474_));
 OAI21_X1 _29693_ (.A(_02010_),
    .B1(_03154_),
    .B2(_03768_),
    .ZN(_04475_));
 OAI211_X2 _29694_ (.A(_02006_),
    .B(_01990_),
    .C1(_02113_),
    .C2(_02106_),
    .ZN(_04476_));
 AND4_X1 _29695_ (.A1(_02000_),
    .A2(_04096_),
    .A3(_02003_),
    .A4(_04476_),
    .ZN(_04477_));
 NAND4_X2 _29696_ (.A1(_04473_),
    .A2(_04474_),
    .A3(_04475_),
    .A4(_04477_),
    .ZN(_04478_));
 NOR2_X1 _29697_ (.A1(_02101_),
    .A2(_03182_),
    .ZN(_04479_));
 INV_X1 _29698_ (.A(_04479_),
    .ZN(_04480_));
 AND2_X1 _29699_ (.A1(_01995_),
    .A2(_01927_),
    .ZN(_04481_));
 AND2_X4 _29700_ (.A1(_01939_),
    .A2(_01927_),
    .ZN(_04482_));
 AND2_X1 _29701_ (.A1(_01968_),
    .A2(_01927_),
    .ZN(_04484_));
 NOR4_X2 _29702_ (.A1(_04481_),
    .A2(_04482_),
    .A3(_04077_),
    .A4(_04484_),
    .ZN(_04485_));
 OAI21_X1 _29703_ (.A(_02084_),
    .B1(_02054_),
    .B2(_02098_),
    .ZN(_04486_));
 AND4_X1 _29704_ (.A1(_04480_),
    .A2(_04485_),
    .A3(_03571_),
    .A4(_04486_),
    .ZN(_04487_));
 AOI211_X2 _29705_ (.A(_03170_),
    .B(_03173_),
    .C1(_01923_),
    .C2(_02123_),
    .ZN(_04488_));
 OAI221_X1 _29706_ (.A(_02123_),
    .B1(_03161_),
    .B2(_03159_),
    .C1(_02025_),
    .C2(_02098_),
    .ZN(_04489_));
 NAND2_X1 _29707_ (.A1(_02069_),
    .A2(_01949_),
    .ZN(_04490_));
 OAI21_X1 _29708_ (.A(_02070_),
    .B1(_03758_),
    .B2(_02061_),
    .ZN(_04491_));
 INV_X1 _29709_ (.A(_03178_),
    .ZN(_04492_));
 NAND4_X1 _29710_ (.A1(_01892_),
    .A2(_02005_),
    .A3(_01925_),
    .A4(_02006_),
    .ZN(_04493_));
 AND4_X1 _29711_ (.A1(_04490_),
    .A2(_04491_),
    .A3(_04492_),
    .A4(_04493_),
    .ZN(_04495_));
 NAND4_X1 _29712_ (.A1(_04487_),
    .A2(_04488_),
    .A3(_04489_),
    .A4(_04495_),
    .ZN(_04496_));
 AOI211_X4 _29713_ (.A(_01931_),
    .B(_03143_),
    .C1(_03161_),
    .C2(_02017_),
    .ZN(_04497_));
 AOI21_X1 _29714_ (.A(_03143_),
    .B1(_03783_),
    .B2(_01950_),
    .ZN(_04498_));
 NOR3_X1 _29715_ (.A1(_04497_),
    .A2(_03785_),
    .A3(_04498_),
    .ZN(_04499_));
 OAI21_X1 _29716_ (.A(_02014_),
    .B1(_01995_),
    .B2(_02081_),
    .ZN(_04500_));
 AND3_X1 _29717_ (.A1(_04500_),
    .A2(_02016_),
    .A3(_02018_),
    .ZN(_04501_));
 INV_X1 _29718_ (.A(_02065_),
    .ZN(_04502_));
 NAND2_X1 _29719_ (.A1(_01960_),
    .A2(_02026_),
    .ZN(_04503_));
 AND4_X1 _29720_ (.A1(_04060_),
    .A2(_03158_),
    .A3(_04502_),
    .A4(_04503_),
    .ZN(_04504_));
 NAND2_X1 _29721_ (.A1(_02080_),
    .A2(_02053_),
    .ZN(_04506_));
 OAI21_X1 _29722_ (.A(_01938_),
    .B1(_01999_),
    .B2(_01940_),
    .ZN(_04507_));
 NAND3_X1 _29723_ (.A1(_02080_),
    .A2(_02005_),
    .A3(_01892_),
    .ZN(_04508_));
 NAND2_X1 _29724_ (.A1(_02080_),
    .A2(_02112_),
    .ZN(_04509_));
 AND4_X1 _29725_ (.A1(_04506_),
    .A2(_04507_),
    .A3(_04508_),
    .A4(_04509_),
    .ZN(_04510_));
 NAND4_X1 _29726_ (.A1(_04499_),
    .A2(_04501_),
    .A3(_04504_),
    .A4(_04510_),
    .ZN(_04511_));
 NOR4_X4 _29727_ (.A1(_04464_),
    .A2(_04478_),
    .A3(_04496_),
    .A4(_04511_),
    .ZN(_04512_));
 NAND2_X2 _29728_ (.A1(_04512_),
    .A2(_02031_),
    .ZN(_04513_));
 XNOR2_X1 _29729_ (.A(_04513_),
    .B(_04246_),
    .ZN(_04514_));
 XNOR2_X1 _29730_ (.A(_04443_),
    .B(_04514_),
    .ZN(_04515_));
 AOI21_X1 _29731_ (.A(_03268_),
    .B1(_02900_),
    .B2(_02779_),
    .ZN(_04517_));
 AND4_X1 _29732_ (.A1(_02800_),
    .A2(_02845_),
    .A3(_02741_),
    .A4(_02753_),
    .ZN(_04518_));
 AND4_X1 _29733_ (.A1(_02755_),
    .A2(_02845_),
    .A3(_02741_),
    .A4(_02709_),
    .ZN(_04519_));
 OR4_X2 _29734_ (.A1(_03985_),
    .A2(_04517_),
    .A3(_04518_),
    .A4(_04519_),
    .ZN(_04520_));
 AND2_X1 _29735_ (.A1(_02898_),
    .A2(_02790_),
    .ZN(_04521_));
 NOR4_X4 _29736_ (.A1(_04520_),
    .A2(_03305_),
    .A3(_03667_),
    .A4(_04521_),
    .ZN(_04522_));
 OAI21_X1 _29737_ (.A(_02835_),
    .B1(_03259_),
    .B2(_03273_),
    .ZN(_04523_));
 OAI21_X1 _29738_ (.A(_02835_),
    .B1(_02881_),
    .B2(_02791_),
    .ZN(_04524_));
 OAI211_X2 _29739_ (.A(_02823_),
    .B(_16855_),
    .C1(_16854_),
    .C2(_02712_),
    .ZN(_04525_));
 AND4_X1 _29740_ (.A1(_03227_),
    .A2(_04523_),
    .A3(_04524_),
    .A4(_04525_),
    .ZN(_04526_));
 NAND3_X1 _29741_ (.A1(_04261_),
    .A2(_02873_),
    .A3(_02874_),
    .ZN(_04528_));
 OAI21_X1 _29742_ (.A(_04267_),
    .B1(_03623_),
    .B2(_02887_),
    .ZN(_04529_));
 NAND2_X1 _29743_ (.A1(_02731_),
    .A2(_03279_),
    .ZN(_04530_));
 NAND2_X1 _29744_ (.A1(_03279_),
    .A2(_02732_),
    .ZN(_04531_));
 OAI211_X2 _29745_ (.A(_04530_),
    .B(_04531_),
    .C1(_04262_),
    .C2(_03588_),
    .ZN(_04532_));
 NOR4_X1 _29746_ (.A1(_04528_),
    .A2(_03993_),
    .A3(_04529_),
    .A4(_04532_),
    .ZN(_04533_));
 OAI21_X1 _29747_ (.A(_02861_),
    .B1(_02784_),
    .B2(_02702_),
    .ZN(_04534_));
 OAI21_X1 _29748_ (.A(_02861_),
    .B1(_02903_),
    .B2(_02749_),
    .ZN(_04535_));
 NOR2_X1 _29749_ (.A1(_03217_),
    .A2(_03269_),
    .ZN(_04536_));
 NOR2_X1 _29750_ (.A1(_04536_),
    .A2(_04278_),
    .ZN(_04537_));
 AND4_X1 _29751_ (.A1(_03291_),
    .A2(_04534_),
    .A3(_04535_),
    .A4(_04537_),
    .ZN(_04539_));
 NAND4_X1 _29752_ (.A1(_04522_),
    .A2(_04526_),
    .A3(_04533_),
    .A4(_04539_),
    .ZN(_04540_));
 NOR2_X1 _29753_ (.A1(_02692_),
    .A2(_02695_),
    .ZN(_04541_));
 OAI21_X1 _29754_ (.A(_02727_),
    .B1(_02902_),
    .B2(_02778_),
    .ZN(_04542_));
 OAI211_X2 _29755_ (.A(_02727_),
    .B(_02858_),
    .C1(_02856_),
    .C2(_02857_),
    .ZN(_04543_));
 AND3_X1 _29756_ (.A1(_04542_),
    .A2(_04296_),
    .A3(_04543_),
    .ZN(_04544_));
 OAI21_X1 _29757_ (.A(_02697_),
    .B1(_02756_),
    .B2(_02732_),
    .ZN(_04545_));
 NAND3_X1 _29758_ (.A1(_02801_),
    .A2(_02683_),
    .A3(_02773_),
    .ZN(_04546_));
 AND3_X1 _29759_ (.A1(_02720_),
    .A2(_03216_),
    .A3(_04546_),
    .ZN(_04547_));
 AND4_X1 _29760_ (.A1(_04541_),
    .A2(_04544_),
    .A3(_04545_),
    .A4(_04547_),
    .ZN(_04548_));
 AOI21_X1 _29761_ (.A(_03611_),
    .B1(_02900_),
    .B2(_03623_),
    .ZN(_04550_));
 NAND2_X1 _29762_ (.A1(_03309_),
    .A2(_02747_),
    .ZN(_04551_));
 OAI211_X2 _29763_ (.A(_02776_),
    .B(_04551_),
    .C1(_02777_),
    .C2(_02886_),
    .ZN(_04552_));
 AOI21_X1 _29764_ (.A(_02777_),
    .B1(_03588_),
    .B2(_04008_),
    .ZN(_04553_));
 NOR4_X1 _29765_ (.A1(_04550_),
    .A2(_04552_),
    .A3(_04553_),
    .A4(_03606_),
    .ZN(_04554_));
 OAI21_X1 _29766_ (.A(_02752_),
    .B1(_02731_),
    .B2(_02797_),
    .ZN(_04555_));
 NAND3_X1 _29767_ (.A1(_02759_),
    .A2(_02735_),
    .A3(_02859_),
    .ZN(_04556_));
 NAND2_X1 _29768_ (.A1(_02767_),
    .A2(_02759_),
    .ZN(_04557_));
 AND3_X1 _29769_ (.A1(_04556_),
    .A2(_04557_),
    .A3(_02760_),
    .ZN(_04558_));
 OAI21_X1 _29770_ (.A(_03222_),
    .B1(_03259_),
    .B2(_02736_),
    .ZN(_04559_));
 OAI21_X1 _29771_ (.A(_02752_),
    .B1(_02864_),
    .B2(_03595_),
    .ZN(_04561_));
 AND4_X1 _29772_ (.A1(_04555_),
    .A2(_04558_),
    .A3(_04559_),
    .A4(_04561_),
    .ZN(_04562_));
 OAI21_X1 _29773_ (.A(_02799_),
    .B1(_02701_),
    .B2(_02831_),
    .ZN(_04563_));
 NAND3_X1 _29774_ (.A1(_02732_),
    .A2(_02724_),
    .A3(_02743_),
    .ZN(_04564_));
 NAND4_X1 _29775_ (.A1(_03246_),
    .A2(_02724_),
    .A3(_02859_),
    .A4(_02743_),
    .ZN(_04565_));
 NAND3_X1 _29776_ (.A1(_04563_),
    .A2(_04564_),
    .A3(_04565_),
    .ZN(_04566_));
 NAND2_X1 _29777_ (.A1(_02731_),
    .A2(_02796_),
    .ZN(_04567_));
 NAND3_X1 _29778_ (.A1(_02796_),
    .A2(_02863_),
    .A3(_03233_),
    .ZN(_04568_));
 NAND2_X1 _29779_ (.A1(_02795_),
    .A2(_02704_),
    .ZN(_04569_));
 NAND3_X1 _29780_ (.A1(_04567_),
    .A2(_04568_),
    .A3(_04569_),
    .ZN(_04570_));
 NOR4_X1 _29781_ (.A1(_03240_),
    .A2(_04566_),
    .A3(_03594_),
    .A4(_04570_),
    .ZN(_04572_));
 NAND4_X1 _29782_ (.A1(_04548_),
    .A2(_04554_),
    .A3(_04562_),
    .A4(_04572_),
    .ZN(_04573_));
 NOR2_X2 _29783_ (.A1(_04540_),
    .A2(_04573_),
    .ZN(_04574_));
 XNOR2_X1 _29784_ (.A(_04515_),
    .B(_04574_),
    .ZN(_04575_));
 XNOR2_X1 _29785_ (.A(_04575_),
    .B(_17235_),
    .ZN(_04576_));
 MUX2_X1 _29786_ (.A(_04324_),
    .B(_04576_),
    .S(_01876_),
    .Z(_00713_));
 XOR2_X1 _29787_ (.A(_17236_),
    .B(_17107_),
    .Z(_04577_));
 OAI21_X1 _29788_ (.A(_02241_),
    .B1(_02264_),
    .B2(_02266_),
    .ZN(_04578_));
 NAND2_X1 _29789_ (.A1(_02247_),
    .A2(_02294_),
    .ZN(_04579_));
 OR2_X4 _29790_ (.A1(_02259_),
    .A2(_03882_),
    .ZN(_04580_));
 AOI211_X2 _29791_ (.A(_04383_),
    .B(_04580_),
    .C1(_03018_),
    .C2(_02258_),
    .ZN(_04582_));
 OAI21_X1 _29792_ (.A(_02246_),
    .B1(_02209_),
    .B2(_02276_),
    .ZN(_04583_));
 AND4_X2 _29793_ (.A1(_04579_),
    .A2(_04582_),
    .A3(_03887_),
    .A4(_04583_),
    .ZN(_04584_));
 INV_X1 _29794_ (.A(_03419_),
    .ZN(_04585_));
 OAI21_X1 _29795_ (.A(_02226_),
    .B1(_02294_),
    .B2(_02185_),
    .ZN(_04586_));
 OAI21_X1 _29796_ (.A(_02226_),
    .B1(_02335_),
    .B2(_02251_),
    .ZN(_04587_));
 AND3_X1 _29797_ (.A1(_04586_),
    .A2(_04587_),
    .A3(_03854_),
    .ZN(_04588_));
 AND4_X4 _29798_ (.A1(_04578_),
    .A2(_04584_),
    .A3(_04585_),
    .A4(_04588_),
    .ZN(_04589_));
 OAI21_X1 _29799_ (.A(_02275_),
    .B1(_04431_),
    .B2(_02153_),
    .ZN(_04590_));
 AND3_X1 _29800_ (.A1(_03081_),
    .A2(_02278_),
    .A3(_02267_),
    .ZN(_04591_));
 AND4_X1 _29801_ (.A1(_02350_),
    .A2(_02278_),
    .A3(_02211_),
    .A4(_02267_),
    .ZN(_04593_));
 NOR4_X1 _29802_ (.A1(_03072_),
    .A2(_04126_),
    .A3(_04591_),
    .A4(_04593_),
    .ZN(_04594_));
 OAI21_X1 _29803_ (.A(_02291_),
    .B1(_02318_),
    .B2(_02189_),
    .ZN(_04595_));
 AND3_X1 _29804_ (.A1(_04595_),
    .A2(_03085_),
    .A3(_03866_),
    .ZN(_04596_));
 NAND3_X1 _29805_ (.A1(_02185_),
    .A2(_02194_),
    .A3(_02279_),
    .ZN(_04597_));
 OAI211_X2 _29806_ (.A(_02194_),
    .B(_02278_),
    .C1(_02306_),
    .C2(_02286_),
    .ZN(_04598_));
 NAND4_X1 _29807_ (.A1(_02278_),
    .A2(_02220_),
    .A3(_02194_),
    .A4(_02191_),
    .ZN(_04599_));
 AND4_X1 _29808_ (.A1(_04597_),
    .A2(_04598_),
    .A3(_02310_),
    .A4(_04599_),
    .ZN(_04600_));
 AND4_X1 _29809_ (.A1(_04590_),
    .A2(_04594_),
    .A3(_04596_),
    .A4(_04600_),
    .ZN(_04601_));
 AND4_X1 _29810_ (.A1(_02146_),
    .A2(_02326_),
    .A3(_02169_),
    .A4(_02267_),
    .ZN(_04602_));
 AND2_X1 _29811_ (.A1(_02342_),
    .A2(_02285_),
    .ZN(_04604_));
 AOI211_X4 _29812_ (.A(_04602_),
    .B(_04604_),
    .C1(_02239_),
    .C2(_03097_),
    .ZN(_04605_));
 OAI21_X1 _29813_ (.A(_02353_),
    .B1(_03371_),
    .B2(_03050_),
    .ZN(_04606_));
 AND3_X1 _29814_ (.A1(_02260_),
    .A2(_02326_),
    .A3(_02164_),
    .ZN(_04607_));
 AND2_X1 _29815_ (.A1(_02352_),
    .A2(_02257_),
    .ZN(_04608_));
 AOI211_X2 _29816_ (.A(_04607_),
    .B(_04608_),
    .C1(_02352_),
    .C2(_03877_),
    .ZN(_04609_));
 OAI211_X2 _29817_ (.A(_03032_),
    .B(_02347_),
    .C1(_02359_),
    .C2(_02230_),
    .ZN(_04610_));
 OAI21_X1 _29818_ (.A(_02328_),
    .B1(_03083_),
    .B2(_02206_),
    .ZN(_04611_));
 AND4_X1 _29819_ (.A1(_04606_),
    .A2(_04609_),
    .A3(_04610_),
    .A4(_04611_),
    .ZN(_04612_));
 OAI211_X2 _29820_ (.A(_03097_),
    .B(_16807_),
    .C1(_03055_),
    .C2(_02135_),
    .ZN(_04613_));
 NAND2_X1 _29821_ (.A1(_02334_),
    .A2(_02251_),
    .ZN(_04615_));
 NAND2_X1 _29822_ (.A1(_02334_),
    .A2(_02359_),
    .ZN(_04616_));
 AND4_X1 _29823_ (.A1(_03110_),
    .A2(_03824_),
    .A3(_04615_),
    .A4(_04616_),
    .ZN(_04617_));
 AND4_X4 _29824_ (.A1(_04605_),
    .A2(_04612_),
    .A3(_04613_),
    .A4(_04617_),
    .ZN(_04618_));
 OAI21_X1 _29825_ (.A(_02134_),
    .B1(_03371_),
    .B2(_03050_),
    .ZN(_04619_));
 OAI21_X1 _29826_ (.A(_02201_),
    .B1(_02221_),
    .B2(_02153_),
    .ZN(_04620_));
 OAI211_X2 _29827_ (.A(_02201_),
    .B(_02237_),
    .C1(_02173_),
    .C2(_02174_),
    .ZN(_04621_));
 AND2_X1 _29828_ (.A1(_04620_),
    .A2(_04621_),
    .ZN(_04622_));
 NAND2_X1 _29829_ (.A1(_02182_),
    .A2(_02286_),
    .ZN(_04623_));
 OAI21_X1 _29830_ (.A(_02182_),
    .B1(_03083_),
    .B2(_02320_),
    .ZN(_04624_));
 AND4_X1 _29831_ (.A1(_02187_),
    .A2(_04622_),
    .A3(_04623_),
    .A4(_04624_),
    .ZN(_04626_));
 OAI21_X1 _29832_ (.A(_02134_),
    .B1(_02153_),
    .B2(_03877_),
    .ZN(_04627_));
 AND2_X1 _29833_ (.A1(_02205_),
    .A2(_02165_),
    .ZN(_04628_));
 INV_X1 _29834_ (.A(_04628_),
    .ZN(_04629_));
 OAI21_X1 _29835_ (.A(_02176_),
    .B1(_02305_),
    .B2(_03081_),
    .ZN(_04630_));
 NAND4_X1 _29836_ (.A1(_02214_),
    .A2(_02243_),
    .A3(_02193_),
    .A4(_02280_),
    .ZN(_04631_));
 AND4_X1 _29837_ (.A1(_03042_),
    .A2(_04629_),
    .A3(_04630_),
    .A4(_04631_),
    .ZN(_04632_));
 AND4_X1 _29838_ (.A1(_04619_),
    .A2(_04626_),
    .A3(_04627_),
    .A4(_04632_),
    .ZN(_04633_));
 NAND4_X4 _29839_ (.A1(_04589_),
    .A2(_04601_),
    .A3(_04618_),
    .A4(_04633_),
    .ZN(_04634_));
 NOR2_X4 _29840_ (.A1(_04634_),
    .A2(_02360_),
    .ZN(_04635_));
 INV_X1 _29841_ (.A(_03938_),
    .ZN(_04637_));
 NAND2_X1 _29842_ (.A1(_02556_),
    .A2(_02419_),
    .ZN(_04638_));
 NAND2_X1 _29843_ (.A1(_02556_),
    .A2(_03437_),
    .ZN(_04639_));
 NAND4_X1 _29844_ (.A1(_04637_),
    .A2(_04638_),
    .A3(_02952_),
    .A4(_04639_),
    .ZN(_04640_));
 AND2_X1 _29845_ (.A1(_02557_),
    .A2(_02445_),
    .ZN(_04641_));
 AOI21_X1 _29846_ (.A(_03465_),
    .B1(_02417_),
    .B2(_02589_),
    .ZN(_04642_));
 NAND2_X1 _29847_ (.A1(_02475_),
    .A2(_03462_),
    .ZN(_04643_));
 AND4_X2 _29848_ (.A1(_02371_),
    .A2(_02509_),
    .A3(_02378_),
    .A4(_02593_),
    .ZN(_04644_));
 OR4_X4 _29849_ (.A1(_04641_),
    .A2(_04642_),
    .A3(_04643_),
    .A4(_04644_),
    .ZN(_04645_));
 OAI21_X1 _29850_ (.A(_02610_),
    .B1(_02421_),
    .B2(_02987_),
    .ZN(_04646_));
 NAND4_X1 _29851_ (.A1(_02991_),
    .A2(_02553_),
    .A3(_02506_),
    .A4(_02944_),
    .ZN(_04648_));
 OAI21_X1 _29852_ (.A(_02610_),
    .B1(_02423_),
    .B2(_02445_),
    .ZN(_04649_));
 NAND3_X1 _29853_ (.A1(_04646_),
    .A2(_04648_),
    .A3(_04649_),
    .ZN(_04650_));
 OAI211_X2 _29854_ (.A(_03431_),
    .B(_02553_),
    .C1(_02419_),
    .C2(_02619_),
    .ZN(_04651_));
 OAI211_X2 _29855_ (.A(_04651_),
    .B(_04206_),
    .C1(_02385_),
    .C2(_02493_),
    .ZN(_04652_));
 NOR4_X4 _29856_ (.A1(_04640_),
    .A2(_04645_),
    .A3(_04650_),
    .A4(_04652_),
    .ZN(_04653_));
 OAI21_X1 _29857_ (.A(_02548_),
    .B1(_02999_),
    .B2(_03893_),
    .ZN(_04654_));
 NAND4_X1 _29858_ (.A1(_02509_),
    .A2(_02672_),
    .A3(_02371_),
    .A4(_02944_),
    .ZN(_04655_));
 AND2_X1 _29859_ (.A1(_04654_),
    .A2(_04655_),
    .ZN(_04656_));
 AOI21_X1 _29860_ (.A(_02469_),
    .B1(_02417_),
    .B2(_02589_),
    .ZN(_04657_));
 NAND3_X4 _29861_ (.A1(_02572_),
    .A2(_02534_),
    .A3(_02429_),
    .ZN(_04659_));
 NAND4_X1 _29862_ (.A1(_02534_),
    .A2(_02429_),
    .A3(_02394_),
    .A4(_02621_),
    .ZN(_04660_));
 OAI211_X2 _29863_ (.A(_04659_),
    .B(_04660_),
    .C1(_02469_),
    .C2(_02493_),
    .ZN(_04661_));
 AOI211_X4 _29864_ (.A(_04657_),
    .B(_04661_),
    .C1(_02527_),
    .C2(_02465_),
    .ZN(_04662_));
 AND2_X1 _29865_ (.A1(_02583_),
    .A2(_02584_),
    .ZN(_04663_));
 AND2_X1 _29866_ (.A1(_02532_),
    .A2(_02439_),
    .ZN(_04664_));
 INV_X1 _29867_ (.A(_04664_),
    .ZN(_04665_));
 AND4_X1 _29868_ (.A1(_04663_),
    .A2(_04665_),
    .A3(_02995_),
    .A4(_03925_),
    .ZN(_04666_));
 INV_X1 _29869_ (.A(_02501_),
    .ZN(_04667_));
 OAI21_X1 _29870_ (.A(_03003_),
    .B1(_02999_),
    .B2(_02466_),
    .ZN(_04668_));
 NAND3_X1 _29871_ (.A1(_02611_),
    .A2(_02672_),
    .A3(_02593_),
    .ZN(_04670_));
 AND4_X1 _29872_ (.A1(_04667_),
    .A2(_04668_),
    .A3(_02568_),
    .A4(_04670_),
    .ZN(_04671_));
 AND4_X4 _29873_ (.A1(_04656_),
    .A2(_04662_),
    .A3(_04666_),
    .A4(_04671_),
    .ZN(_04672_));
 AND2_X1 _29874_ (.A1(_02505_),
    .A2(_02614_),
    .ZN(_04673_));
 AND2_X1 _29875_ (.A1(_02549_),
    .A2(_02614_),
    .ZN(_04674_));
 AND2_X1 _29876_ (.A1(_02494_),
    .A2(_02444_),
    .ZN(_04675_));
 OR4_X2 _29877_ (.A1(_04673_),
    .A2(_02519_),
    .A3(_04674_),
    .A4(_04675_),
    .ZN(_04676_));
 OAI21_X1 _29878_ (.A(_02516_),
    .B1(_02390_),
    .B2(_02527_),
    .ZN(_04677_));
 OAI21_X1 _29879_ (.A(_02516_),
    .B1(_02560_),
    .B2(_03437_),
    .ZN(_04678_));
 NAND3_X1 _29880_ (.A1(_04677_),
    .A2(_04678_),
    .A3(_03908_),
    .ZN(_04679_));
 OAI21_X1 _29881_ (.A(_02449_),
    .B1(_02390_),
    .B2(_02527_),
    .ZN(_04681_));
 NAND4_X1 _29882_ (.A1(_02991_),
    .A2(_02598_),
    .A3(_02446_),
    .A4(_02944_),
    .ZN(_04682_));
 NAND4_X1 _29883_ (.A1(_04225_),
    .A2(_03482_),
    .A3(_04681_),
    .A4(_04682_),
    .ZN(_04683_));
 NAND2_X1 _29884_ (.A1(_02522_),
    .A2(_02528_),
    .ZN(_04684_));
 NAND4_X1 _29885_ (.A1(_02983_),
    .A2(_03914_),
    .A3(_02627_),
    .A4(_04684_),
    .ZN(_04685_));
 NOR4_X1 _29886_ (.A1(_04676_),
    .A2(_04679_),
    .A3(_04683_),
    .A4(_04685_),
    .ZN(_04686_));
 OAI21_X1 _29887_ (.A(_02662_),
    .B1(_02421_),
    .B2(_02987_),
    .ZN(_04687_));
 OAI21_X1 _29888_ (.A(_02525_),
    .B1(_02650_),
    .B2(_02564_),
    .ZN(_04688_));
 OAI211_X2 _29889_ (.A(_02524_),
    .B(_02581_),
    .C1(_02388_),
    .C2(_02535_),
    .ZN(_04689_));
 AND2_X1 _29890_ (.A1(_04688_),
    .A2(_04689_),
    .ZN(_04690_));
 NAND2_X1 _29891_ (.A1(_02572_),
    .A2(_02431_),
    .ZN(_04692_));
 OAI21_X1 _29892_ (.A(_02431_),
    .B1(_02527_),
    .B2(_02441_),
    .ZN(_04693_));
 AND4_X1 _29893_ (.A1(_03451_),
    .A2(_04690_),
    .A3(_04692_),
    .A4(_04693_),
    .ZN(_04694_));
 OAI21_X1 _29894_ (.A(_02662_),
    .B1(_02999_),
    .B2(_03893_),
    .ZN(_04695_));
 AOI21_X1 _29895_ (.A(_03441_),
    .B1(_02550_),
    .B2(_02484_),
    .ZN(_04696_));
 AND4_X1 _29896_ (.A1(_02499_),
    .A2(_02598_),
    .A3(_02472_),
    .A4(_02411_),
    .ZN(_04697_));
 NOR4_X1 _29897_ (.A1(_04696_),
    .A2(_03963_),
    .A3(_02957_),
    .A4(_04697_),
    .ZN(_04698_));
 AND4_X2 _29898_ (.A1(_04687_),
    .A2(_04694_),
    .A3(_04695_),
    .A4(_04698_),
    .ZN(_04699_));
 NAND4_X1 _29899_ (.A1(_04653_),
    .A2(_04672_),
    .A3(_04686_),
    .A4(_04699_),
    .ZN(_04700_));
 NOR2_X2 _29900_ (.A1(_04700_),
    .A2(_02670_),
    .ZN(_04701_));
 XOR2_X2 _29901_ (.A(_04635_),
    .B(_04701_),
    .Z(_04703_));
 AND4_X1 _29902_ (.A1(_01924_),
    .A2(_01894_),
    .A3(_01913_),
    .A4(_01907_),
    .ZN(_04704_));
 AND2_X1 _29903_ (.A1(_01983_),
    .A2(_02039_),
    .ZN(_04705_));
 AOI211_X4 _29904_ (.A(_04704_),
    .B(_04705_),
    .C1(_02072_),
    .C2(_01984_),
    .ZN(_04706_));
 OAI21_X1 _29905_ (.A(_03130_),
    .B1(_03154_),
    .B2(_03202_),
    .ZN(_04707_));
 OAI21_X1 _29906_ (.A(_03130_),
    .B1(_01999_),
    .B2(_02122_),
    .ZN(_04708_));
 AND3_X1 _29907_ (.A1(_04706_),
    .A2(_04707_),
    .A3(_04708_),
    .ZN(_04709_));
 NAND3_X1 _29908_ (.A1(_02093_),
    .A2(_01972_),
    .A3(_01973_),
    .ZN(_04710_));
 AND2_X1 _29909_ (.A1(_03731_),
    .A2(_04710_),
    .ZN(_04711_));
 NAND2_X1 _29910_ (.A1(_01966_),
    .A2(_02015_),
    .ZN(_04712_));
 AND4_X1 _29911_ (.A1(_03728_),
    .A2(_04711_),
    .A3(_03123_),
    .A4(_04712_),
    .ZN(_04714_));
 NAND2_X1 _29912_ (.A1(_02033_),
    .A2(_01898_),
    .ZN(_04715_));
 NAND4_X1 _29913_ (.A1(_01986_),
    .A2(_01973_),
    .A3(_01910_),
    .A4(_01896_),
    .ZN(_04716_));
 NAND4_X1 _29914_ (.A1(_01971_),
    .A2(_01973_),
    .A3(_01910_),
    .A4(_01896_),
    .ZN(_04717_));
 OAI21_X1 _29915_ (.A(_01897_),
    .B1(_01967_),
    .B2(_01969_),
    .ZN(_04718_));
 AND4_X1 _29916_ (.A1(_04715_),
    .A2(_04716_),
    .A3(_04717_),
    .A4(_04718_),
    .ZN(_04719_));
 NAND3_X1 _29917_ (.A1(_02093_),
    .A2(_01918_),
    .A3(_01973_),
    .ZN(_04720_));
 NAND2_X1 _29918_ (.A1(_03538_),
    .A2(_04720_),
    .ZN(_04721_));
 AOI211_X4 _29919_ (.A(_03138_),
    .B(_04721_),
    .C1(_01985_),
    .C2(_03136_),
    .ZN(_04722_));
 AND4_X1 _29920_ (.A1(_04709_),
    .A2(_04714_),
    .A3(_04719_),
    .A4(_04722_),
    .ZN(_04723_));
 AND2_X1 _29921_ (.A1(_02069_),
    .A2(_01961_),
    .ZN(_04725_));
 AOI211_X2 _29922_ (.A(_03179_),
    .B(_04725_),
    .C1(_02070_),
    .C2(_01967_),
    .ZN(_04726_));
 OAI21_X1 _29923_ (.A(_02070_),
    .B1(_02064_),
    .B2(_02090_),
    .ZN(_04727_));
 NAND4_X1 _29924_ (.A1(_04726_),
    .A2(_03792_),
    .A3(_03793_),
    .A4(_04727_),
    .ZN(_04728_));
 AOI221_X1 _29925_ (.A(_04482_),
    .B1(_01914_),
    .B2(_01927_),
    .C1(_01910_),
    .C2(_04484_),
    .ZN(_04729_));
 AND2_X1 _29926_ (.A1(_02103_),
    .A2(_02082_),
    .ZN(_04730_));
 INV_X1 _29927_ (.A(_04730_),
    .ZN(_04731_));
 OAI21_X1 _29928_ (.A(_02084_),
    .B1(_02053_),
    .B2(_02112_),
    .ZN(_04732_));
 OAI21_X1 _29929_ (.A(_02084_),
    .B1(_02122_),
    .B2(_01969_),
    .ZN(_04733_));
 NAND4_X1 _29930_ (.A1(_04729_),
    .A2(_04731_),
    .A3(_04732_),
    .A4(_04733_),
    .ZN(_04734_));
 NOR2_X1 _29931_ (.A1(_02119_),
    .A2(_02028_),
    .ZN(_04736_));
 NOR4_X2 _29932_ (.A1(_04728_),
    .A2(_04734_),
    .A3(_04736_),
    .A4(_03559_),
    .ZN(_04737_));
 AND2_X1 _29933_ (.A1(_02013_),
    .A2(_01945_),
    .ZN(_04738_));
 AOI211_X4 _29934_ (.A(_04738_),
    .B(_03150_),
    .C1(_02014_),
    .C2(_03768_),
    .ZN(_04739_));
 AND2_X1 _29935_ (.A1(_01957_),
    .A2(_01959_),
    .ZN(_04740_));
 NOR4_X1 _29936_ (.A1(_03781_),
    .A2(_04740_),
    .A3(_03142_),
    .A4(_03786_),
    .ZN(_04741_));
 AND2_X1 _29937_ (.A1(_01954_),
    .A2(_03202_),
    .ZN(_04742_));
 INV_X1 _29938_ (.A(_04742_),
    .ZN(_04743_));
 OAI21_X1 _29939_ (.A(_01954_),
    .B1(_01999_),
    .B2(_01940_),
    .ZN(_04744_));
 OAI211_X2 _29940_ (.A(_01916_),
    .B(_01972_),
    .C1(_02060_),
    .C2(_02113_),
    .ZN(_04745_));
 AND4_X1 _29941_ (.A1(_02115_),
    .A2(_04743_),
    .A3(_04744_),
    .A4(_04745_),
    .ZN(_04747_));
 OAI21_X1 _29942_ (.A(_01938_),
    .B1(_02090_),
    .B2(_01911_),
    .ZN(_04748_));
 NAND2_X1 _29943_ (.A1(_01938_),
    .A2(_02001_),
    .ZN(_04749_));
 AND3_X1 _29944_ (.A1(_03165_),
    .A2(_04748_),
    .A3(_04749_),
    .ZN(_04750_));
 AND4_X1 _29945_ (.A1(_04739_),
    .A2(_04741_),
    .A3(_04747_),
    .A4(_04750_),
    .ZN(_04751_));
 OAI21_X1 _29946_ (.A(_01992_),
    .B1(_03154_),
    .B2(_03768_),
    .ZN(_04752_));
 NAND4_X1 _29947_ (.A1(_02032_),
    .A2(_01985_),
    .A3(_02006_),
    .A4(_01990_),
    .ZN(_04753_));
 NAND4_X1 _29948_ (.A1(_02006_),
    .A2(_03159_),
    .A3(_01986_),
    .A4(_01990_),
    .ZN(_04754_));
 AND3_X1 _29949_ (.A1(_04752_),
    .A2(_04753_),
    .A3(_04754_),
    .ZN(_04755_));
 NAND2_X1 _29950_ (.A1(_03202_),
    .A2(_02009_),
    .ZN(_04756_));
 AND2_X1 _29951_ (.A1(_01999_),
    .A2(_02009_),
    .ZN(_04758_));
 INV_X1 _29952_ (.A(_04758_),
    .ZN(_04759_));
 NAND2_X1 _29953_ (.A1(_02001_),
    .A2(_02009_),
    .ZN(_04760_));
 OAI21_X1 _29954_ (.A(_02009_),
    .B1(_02053_),
    .B2(_02090_),
    .ZN(_04761_));
 AND4_X1 _29955_ (.A1(_04756_),
    .A2(_04759_),
    .A3(_04760_),
    .A4(_04761_),
    .ZN(_04762_));
 OAI21_X1 _29956_ (.A(_01980_),
    .B1(_03517_),
    .B2(_01940_),
    .ZN(_04763_));
 AND4_X1 _29957_ (.A1(_03745_),
    .A2(_04763_),
    .A3(_03747_),
    .A4(_04470_),
    .ZN(_04764_));
 OAI21_X1 _29958_ (.A(_03195_),
    .B1(_01949_),
    .B2(_03154_),
    .ZN(_04765_));
 OAI211_X2 _29959_ (.A(_03195_),
    .B(_02099_),
    .C1(_03161_),
    .C2(_02017_),
    .ZN(_04766_));
 AND2_X1 _29960_ (.A1(_04765_),
    .A2(_04766_),
    .ZN(_04767_));
 AND4_X1 _29961_ (.A1(_04755_),
    .A2(_04762_),
    .A3(_04764_),
    .A4(_04767_),
    .ZN(_04769_));
 NAND4_X2 _29962_ (.A1(_04723_),
    .A2(_04737_),
    .A3(_04751_),
    .A4(_04769_),
    .ZN(_04770_));
 NOR2_X4 _29963_ (.A1(_04770_),
    .A2(_02030_),
    .ZN(_04771_));
 XNOR2_X1 _29964_ (.A(_04380_),
    .B(_04771_),
    .ZN(_04772_));
 XNOR2_X2 _29965_ (.A(_04703_),
    .B(_04772_),
    .ZN(_04773_));
 AND2_X1 _29966_ (.A1(_02897_),
    .A2(_03595_),
    .ZN(_04774_));
 AND2_X1 _29967_ (.A1(_03616_),
    .A2(_02818_),
    .ZN(_04775_));
 NOR4_X1 _29968_ (.A1(_04774_),
    .A2(_04775_),
    .A3(_03238_),
    .A4(_04291_),
    .ZN(_04776_));
 AOI22_X1 _29969_ (.A1(_02778_),
    .A2(_02847_),
    .B1(_02861_),
    .B2(_03230_),
    .ZN(_04777_));
 NAND4_X1 _29970_ (.A1(_04776_),
    .A2(_03653_),
    .A3(_03601_),
    .A4(_04777_),
    .ZN(_04778_));
 NAND2_X1 _29971_ (.A1(_03616_),
    .A2(_02847_),
    .ZN(_04780_));
 AND3_X1 _29972_ (.A1(_02872_),
    .A2(_02849_),
    .A3(_04780_),
    .ZN(_04781_));
 AOI22_X1 _29973_ (.A1(_03595_),
    .A2(_02752_),
    .B1(_02749_),
    .B2(_02795_),
    .ZN(_04782_));
 AOI22_X1 _29974_ (.A1(_02835_),
    .A2(_02736_),
    .B1(_02861_),
    .B2(_02710_),
    .ZN(_04783_));
 NAND4_X1 _29975_ (.A1(_04781_),
    .A2(_02874_),
    .A3(_04782_),
    .A4(_04783_),
    .ZN(_04784_));
 OAI221_X1 _29976_ (.A(_02854_),
    .B1(_03268_),
    .B2(_02901_),
    .C1(_03214_),
    .C2(_04008_),
    .ZN(_04785_));
 AOI22_X1 _29977_ (.A1(_02726_),
    .A2(_02778_),
    .B1(_02710_),
    .B2(_02823_),
    .ZN(_04786_));
 NAND2_X1 _29978_ (.A1(_03259_),
    .A2(_02759_),
    .ZN(_04787_));
 OAI211_X2 _29979_ (.A(_04786_),
    .B(_04787_),
    .C1(_02842_),
    .C2(_02765_),
    .ZN(_04788_));
 NOR4_X1 _29980_ (.A1(_04778_),
    .A2(_04784_),
    .A3(_04785_),
    .A4(_04788_),
    .ZN(_04789_));
 AND2_X1 _29981_ (.A1(_02868_),
    .A2(_02881_),
    .ZN(_04791_));
 AND2_X1 _29982_ (.A1(_02726_),
    .A2(_03271_),
    .ZN(_04792_));
 AND3_X1 _29983_ (.A1(_03254_),
    .A2(_02722_),
    .A3(_02817_),
    .ZN(_04793_));
 OR4_X4 _29984_ (.A1(_04791_),
    .A2(_04792_),
    .A3(_03659_),
    .A4(_04793_),
    .ZN(_04794_));
 OAI211_X2 _29985_ (.A(_04267_),
    .B(_04546_),
    .C1(_02783_),
    .C2(_03268_),
    .ZN(_04795_));
 NAND4_X1 _29986_ (.A1(_02696_),
    .A2(_02824_),
    .A3(_03991_),
    .A4(_02716_),
    .ZN(_04796_));
 NAND4_X1 _29987_ (.A1(_02822_),
    .A2(_02763_),
    .A3(_02837_),
    .A4(_04557_),
    .ZN(_04797_));
 NOR4_X1 _29988_ (.A1(_04794_),
    .A2(_04795_),
    .A3(_04796_),
    .A4(_04797_),
    .ZN(_04798_));
 OAI21_X1 _29989_ (.A(_02835_),
    .B1(_02761_),
    .B2(_02870_),
    .ZN(_04799_));
 AOI221_X4 _29990_ (.A(_04260_),
    .B1(_02791_),
    .B2(_02725_),
    .C1(_02704_),
    .C2(_02795_),
    .ZN(_04800_));
 AND2_X1 _29991_ (.A1(_02846_),
    .A2(_02704_),
    .ZN(_04802_));
 AND3_X1 _29992_ (.A1(_02756_),
    .A2(_02845_),
    .A3(_02683_),
    .ZN(_04803_));
 NOR2_X1 _29993_ (.A1(_04802_),
    .A2(_04803_),
    .ZN(_04804_));
 AOI21_X1 _29994_ (.A(_03244_),
    .B1(_02739_),
    .B2(_02752_),
    .ZN(_04805_));
 AND4_X1 _29995_ (.A1(_04799_),
    .A2(_04800_),
    .A3(_04804_),
    .A4(_04805_),
    .ZN(_04806_));
 OAI21_X1 _29996_ (.A(_03309_),
    .B1(_03261_),
    .B2(_03608_),
    .ZN(_04807_));
 INV_X1 _29997_ (.A(_03230_),
    .ZN(_04808_));
 AOI21_X1 _29998_ (.A(_02769_),
    .B1(_03588_),
    .B2(_04808_),
    .ZN(_04809_));
 AND2_X1 _29999_ (.A1(_03248_),
    .A2(_02744_),
    .ZN(_04810_));
 NOR4_X1 _30000_ (.A1(_03285_),
    .A2(_04809_),
    .A3(_04536_),
    .A4(_04810_),
    .ZN(_04811_));
 OAI21_X1 _30001_ (.A(_02898_),
    .B1(_02895_),
    .B2(_02809_),
    .ZN(_04813_));
 AND2_X1 _30002_ (.A1(_02774_),
    .A2(_03595_),
    .ZN(_04814_));
 INV_X1 _30003_ (.A(_04814_),
    .ZN(_04815_));
 OAI21_X1 _30004_ (.A(_02806_),
    .B1(_02797_),
    .B2(_02753_),
    .ZN(_04816_));
 AND3_X1 _30005_ (.A1(_04815_),
    .A2(_03670_),
    .A3(_04816_),
    .ZN(_04817_));
 AND4_X1 _30006_ (.A1(_04807_),
    .A2(_04811_),
    .A3(_04813_),
    .A4(_04817_),
    .ZN(_04818_));
 AND4_X1 _30007_ (.A1(_04789_),
    .A2(_04798_),
    .A3(_04806_),
    .A4(_04818_),
    .ZN(_04819_));
 OAI211_X2 _30008_ (.A(_03298_),
    .B(_03299_),
    .C1(_03294_),
    .C2(_03214_),
    .ZN(_04820_));
 AND2_X1 _30009_ (.A1(_02690_),
    .A2(_02698_),
    .ZN(_04821_));
 OAI21_X1 _30010_ (.A(_02883_),
    .B1(_03253_),
    .B2(_04821_),
    .ZN(_04822_));
 NOR2_X1 _30011_ (.A1(_03592_),
    .A2(_03982_),
    .ZN(_04824_));
 INV_X1 _30012_ (.A(_04824_),
    .ZN(_04825_));
 OAI21_X1 _30013_ (.A(_02787_),
    .B1(_02749_),
    .B2(_03273_),
    .ZN(_04826_));
 NAND4_X1 _30014_ (.A1(_04822_),
    .A2(_03620_),
    .A3(_04825_),
    .A4(_04826_),
    .ZN(_04827_));
 AND3_X1 _30015_ (.A1(_02825_),
    .A2(_03233_),
    .A3(_02743_),
    .ZN(_04828_));
 AOI211_X4 _30016_ (.A(_04820_),
    .B(_04827_),
    .C1(_02740_),
    .C2(_04828_),
    .ZN(_04829_));
 NAND2_X1 _30017_ (.A1(_04819_),
    .A2(_04829_),
    .ZN(_04830_));
 XNOR2_X2 _30018_ (.A(_04773_),
    .B(_04830_),
    .ZN(_04831_));
 XNOR2_X2 _30019_ (.A(_04831_),
    .B(_17236_),
    .ZN(_04832_));
 MUX2_X2 _30020_ (.A(_04577_),
    .B(_04832_),
    .S(_01876_),
    .Z(_00714_));
 XOR2_X1 _30021_ (.A(_17237_),
    .B(_17108_),
    .Z(_04834_));
 XOR2_X1 _30022_ (.A(_02580_),
    .B(_04701_),
    .Z(_04835_));
 AOI21_X1 _30023_ (.A(_03664_),
    .B1(_02893_),
    .B2(_02770_),
    .ZN(_04836_));
 AOI21_X1 _30024_ (.A(_04836_),
    .B1(_02898_),
    .B2(_04821_),
    .ZN(_04837_));
 OAI221_X1 _30025_ (.A(_04837_),
    .B1(_02712_),
    .B2(_03983_),
    .C1(_03664_),
    .C2(_03623_),
    .ZN(_04838_));
 AOI21_X1 _30026_ (.A(_03268_),
    .B1(_04281_),
    .B2(_02901_),
    .ZN(_04839_));
 OR4_X2 _30027_ (.A1(_03985_),
    .A2(_04839_),
    .A3(_03662_),
    .A4(_04519_),
    .ZN(_04840_));
 INV_X1 _30028_ (.A(_04802_),
    .ZN(_04841_));
 NAND4_X1 _30029_ (.A1(_03655_),
    .A2(_02849_),
    .A3(_04841_),
    .A4(_04279_),
    .ZN(_04842_));
 OAI211_X2 _30030_ (.A(_02861_),
    .B(_16855_),
    .C1(_02857_),
    .C2(_02707_),
    .ZN(_04843_));
 OAI21_X1 _30031_ (.A(_02861_),
    .B1(_03595_),
    .B2(_02747_),
    .ZN(_04845_));
 OAI211_X2 _30032_ (.A(_04843_),
    .B(_04845_),
    .C1(_03252_),
    .C2(_03214_),
    .ZN(_04846_));
 NOR4_X2 _30033_ (.A1(_04838_),
    .A2(_04840_),
    .A3(_04842_),
    .A4(_04846_),
    .ZN(_04847_));
 AND2_X1 _30034_ (.A1(_02795_),
    .A2(_02781_),
    .ZN(_04848_));
 OAI21_X1 _30035_ (.A(_04563_),
    .B1(_03588_),
    .B2(_03592_),
    .ZN(_04849_));
 OAI211_X2 _30036_ (.A(_03601_),
    .B(_04312_),
    .C1(_04569_),
    .C2(_02698_),
    .ZN(_04850_));
 NAND2_X1 _30037_ (.A1(_02715_),
    .A2(_02799_),
    .ZN(_04851_));
 NAND2_X1 _30038_ (.A1(_02802_),
    .A2(_04851_),
    .ZN(_04852_));
 OR4_X4 _30039_ (.A1(_04848_),
    .A2(_04849_),
    .A3(_04850_),
    .A4(_04852_),
    .ZN(_04853_));
 AND2_X1 _30040_ (.A1(_02744_),
    .A2(_02719_),
    .ZN(_04854_));
 NAND2_X1 _30041_ (.A1(_02730_),
    .A2(_02744_),
    .ZN(_04856_));
 NAND3_X1 _30042_ (.A1(_04856_),
    .A2(_03587_),
    .A3(_02768_),
    .ZN(_04857_));
 AOI21_X1 _30043_ (.A(_02769_),
    .B1(_02779_),
    .B2(_02738_),
    .ZN(_04858_));
 NOR2_X1 _30044_ (.A1(_02769_),
    .A2(_03294_),
    .ZN(_04859_));
 OR4_X2 _30045_ (.A1(_04854_),
    .A2(_04857_),
    .A3(_04858_),
    .A4(_04859_),
    .ZN(_04860_));
 AND2_X1 _30046_ (.A1(_03222_),
    .A2(_03265_),
    .ZN(_04861_));
 NOR4_X4 _30047_ (.A1(_04853_),
    .A2(_04860_),
    .A3(_04861_),
    .A4(_04037_),
    .ZN(_04862_));
 INV_X1 _30048_ (.A(_03613_),
    .ZN(_04863_));
 NAND2_X1 _30049_ (.A1(_03309_),
    .A2(_03273_),
    .ZN(_04864_));
 NAND4_X1 _30050_ (.A1(_04863_),
    .A2(_04864_),
    .A3(_03312_),
    .A4(_04304_),
    .ZN(_04865_));
 AND2_X1 _30051_ (.A1(_02726_),
    .A2(_02831_),
    .ZN(_04867_));
 INV_X1 _30052_ (.A(_04867_),
    .ZN(_04868_));
 NAND2_X1 _30053_ (.A1(_02727_),
    .A2(_02719_),
    .ZN(_04869_));
 OAI211_X2 _30054_ (.A(_02724_),
    .B(_02773_),
    .C1(_03595_),
    .C2(_02747_),
    .ZN(_04870_));
 NAND4_X1 _30055_ (.A1(_04868_),
    .A2(_03313_),
    .A3(_04869_),
    .A4(_04870_),
    .ZN(_04871_));
 NAND2_X1 _30056_ (.A1(_02697_),
    .A2(_03301_),
    .ZN(_04872_));
 NAND4_X1 _30057_ (.A1(_02693_),
    .A2(_02711_),
    .A3(_02705_),
    .A4(_04872_),
    .ZN(_04873_));
 OAI21_X1 _30058_ (.A(_02787_),
    .B1(_02702_),
    .B2(_04821_),
    .ZN(_04874_));
 OAI21_X1 _30059_ (.A(_04874_),
    .B1(_03252_),
    .B2(_03611_),
    .ZN(_04875_));
 NOR4_X1 _30060_ (.A1(_04865_),
    .A2(_04871_),
    .A3(_04873_),
    .A4(_04875_),
    .ZN(_04876_));
 OAI21_X1 _30061_ (.A(_02868_),
    .B1(_02702_),
    .B2(_04821_),
    .ZN(_04878_));
 OAI21_X1 _30062_ (.A(_02868_),
    .B1(_03595_),
    .B2(_02848_),
    .ZN(_04879_));
 NAND4_X1 _30063_ (.A1(_02741_),
    .A2(_02812_),
    .A3(_02856_),
    .A4(_02817_),
    .ZN(_04880_));
 AND3_X1 _30064_ (.A1(_04878_),
    .A2(_04879_),
    .A3(_04880_),
    .ZN(_04881_));
 AOI21_X1 _30065_ (.A(_03634_),
    .B1(_04015_),
    .B2(_04808_),
    .ZN(_04882_));
 AOI21_X1 _30066_ (.A(_03634_),
    .B1(_02779_),
    .B2(_02738_),
    .ZN(_04883_));
 AOI211_X4 _30067_ (.A(_04882_),
    .B(_04883_),
    .C1(_02903_),
    .C2(_02823_),
    .ZN(_04884_));
 NAND2_X1 _30068_ (.A1(_02870_),
    .A2(_02829_),
    .ZN(_04885_));
 AND4_X1 _30069_ (.A1(_03974_),
    .A2(_02837_),
    .A3(_04885_),
    .A4(_04252_),
    .ZN(_04886_));
 OAI21_X1 _30070_ (.A(_02883_),
    .B1(_02710_),
    .B2(_02715_),
    .ZN(_04887_));
 OAI211_X2 _30071_ (.A(_02877_),
    .B(_02753_),
    .C1(_02856_),
    .C2(_02857_),
    .ZN(_04889_));
 AND3_X1 _30072_ (.A1(_04887_),
    .A2(_03642_),
    .A3(_04889_),
    .ZN(_04890_));
 AND4_X2 _30073_ (.A1(_04881_),
    .A2(_04884_),
    .A3(_04886_),
    .A4(_04890_),
    .ZN(_04891_));
 NAND4_X2 _30074_ (.A1(_04847_),
    .A2(_04862_),
    .A3(_04876_),
    .A4(_04891_),
    .ZN(_04892_));
 NOR2_X4 _30075_ (.A1(_04892_),
    .A2(_03267_),
    .ZN(_04893_));
 XNOR2_X1 _30076_ (.A(_04835_),
    .B(_04893_),
    .ZN(_04894_));
 NAND2_X1 _30077_ (.A1(_01938_),
    .A2(_02082_),
    .ZN(_04895_));
 OAI21_X1 _30078_ (.A(_01938_),
    .B1(_02090_),
    .B2(_02034_),
    .ZN(_04896_));
 AND4_X1 _30079_ (.A1(_04895_),
    .A2(_04896_),
    .A3(_03165_),
    .A4(_04064_),
    .ZN(_04897_));
 OAI211_X2 _30080_ (.A(_01916_),
    .B(_01972_),
    .C1(_02113_),
    .C2(_02106_),
    .ZN(_04898_));
 OAI21_X1 _30081_ (.A(_01960_),
    .B1(_01961_),
    .B2(_02077_),
    .ZN(_04900_));
 NAND4_X1 _30082_ (.A1(_04897_),
    .A2(_02091_),
    .A3(_04898_),
    .A4(_04900_),
    .ZN(_04901_));
 AND2_X1 _30083_ (.A1(_01941_),
    .A2(_02096_),
    .ZN(_04902_));
 AND2_X4 _30084_ (.A1(_03758_),
    .A2(_02096_),
    .ZN(_04903_));
 AOI211_X2 _30085_ (.A(_04902_),
    .B(_04903_),
    .C1(_01968_),
    .C2(_02097_),
    .ZN(_04904_));
 AND3_X1 _30086_ (.A1(_01994_),
    .A2(_01925_),
    .A3(_01918_),
    .ZN(_04905_));
 AOI211_X2 _30087_ (.A(_04905_),
    .B(_03180_),
    .C1(_02069_),
    .C2(_03758_),
    .ZN(_04906_));
 AND3_X1 _30088_ (.A1(_04492_),
    .A2(_04490_),
    .A3(_04068_),
    .ZN(_04907_));
 OAI21_X1 _30089_ (.A(_02069_),
    .B1(_01968_),
    .B2(_01967_),
    .ZN(_04908_));
 NAND4_X1 _30090_ (.A1(_04904_),
    .A2(_04906_),
    .A3(_04907_),
    .A4(_04908_),
    .ZN(_04909_));
 AND3_X1 _30091_ (.A1(_02063_),
    .A2(_01915_),
    .A3(_01918_),
    .ZN(_04911_));
 AOI211_X2 _30092_ (.A(_04911_),
    .B(_04053_),
    .C1(_02082_),
    .C2(_01920_),
    .ZN(_04912_));
 OAI21_X1 _30093_ (.A(_01920_),
    .B1(_03134_),
    .B2(_01967_),
    .ZN(_04913_));
 OAI21_X1 _30094_ (.A(_02013_),
    .B1(_02053_),
    .B2(_02090_),
    .ZN(_04914_));
 OAI21_X1 _30095_ (.A(_02013_),
    .B1(_02121_),
    .B2(_02026_),
    .ZN(_04915_));
 NAND4_X1 _30096_ (.A1(_04912_),
    .A2(_04913_),
    .A3(_04914_),
    .A4(_04915_),
    .ZN(_04916_));
 AND4_X2 _30097_ (.A1(_02041_),
    .A2(_02049_),
    .A3(_03570_),
    .A4(_03801_),
    .ZN(_04917_));
 OAI21_X1 _30098_ (.A(_01927_),
    .B1(_02122_),
    .B2(_02054_),
    .ZN(_04918_));
 OAI211_X2 _30099_ (.A(_01927_),
    .B(_01904_),
    .C1(_01908_),
    .C2(_01986_),
    .ZN(_04919_));
 NAND3_X2 _30100_ (.A1(_04917_),
    .A2(_04918_),
    .A3(_04919_),
    .ZN(_04920_));
 OR4_X4 _30101_ (.A1(_04901_),
    .A2(_04909_),
    .A3(_04916_),
    .A4(_04920_),
    .ZN(_04922_));
 NAND3_X1 _30102_ (.A1(_01995_),
    .A2(_02006_),
    .A3(_01990_),
    .ZN(_04923_));
 OAI21_X1 _30103_ (.A(_01991_),
    .B1(_01968_),
    .B2(_01914_),
    .ZN(_04924_));
 AND4_X1 _30104_ (.A1(_04923_),
    .A2(_04096_),
    .A3(_02003_),
    .A4(_04924_),
    .ZN(_04925_));
 OAI21_X1 _30105_ (.A(_02009_),
    .B1(_02071_),
    .B2(_02093_),
    .ZN(_04926_));
 OAI211_X2 _30106_ (.A(_02009_),
    .B(_02025_),
    .C1(_03161_),
    .C2(_02017_),
    .ZN(_04927_));
 AND4_X2 _30107_ (.A1(_04759_),
    .A2(_04925_),
    .A3(_04926_),
    .A4(_04927_),
    .ZN(_04928_));
 OAI21_X1 _30108_ (.A(_03195_),
    .B1(_01961_),
    .B2(_02054_),
    .ZN(_04929_));
 NAND2_X1 _30109_ (.A1(_01994_),
    .A2(_01980_),
    .ZN(_04930_));
 AND4_X1 _30110_ (.A1(_03747_),
    .A2(_03520_),
    .A3(_04930_),
    .A4(_04470_),
    .ZN(_04931_));
 AND2_X4 _30111_ (.A1(_02020_),
    .A2(_02093_),
    .ZN(_04933_));
 AND4_X1 _30112_ (.A1(_01924_),
    .A2(_01933_),
    .A3(_01907_),
    .A4(_01990_),
    .ZN(_04934_));
 NOR4_X2 _30113_ (.A1(_04466_),
    .A2(_03198_),
    .A3(_04933_),
    .A4(_04934_),
    .ZN(_04935_));
 OAI221_X1 _30114_ (.A(_01980_),
    .B1(_02022_),
    .B2(_01910_),
    .C1(_03517_),
    .C2(_01971_),
    .ZN(_04936_));
 AND4_X1 _30115_ (.A1(_04929_),
    .A2(_04931_),
    .A3(_04935_),
    .A4(_04936_),
    .ZN(_04937_));
 AND2_X1 _30116_ (.A1(_01999_),
    .A2(_01897_),
    .ZN(_04938_));
 INV_X1 _30117_ (.A(_04938_),
    .ZN(_04939_));
 OAI21_X1 _30118_ (.A(_02078_),
    .B1(_04447_),
    .B2(_03134_),
    .ZN(_04940_));
 OAI21_X1 _30119_ (.A(_01897_),
    .B1(_02033_),
    .B2(_01993_),
    .ZN(_04941_));
 OAI21_X1 _30120_ (.A(_02078_),
    .B1(_02112_),
    .B2(_02082_),
    .ZN(_04942_));
 AND4_X1 _30121_ (.A1(_04939_),
    .A2(_04940_),
    .A3(_04941_),
    .A4(_04942_),
    .ZN(_04944_));
 NOR2_X1 _30122_ (.A1(_03124_),
    .A2(_04459_),
    .ZN(_04945_));
 OAI221_X1 _30123_ (.A(_01966_),
    .B1(_02118_),
    .B2(_01910_),
    .C1(_02025_),
    .C2(_01971_),
    .ZN(_04946_));
 OAI21_X1 _30124_ (.A(_01984_),
    .B1(_01935_),
    .B2(_02113_),
    .ZN(_04947_));
 AND4_X1 _30125_ (.A1(_04945_),
    .A2(_04710_),
    .A3(_04946_),
    .A4(_04947_),
    .ZN(_04948_));
 NAND4_X4 _30126_ (.A1(_04928_),
    .A2(_04937_),
    .A3(_04944_),
    .A4(_04948_),
    .ZN(_04949_));
 NOR2_X4 _30127_ (.A1(_04922_),
    .A2(_04949_),
    .ZN(_04950_));
 OAI21_X1 _30128_ (.A(_02233_),
    .B1(_03884_),
    .B2(_02242_),
    .ZN(_04951_));
 AND4_X1 _30129_ (.A1(_02324_),
    .A2(_02143_),
    .A3(_02146_),
    .A4(_02223_),
    .ZN(_04952_));
 AND2_X2 _30130_ (.A1(_02225_),
    .A2(_02285_),
    .ZN(_04953_));
 AOI211_X2 _30131_ (.A(_04952_),
    .B(_04953_),
    .C1(_02225_),
    .C2(_03884_),
    .ZN(_04955_));
 OAI21_X1 _30132_ (.A(_02225_),
    .B1(_02206_),
    .B2(_02208_),
    .ZN(_04956_));
 OAI21_X1 _30133_ (.A(_02225_),
    .B1(_02257_),
    .B2(_02260_),
    .ZN(_04957_));
 AND4_X1 _30134_ (.A1(_04951_),
    .A2(_04955_),
    .A3(_04956_),
    .A4(_04957_),
    .ZN(_04958_));
 OAI21_X1 _30135_ (.A(_02290_),
    .B1(_03078_),
    .B2(_02257_),
    .ZN(_04959_));
 NAND4_X1 _30136_ (.A1(_02273_),
    .A2(_02324_),
    .A3(_02317_),
    .A4(_02135_),
    .ZN(_04960_));
 OAI21_X1 _30137_ (.A(_02290_),
    .B1(_02140_),
    .B2(_03096_),
    .ZN(_04961_));
 AND3_X1 _30138_ (.A1(_04959_),
    .A2(_04960_),
    .A3(_04961_),
    .ZN(_04962_));
 OAI21_X1 _30139_ (.A(_02275_),
    .B1(_02305_),
    .B2(_03081_),
    .ZN(_04963_));
 OAI21_X1 _30140_ (.A(_02275_),
    .B1(_02208_),
    .B2(_02192_),
    .ZN(_04964_));
 AND3_X1 _30141_ (.A1(_04962_),
    .A2(_04963_),
    .A3(_04964_),
    .ZN(_04966_));
 OAI21_X1 _30142_ (.A(_02301_),
    .B1(_02335_),
    .B2(_02250_),
    .ZN(_04967_));
 OAI211_X2 _30143_ (.A(_02179_),
    .B(_02278_),
    .C1(_02285_),
    .C2(_02230_),
    .ZN(_04968_));
 NAND3_X1 _30144_ (.A1(_04967_),
    .A2(_04968_),
    .A3(_03406_),
    .ZN(_04969_));
 NAND2_X1 _30145_ (.A1(_02341_),
    .A2(_02313_),
    .ZN(_04970_));
 NAND3_X1 _30146_ (.A1(_04970_),
    .A2(_03073_),
    .A3(_03074_),
    .ZN(_04971_));
 NOR4_X1 _30147_ (.A1(_04127_),
    .A2(_03072_),
    .A3(_04969_),
    .A4(_04971_),
    .ZN(_04972_));
 OAI21_X1 _30148_ (.A(_02262_),
    .B1(_02208_),
    .B2(_03871_),
    .ZN(_04973_));
 OAI21_X1 _30149_ (.A(_02246_),
    .B1(_03077_),
    .B2(_02153_),
    .ZN(_04974_));
 NOR2_X1 _30150_ (.A1(_02188_),
    .A2(_02169_),
    .ZN(_04975_));
 OAI21_X1 _30151_ (.A(_02246_),
    .B1(_02294_),
    .B2(_04975_),
    .ZN(_04977_));
 OAI211_X2 _30152_ (.A(_02262_),
    .B(_02212_),
    .C1(_02146_),
    .C2(_02237_),
    .ZN(_04978_));
 AND4_X1 _30153_ (.A1(_04973_),
    .A2(_04974_),
    .A3(_04977_),
    .A4(_04978_),
    .ZN(_04979_));
 NAND4_X1 _30154_ (.A1(_04958_),
    .A2(_04966_),
    .A3(_04972_),
    .A4(_04979_),
    .ZN(_04980_));
 NAND2_X1 _30155_ (.A1(_02238_),
    .A2(_02181_),
    .ZN(_04981_));
 NAND2_X1 _30156_ (.A1(_04975_),
    .A2(_02201_),
    .ZN(_04982_));
 AND4_X1 _30157_ (.A1(_03021_),
    .A2(_03835_),
    .A3(_04413_),
    .A4(_04982_),
    .ZN(_04983_));
 OAI21_X1 _30158_ (.A(_02181_),
    .B1(_02147_),
    .B2(_02285_),
    .ZN(_04984_));
 OAI211_X2 _30159_ (.A(_02167_),
    .B(_02181_),
    .C1(_03083_),
    .C2(_02219_),
    .ZN(_04985_));
 AND4_X1 _30160_ (.A1(_04981_),
    .A2(_04983_),
    .A3(_04984_),
    .A4(_04985_),
    .ZN(_04986_));
 AND2_X1 _30161_ (.A1(_04168_),
    .A2(_04169_),
    .ZN(_04988_));
 AND3_X1 _30162_ (.A1(_04629_),
    .A2(_03043_),
    .A3(_03365_),
    .ZN(_04989_));
 OAI21_X1 _30163_ (.A(_02176_),
    .B1(_02238_),
    .B2(_02359_),
    .ZN(_04990_));
 OAI21_X1 _30164_ (.A(_02134_),
    .B1(_03083_),
    .B2(_02320_),
    .ZN(_04991_));
 AND4_X1 _30165_ (.A1(_04988_),
    .A2(_04989_),
    .A3(_04990_),
    .A4(_04991_),
    .ZN(_04992_));
 NAND2_X1 _30166_ (.A1(_02352_),
    .A2(_02206_),
    .ZN(_04993_));
 AND3_X2 _30167_ (.A1(_02327_),
    .A2(_03083_),
    .A3(_02167_),
    .ZN(_04994_));
 AOI21_X2 _30168_ (.A(_04994_),
    .B1(_02328_),
    .B2(_03078_),
    .ZN(_04995_));
 OAI21_X1 _30169_ (.A(_02352_),
    .B1(_03371_),
    .B2(_02141_),
    .ZN(_04996_));
 OAI21_X1 _30170_ (.A(_02328_),
    .B1(_02294_),
    .B2(_03018_),
    .ZN(_04997_));
 AND4_X2 _30171_ (.A1(_04993_),
    .A2(_04995_),
    .A3(_04996_),
    .A4(_04997_),
    .ZN(_04999_));
 OAI21_X1 _30172_ (.A(_02331_),
    .B1(_03037_),
    .B2(_02206_),
    .ZN(_05000_));
 OAI21_X1 _30173_ (.A(_02331_),
    .B1(_02156_),
    .B2(_02260_),
    .ZN(_05001_));
 NAND3_X1 _30174_ (.A1(_05000_),
    .A2(_04616_),
    .A3(_05001_),
    .ZN(_05002_));
 NOR4_X4 _30175_ (.A1(_05002_),
    .A2(_04390_),
    .A3(_02343_),
    .A4(_04604_),
    .ZN(_05003_));
 NAND4_X2 _30176_ (.A1(_04986_),
    .A2(_04992_),
    .A3(_04999_),
    .A4(_05003_),
    .ZN(_05004_));
 NOR2_X2 _30177_ (.A1(_04980_),
    .A2(_05004_),
    .ZN(_05005_));
 INV_X4 _30178_ (.A(_05005_),
    .ZN(_05006_));
 XNOR2_X1 _30179_ (.A(_04950_),
    .B(_05006_),
    .ZN(_05007_));
 XNOR2_X1 _30180_ (.A(_04894_),
    .B(_05007_),
    .ZN(_05008_));
 XNOR2_X1 _30181_ (.A(_05008_),
    .B(_17237_),
    .ZN(_05010_));
 MUX2_X1 _30182_ (.A(_04834_),
    .B(_05010_),
    .S(_01876_),
    .Z(_00715_));
 XOR2_X1 _30183_ (.A(_17238_),
    .B(_17109_),
    .Z(_05011_));
 XNOR2_X1 _30184_ (.A(_04950_),
    .B(_01037_),
    .ZN(_05012_));
 XOR2_X1 _30185_ (.A(_05012_),
    .B(_03317_),
    .Z(_05013_));
 XNOR2_X1 _30186_ (.A(_02677_),
    .B(_02361_),
    .ZN(_05014_));
 XNOR2_X1 _30187_ (.A(_05013_),
    .B(_05014_),
    .ZN(_05015_));
 BUF_X4 _30188_ (.A(_09098_),
    .Z(_05016_));
 MUX2_X1 _30189_ (.A(_05011_),
    .B(_05015_),
    .S(_05016_),
    .Z(_00676_));
 XOR2_X1 _30190_ (.A(_17239_),
    .B(_17110_),
    .Z(_05017_));
 INV_X1 _30191_ (.A(_04950_),
    .ZN(_05019_));
 XNOR2_X2 _30192_ (.A(_05019_),
    .B(_02128_),
    .ZN(_05020_));
 XNOR2_X2 _30193_ (.A(_05020_),
    .B(_03671_),
    .ZN(_05021_));
 XNOR2_X1 _30194_ (.A(_03117_),
    .B(_03317_),
    .ZN(_05022_));
 XNOR2_X1 _30195_ (.A(_05021_),
    .B(_05022_),
    .ZN(_05023_));
 XOR2_X1 _30196_ (.A(_05023_),
    .B(_17239_),
    .Z(_05024_));
 MUX2_X1 _30197_ (.A(_05017_),
    .B(_05024_),
    .S(_05016_),
    .Z(_00677_));
 XOR2_X1 _30198_ (.A(_17209_),
    .B(_17111_),
    .Z(_05025_));
 XNOR2_X1 _30199_ (.A(_03504_),
    .B(_04045_),
    .ZN(_05026_));
 XOR2_X2 _30200_ (.A(_03671_),
    .B(_03212_),
    .Z(_05027_));
 XNOR2_X1 _30201_ (.A(_05026_),
    .B(_05027_),
    .ZN(_05029_));
 INV_X1 _30202_ (.A(_17209_),
    .ZN(_05030_));
 XNOR2_X1 _30203_ (.A(_05029_),
    .B(_05030_),
    .ZN(_05031_));
 MUX2_X1 _30204_ (.A(_05025_),
    .B(_05031_),
    .S(_05016_),
    .Z(_00678_));
 XOR2_X1 _30205_ (.A(_17210_),
    .B(_17112_),
    .Z(_05032_));
 XNOR2_X1 _30206_ (.A(_04950_),
    .B(_03577_),
    .ZN(_05033_));
 XNOR2_X1 _30207_ (.A(_05033_),
    .B(_04318_),
    .ZN(_05034_));
 XOR2_X1 _30208_ (.A(_05034_),
    .B(_04047_),
    .Z(_05035_));
 XNOR2_X1 _30209_ (.A(_05035_),
    .B(_17210_),
    .ZN(_05036_));
 MUX2_X1 _30210_ (.A(_05032_),
    .B(_05036_),
    .S(_05016_),
    .Z(_00679_));
 XOR2_X1 _30211_ (.A(_17211_),
    .B(_17113_),
    .Z(_05038_));
 XOR2_X2 _30212_ (.A(_04950_),
    .B(_03805_),
    .Z(_05039_));
 XNOR2_X1 _30213_ (.A(_05039_),
    .B(_04574_),
    .ZN(_05040_));
 XOR2_X1 _30214_ (.A(_05040_),
    .B(_04321_),
    .Z(_05041_));
 XOR2_X1 _30215_ (.A(_05041_),
    .B(_17211_),
    .Z(_05042_));
 MUX2_X1 _30216_ (.A(_05038_),
    .B(_05042_),
    .S(_05016_),
    .Z(_00680_));
 XOR2_X1 _30217_ (.A(_17212_),
    .B(_17114_),
    .Z(_05043_));
 XNOR2_X1 _30218_ (.A(_04574_),
    .B(_04108_),
    .ZN(_05044_));
 XNOR2_X1 _30219_ (.A(_04443_),
    .B(_05044_),
    .ZN(_05045_));
 XNOR2_X1 _30220_ (.A(_05045_),
    .B(_04830_),
    .ZN(_05046_));
 INV_X1 _30221_ (.A(_17212_),
    .ZN(_05048_));
 XNOR2_X1 _30222_ (.A(_05046_),
    .B(_05048_),
    .ZN(_05049_));
 MUX2_X1 _30223_ (.A(_05043_),
    .B(_05049_),
    .S(_05016_),
    .Z(_00681_));
 XOR2_X1 _30224_ (.A(_17213_),
    .B(_17115_),
    .Z(_05050_));
 XOR2_X1 _30225_ (.A(_04513_),
    .B(_04830_),
    .Z(_05051_));
 XNOR2_X2 _30226_ (.A(_04703_),
    .B(_05051_),
    .ZN(_05052_));
 XNOR2_X2 _30227_ (.A(_05052_),
    .B(_04893_),
    .ZN(_05053_));
 XNOR2_X2 _30228_ (.A(_05053_),
    .B(_17213_),
    .ZN(_05054_));
 MUX2_X2 _30229_ (.A(_05050_),
    .B(_05054_),
    .S(_05016_),
    .Z(_00682_));
 XOR2_X1 _30230_ (.A(_17214_),
    .B(_17116_),
    .Z(_05055_));
 XNOR2_X1 _30231_ (.A(_02580_),
    .B(_05006_),
    .ZN(_05057_));
 XOR2_X2 _30232_ (.A(_04771_),
    .B(_04893_),
    .Z(_05058_));
 XOR2_X1 _30233_ (.A(_05057_),
    .B(_05058_),
    .Z(_05059_));
 XNOR2_X1 _30234_ (.A(_05059_),
    .B(_02907_),
    .ZN(_05060_));
 XNOR2_X1 _30235_ (.A(_05060_),
    .B(_17214_),
    .ZN(_05061_));
 MUX2_X1 _30236_ (.A(_05055_),
    .B(_05061_),
    .S(_05016_),
    .Z(_00683_));
 XOR2_X1 _30237_ (.A(_17215_),
    .B(_17118_),
    .Z(_05062_));
 XNOR2_X1 _30238_ (.A(_05020_),
    .B(_01038_),
    .ZN(_05063_));
 XNOR2_X1 _30239_ (.A(_02677_),
    .B(_03316_),
    .ZN(_05064_));
 XNOR2_X1 _30240_ (.A(_05064_),
    .B(_05006_),
    .ZN(_05065_));
 XNOR2_X1 _30241_ (.A(_05063_),
    .B(_05065_),
    .ZN(_05067_));
 MUX2_X1 _30242_ (.A(_05062_),
    .B(_05067_),
    .S(_05016_),
    .Z(_00644_));
 XOR2_X1 _30243_ (.A(_17216_),
    .B(_17119_),
    .Z(_05068_));
 XNOR2_X1 _30244_ (.A(_05020_),
    .B(_05027_),
    .ZN(_05069_));
 XNOR2_X1 _30245_ (.A(_02361_),
    .B(_05006_),
    .ZN(_05070_));
 INV_X1 _30246_ (.A(_01039_),
    .ZN(_05071_));
 XNOR2_X1 _30247_ (.A(_03015_),
    .B(_05071_),
    .ZN(_05072_));
 XOR2_X1 _30248_ (.A(_05070_),
    .B(_05072_),
    .Z(_05073_));
 XNOR2_X1 _30249_ (.A(_05069_),
    .B(_05073_),
    .ZN(_05074_));
 MUX2_X1 _30250_ (.A(_05068_),
    .B(_05074_),
    .S(_05016_),
    .Z(_00645_));
 XNOR2_X1 _30251_ (.A(_03577_),
    .B(_03503_),
    .ZN(_05076_));
 XNOR2_X1 _30252_ (.A(_05076_),
    .B(_04045_),
    .ZN(_05077_));
 XNOR2_X1 _30253_ (.A(_03212_),
    .B(_03116_),
    .ZN(_05078_));
 OAI21_X1 _30254_ (.A(_09098_),
    .B1(_05077_),
    .B2(_05078_),
    .ZN(_05079_));
 AOI21_X1 _30255_ (.A(_05079_),
    .B1(_05077_),
    .B2(_05078_),
    .ZN(_05080_));
 AND2_X1 _30256_ (.A1(_01331_),
    .A2(_17120_),
    .ZN(_05081_));
 NOR2_X1 _30257_ (.A1(_05080_),
    .A2(_05081_),
    .ZN(_05082_));
 XNOR2_X1 _30258_ (.A(_05082_),
    .B(_17217_),
    .ZN(_00646_));
 XOR2_X1 _30259_ (.A(_17218_),
    .B(_17121_),
    .Z(_05083_));
 XNOR2_X1 _30260_ (.A(_03577_),
    .B(_04318_),
    .ZN(_05084_));
 XNOR2_X1 _30261_ (.A(_05039_),
    .B(_05084_),
    .ZN(_05086_));
 XNOR2_X1 _30262_ (.A(_03427_),
    .B(_05005_),
    .ZN(_05087_));
 XOR2_X1 _30263_ (.A(_05087_),
    .B(_03971_),
    .Z(_05088_));
 XNOR2_X1 _30264_ (.A(_05086_),
    .B(_05088_),
    .ZN(_05089_));
 XNOR2_X1 _30265_ (.A(_05089_),
    .B(_17218_),
    .ZN(_05090_));
 BUF_X4 _30266_ (.A(_09098_),
    .Z(_05091_));
 MUX2_X1 _30267_ (.A(_05083_),
    .B(_05090_),
    .S(_05091_),
    .Z(_00647_));
 XOR2_X1 _30268_ (.A(_17220_),
    .B(_17122_),
    .Z(_05092_));
 XNOR2_X1 _30269_ (.A(_05039_),
    .B(_04108_),
    .ZN(_05093_));
 XNOR2_X1 _30270_ (.A(_03892_),
    .B(_05006_),
    .ZN(_05094_));
 XOR2_X1 _30271_ (.A(_05094_),
    .B(_04246_),
    .Z(_05096_));
 XNOR2_X1 _30272_ (.A(_05093_),
    .B(_05096_),
    .ZN(_05097_));
 XNOR2_X1 _30273_ (.A(_05097_),
    .B(_04574_),
    .ZN(_05098_));
 XOR2_X1 _30274_ (.A(_05098_),
    .B(_17220_),
    .Z(_05099_));
 MUX2_X1 _30275_ (.A(_05092_),
    .B(_05099_),
    .S(_05091_),
    .Z(_00648_));
 XOR2_X1 _30276_ (.A(_17221_),
    .B(_17123_),
    .Z(_05100_));
 XOR2_X1 _30277_ (.A(_05051_),
    .B(_04178_),
    .Z(_05101_));
 INV_X1 _30278_ (.A(_01040_),
    .ZN(_05102_));
 XNOR2_X1 _30279_ (.A(_04380_),
    .B(_05102_),
    .ZN(_05103_));
 XNOR2_X1 _30280_ (.A(_05103_),
    .B(_04108_),
    .ZN(_05104_));
 XNOR2_X1 _30281_ (.A(_05101_),
    .B(_05104_),
    .ZN(_05106_));
 MUX2_X1 _30282_ (.A(_05100_),
    .B(_05106_),
    .S(_05091_),
    .Z(_00649_));
 XOR2_X1 _30283_ (.A(_17222_),
    .B(_17124_),
    .Z(_05107_));
 XNOR2_X1 _30284_ (.A(_04513_),
    .B(_01041_),
    .ZN(_05108_));
 XOR2_X1 _30285_ (.A(_05108_),
    .B(_04701_),
    .Z(_05109_));
 XNOR2_X1 _30286_ (.A(_05058_),
    .B(_04442_),
    .ZN(_05110_));
 XNOR2_X1 _30287_ (.A(_05109_),
    .B(_05110_),
    .ZN(_05111_));
 MUX2_X1 _30288_ (.A(_05107_),
    .B(_05111_),
    .S(_05091_),
    .Z(_00650_));
 XOR2_X1 _30289_ (.A(_17223_),
    .B(_17125_),
    .Z(_05112_));
 XNOR2_X1 _30290_ (.A(_04635_),
    .B(_02580_),
    .ZN(_05113_));
 XOR2_X1 _30291_ (.A(_04950_),
    .B(_04771_),
    .Z(_05115_));
 XNOR2_X1 _30292_ (.A(_05113_),
    .B(_05115_),
    .ZN(_05116_));
 XNOR2_X1 _30293_ (.A(_05116_),
    .B(_02907_),
    .ZN(_05117_));
 XNOR2_X1 _30294_ (.A(_05117_),
    .B(_17223_),
    .ZN(_05118_));
 MUX2_X1 _30295_ (.A(_05112_),
    .B(_05118_),
    .S(_05091_),
    .Z(_00651_));
 XOR2_X1 _30296_ (.A(_17224_),
    .B(_17126_),
    .Z(_05119_));
 XNOR2_X1 _30297_ (.A(_02361_),
    .B(_01042_),
    .ZN(_05120_));
 XNOR2_X1 _30298_ (.A(_05057_),
    .B(_05120_),
    .ZN(_05121_));
 XNOR2_X1 _30299_ (.A(_02128_),
    .B(_03316_),
    .ZN(_05122_));
 XNOR2_X1 _30300_ (.A(_05121_),
    .B(_05122_),
    .ZN(_05123_));
 MUX2_X1 _30301_ (.A(_05119_),
    .B(_05123_),
    .S(_05091_),
    .Z(_00612_));
 XOR2_X1 _30302_ (.A(_17225_),
    .B(_17127_),
    .Z(_05125_));
 XOR2_X1 _30303_ (.A(_02678_),
    .B(_05070_),
    .Z(_05126_));
 XNOR2_X2 _30304_ (.A(_05078_),
    .B(_03671_),
    .ZN(_05127_));
 XNOR2_X1 _30305_ (.A(_05126_),
    .B(_05127_),
    .ZN(_05128_));
 INV_X1 _30306_ (.A(_01043_),
    .ZN(_05129_));
 XNOR2_X1 _30307_ (.A(_05128_),
    .B(_05129_),
    .ZN(_05130_));
 MUX2_X1 _30308_ (.A(_05125_),
    .B(_05130_),
    .S(_05091_),
    .Z(_00613_));
 XOR2_X1 _30309_ (.A(_17226_),
    .B(_17129_),
    .Z(_05131_));
 XNOR2_X2 _30310_ (.A(_03577_),
    .B(_03427_),
    .ZN(_05132_));
 XNOR2_X1 _30311_ (.A(_03117_),
    .B(_05132_),
    .ZN(_05134_));
 XNOR2_X1 _30312_ (.A(_05134_),
    .B(_04045_),
    .ZN(_05135_));
 XNOR2_X1 _30313_ (.A(_05135_),
    .B(_17226_),
    .ZN(_05136_));
 MUX2_X1 _30314_ (.A(_05131_),
    .B(_05136_),
    .S(_05091_),
    .Z(_00614_));
 XOR2_X1 _30315_ (.A(_17227_),
    .B(_17130_),
    .Z(_05137_));
 XNOR2_X1 _30316_ (.A(_03892_),
    .B(_04318_),
    .ZN(_05138_));
 XNOR2_X1 _30317_ (.A(_03725_),
    .B(_05138_),
    .ZN(_05139_));
 XNOR2_X1 _30318_ (.A(_05087_),
    .B(_03805_),
    .ZN(_05140_));
 XNOR2_X1 _30319_ (.A(_05139_),
    .B(_05140_),
    .ZN(_05141_));
 XNOR2_X1 _30320_ (.A(_05141_),
    .B(_17227_),
    .ZN(_05142_));
 MUX2_X1 _30321_ (.A(_05137_),
    .B(_05142_),
    .S(_05091_),
    .Z(_00615_));
 XOR2_X1 _30322_ (.A(_17228_),
    .B(_17131_),
    .Z(_05144_));
 XNOR2_X1 _30323_ (.A(_04051_),
    .B(_05094_),
    .ZN(_05145_));
 XNOR2_X1 _30324_ (.A(_04178_),
    .B(_04108_),
    .ZN(_05146_));
 XNOR2_X1 _30325_ (.A(_05146_),
    .B(_04574_),
    .ZN(_05147_));
 XNOR2_X1 _30326_ (.A(_05145_),
    .B(_05147_),
    .ZN(_05148_));
 XNOR2_X1 _30327_ (.A(_05148_),
    .B(_17228_),
    .ZN(_05149_));
 MUX2_X1 _30328_ (.A(_05144_),
    .B(_05149_),
    .S(_05091_),
    .Z(_00616_));
 XOR2_X1 _30329_ (.A(_17229_),
    .B(_17132_),
    .Z(_05150_));
 XOR2_X1 _30330_ (.A(_04247_),
    .B(_04830_),
    .Z(_05151_));
 XOR2_X1 _30331_ (.A(_04442_),
    .B(_01044_),
    .Z(_05153_));
 XNOR2_X1 _30332_ (.A(_05153_),
    .B(_04513_),
    .ZN(_05154_));
 XNOR2_X1 _30333_ (.A(_05151_),
    .B(_05154_),
    .ZN(_05155_));
 BUF_X4 _30334_ (.A(_09098_),
    .Z(_05156_));
 MUX2_X1 _30335_ (.A(_05150_),
    .B(_05155_),
    .S(_05156_),
    .Z(_00617_));
 INV_X1 _30336_ (.A(_16755_),
    .ZN(_05157_));
 NOR2_X1 _30337_ (.A1(_01200_),
    .A2(_01201_),
    .ZN(_05158_));
 NOR2_X1 _30338_ (.A1(_01330_),
    .A2(_01199_),
    .ZN(_05159_));
 AOI221_X4 _30339_ (.A(_05157_),
    .B1(_03933_),
    .B2(_01198_),
    .C1(_05158_),
    .C2(_05159_),
    .ZN(_00599_));
 NOR3_X1 _30340_ (.A1(_01198_),
    .A2(_01199_),
    .A3(_01045_),
    .ZN(_05160_));
 INV_X1 _30341_ (.A(_05158_),
    .ZN(_05162_));
 NOR2_X1 _30342_ (.A1(_01198_),
    .A2(_01199_),
    .ZN(_05163_));
 AOI21_X1 _30343_ (.A(_05160_),
    .B1(_05162_),
    .B2(_05163_),
    .ZN(_05164_));
 AOI21_X1 _30344_ (.A(_03847_),
    .B1(_01198_),
    .B2(_01199_),
    .ZN(_05165_));
 AOI21_X1 _30345_ (.A(_05157_),
    .B1(_05164_),
    .B2(_05165_),
    .ZN(_00600_));
 AND2_X1 _30346_ (.A1(_05162_),
    .A2(_05163_),
    .ZN(_05166_));
 INV_X1 _30347_ (.A(_01046_),
    .ZN(_05167_));
 OAI211_X2 _30348_ (.A(_03749_),
    .B(_16755_),
    .C1(_05166_),
    .C2(_05167_),
    .ZN(_05168_));
 AOI21_X1 _30349_ (.A(_05168_),
    .B1(_05167_),
    .B2(_05166_),
    .ZN(_00601_));
 INV_X1 _30350_ (.A(_01200_),
    .ZN(_05169_));
 NAND3_X1 _30351_ (.A1(_05163_),
    .A2(_05169_),
    .A3(_01201_),
    .ZN(_05171_));
 INV_X1 _30352_ (.A(_01047_),
    .ZN(_05172_));
 OR2_X1 _30353_ (.A1(_05171_),
    .A2(_05172_),
    .ZN(_05173_));
 AOI21_X1 _30354_ (.A(_03847_),
    .B1(_05171_),
    .B2(_05172_),
    .ZN(_05174_));
 AOI21_X1 _30355_ (.A(_05157_),
    .B1(_05173_),
    .B2(_05174_),
    .ZN(_00602_));
 XOR2_X1 _30356_ (.A(_17231_),
    .B(_17133_),
    .Z(_05175_));
 XNOR2_X1 _30357_ (.A(_04893_),
    .B(_01048_),
    .ZN(_05176_));
 XNOR2_X1 _30358_ (.A(_04443_),
    .B(_05176_),
    .ZN(_05177_));
 XOR2_X1 _30359_ (.A(_04635_),
    .B(_04771_),
    .Z(_05178_));
 XNOR2_X1 _30360_ (.A(_05177_),
    .B(_05178_),
    .ZN(_05179_));
 MUX2_X1 _30361_ (.A(_05175_),
    .B(_05179_),
    .S(_05156_),
    .Z(_00618_));
 MUX2_X1 _30362_ (.A(_17012_),
    .B(_16884_),
    .S(_03847_),
    .Z(_00732_));
 BUF_X4 _30363_ (.A(_03836_),
    .Z(_05181_));
 MUX2_X1 _30364_ (.A(_17051_),
    .B(_16923_),
    .S(_05181_),
    .Z(_00771_));
 MUX2_X1 _30365_ (.A(_17062_),
    .B(_16934_),
    .S(_05181_),
    .Z(_00782_));
 MUX2_X1 _30366_ (.A(_17073_),
    .B(_16945_),
    .S(_05181_),
    .Z(_00793_));
 MUX2_X1 _30367_ (.A(_17084_),
    .B(_16956_),
    .S(_05181_),
    .Z(_00804_));
 MUX2_X1 _30368_ (.A(_17095_),
    .B(_16967_),
    .S(_05181_),
    .Z(_00815_));
 XOR2_X1 _30369_ (.A(_17232_),
    .B(_17134_),
    .Z(_05182_));
 XNOR2_X1 _30370_ (.A(_05007_),
    .B(_02907_),
    .ZN(_05183_));
 XOR2_X1 _30371_ (.A(_05183_),
    .B(_04703_),
    .Z(_05185_));
 XNOR2_X1 _30372_ (.A(_05185_),
    .B(_17232_),
    .ZN(_05186_));
 MUX2_X1 _30373_ (.A(_05182_),
    .B(_05186_),
    .S(_05156_),
    .Z(_00619_));
 MUX2_X1 _30374_ (.A(_17106_),
    .B(_16978_),
    .S(_05181_),
    .Z(_00826_));
 MUX2_X1 _30375_ (.A(_17117_),
    .B(_16989_),
    .S(_05181_),
    .Z(_00837_));
 MUX2_X1 _30376_ (.A(_17128_),
    .B(_17000_),
    .S(_05181_),
    .Z(_00848_));
 MUX2_X1 _30377_ (.A(_17139_),
    .B(_17011_),
    .S(_05181_),
    .Z(_00859_));
 MUX2_X1 _30378_ (.A(_17023_),
    .B(_16895_),
    .S(_05181_),
    .Z(_00743_));
 BUF_X4 _30379_ (.A(_03836_),
    .Z(_05187_));
 MUX2_X1 _30380_ (.A(_17034_),
    .B(_16906_),
    .S(_05187_),
    .Z(_00754_));
 MUX2_X1 _30381_ (.A(_17043_),
    .B(_16915_),
    .S(_05187_),
    .Z(_00763_));
 MUX2_X1 _30382_ (.A(_17044_),
    .B(_16916_),
    .S(_05187_),
    .Z(_00764_));
 MUX2_X1 _30383_ (.A(_17045_),
    .B(_16917_),
    .S(_05187_),
    .Z(_00765_));
 MUX2_X1 _30384_ (.A(_17046_),
    .B(_16918_),
    .S(_05187_),
    .Z(_00766_));
 MUX2_X1 _30385_ (.A(_17047_),
    .B(_16919_),
    .S(_05187_),
    .Z(_00767_));
 MUX2_X1 _30386_ (.A(_17048_),
    .B(_16920_),
    .S(_05187_),
    .Z(_00768_));
 MUX2_X1 _30387_ (.A(_17049_),
    .B(_16921_),
    .S(_05187_),
    .Z(_00769_));
 MUX2_X1 _30388_ (.A(_17050_),
    .B(_16922_),
    .S(_05187_),
    .Z(_00770_));
 MUX2_X1 _30389_ (.A(_17052_),
    .B(_16924_),
    .S(_05187_),
    .Z(_00772_));
 BUF_X8 _30390_ (.A(_01330_),
    .Z(_05189_));
 BUF_X4 _30391_ (.A(_05189_),
    .Z(_05191_));
 MUX2_X1 _30392_ (.A(_17053_),
    .B(_16925_),
    .S(_05191_),
    .Z(_00773_));
 MUX2_X1 _30393_ (.A(_17054_),
    .B(_16926_),
    .S(_05191_),
    .Z(_00774_));
 MUX2_X1 _30394_ (.A(_17055_),
    .B(_16927_),
    .S(_05191_),
    .Z(_00775_));
 MUX2_X1 _30395_ (.A(_17056_),
    .B(_16928_),
    .S(_05191_),
    .Z(_00776_));
 MUX2_X1 _30396_ (.A(_17057_),
    .B(_16929_),
    .S(_05191_),
    .Z(_00777_));
 MUX2_X1 _30397_ (.A(_17058_),
    .B(_16930_),
    .S(_05191_),
    .Z(_00778_));
 MUX2_X1 _30398_ (.A(_17059_),
    .B(_16931_),
    .S(_05191_),
    .Z(_00779_));
 MUX2_X1 _30399_ (.A(_17060_),
    .B(_16932_),
    .S(_05191_),
    .Z(_00780_));
 MUX2_X1 _30400_ (.A(_17061_),
    .B(_16933_),
    .S(_05191_),
    .Z(_00781_));
 MUX2_X1 _30401_ (.A(_17063_),
    .B(_16935_),
    .S(_05191_),
    .Z(_00783_));
 BUF_X4 _30402_ (.A(_05189_),
    .Z(_05193_));
 MUX2_X1 _30403_ (.A(_17064_),
    .B(_16936_),
    .S(_05193_),
    .Z(_00784_));
 MUX2_X1 _30404_ (.A(_17065_),
    .B(_16937_),
    .S(_05193_),
    .Z(_00785_));
 MUX2_X1 _30405_ (.A(_17066_),
    .B(_16938_),
    .S(_05193_),
    .Z(_00786_));
 MUX2_X1 _30406_ (.A(_17067_),
    .B(_16939_),
    .S(_05193_),
    .Z(_00787_));
 MUX2_X1 _30407_ (.A(_17068_),
    .B(_16940_),
    .S(_05193_),
    .Z(_00788_));
 MUX2_X1 _30408_ (.A(_17069_),
    .B(_16941_),
    .S(_05193_),
    .Z(_00789_));
 MUX2_X1 _30409_ (.A(_17070_),
    .B(_16942_),
    .S(_05193_),
    .Z(_00790_));
 MUX2_X1 _30410_ (.A(_17071_),
    .B(_16943_),
    .S(_05193_),
    .Z(_00791_));
 MUX2_X1 _30411_ (.A(_17072_),
    .B(_16944_),
    .S(_05193_),
    .Z(_00792_));
 MUX2_X1 _30412_ (.A(_17074_),
    .B(_16946_),
    .S(_05193_),
    .Z(_00794_));
 BUF_X4 _30413_ (.A(_05189_),
    .Z(_05195_));
 MUX2_X1 _30414_ (.A(_17075_),
    .B(_16947_),
    .S(_05195_),
    .Z(_00795_));
 MUX2_X1 _30415_ (.A(_17076_),
    .B(_16948_),
    .S(_05195_),
    .Z(_00796_));
 MUX2_X1 _30416_ (.A(_17077_),
    .B(_16949_),
    .S(_05195_),
    .Z(_00797_));
 MUX2_X1 _30417_ (.A(_17078_),
    .B(_16950_),
    .S(_05195_),
    .Z(_00798_));
 MUX2_X1 _30418_ (.A(_17079_),
    .B(_16951_),
    .S(_05195_),
    .Z(_00799_));
 MUX2_X1 _30419_ (.A(_17080_),
    .B(_16952_),
    .S(_05195_),
    .Z(_00800_));
 MUX2_X1 _30420_ (.A(_17081_),
    .B(_16953_),
    .S(_05195_),
    .Z(_00801_));
 MUX2_X1 _30421_ (.A(_17082_),
    .B(_16954_),
    .S(_05195_),
    .Z(_00802_));
 MUX2_X1 _30422_ (.A(_17083_),
    .B(_16955_),
    .S(_05195_),
    .Z(_00803_));
 MUX2_X1 _30423_ (.A(_17085_),
    .B(_16957_),
    .S(_05195_),
    .Z(_00805_));
 BUF_X4 _30424_ (.A(_05189_),
    .Z(_05197_));
 MUX2_X1 _30425_ (.A(_17086_),
    .B(_16958_),
    .S(_05197_),
    .Z(_00806_));
 MUX2_X1 _30426_ (.A(_17087_),
    .B(_16959_),
    .S(_05197_),
    .Z(_00807_));
 MUX2_X1 _30427_ (.A(_17088_),
    .B(_16960_),
    .S(_05197_),
    .Z(_00808_));
 MUX2_X1 _30428_ (.A(_17089_),
    .B(_16961_),
    .S(_05197_),
    .Z(_00809_));
 MUX2_X1 _30429_ (.A(_17090_),
    .B(_16962_),
    .S(_05197_),
    .Z(_00810_));
 MUX2_X1 _30430_ (.A(_17091_),
    .B(_16963_),
    .S(_05197_),
    .Z(_00811_));
 MUX2_X1 _30431_ (.A(_17092_),
    .B(_16964_),
    .S(_05197_),
    .Z(_00812_));
 MUX2_X1 _30432_ (.A(_17093_),
    .B(_16965_),
    .S(_05197_),
    .Z(_00813_));
 MUX2_X1 _30433_ (.A(_17094_),
    .B(_16966_),
    .S(_05197_),
    .Z(_00814_));
 MUX2_X1 _30434_ (.A(_17096_),
    .B(_16968_),
    .S(_05197_),
    .Z(_00816_));
 BUF_X4 _30435_ (.A(_05189_),
    .Z(_05199_));
 MUX2_X1 _30436_ (.A(_17097_),
    .B(_16969_),
    .S(_05199_),
    .Z(_00817_));
 MUX2_X1 _30437_ (.A(_17098_),
    .B(_16970_),
    .S(_05199_),
    .Z(_00818_));
 MUX2_X1 _30438_ (.A(_17099_),
    .B(_16971_),
    .S(_05199_),
    .Z(_00819_));
 MUX2_X1 _30439_ (.A(_17100_),
    .B(_16972_),
    .S(_05199_),
    .Z(_00820_));
 MUX2_X1 _30440_ (.A(_17101_),
    .B(_16973_),
    .S(_05199_),
    .Z(_00821_));
 MUX2_X1 _30441_ (.A(_17102_),
    .B(_16974_),
    .S(_05199_),
    .Z(_00822_));
 MUX2_X1 _30442_ (.A(_17103_),
    .B(_16975_),
    .S(_05199_),
    .Z(_00823_));
 MUX2_X1 _30443_ (.A(_17104_),
    .B(_16976_),
    .S(_05199_),
    .Z(_00824_));
 MUX2_X1 _30444_ (.A(_17105_),
    .B(_16977_),
    .S(_05199_),
    .Z(_00825_));
 MUX2_X1 _30445_ (.A(_17107_),
    .B(_16979_),
    .S(_05199_),
    .Z(_00827_));
 BUF_X4 _30446_ (.A(_05189_),
    .Z(_05201_));
 MUX2_X1 _30447_ (.A(_17108_),
    .B(_16980_),
    .S(_05201_),
    .Z(_00828_));
 MUX2_X1 _30448_ (.A(_17109_),
    .B(_16981_),
    .S(_05201_),
    .Z(_00829_));
 MUX2_X1 _30449_ (.A(_17110_),
    .B(_16982_),
    .S(_05201_),
    .Z(_00830_));
 MUX2_X1 _30450_ (.A(_17111_),
    .B(_16983_),
    .S(_05201_),
    .Z(_00831_));
 MUX2_X1 _30451_ (.A(_17112_),
    .B(_16984_),
    .S(_05201_),
    .Z(_00832_));
 MUX2_X1 _30452_ (.A(_17113_),
    .B(_16985_),
    .S(_05201_),
    .Z(_00833_));
 MUX2_X1 _30453_ (.A(_17114_),
    .B(_16986_),
    .S(_05201_),
    .Z(_00834_));
 MUX2_X1 _30454_ (.A(_17115_),
    .B(_16987_),
    .S(_05201_),
    .Z(_00835_));
 MUX2_X1 _30455_ (.A(_17116_),
    .B(_16988_),
    .S(_05201_),
    .Z(_00836_));
 MUX2_X1 _30456_ (.A(_17118_),
    .B(_16990_),
    .S(_05201_),
    .Z(_00838_));
 BUF_X4 _30457_ (.A(_05189_),
    .Z(_05203_));
 MUX2_X1 _30458_ (.A(_17119_),
    .B(_16991_),
    .S(_05203_),
    .Z(_00839_));
 MUX2_X1 _30459_ (.A(_17120_),
    .B(_16992_),
    .S(_05203_),
    .Z(_00840_));
 MUX2_X1 _30460_ (.A(_17121_),
    .B(_16993_),
    .S(_05203_),
    .Z(_00841_));
 MUX2_X1 _30461_ (.A(_17122_),
    .B(_16994_),
    .S(_05203_),
    .Z(_00842_));
 MUX2_X1 _30462_ (.A(_17123_),
    .B(_16995_),
    .S(_05203_),
    .Z(_00843_));
 MUX2_X1 _30463_ (.A(_17124_),
    .B(_16996_),
    .S(_05203_),
    .Z(_00844_));
 MUX2_X1 _30464_ (.A(_17125_),
    .B(_16997_),
    .S(_05203_),
    .Z(_00845_));
 MUX2_X1 _30465_ (.A(_17126_),
    .B(_16998_),
    .S(_05203_),
    .Z(_00846_));
 MUX2_X1 _30466_ (.A(_17127_),
    .B(_16999_),
    .S(_05203_),
    .Z(_00847_));
 MUX2_X1 _30467_ (.A(_17129_),
    .B(_17001_),
    .S(_05203_),
    .Z(_00849_));
 BUF_X4 _30468_ (.A(_05189_),
    .Z(_05205_));
 MUX2_X1 _30469_ (.A(_17130_),
    .B(_17002_),
    .S(_05205_),
    .Z(_00850_));
 MUX2_X1 _30470_ (.A(_17131_),
    .B(_17003_),
    .S(_05205_),
    .Z(_00851_));
 MUX2_X1 _30471_ (.A(_17132_),
    .B(_17004_),
    .S(_05205_),
    .Z(_00852_));
 MUX2_X1 _30472_ (.A(_17133_),
    .B(_17005_),
    .S(_05205_),
    .Z(_00853_));
 MUX2_X1 _30473_ (.A(_17134_),
    .B(_17006_),
    .S(_05205_),
    .Z(_00854_));
 XOR2_X1 _30474_ (.A(_17176_),
    .B(_17135_),
    .Z(_05207_));
 BUF_X32 _30475_ (.A(_16757_),
    .Z(_05208_));
 AND2_X4 _30476_ (.A1(_05208_),
    .A2(_16756_),
    .ZN(_05209_));
 AND2_X4 _30477_ (.A1(_16758_),
    .A2(_16759_),
    .ZN(_05210_));
 AND2_X2 _30478_ (.A1(_05209_),
    .A2(_05210_),
    .ZN(_05211_));
 AND2_X4 _30479_ (.A1(_16761_),
    .A2(_16760_),
    .ZN(_05212_));
 NOR2_X1 _30480_ (.A1(_16763_),
    .A2(_16762_),
    .ZN(_05213_));
 BUF_X2 _30481_ (.A(_05213_),
    .Z(_05215_));
 AND2_X2 _30482_ (.A1(_05212_),
    .A2(_05215_),
    .ZN(_05216_));
 AND2_X1 _30483_ (.A1(_05211_),
    .A2(_05216_),
    .ZN(_05217_));
 INV_X32 _30484_ (.A(_16759_),
    .ZN(_05218_));
 NOR2_X4 _30485_ (.A1(_05218_),
    .A2(_16758_),
    .ZN(_05219_));
 NOR2_X4 _30486_ (.A1(_05208_),
    .A2(_16756_),
    .ZN(_05220_));
 AND3_X1 _30487_ (.A1(_05216_),
    .A2(_05219_),
    .A3(_05220_),
    .ZN(_05221_));
 INV_X32 _30488_ (.A(_16757_),
    .ZN(_05222_));
 AND2_X4 _30489_ (.A1(_05210_),
    .A2(_05222_),
    .ZN(_05223_));
 BUF_X8 _30490_ (.A(_05223_),
    .Z(_05224_));
 AOI211_X2 _30491_ (.A(_05217_),
    .B(_05221_),
    .C1(_05224_),
    .C2(_05216_),
    .ZN(_05226_));
 AND2_X4 _30492_ (.A1(_05218_),
    .A2(_16758_),
    .ZN(_05227_));
 BUF_X8 _30493_ (.A(_05227_),
    .Z(_05228_));
 BUF_X4 _30494_ (.A(_05228_),
    .Z(_05229_));
 BUF_X4 _30495_ (.A(_05229_),
    .Z(_05230_));
 NOR2_X4 _30496_ (.A1(_05222_),
    .A2(_16756_),
    .ZN(_05231_));
 BUF_X4 _30497_ (.A(_05231_),
    .Z(_05232_));
 BUF_X2 _30498_ (.A(_05212_),
    .Z(_05233_));
 NAND4_X1 _30499_ (.A1(_05230_),
    .A2(_05232_),
    .A3(_05233_),
    .A4(_05215_),
    .ZN(_05234_));
 INV_X1 _30500_ (.A(_05216_),
    .ZN(_05235_));
 INV_X1 _30501_ (.A(_05220_),
    .ZN(_05237_));
 NOR2_X4 _30502_ (.A1(_16758_),
    .A2(_16759_),
    .ZN(_05238_));
 BUF_X2 _30503_ (.A(_05238_),
    .Z(_05239_));
 BUF_X4 _30504_ (.A(_05239_),
    .Z(_05240_));
 NAND2_X1 _30505_ (.A1(_05237_),
    .A2(_05240_),
    .ZN(_05241_));
 OAI211_X2 _30506_ (.A(_05226_),
    .B(_05234_),
    .C1(_05235_),
    .C2(_05241_),
    .ZN(_05242_));
 NOR2_X4 _30507_ (.A1(_16761_),
    .A2(_16760_),
    .ZN(_05243_));
 AND2_X1 _30508_ (.A1(_05243_),
    .A2(_05215_),
    .ZN(_05244_));
 BUF_X4 _30509_ (.A(_05244_),
    .Z(_05245_));
 BUF_X4 _30510_ (.A(_05208_),
    .Z(_05246_));
 BUF_X4 _30511_ (.A(_16756_),
    .Z(_05248_));
 OAI211_X2 _30512_ (.A(_05245_),
    .B(_05230_),
    .C1(_05246_),
    .C2(_05248_),
    .ZN(_05249_));
 BUF_X4 _30513_ (.A(_05219_),
    .Z(_05250_));
 OAI211_X2 _30514_ (.A(_05245_),
    .B(_05250_),
    .C1(_05246_),
    .C2(_05248_),
    .ZN(_05251_));
 BUF_X4 _30515_ (.A(_05210_),
    .Z(_05252_));
 INV_X4 _30516_ (.A(_16756_),
    .ZN(_05253_));
 NOR2_X4 _30517_ (.A1(_05253_),
    .A2(_05208_),
    .ZN(_05254_));
 BUF_X4 _30518_ (.A(_05254_),
    .Z(_05255_));
 OAI211_X2 _30519_ (.A(_05245_),
    .B(_05252_),
    .C1(_05232_),
    .C2(_05255_),
    .ZN(_05256_));
 AND2_X4 _30520_ (.A1(_05239_),
    .A2(_05208_),
    .ZN(_05257_));
 NAND2_X1 _30521_ (.A1(_05245_),
    .A2(_05257_),
    .ZN(_05259_));
 NAND4_X1 _30522_ (.A1(_05249_),
    .A2(_05251_),
    .A3(_05256_),
    .A4(_05259_),
    .ZN(_05260_));
 NOR3_X1 _30523_ (.A1(_05231_),
    .A2(_16758_),
    .A3(_05218_),
    .ZN(_05261_));
 INV_X1 _30524_ (.A(_05255_),
    .ZN(_05262_));
 AND2_X1 _30525_ (.A1(_05261_),
    .A2(_05262_),
    .ZN(_05263_));
 INV_X32 _30526_ (.A(_16760_),
    .ZN(_05264_));
 NOR2_X4 _30527_ (.A1(_05264_),
    .A2(_16761_),
    .ZN(_05265_));
 AND2_X1 _30528_ (.A1(_05265_),
    .A2(_05213_),
    .ZN(_05266_));
 BUF_X4 _30529_ (.A(_05266_),
    .Z(_05267_));
 NAND2_X1 _30530_ (.A1(_05263_),
    .A2(_05267_),
    .ZN(_05268_));
 BUF_X4 _30531_ (.A(_05267_),
    .Z(_05270_));
 NAND2_X1 _30532_ (.A1(_05270_),
    .A2(_05257_),
    .ZN(_05271_));
 BUF_X8 _30533_ (.A(_05209_),
    .Z(_05272_));
 INV_X1 _30534_ (.A(_05272_),
    .ZN(_05273_));
 NAND2_X1 _30535_ (.A1(_05273_),
    .A2(_05229_),
    .ZN(_05274_));
 BUF_X4 _30536_ (.A(_05220_),
    .Z(_05275_));
 NOR2_X1 _30537_ (.A1(_05274_),
    .A2(_05275_),
    .ZN(_05276_));
 INV_X1 _30538_ (.A(_05276_),
    .ZN(_05277_));
 INV_X2 _30539_ (.A(_05266_),
    .ZN(_05278_));
 OAI211_X2 _30540_ (.A(_05268_),
    .B(_05271_),
    .C1(_05277_),
    .C2(_05278_),
    .ZN(_05279_));
 AND2_X1 _30541_ (.A1(_05238_),
    .A2(_05222_),
    .ZN(_05281_));
 AND2_X4 _30542_ (.A1(_05264_),
    .A2(_16761_),
    .ZN(_05282_));
 BUF_X4 _30543_ (.A(_05282_),
    .Z(_05283_));
 NAND3_X1 _30544_ (.A1(_05281_),
    .A2(_05283_),
    .A3(_05215_),
    .ZN(_05284_));
 NAND4_X1 _30545_ (.A1(_05282_),
    .A2(_05231_),
    .A3(_05239_),
    .A4(_05215_),
    .ZN(_05285_));
 NAND2_X1 _30546_ (.A1(_05284_),
    .A2(_05285_),
    .ZN(_05286_));
 INV_X1 _30547_ (.A(_05286_),
    .ZN(_05287_));
 AND2_X1 _30548_ (.A1(_05282_),
    .A2(_05215_),
    .ZN(_05288_));
 BUF_X4 _30549_ (.A(_05288_),
    .Z(_05289_));
 AND2_X4 _30550_ (.A1(_05237_),
    .A2(_05219_),
    .ZN(_05290_));
 NAND2_X1 _30551_ (.A1(_05289_),
    .A2(_05290_),
    .ZN(_05292_));
 AND2_X1 _30552_ (.A1(_05229_),
    .A2(_05237_),
    .ZN(_05293_));
 NAND3_X1 _30553_ (.A1(_05293_),
    .A2(_05289_),
    .A3(_05273_),
    .ZN(_05294_));
 AND2_X2 _30554_ (.A1(_05210_),
    .A2(_05220_),
    .ZN(_05295_));
 BUF_X4 _30555_ (.A(_05295_),
    .Z(_05296_));
 AND2_X2 _30556_ (.A1(_05252_),
    .A2(_05208_),
    .ZN(_05297_));
 OAI21_X1 _30557_ (.A(_05289_),
    .B1(_05296_),
    .B2(_05297_),
    .ZN(_05298_));
 NAND4_X1 _30558_ (.A1(_05287_),
    .A2(_05292_),
    .A3(_05294_),
    .A4(_05298_),
    .ZN(_05299_));
 NOR4_X1 _30559_ (.A1(_05242_),
    .A2(_05260_),
    .A3(_05279_),
    .A4(_05299_),
    .ZN(_05300_));
 AND2_X4 _30560_ (.A1(_16763_),
    .A2(_16762_),
    .ZN(_05301_));
 BUF_X8 _30561_ (.A(_05301_),
    .Z(_05303_));
 AND2_X4 _30562_ (.A1(_05265_),
    .A2(_05303_),
    .ZN(_05304_));
 BUF_X8 _30563_ (.A(_05304_),
    .Z(_05305_));
 NAND3_X1 _30564_ (.A1(_05305_),
    .A2(_05255_),
    .A3(_05229_),
    .ZN(_05306_));
 AND2_X2 _30565_ (.A1(_05231_),
    .A2(_05238_),
    .ZN(_05307_));
 NAND2_X1 _30566_ (.A1(_05307_),
    .A2(_05305_),
    .ZN(_05308_));
 NAND2_X1 _30567_ (.A1(_05306_),
    .A2(_05308_),
    .ZN(_05309_));
 BUF_X4 _30568_ (.A(_05222_),
    .Z(_05310_));
 AND2_X2 _30569_ (.A1(_05219_),
    .A2(_05310_),
    .ZN(_05311_));
 NAND2_X2 _30570_ (.A1(_05311_),
    .A2(_05305_),
    .ZN(_05312_));
 AND2_X2 _30571_ (.A1(_05219_),
    .A2(_05208_),
    .ZN(_05314_));
 NAND2_X2 _30572_ (.A1(_05314_),
    .A2(_05305_),
    .ZN(_05315_));
 AND2_X2 _30573_ (.A1(_05231_),
    .A2(_05210_),
    .ZN(_05316_));
 AND2_X4 _30574_ (.A1(_05254_),
    .A2(_05210_),
    .ZN(_05317_));
 BUF_X4 _30575_ (.A(_05317_),
    .Z(_05318_));
 NOR2_X2 _30576_ (.A1(_05316_),
    .A2(_05318_),
    .ZN(_05319_));
 INV_X2 _30577_ (.A(_05305_),
    .ZN(_05320_));
 OAI211_X2 _30578_ (.A(_05312_),
    .B(_05315_),
    .C1(_05319_),
    .C2(_05320_),
    .ZN(_05321_));
 AND2_X4 _30579_ (.A1(_05303_),
    .A2(_05243_),
    .ZN(_05322_));
 NAND3_X1 _30580_ (.A1(_05322_),
    .A2(_05248_),
    .A3(_05250_),
    .ZN(_05323_));
 NAND2_X1 _30581_ (.A1(_05322_),
    .A2(_05224_),
    .ZN(_05325_));
 INV_X1 _30582_ (.A(_05316_),
    .ZN(_05326_));
 INV_X2 _30583_ (.A(_05322_),
    .ZN(_05327_));
 OAI211_X2 _30584_ (.A(_05323_),
    .B(_05325_),
    .C1(_05326_),
    .C2(_05327_),
    .ZN(_05328_));
 BUF_X4 _30585_ (.A(_05243_),
    .Z(_05329_));
 AND4_X1 _30586_ (.A1(_05231_),
    .A2(_05239_),
    .A3(_05329_),
    .A4(_05303_),
    .ZN(_05330_));
 OR4_X4 _30587_ (.A1(_05309_),
    .A2(_05321_),
    .A3(_05328_),
    .A4(_05330_),
    .ZN(_05331_));
 AND2_X4 _30588_ (.A1(_05282_),
    .A2(_05301_),
    .ZN(_05332_));
 BUF_X4 _30589_ (.A(_05332_),
    .Z(_05333_));
 AND2_X4 _30590_ (.A1(_05272_),
    .A2(_05238_),
    .ZN(_05334_));
 INV_X4 _30591_ (.A(_05334_),
    .ZN(_05336_));
 AND2_X2 _30592_ (.A1(_05220_),
    .A2(_05238_),
    .ZN(_05337_));
 INV_X1 _30593_ (.A(_05337_),
    .ZN(_05338_));
 NAND2_X2 _30594_ (.A1(_05336_),
    .A2(_05338_),
    .ZN(_05339_));
 AND2_X1 _30595_ (.A1(_05228_),
    .A2(_05310_),
    .ZN(_05340_));
 BUF_X2 _30596_ (.A(_05340_),
    .Z(_05341_));
 OAI21_X1 _30597_ (.A(_05333_),
    .B1(_05339_),
    .B2(_05341_),
    .ZN(_05342_));
 NAND3_X1 _30598_ (.A1(_05333_),
    .A2(_05250_),
    .A3(_05262_),
    .ZN(_05343_));
 INV_X1 _30599_ (.A(_05333_),
    .ZN(_05344_));
 AND2_X2 _30600_ (.A1(_05210_),
    .A2(_16756_),
    .ZN(_05345_));
 INV_X1 _30601_ (.A(_05345_),
    .ZN(_05347_));
 OAI211_X2 _30602_ (.A(_05342_),
    .B(_05343_),
    .C1(_05344_),
    .C2(_05347_),
    .ZN(_05348_));
 AND2_X2 _30603_ (.A1(_05228_),
    .A2(_05275_),
    .ZN(_05349_));
 AND2_X2 _30604_ (.A1(_05212_),
    .A2(_05301_),
    .ZN(_05350_));
 NAND2_X1 _30605_ (.A1(_05349_),
    .A2(_05350_),
    .ZN(_05351_));
 AND2_X2 _30606_ (.A1(_05254_),
    .A2(_05238_),
    .ZN(_05352_));
 BUF_X4 _30607_ (.A(_05352_),
    .Z(_05353_));
 BUF_X4 _30608_ (.A(_05350_),
    .Z(_05354_));
 NAND2_X1 _30609_ (.A1(_05353_),
    .A2(_05354_),
    .ZN(_05355_));
 BUF_X4 _30610_ (.A(_05257_),
    .Z(_05356_));
 NAND3_X1 _30611_ (.A1(_05356_),
    .A2(_05233_),
    .A3(_05303_),
    .ZN(_05358_));
 NAND3_X1 _30612_ (.A1(_05351_),
    .A2(_05355_),
    .A3(_05358_),
    .ZN(_05359_));
 BUF_X4 _30613_ (.A(_05314_),
    .Z(_05360_));
 NAND2_X1 _30614_ (.A1(_05360_),
    .A2(_05350_),
    .ZN(_05361_));
 NAND3_X1 _30615_ (.A1(_05350_),
    .A2(_05232_),
    .A3(_05252_),
    .ZN(_05362_));
 INV_X1 _30616_ (.A(_05311_),
    .ZN(_05363_));
 INV_X4 _30617_ (.A(_05350_),
    .ZN(_05364_));
 OAI211_X2 _30618_ (.A(_05361_),
    .B(_05362_),
    .C1(_05363_),
    .C2(_05364_),
    .ZN(_05365_));
 NOR4_X4 _30619_ (.A1(_05331_),
    .A2(_05348_),
    .A3(_05359_),
    .A4(_05365_),
    .ZN(_05366_));
 INV_X32 _30620_ (.A(_16763_),
    .ZN(_05367_));
 AND2_X2 _30621_ (.A1(_05367_),
    .A2(_16762_),
    .ZN(_05369_));
 AND2_X2 _30622_ (.A1(_05369_),
    .A2(_05212_),
    .ZN(_05370_));
 BUF_X4 _30623_ (.A(_05316_),
    .Z(_05371_));
 AND2_X4 _30624_ (.A1(_05219_),
    .A2(_05272_),
    .ZN(_05372_));
 BUF_X8 _30625_ (.A(_05372_),
    .Z(_05373_));
 OAI21_X1 _30626_ (.A(_05370_),
    .B1(_05371_),
    .B2(_05373_),
    .ZN(_05374_));
 BUF_X4 _30627_ (.A(_05370_),
    .Z(_05375_));
 NAND3_X1 _30628_ (.A1(_05375_),
    .A2(_05248_),
    .A3(_05224_),
    .ZN(_05376_));
 AND2_X1 _30629_ (.A1(_05374_),
    .A2(_05376_),
    .ZN(_05377_));
 BUF_X2 _30630_ (.A(_05334_),
    .Z(_05378_));
 NAND2_X1 _30631_ (.A1(_05375_),
    .A2(_05378_),
    .ZN(_05380_));
 AND2_X2 _30632_ (.A1(_05228_),
    .A2(_16756_),
    .ZN(_05381_));
 NAND2_X1 _30633_ (.A1(_05381_),
    .A2(_05375_),
    .ZN(_05382_));
 BUF_X2 _30634_ (.A(_05281_),
    .Z(_05383_));
 BUF_X4 _30635_ (.A(_05369_),
    .Z(_05384_));
 NAND3_X1 _30636_ (.A1(_05383_),
    .A2(_05384_),
    .A3(_05233_),
    .ZN(_05385_));
 NAND4_X1 _30637_ (.A1(_05377_),
    .A2(_05380_),
    .A3(_05382_),
    .A4(_05385_),
    .ZN(_05386_));
 AND2_X1 _30638_ (.A1(_05369_),
    .A2(_05329_),
    .ZN(_05387_));
 OAI21_X1 _30639_ (.A(_05387_),
    .B1(_05371_),
    .B2(_05224_),
    .ZN(_05388_));
 NAND4_X1 _30640_ (.A1(_05384_),
    .A2(_05250_),
    .A3(_05248_),
    .A4(_05329_),
    .ZN(_05389_));
 AND2_X1 _30641_ (.A1(_05388_),
    .A2(_05389_),
    .ZN(_05391_));
 BUF_X4 _30642_ (.A(_05387_),
    .Z(_05392_));
 OAI21_X1 _30643_ (.A(_05392_),
    .B1(_05349_),
    .B2(_05383_),
    .ZN(_05393_));
 AND2_X2 _30644_ (.A1(_05369_),
    .A2(_05265_),
    .ZN(_05394_));
 BUF_X2 _30645_ (.A(_05394_),
    .Z(_05395_));
 INV_X1 _30646_ (.A(_05231_),
    .ZN(_05396_));
 NAND2_X1 _30647_ (.A1(_05396_),
    .A2(_05239_),
    .ZN(_05397_));
 INV_X1 _30648_ (.A(_05397_),
    .ZN(_05398_));
 AND2_X4 _30649_ (.A1(_05228_),
    .A2(_05208_),
    .ZN(_05399_));
 OAI21_X1 _30650_ (.A(_05395_),
    .B1(_05398_),
    .B2(_05399_),
    .ZN(_05400_));
 AND2_X1 _30651_ (.A1(_05250_),
    .A2(_05248_),
    .ZN(_05402_));
 OAI21_X1 _30652_ (.A(_05395_),
    .B1(_05402_),
    .B2(_05211_),
    .ZN(_05403_));
 NAND4_X1 _30653_ (.A1(_05391_),
    .A2(_05393_),
    .A3(_05400_),
    .A4(_05403_),
    .ZN(_05404_));
 AND2_X2 _30654_ (.A1(_05282_),
    .A2(_05369_),
    .ZN(_05405_));
 INV_X1 _30655_ (.A(_05405_),
    .ZN(_05406_));
 AND2_X1 _30656_ (.A1(_05239_),
    .A2(_16756_),
    .ZN(_05407_));
 INV_X1 _30657_ (.A(_05407_),
    .ZN(_05408_));
 INV_X1 _30658_ (.A(_05230_),
    .ZN(_05409_));
 AOI21_X1 _30659_ (.A(_05406_),
    .B1(_05408_),
    .B2(_05409_),
    .ZN(_05410_));
 NAND2_X1 _30660_ (.A1(_05405_),
    .A2(_05261_),
    .ZN(_05411_));
 BUF_X4 _30661_ (.A(_05405_),
    .Z(_05413_));
 NAND2_X1 _30662_ (.A1(_05413_),
    .A2(_05371_),
    .ZN(_05414_));
 NAND2_X1 _30663_ (.A1(_05411_),
    .A2(_05414_),
    .ZN(_05415_));
 NOR4_X1 _30664_ (.A1(_05386_),
    .A2(_05404_),
    .A3(_05410_),
    .A4(_05415_),
    .ZN(_05416_));
 NOR2_X4 _30665_ (.A1(_05367_),
    .A2(_16762_),
    .ZN(_05417_));
 AND2_X2 _30666_ (.A1(_05265_),
    .A2(_05417_),
    .ZN(_05418_));
 BUF_X2 _30667_ (.A(_05418_),
    .Z(_05419_));
 INV_X1 _30668_ (.A(_05239_),
    .ZN(_05420_));
 NOR3_X1 _30669_ (.A1(_05420_),
    .A2(_05272_),
    .A3(_05275_),
    .ZN(_05421_));
 OAI21_X1 _30670_ (.A(_05419_),
    .B1(_05421_),
    .B2(_05297_),
    .ZN(_05422_));
 AND2_X1 _30671_ (.A1(_05282_),
    .A2(_05417_),
    .ZN(_05424_));
 OAI21_X1 _30672_ (.A(_05424_),
    .B1(_05211_),
    .B2(_05224_),
    .ZN(_05425_));
 NAND4_X1 _30673_ (.A1(_05282_),
    .A2(_05250_),
    .A3(_05255_),
    .A4(_05417_),
    .ZN(_05426_));
 INV_X1 _30674_ (.A(_05349_),
    .ZN(_05427_));
 INV_X1 _30675_ (.A(_05424_),
    .ZN(_05428_));
 OAI211_X2 _30676_ (.A(_05425_),
    .B(_05426_),
    .C1(_05427_),
    .C2(_05428_),
    .ZN(_05429_));
 AND2_X2 _30677_ (.A1(_05417_),
    .A2(_05212_),
    .ZN(_05430_));
 INV_X2 _30678_ (.A(_05430_),
    .ZN(_05431_));
 NAND2_X1 _30679_ (.A1(_05396_),
    .A2(_05228_),
    .ZN(_05432_));
 NOR2_X1 _30680_ (.A1(_05431_),
    .A2(_05432_),
    .ZN(_05433_));
 NOR2_X2 _30681_ (.A1(_05420_),
    .A2(_05255_),
    .ZN(_05435_));
 AND2_X1 _30682_ (.A1(_05430_),
    .A2(_05435_),
    .ZN(_05436_));
 AND3_X1 _30683_ (.A1(_05295_),
    .A2(_05212_),
    .A3(_05417_),
    .ZN(_05437_));
 NOR4_X1 _30684_ (.A1(_05429_),
    .A2(_05433_),
    .A3(_05436_),
    .A4(_05437_),
    .ZN(_05438_));
 AND2_X2 _30685_ (.A1(_05417_),
    .A2(_05243_),
    .ZN(_05439_));
 NAND3_X1 _30686_ (.A1(_05439_),
    .A2(_05310_),
    .A3(_05229_),
    .ZN(_05440_));
 BUF_X2 _30687_ (.A(_05417_),
    .Z(_05441_));
 NAND4_X1 _30688_ (.A1(_05229_),
    .A2(_05272_),
    .A3(_05441_),
    .A4(_05329_),
    .ZN(_05442_));
 NAND2_X1 _30689_ (.A1(_05440_),
    .A2(_05442_),
    .ZN(_05443_));
 BUF_X2 _30690_ (.A(_05439_),
    .Z(_05444_));
 BUF_X4 _30691_ (.A(_05253_),
    .Z(_05446_));
 AND2_X1 _30692_ (.A1(_05240_),
    .A2(_05446_),
    .ZN(_05447_));
 AOI21_X1 _30693_ (.A(_05443_),
    .B1(_05444_),
    .B2(_05447_),
    .ZN(_05448_));
 OAI21_X1 _30694_ (.A(_05210_),
    .B1(_05208_),
    .B2(_16756_),
    .ZN(_05449_));
 INV_X1 _30695_ (.A(_05449_),
    .ZN(_05450_));
 OAI21_X1 _30696_ (.A(_05444_),
    .B1(_05450_),
    .B2(_05402_),
    .ZN(_05451_));
 AND4_X1 _30697_ (.A1(_05422_),
    .A2(_05438_),
    .A3(_05448_),
    .A4(_05451_),
    .ZN(_05452_));
 AND4_X2 _30698_ (.A1(_05300_),
    .A2(_05366_),
    .A3(_05416_),
    .A4(_05452_),
    .ZN(_05453_));
 AND2_X1 _30699_ (.A1(_05337_),
    .A2(_05245_),
    .ZN(_05454_));
 INV_X1 _30700_ (.A(_05454_),
    .ZN(_05455_));
 NAND2_X2 _30701_ (.A1(_05453_),
    .A2(_05455_),
    .ZN(_05457_));
 INV_X4 _30702_ (.A(_05211_),
    .ZN(_05458_));
 INV_X1 _30703_ (.A(_05295_),
    .ZN(_05459_));
 NAND2_X2 _30704_ (.A1(_05458_),
    .A2(_05459_),
    .ZN(_05460_));
 AND2_X1 _30705_ (.A1(_05460_),
    .A2(_05333_),
    .ZN(_05461_));
 NAND2_X1 _30706_ (.A1(_05381_),
    .A2(_05332_),
    .ZN(_05462_));
 INV_X1 _30707_ (.A(_05281_),
    .ZN(_05463_));
 OAI21_X1 _30708_ (.A(_05462_),
    .B1(_05344_),
    .B2(_05463_),
    .ZN(_05464_));
 AND2_X1 _30709_ (.A1(_05311_),
    .A2(_05322_),
    .ZN(_05465_));
 AND2_X1 _30710_ (.A1(_05439_),
    .A2(_05311_),
    .ZN(_05466_));
 OR4_X4 _30711_ (.A1(_05461_),
    .A2(_05464_),
    .A3(_05465_),
    .A4(_05466_),
    .ZN(_05468_));
 AND2_X1 _30712_ (.A1(_05399_),
    .A2(_05289_),
    .ZN(_05469_));
 NAND2_X1 _30713_ (.A1(_05339_),
    .A2(_05439_),
    .ZN(_05470_));
 AND2_X1 _30714_ (.A1(_05297_),
    .A2(_05322_),
    .ZN(_05471_));
 INV_X1 _30715_ (.A(_05471_),
    .ZN(_05472_));
 AND2_X2 _30716_ (.A1(_05228_),
    .A2(_05231_),
    .ZN(_05473_));
 NAND2_X1 _30717_ (.A1(_05473_),
    .A2(_05305_),
    .ZN(_05474_));
 NAND4_X4 _30718_ (.A1(_05470_),
    .A2(_05472_),
    .A3(_05308_),
    .A4(_05474_),
    .ZN(_05475_));
 NAND2_X1 _30719_ (.A1(_05267_),
    .A2(_05281_),
    .ZN(_05476_));
 OAI21_X1 _30720_ (.A(_05476_),
    .B1(_05363_),
    .B2(_05278_),
    .ZN(_05477_));
 NOR4_X4 _30721_ (.A1(_05468_),
    .A2(_05469_),
    .A3(_05475_),
    .A4(_05477_),
    .ZN(_05479_));
 AND2_X4 _30722_ (.A1(_05290_),
    .A2(_05273_),
    .ZN(_05480_));
 AND2_X1 _30723_ (.A1(_05480_),
    .A2(_05418_),
    .ZN(_05481_));
 INV_X1 _30724_ (.A(_05418_),
    .ZN(_05482_));
 INV_X1 _30725_ (.A(_05399_),
    .ZN(_05483_));
 AOI21_X1 _30726_ (.A(_05482_),
    .B1(_05483_),
    .B2(_05408_),
    .ZN(_05484_));
 AOI21_X1 _30727_ (.A(_05482_),
    .B1(_05458_),
    .B2(_05459_),
    .ZN(_05485_));
 AND3_X1 _30728_ (.A1(_05224_),
    .A2(_05441_),
    .A3(_05283_),
    .ZN(_05486_));
 NOR4_X1 _30729_ (.A1(_05481_),
    .A2(_05484_),
    .A3(_05485_),
    .A4(_05486_),
    .ZN(_05487_));
 OAI21_X1 _30730_ (.A(_05394_),
    .B1(_05480_),
    .B2(_05211_),
    .ZN(_05488_));
 NAND4_X1 _30731_ (.A1(_05384_),
    .A2(_05265_),
    .A3(_05248_),
    .A4(_05239_),
    .ZN(_05490_));
 OAI211_X2 _30732_ (.A(_05394_),
    .B(_05229_),
    .C1(_05232_),
    .C2(_05255_),
    .ZN(_05491_));
 AND3_X1 _30733_ (.A1(_05488_),
    .A2(_05490_),
    .A3(_05491_),
    .ZN(_05492_));
 AND2_X4 _30734_ (.A1(_05228_),
    .A2(_05272_),
    .ZN(_05493_));
 OAI21_X1 _30735_ (.A(_05392_),
    .B1(_05493_),
    .B2(_05352_),
    .ZN(_05494_));
 OAI21_X1 _30736_ (.A(_05387_),
    .B1(_05360_),
    .B2(_05345_),
    .ZN(_05495_));
 BUF_X4 _30737_ (.A(_05424_),
    .Z(_05496_));
 BUF_X2 _30738_ (.A(_05311_),
    .Z(_05497_));
 BUF_X2 _30739_ (.A(_05430_),
    .Z(_05498_));
 AOI22_X1 _30740_ (.A1(_05496_),
    .A2(_05497_),
    .B1(_05498_),
    .B2(_05281_),
    .ZN(_05499_));
 AND4_X1 _30741_ (.A1(_05492_),
    .A2(_05494_),
    .A3(_05495_),
    .A4(_05499_),
    .ZN(_05501_));
 NOR2_X1 _30742_ (.A1(_05432_),
    .A2(_05255_),
    .ZN(_05502_));
 AND2_X1 _30743_ (.A1(_05502_),
    .A2(_05267_),
    .ZN(_05503_));
 INV_X1 _30744_ (.A(_05340_),
    .ZN(_05504_));
 OAI22_X1 _30745_ (.A1(_05504_),
    .A2(_05364_),
    .B1(_05408_),
    .B2(_05235_),
    .ZN(_05505_));
 AND2_X1 _30746_ (.A1(_05381_),
    .A2(_05216_),
    .ZN(_05506_));
 AND2_X1 _30747_ (.A1(_05252_),
    .A2(_05446_),
    .ZN(_05507_));
 AND2_X1 _30748_ (.A1(_05350_),
    .A2(_05507_),
    .ZN(_05508_));
 NOR4_X1 _30749_ (.A1(_05503_),
    .A2(_05505_),
    .A3(_05506_),
    .A4(_05508_),
    .ZN(_05509_));
 NAND4_X2 _30750_ (.A1(_05479_),
    .A2(_05487_),
    .A3(_05501_),
    .A4(_05509_),
    .ZN(_05510_));
 NAND2_X1 _30751_ (.A1(_05413_),
    .A2(_05240_),
    .ZN(_05512_));
 AND2_X1 _30752_ (.A1(_05314_),
    .A2(_05266_),
    .ZN(_05513_));
 INV_X1 _30753_ (.A(_05307_),
    .ZN(_05514_));
 AOI21_X1 _30754_ (.A(_05278_),
    .B1(_05458_),
    .B2(_05514_),
    .ZN(_05515_));
 AOI211_X2 _30755_ (.A(_05513_),
    .B(_05515_),
    .C1(_05267_),
    .C2(_05224_),
    .ZN(_05516_));
 BUF_X4 _30756_ (.A(_05224_),
    .Z(_05517_));
 NAND2_X1 _30757_ (.A1(_05517_),
    .A2(_05245_),
    .ZN(_05518_));
 AOI22_X1 _30758_ (.A1(_05341_),
    .A2(_05375_),
    .B1(_05405_),
    .B2(_05297_),
    .ZN(_05519_));
 AND4_X1 _30759_ (.A1(_05512_),
    .A2(_05516_),
    .A3(_05518_),
    .A4(_05519_),
    .ZN(_05520_));
 AND2_X2 _30760_ (.A1(_05219_),
    .A2(_05231_),
    .ZN(_05521_));
 AND2_X1 _30761_ (.A1(_05370_),
    .A2(_05521_),
    .ZN(_05523_));
 INV_X1 _30762_ (.A(_05523_),
    .ZN(_05524_));
 NAND2_X1 _30763_ (.A1(_05316_),
    .A2(_05430_),
    .ZN(_05525_));
 NAND2_X1 _30764_ (.A1(_05314_),
    .A2(_05430_),
    .ZN(_05526_));
 NAND2_X1 _30765_ (.A1(_05525_),
    .A2(_05526_),
    .ZN(_05527_));
 NOR2_X1 _30766_ (.A1(_05345_),
    .A2(_05224_),
    .ZN(_05528_));
 INV_X1 _30767_ (.A(_05528_),
    .ZN(_05529_));
 AOI211_X2 _30768_ (.A(_05433_),
    .B(_05527_),
    .C1(_05305_),
    .C2(_05529_),
    .ZN(_05530_));
 AND2_X1 _30769_ (.A1(_05370_),
    .A2(_05311_),
    .ZN(_05531_));
 INV_X1 _30770_ (.A(_05531_),
    .ZN(_05532_));
 AND4_X1 _30771_ (.A1(_05524_),
    .A2(_05530_),
    .A3(_05532_),
    .A4(_05287_),
    .ZN(_05534_));
 AND2_X1 _30772_ (.A1(_05424_),
    .A2(_05521_),
    .ZN(_05535_));
 INV_X1 _30773_ (.A(_05535_),
    .ZN(_05536_));
 NAND3_X1 _30774_ (.A1(_05439_),
    .A2(_05255_),
    .A3(_05229_),
    .ZN(_05537_));
 NAND2_X1 _30775_ (.A1(_05373_),
    .A2(_05305_),
    .ZN(_05538_));
 NAND4_X1 _30776_ (.A1(_05283_),
    .A2(_05218_),
    .A3(_05232_),
    .A4(_05303_),
    .ZN(_05539_));
 NAND4_X1 _30777_ (.A1(_05536_),
    .A2(_05537_),
    .A3(_05538_),
    .A4(_05539_),
    .ZN(_05540_));
 AND2_X2 _30778_ (.A1(_05219_),
    .A2(_05255_),
    .ZN(_05541_));
 AND2_X1 _30779_ (.A1(_05541_),
    .A2(_05350_),
    .ZN(_05542_));
 INV_X1 _30780_ (.A(_05542_),
    .ZN(_05543_));
 NAND2_X1 _30781_ (.A1(_05405_),
    .A2(_05541_),
    .ZN(_05545_));
 NAND3_X1 _30782_ (.A1(_05350_),
    .A2(_05273_),
    .A3(_05239_),
    .ZN(_05546_));
 NAND2_X1 _30783_ (.A1(_05289_),
    .A2(_05318_),
    .ZN(_05547_));
 NAND4_X1 _30784_ (.A1(_05543_),
    .A2(_05545_),
    .A3(_05546_),
    .A4(_05547_),
    .ZN(_05548_));
 NAND3_X1 _30785_ (.A1(_05371_),
    .A2(_05441_),
    .A3(_05283_),
    .ZN(_05549_));
 INV_X1 _30786_ (.A(_05318_),
    .ZN(_05550_));
 OAI221_X1 _30787_ (.A(_05549_),
    .B1(_05550_),
    .B2(_05327_),
    .C1(_05428_),
    .C2(_05338_),
    .ZN(_05551_));
 NAND2_X2 _30788_ (.A1(_05405_),
    .A2(_05493_),
    .ZN(_05552_));
 NAND2_X1 _30789_ (.A1(_05370_),
    .A2(_05407_),
    .ZN(_05553_));
 INV_X1 _30790_ (.A(_05493_),
    .ZN(_05554_));
 INV_X1 _30791_ (.A(_05370_),
    .ZN(_05556_));
 OAI211_X2 _30792_ (.A(_05552_),
    .B(_05553_),
    .C1(_05554_),
    .C2(_05556_),
    .ZN(_05557_));
 NOR4_X1 _30793_ (.A1(_05540_),
    .A2(_05548_),
    .A3(_05551_),
    .A4(_05557_),
    .ZN(_05558_));
 AND2_X1 _30794_ (.A1(_05343_),
    .A2(_05292_),
    .ZN(_05559_));
 OAI21_X1 _30795_ (.A(_05244_),
    .B1(_05502_),
    .B2(_05371_),
    .ZN(_05560_));
 AND2_X1 _30796_ (.A1(_05370_),
    .A2(_05450_),
    .ZN(_05561_));
 INV_X1 _30797_ (.A(_05561_),
    .ZN(_05562_));
 AND2_X1 _30798_ (.A1(_05560_),
    .A2(_05562_),
    .ZN(_05563_));
 BUF_X4 _30799_ (.A(_05322_),
    .Z(_05564_));
 OAI21_X1 _30800_ (.A(_05564_),
    .B1(_05293_),
    .B2(_05337_),
    .ZN(_05565_));
 OAI21_X1 _30801_ (.A(_05216_),
    .B1(_05314_),
    .B2(_05507_),
    .ZN(_05567_));
 AND4_X1 _30802_ (.A1(_05559_),
    .A2(_05563_),
    .A3(_05565_),
    .A4(_05567_),
    .ZN(_05568_));
 NAND4_X1 _30803_ (.A1(_05520_),
    .A2(_05534_),
    .A3(_05558_),
    .A4(_05568_),
    .ZN(_05569_));
 NOR2_X4 _30804_ (.A1(_05510_),
    .A2(_05569_),
    .ZN(_05570_));
 XOR2_X1 _30805_ (.A(_05457_),
    .B(_05570_),
    .Z(_05571_));
 INV_X1 _30806_ (.A(_16802_),
    .ZN(_05572_));
 NOR2_X2 _30807_ (.A1(_05572_),
    .A2(_16803_),
    .ZN(_05573_));
 NOR2_X1 _30808_ (.A1(_16801_),
    .A2(_16800_),
    .ZN(_05574_));
 AND2_X1 _30809_ (.A1(_05573_),
    .A2(_05574_),
    .ZN(_05575_));
 BUF_X2 _30810_ (.A(_05575_),
    .Z(_05576_));
 BUF_X32 _30811_ (.A(_16798_),
    .Z(_05578_));
 BUF_X32 _30812_ (.A(_16799_),
    .Z(_05579_));
 NOR2_X4 _30813_ (.A1(_05578_),
    .A2(_05579_),
    .ZN(_05580_));
 BUF_X8 _30814_ (.A(_05580_),
    .Z(_05581_));
 INV_X32 _30815_ (.A(_16797_),
    .ZN(_05582_));
 AND2_X2 _30816_ (.A1(_05581_),
    .A2(_05582_),
    .ZN(_05583_));
 INV_X1 _30817_ (.A(_05583_),
    .ZN(_05584_));
 INV_X8 _30818_ (.A(_16798_),
    .ZN(_05585_));
 NOR2_X4 _30819_ (.A1(_05585_),
    .A2(_05579_),
    .ZN(_05586_));
 BUF_X8 _30820_ (.A(_05586_),
    .Z(_05587_));
 BUF_X2 _30821_ (.A(_05587_),
    .Z(_05589_));
 INV_X1 _30822_ (.A(_05589_),
    .ZN(_05590_));
 NOR2_X4 _30823_ (.A1(_16797_),
    .A2(_16796_),
    .ZN(_05591_));
 INV_X4 _30824_ (.A(_05591_),
    .ZN(_05592_));
 OAI21_X1 _30825_ (.A(_05584_),
    .B1(_05590_),
    .B2(_05592_),
    .ZN(_05593_));
 AND2_X4 _30826_ (.A1(_16798_),
    .A2(_16799_),
    .ZN(_05594_));
 BUF_X8 _30827_ (.A(_05594_),
    .Z(_05595_));
 INV_X32 _30828_ (.A(_16796_),
    .ZN(_05596_));
 OAI21_X1 _30829_ (.A(_05595_),
    .B1(_05582_),
    .B2(_05596_),
    .ZN(_05597_));
 INV_X1 _30830_ (.A(_16799_),
    .ZN(_05598_));
 NOR2_X4 _30831_ (.A1(_05598_),
    .A2(_05578_),
    .ZN(_05600_));
 BUF_X4 _30832_ (.A(_05600_),
    .Z(_05601_));
 INV_X1 _30833_ (.A(_05601_),
    .ZN(_05602_));
 BUF_X4 _30834_ (.A(_05596_),
    .Z(_05603_));
 OAI21_X1 _30835_ (.A(_05597_),
    .B1(_05602_),
    .B2(_05603_),
    .ZN(_05604_));
 OAI21_X1 _30836_ (.A(_05576_),
    .B1(_05593_),
    .B2(_05604_),
    .ZN(_05605_));
 INV_X16 _30837_ (.A(_16801_),
    .ZN(_05606_));
 NOR2_X4 _30838_ (.A1(_05606_),
    .A2(_16800_),
    .ZN(_05607_));
 AND2_X2 _30839_ (.A1(_05607_),
    .A2(_05573_),
    .ZN(_05608_));
 AND2_X4 _30840_ (.A1(_05587_),
    .A2(_05582_),
    .ZN(_05609_));
 BUF_X8 _30841_ (.A(_05609_),
    .Z(_05611_));
 AND2_X2 _30842_ (.A1(_05587_),
    .A2(_16797_),
    .ZN(_05612_));
 BUF_X4 _30843_ (.A(_05612_),
    .Z(_05613_));
 OAI21_X1 _30844_ (.A(_05608_),
    .B1(_05611_),
    .B2(_05613_),
    .ZN(_05614_));
 NOR2_X4 _30845_ (.A1(_05596_),
    .A2(_16797_),
    .ZN(_05615_));
 AND2_X1 _30846_ (.A1(_05615_),
    .A2(_05581_),
    .ZN(_05616_));
 AND2_X1 _30847_ (.A1(_05608_),
    .A2(_05616_),
    .ZN(_05617_));
 INV_X1 _30848_ (.A(_05617_),
    .ZN(_05618_));
 AND2_X4 _30849_ (.A1(_16797_),
    .A2(_16796_),
    .ZN(_05619_));
 BUF_X8 _30850_ (.A(_05619_),
    .Z(_05620_));
 AND2_X4 _30851_ (.A1(_05620_),
    .A2(_05581_),
    .ZN(_05622_));
 BUF_X2 _30852_ (.A(_05622_),
    .Z(_05623_));
 BUF_X2 _30853_ (.A(_05607_),
    .Z(_05624_));
 NAND3_X1 _30854_ (.A1(_05623_),
    .A2(_05624_),
    .A3(_05573_),
    .ZN(_05625_));
 INV_X1 _30855_ (.A(_05608_),
    .ZN(_05626_));
 OAI21_X1 _30856_ (.A(_05600_),
    .B1(_05582_),
    .B2(_16796_),
    .ZN(_05627_));
 NOR2_X1 _30857_ (.A1(_05626_),
    .A2(_05627_),
    .ZN(_05628_));
 NOR2_X4 _30858_ (.A1(_05582_),
    .A2(_16796_),
    .ZN(_05629_));
 BUF_X4 _30859_ (.A(_05629_),
    .Z(_05630_));
 AND2_X4 _30860_ (.A1(_05630_),
    .A2(_05595_),
    .ZN(_05631_));
 AOI21_X1 _30861_ (.A(_05628_),
    .B1(_05631_),
    .B2(_05608_),
    .ZN(_05633_));
 AND4_X1 _30862_ (.A1(_05614_),
    .A2(_05618_),
    .A3(_05625_),
    .A4(_05633_),
    .ZN(_05634_));
 AND2_X1 _30863_ (.A1(_05606_),
    .A2(_16800_),
    .ZN(_05635_));
 BUF_X4 _30864_ (.A(_05635_),
    .Z(_05636_));
 AND2_X2 _30865_ (.A1(_05636_),
    .A2(_05573_),
    .ZN(_05637_));
 BUF_X4 _30866_ (.A(_16796_),
    .Z(_05638_));
 AND2_X2 _30867_ (.A1(_05601_),
    .A2(_05638_),
    .ZN(_05639_));
 AND2_X1 _30868_ (.A1(_05594_),
    .A2(_05619_),
    .ZN(_05640_));
 BUF_X2 _30869_ (.A(_05640_),
    .Z(_05641_));
 OAI21_X1 _30870_ (.A(_05637_),
    .B1(_05639_),
    .B2(_05641_),
    .ZN(_05642_));
 AND2_X1 _30871_ (.A1(_05637_),
    .A2(_05612_),
    .ZN(_05644_));
 INV_X1 _30872_ (.A(_05644_),
    .ZN(_05645_));
 BUF_X4 _30873_ (.A(_05583_),
    .Z(_05646_));
 NAND2_X1 _30874_ (.A1(_05637_),
    .A2(_05646_),
    .ZN(_05647_));
 NAND2_X1 _30875_ (.A1(_05637_),
    .A2(_05623_),
    .ZN(_05648_));
 AND4_X1 _30876_ (.A1(_05642_),
    .A2(_05645_),
    .A3(_05647_),
    .A4(_05648_),
    .ZN(_05649_));
 AND2_X4 _30877_ (.A1(_16801_),
    .A2(_16800_),
    .ZN(_05650_));
 BUF_X4 _30878_ (.A(_05650_),
    .Z(_05651_));
 BUF_X2 _30879_ (.A(_05651_),
    .Z(_05652_));
 NAND3_X1 _30880_ (.A1(_05646_),
    .A2(_05573_),
    .A3(_05652_),
    .ZN(_05653_));
 AND2_X2 _30881_ (.A1(_05573_),
    .A2(_05651_),
    .ZN(_05655_));
 BUF_X8 _30882_ (.A(_05655_),
    .Z(_05656_));
 AND2_X4 _30883_ (.A1(_05615_),
    .A2(_05595_),
    .ZN(_05657_));
 NOR2_X4 _30884_ (.A1(_05631_),
    .A2(_05657_),
    .ZN(_05658_));
 INV_X1 _30885_ (.A(_05658_),
    .ZN(_05659_));
 AND2_X1 _30886_ (.A1(_05600_),
    .A2(_05620_),
    .ZN(_05660_));
 BUF_X4 _30887_ (.A(_05660_),
    .Z(_05661_));
 OAI21_X1 _30888_ (.A(_05656_),
    .B1(_05659_),
    .B2(_05661_),
    .ZN(_05662_));
 NAND2_X1 _30889_ (.A1(_05655_),
    .A2(_05622_),
    .ZN(_05663_));
 NOR2_X1 _30890_ (.A1(_05596_),
    .A2(_05579_),
    .ZN(_05664_));
 AND2_X2 _30891_ (.A1(_05664_),
    .A2(_05578_),
    .ZN(_05666_));
 NAND2_X1 _30892_ (.A1(_05666_),
    .A2(_05655_),
    .ZN(_05667_));
 AND4_X1 _30893_ (.A1(_05653_),
    .A2(_05662_),
    .A3(_05663_),
    .A4(_05667_),
    .ZN(_05668_));
 AND4_X1 _30894_ (.A1(_05605_),
    .A2(_05634_),
    .A3(_05649_),
    .A4(_05668_),
    .ZN(_05669_));
 NOR2_X1 _30895_ (.A1(_16803_),
    .A2(_16802_),
    .ZN(_05670_));
 AND2_X2 _30896_ (.A1(_05670_),
    .A2(_05574_),
    .ZN(_05671_));
 BUF_X4 _30897_ (.A(_05595_),
    .Z(_05672_));
 BUF_X4 _30898_ (.A(_05615_),
    .Z(_05673_));
 OAI211_X2 _30899_ (.A(_05671_),
    .B(_05672_),
    .C1(_05630_),
    .C2(_05673_),
    .ZN(_05674_));
 CLKBUF_X2 _30900_ (.A(_05670_),
    .Z(_05675_));
 BUF_X2 _30901_ (.A(_05574_),
    .Z(_05677_));
 NAND4_X1 _30902_ (.A1(_05601_),
    .A2(_05673_),
    .A3(_05675_),
    .A4(_05677_),
    .ZN(_05678_));
 AND2_X2 _30903_ (.A1(_05600_),
    .A2(_16797_),
    .ZN(_05679_));
 INV_X4 _30904_ (.A(_05679_),
    .ZN(_05680_));
 INV_X1 _30905_ (.A(_05671_),
    .ZN(_05681_));
 OAI211_X2 _30906_ (.A(_05674_),
    .B(_05678_),
    .C1(_05680_),
    .C2(_05681_),
    .ZN(_05682_));
 BUF_X2 _30907_ (.A(_05671_),
    .Z(_05683_));
 AND2_X1 _30908_ (.A1(_05581_),
    .A2(_16797_),
    .ZN(_05684_));
 BUF_X4 _30909_ (.A(_05684_),
    .Z(_05685_));
 AND2_X1 _30910_ (.A1(_05683_),
    .A2(_05685_),
    .ZN(_05686_));
 AND2_X1 _30911_ (.A1(_05612_),
    .A2(_05671_),
    .ZN(_05688_));
 AND3_X1 _30912_ (.A1(_05671_),
    .A2(_05587_),
    .A3(_05673_),
    .ZN(_05689_));
 NOR4_X1 _30913_ (.A1(_05682_),
    .A2(_05686_),
    .A3(_05688_),
    .A4(_05689_),
    .ZN(_05690_));
 AND2_X2 _30914_ (.A1(_05635_),
    .A2(_05670_),
    .ZN(_05691_));
 AND2_X2 _30915_ (.A1(_05592_),
    .A2(_05586_),
    .ZN(_05692_));
 INV_X1 _30916_ (.A(_05620_),
    .ZN(_05693_));
 BUF_X2 _30917_ (.A(_05693_),
    .Z(_05694_));
 AND3_X1 _30918_ (.A1(_05691_),
    .A2(_05692_),
    .A3(_05694_),
    .ZN(_05695_));
 NOR2_X1 _30919_ (.A1(_05627_),
    .A2(_05615_),
    .ZN(_05696_));
 AND2_X1 _30920_ (.A1(_05696_),
    .A2(_05691_),
    .ZN(_05697_));
 BUF_X2 _30921_ (.A(_05691_),
    .Z(_05699_));
 AOI211_X2 _30922_ (.A(_05695_),
    .B(_05697_),
    .C1(_05699_),
    .C2(_05685_),
    .ZN(_05700_));
 NAND3_X1 _30923_ (.A1(_05583_),
    .A2(_05670_),
    .A3(_05607_),
    .ZN(_05701_));
 NAND4_X1 _30924_ (.A1(_05630_),
    .A2(_05607_),
    .A3(_05581_),
    .A4(_05670_),
    .ZN(_05702_));
 NAND2_X1 _30925_ (.A1(_05701_),
    .A2(_05702_),
    .ZN(_05703_));
 INV_X1 _30926_ (.A(_05703_),
    .ZN(_05704_));
 AND2_X1 _30927_ (.A1(_05607_),
    .A2(_05670_),
    .ZN(_05705_));
 AND3_X1 _30928_ (.A1(_05705_),
    .A2(_05601_),
    .A3(_05592_),
    .ZN(_05706_));
 INV_X1 _30929_ (.A(_05706_),
    .ZN(_05707_));
 BUF_X4 _30930_ (.A(_05705_),
    .Z(_05708_));
 NAND3_X1 _30931_ (.A1(_05692_),
    .A2(_05708_),
    .A3(_05694_),
    .ZN(_05710_));
 AND2_X2 _30932_ (.A1(_05595_),
    .A2(_05591_),
    .ZN(_05711_));
 BUF_X4 _30933_ (.A(_16797_),
    .Z(_05712_));
 AND2_X2 _30934_ (.A1(_05595_),
    .A2(_05712_),
    .ZN(_05713_));
 OAI21_X1 _30935_ (.A(_05708_),
    .B1(_05711_),
    .B2(_05713_),
    .ZN(_05714_));
 AND4_X1 _30936_ (.A1(_05704_),
    .A2(_05707_),
    .A3(_05710_),
    .A4(_05714_),
    .ZN(_05715_));
 AND2_X2 _30937_ (.A1(_05651_),
    .A2(_05670_),
    .ZN(_05716_));
 INV_X1 _30938_ (.A(_05716_),
    .ZN(_05717_));
 AND2_X1 _30939_ (.A1(_05629_),
    .A2(_05586_),
    .ZN(_05718_));
 BUF_X2 _30940_ (.A(_05718_),
    .Z(_05719_));
 INV_X1 _30941_ (.A(_05719_),
    .ZN(_05721_));
 BUF_X8 _30942_ (.A(_05581_),
    .Z(_05722_));
 NAND2_X1 _30943_ (.A1(_05592_),
    .A2(_05722_),
    .ZN(_05723_));
 AOI21_X1 _30944_ (.A(_05717_),
    .B1(_05721_),
    .B2(_05723_),
    .ZN(_05724_));
 AND2_X1 _30945_ (.A1(_05641_),
    .A2(_05716_),
    .ZN(_05725_));
 BUF_X2 _30946_ (.A(_05591_),
    .Z(_05726_));
 AND3_X1 _30947_ (.A1(_05716_),
    .A2(_05601_),
    .A3(_05726_),
    .ZN(_05727_));
 NAND2_X1 _30948_ (.A1(_05582_),
    .A2(_05579_),
    .ZN(_05728_));
 NOR2_X2 _30949_ (.A1(_05728_),
    .A2(_05585_),
    .ZN(_05729_));
 AND2_X1 _30950_ (.A1(_05716_),
    .A2(_05729_),
    .ZN(_05730_));
 NOR4_X1 _30951_ (.A1(_05724_),
    .A2(_05725_),
    .A3(_05727_),
    .A4(_05730_),
    .ZN(_05732_));
 AND4_X1 _30952_ (.A1(_05690_),
    .A2(_05700_),
    .A3(_05715_),
    .A4(_05732_),
    .ZN(_05733_));
 AND2_X1 _30953_ (.A1(_05572_),
    .A2(_16803_),
    .ZN(_05734_));
 BUF_X2 _30954_ (.A(_05734_),
    .Z(_05735_));
 BUF_X4 _30955_ (.A(_05735_),
    .Z(_05736_));
 OAI211_X2 _30956_ (.A(_05624_),
    .B(_05736_),
    .C1(_05641_),
    .C2(_05729_),
    .ZN(_05737_));
 BUF_X8 _30957_ (.A(_05601_),
    .Z(_05738_));
 NAND4_X1 _30958_ (.A1(_05736_),
    .A2(_05738_),
    .A3(_05673_),
    .A4(_05624_),
    .ZN(_05739_));
 AND2_X1 _30959_ (.A1(_05737_),
    .A2(_05739_),
    .ZN(_05740_));
 AND2_X1 _30960_ (.A1(_05734_),
    .A2(_05650_),
    .ZN(_05741_));
 INV_X1 _30961_ (.A(_05741_),
    .ZN(_05743_));
 INV_X1 _30962_ (.A(_05615_),
    .ZN(_05744_));
 BUF_X2 _30963_ (.A(_05744_),
    .Z(_05745_));
 NAND2_X1 _30964_ (.A1(_05745_),
    .A2(_05581_),
    .ZN(_05746_));
 NOR2_X1 _30965_ (.A1(_05743_),
    .A2(_05746_),
    .ZN(_05747_));
 INV_X4 _30966_ (.A(_05630_),
    .ZN(_05748_));
 NAND2_X1 _30967_ (.A1(_05748_),
    .A2(_05586_),
    .ZN(_05749_));
 NOR2_X1 _30968_ (.A1(_05743_),
    .A2(_05749_),
    .ZN(_05750_));
 BUF_X4 _30969_ (.A(_05741_),
    .Z(_05751_));
 AOI211_X2 _30970_ (.A(_05747_),
    .B(_05750_),
    .C1(_05711_),
    .C2(_05751_),
    .ZN(_05752_));
 AND2_X1 _30971_ (.A1(_05734_),
    .A2(_05635_),
    .ZN(_05754_));
 BUF_X2 _30972_ (.A(_05754_),
    .Z(_05755_));
 NAND2_X1 _30973_ (.A1(_05755_),
    .A2(_05713_),
    .ZN(_05756_));
 AND2_X1 _30974_ (.A1(_05734_),
    .A2(_05574_),
    .ZN(_05757_));
 BUF_X4 _30975_ (.A(_05757_),
    .Z(_05758_));
 INV_X1 _30976_ (.A(_05749_),
    .ZN(_05759_));
 AND2_X1 _30977_ (.A1(_05722_),
    .A2(_05596_),
    .ZN(_05760_));
 OAI21_X1 _30978_ (.A(_05758_),
    .B1(_05759_),
    .B2(_05760_),
    .ZN(_05761_));
 AND2_X2 _30979_ (.A1(_05630_),
    .A2(_05581_),
    .ZN(_05762_));
 BUF_X4 _30980_ (.A(_05616_),
    .Z(_05763_));
 OAI21_X1 _30981_ (.A(_05755_),
    .B1(_05762_),
    .B2(_05763_),
    .ZN(_05765_));
 NAND2_X1 _30982_ (.A1(_05592_),
    .A2(_05595_),
    .ZN(_05766_));
 INV_X1 _30983_ (.A(_05766_),
    .ZN(_05767_));
 OAI21_X1 _30984_ (.A(_05758_),
    .B1(_05767_),
    .B2(_05639_),
    .ZN(_05768_));
 AND4_X1 _30985_ (.A1(_05756_),
    .A2(_05761_),
    .A3(_05765_),
    .A4(_05768_),
    .ZN(_05769_));
 AND2_X1 _30986_ (.A1(_05734_),
    .A2(_05607_),
    .ZN(_05770_));
 BUF_X2 _30987_ (.A(_05770_),
    .Z(_05771_));
 AND2_X1 _30988_ (.A1(_05587_),
    .A2(_05591_),
    .ZN(_05772_));
 AND2_X1 _30989_ (.A1(_05771_),
    .A2(_05772_),
    .ZN(_05773_));
 INV_X1 _30990_ (.A(_05773_),
    .ZN(_05774_));
 AND4_X1 _30991_ (.A1(_05740_),
    .A2(_05752_),
    .A3(_05769_),
    .A4(_05774_),
    .ZN(_05776_));
 AND2_X4 _30992_ (.A1(_16803_),
    .A2(_16802_),
    .ZN(_05777_));
 AND2_X4 _30993_ (.A1(_05607_),
    .A2(_05777_),
    .ZN(_05778_));
 BUF_X8 _30994_ (.A(_05778_),
    .Z(_05779_));
 INV_X2 _30995_ (.A(_05779_),
    .ZN(_05780_));
 OAI21_X1 _30996_ (.A(_05600_),
    .B1(_16797_),
    .B2(_05596_),
    .ZN(_05781_));
 NOR2_X1 _30997_ (.A1(_05780_),
    .A2(_05781_),
    .ZN(_05782_));
 INV_X1 _30998_ (.A(_05580_),
    .ZN(_05783_));
 NOR2_X2 _30999_ (.A1(_05783_),
    .A2(_05630_),
    .ZN(_05784_));
 AND3_X1 _31000_ (.A1(_05779_),
    .A2(_05784_),
    .A3(_05745_),
    .ZN(_05785_));
 AND2_X1 _31001_ (.A1(_05609_),
    .A2(_05779_),
    .ZN(_05787_));
 AND2_X4 _31002_ (.A1(_05595_),
    .A2(_05638_),
    .ZN(_05788_));
 BUF_X4 _31003_ (.A(_05777_),
    .Z(_05789_));
 AND3_X2 _31004_ (.A1(_05788_),
    .A2(_05789_),
    .A3(_05624_),
    .ZN(_05790_));
 OR4_X2 _31005_ (.A1(_05782_),
    .A2(_05785_),
    .A3(_05787_),
    .A4(_05790_),
    .ZN(_05791_));
 AND2_X2 _31006_ (.A1(_05635_),
    .A2(_05777_),
    .ZN(_05792_));
 AND2_X1 _31007_ (.A1(_05586_),
    .A2(_05615_),
    .ZN(_05793_));
 BUF_X2 _31008_ (.A(_05793_),
    .Z(_05794_));
 OAI21_X1 _31009_ (.A(_05792_),
    .B1(_05794_),
    .B2(_05762_),
    .ZN(_05795_));
 BUF_X4 _31010_ (.A(_05657_),
    .Z(_05796_));
 OAI21_X1 _31011_ (.A(_05792_),
    .B1(_05631_),
    .B2(_05796_),
    .ZN(_05798_));
 NOR2_X1 _31012_ (.A1(_05728_),
    .A2(_05578_),
    .ZN(_05799_));
 BUF_X4 _31013_ (.A(_05799_),
    .Z(_05800_));
 OAI21_X1 _31014_ (.A(_05792_),
    .B1(_05679_),
    .B2(_05800_),
    .ZN(_05801_));
 NAND3_X1 _31015_ (.A1(_05795_),
    .A2(_05798_),
    .A3(_05801_),
    .ZN(_05802_));
 AND2_X1 _31016_ (.A1(_05789_),
    .A2(_05574_),
    .ZN(_05803_));
 BUF_X4 _31017_ (.A(_05803_),
    .Z(_05804_));
 BUF_X4 _31018_ (.A(_05582_),
    .Z(_05805_));
 OAI211_X2 _31019_ (.A(_05804_),
    .B(_05672_),
    .C1(_05805_),
    .C2(_05603_),
    .ZN(_05806_));
 BUF_X2 _31020_ (.A(_05630_),
    .Z(_05807_));
 BUF_X2 _31021_ (.A(_05789_),
    .Z(_05809_));
 NAND4_X1 _31022_ (.A1(_05807_),
    .A2(_05809_),
    .A3(_05722_),
    .A4(_05677_),
    .ZN(_05810_));
 INV_X1 _31023_ (.A(_05804_),
    .ZN(_05811_));
 INV_X1 _31024_ (.A(_05639_),
    .ZN(_05812_));
 OAI211_X2 _31025_ (.A(_05806_),
    .B(_05810_),
    .C1(_05811_),
    .C2(_05812_),
    .ZN(_05813_));
 AND2_X1 _31026_ (.A1(_05789_),
    .A2(_05651_),
    .ZN(_05814_));
 BUF_X4 _31027_ (.A(_05814_),
    .Z(_05815_));
 OAI21_X1 _31028_ (.A(_05815_),
    .B1(_05679_),
    .B2(_05800_),
    .ZN(_05816_));
 BUF_X4 _31029_ (.A(_05722_),
    .Z(_05817_));
 BUF_X4 _31030_ (.A(_05638_),
    .Z(_05818_));
 OAI211_X2 _31031_ (.A(_05815_),
    .B(_05817_),
    .C1(_05712_),
    .C2(_05818_),
    .ZN(_05820_));
 NAND2_X1 _31032_ (.A1(_05772_),
    .A2(_05815_),
    .ZN(_05821_));
 NAND3_X1 _31033_ (.A1(_05815_),
    .A2(_05672_),
    .A3(_05807_),
    .ZN(_05822_));
 NAND4_X1 _31034_ (.A1(_05816_),
    .A2(_05820_),
    .A3(_05821_),
    .A4(_05822_),
    .ZN(_05823_));
 NOR4_X2 _31035_ (.A1(_05791_),
    .A2(_05802_),
    .A3(_05813_),
    .A4(_05823_),
    .ZN(_05824_));
 NAND4_X1 _31036_ (.A1(_05669_),
    .A2(_05733_),
    .A3(_05776_),
    .A4(_05824_),
    .ZN(_05825_));
 OAI21_X1 _31037_ (.A(_05598_),
    .B1(_05592_),
    .B2(_05578_),
    .ZN(_05826_));
 CLKBUF_X2 _31038_ (.A(_05677_),
    .Z(_05827_));
 AND3_X1 _31039_ (.A1(_05675_),
    .A2(_05827_),
    .A3(_05598_),
    .ZN(_05828_));
 AND2_X1 _31040_ (.A1(_05826_),
    .A2(_05828_),
    .ZN(_05829_));
 OR2_X2 _31041_ (.A1(_05825_),
    .A2(_05829_),
    .ZN(_05831_));
 XNOR2_X1 _31042_ (.A(_05831_),
    .B(_14297_),
    .ZN(_05832_));
 XNOR2_X1 _31043_ (.A(_05571_),
    .B(_05832_),
    .ZN(_05833_));
 INV_X16 _31044_ (.A(_16843_),
    .ZN(_05834_));
 AND2_X4 _31045_ (.A1(_05834_),
    .A2(_16842_),
    .ZN(_05835_));
 BUF_X4 _31046_ (.A(_05835_),
    .Z(_05836_));
 NOR2_X1 _31047_ (.A1(_16841_),
    .A2(_16840_),
    .ZN(_05837_));
 AND2_X1 _31048_ (.A1(_05836_),
    .A2(_05837_),
    .ZN(_05838_));
 INV_X1 _31049_ (.A(_16838_),
    .ZN(_05839_));
 NOR2_X2 _31050_ (.A1(_05839_),
    .A2(_16839_),
    .ZN(_05840_));
 BUF_X4 _31051_ (.A(_05840_),
    .Z(_05842_));
 NOR2_X4 _31052_ (.A1(_16837_),
    .A2(_16836_),
    .ZN(_05843_));
 AND2_X2 _31053_ (.A1(_05842_),
    .A2(_05843_),
    .ZN(_05844_));
 AND2_X1 _31054_ (.A1(_05838_),
    .A2(_05844_),
    .ZN(_05845_));
 INV_X16 _31055_ (.A(_16841_),
    .ZN(_05846_));
 NOR2_X4 _31056_ (.A1(_05846_),
    .A2(_16840_),
    .ZN(_05847_));
 AND2_X1 _31057_ (.A1(_05835_),
    .A2(_05847_),
    .ZN(_05848_));
 BUF_X4 _31058_ (.A(_05848_),
    .Z(_05849_));
 INV_X32 _31059_ (.A(_16836_),
    .ZN(_05850_));
 NOR2_X4 _31060_ (.A1(_05850_),
    .A2(_16837_),
    .ZN(_05851_));
 NOR2_X4 _31061_ (.A1(_16838_),
    .A2(_16839_),
    .ZN(_05853_));
 BUF_X4 _31062_ (.A(_05853_),
    .Z(_05854_));
 AND2_X2 _31063_ (.A1(_05851_),
    .A2(_05854_),
    .ZN(_05855_));
 AND2_X1 _31064_ (.A1(_05849_),
    .A2(_05855_),
    .ZN(_05856_));
 AND2_X4 _31065_ (.A1(_16837_),
    .A2(_16836_),
    .ZN(_05857_));
 BUF_X4 _31066_ (.A(_05857_),
    .Z(_05858_));
 AND2_X4 _31067_ (.A1(_05858_),
    .A2(_05853_),
    .ZN(_05859_));
 BUF_X4 _31068_ (.A(_05859_),
    .Z(_05860_));
 AND2_X4 _31069_ (.A1(_05849_),
    .A2(_05860_),
    .ZN(_05861_));
 INV_X32 _31070_ (.A(_16837_),
    .ZN(_05862_));
 NOR2_X2 _31071_ (.A1(_05862_),
    .A2(_16836_),
    .ZN(_05864_));
 AND2_X2 _31072_ (.A1(_05842_),
    .A2(_05864_),
    .ZN(_05865_));
 AND2_X1 _31073_ (.A1(_05849_),
    .A2(_05865_),
    .ZN(_05866_));
 OR4_X4 _31074_ (.A1(_05845_),
    .A2(_05856_),
    .A3(_05861_),
    .A4(_05866_),
    .ZN(_05867_));
 BUF_X4 _31075_ (.A(_05850_),
    .Z(_05868_));
 AND2_X4 _31076_ (.A1(_16838_),
    .A2(_16839_),
    .ZN(_05869_));
 BUF_X4 _31077_ (.A(_05869_),
    .Z(_05870_));
 BUF_X4 _31078_ (.A(_16837_),
    .Z(_05871_));
 AND2_X4 _31079_ (.A1(_05870_),
    .A2(_05871_),
    .ZN(_05872_));
 BUF_X2 _31080_ (.A(_05872_),
    .Z(_05873_));
 AND2_X2 _31081_ (.A1(_16843_),
    .A2(_16842_),
    .ZN(_05875_));
 AND2_X1 _31082_ (.A1(_05875_),
    .A2(_05837_),
    .ZN(_05876_));
 AND2_X1 _31083_ (.A1(_05873_),
    .A2(_05876_),
    .ZN(_05877_));
 NOR2_X1 _31084_ (.A1(_05834_),
    .A2(_16842_),
    .ZN(_05878_));
 AND2_X4 _31085_ (.A1(_16841_),
    .A2(_16840_),
    .ZN(_05879_));
 BUF_X2 _31086_ (.A(_05879_),
    .Z(_05880_));
 AND2_X1 _31087_ (.A1(_05878_),
    .A2(_05880_),
    .ZN(_05881_));
 BUF_X2 _31088_ (.A(_05881_),
    .Z(_05882_));
 BUF_X4 _31089_ (.A(_05882_),
    .Z(_05883_));
 BUF_X4 _31090_ (.A(_05870_),
    .Z(_05884_));
 INV_X1 _31091_ (.A(_05884_),
    .ZN(_05886_));
 INV_X4 _31092_ (.A(_05843_),
    .ZN(_05887_));
 INV_X1 _31093_ (.A(_05854_),
    .ZN(_05888_));
 BUF_X4 _31094_ (.A(_05851_),
    .Z(_05889_));
 OAI22_X1 _31095_ (.A1(_05886_),
    .A2(_05887_),
    .B1(_05888_),
    .B2(_05889_),
    .ZN(_05890_));
 AOI221_X2 _31096_ (.A(_05867_),
    .B1(_05868_),
    .B2(_05877_),
    .C1(_05883_),
    .C2(_05890_),
    .ZN(_05891_));
 AND2_X4 _31097_ (.A1(_05846_),
    .A2(_16840_),
    .ZN(_05892_));
 BUF_X2 _31098_ (.A(_05878_),
    .Z(_05893_));
 AND2_X2 _31099_ (.A1(_05892_),
    .A2(_05893_),
    .ZN(_05894_));
 BUF_X4 _31100_ (.A(_05894_),
    .Z(_05895_));
 OAI21_X1 _31101_ (.A(_05854_),
    .B1(_05889_),
    .B2(_05864_),
    .ZN(_05897_));
 INV_X1 _31102_ (.A(_05897_),
    .ZN(_05898_));
 OAI21_X1 _31103_ (.A(_05895_),
    .B1(_05898_),
    .B2(_05873_),
    .ZN(_05899_));
 BUF_X4 _31104_ (.A(_05862_),
    .Z(_05900_));
 AND2_X2 _31105_ (.A1(_05870_),
    .A2(_05900_),
    .ZN(_05901_));
 NOR2_X1 _31106_ (.A1(_16843_),
    .A2(_16842_),
    .ZN(_05902_));
 AND2_X2 _31107_ (.A1(_05880_),
    .A2(_05902_),
    .ZN(_05903_));
 AND2_X1 _31108_ (.A1(_05901_),
    .A2(_05903_),
    .ZN(_05904_));
 INV_X1 _31109_ (.A(_05904_),
    .ZN(_05905_));
 AND2_X1 _31110_ (.A1(_05836_),
    .A2(_05892_),
    .ZN(_05906_));
 BUF_X2 _31111_ (.A(_05906_),
    .Z(_05908_));
 AND2_X2 _31112_ (.A1(_05842_),
    .A2(_05871_),
    .ZN(_05909_));
 NAND2_X1 _31113_ (.A1(_05908_),
    .A2(_05909_),
    .ZN(_05910_));
 AND2_X1 _31114_ (.A1(_05853_),
    .A2(_05862_),
    .ZN(_05911_));
 BUF_X4 _31115_ (.A(_05911_),
    .Z(_05912_));
 NAND3_X1 _31116_ (.A1(_05912_),
    .A2(_05837_),
    .A3(_05836_),
    .ZN(_05913_));
 BUF_X4 _31117_ (.A(_05849_),
    .Z(_05914_));
 AND2_X2 _31118_ (.A1(_05842_),
    .A2(_05900_),
    .ZN(_05915_));
 NAND2_X1 _31119_ (.A1(_05914_),
    .A2(_05915_),
    .ZN(_05916_));
 AND4_X1 _31120_ (.A1(_05905_),
    .A2(_05910_),
    .A3(_05913_),
    .A4(_05916_),
    .ZN(_05917_));
 AND2_X1 _31121_ (.A1(_05835_),
    .A2(_05879_),
    .ZN(_05919_));
 BUF_X2 _31122_ (.A(_05919_),
    .Z(_05920_));
 BUF_X2 _31123_ (.A(_05920_),
    .Z(_05921_));
 AND2_X2 _31124_ (.A1(_05842_),
    .A2(_16836_),
    .ZN(_05922_));
 AND2_X1 _31125_ (.A1(_05853_),
    .A2(_16836_),
    .ZN(_05923_));
 OAI21_X1 _31126_ (.A(_05921_),
    .B1(_05922_),
    .B2(_05923_),
    .ZN(_05924_));
 AND2_X2 _31127_ (.A1(_05902_),
    .A2(_05837_),
    .ZN(_05925_));
 BUF_X2 _31128_ (.A(_05925_),
    .Z(_05926_));
 NAND2_X1 _31129_ (.A1(_05887_),
    .A2(_05870_),
    .ZN(_05927_));
 NOR2_X1 _31130_ (.A1(_05927_),
    .A2(_05858_),
    .ZN(_05928_));
 NOR2_X1 _31131_ (.A1(_05900_),
    .A2(_16838_),
    .ZN(_05930_));
 OAI21_X1 _31132_ (.A(_05926_),
    .B1(_05928_),
    .B2(_05930_),
    .ZN(_05931_));
 AND4_X1 _31133_ (.A1(_05899_),
    .A2(_05917_),
    .A3(_05924_),
    .A4(_05931_),
    .ZN(_05932_));
 AND2_X1 _31134_ (.A1(_05864_),
    .A2(_05870_),
    .ZN(_05933_));
 BUF_X2 _31135_ (.A(_05933_),
    .Z(_05934_));
 AND2_X2 _31136_ (.A1(_05875_),
    .A2(_05880_),
    .ZN(_05935_));
 BUF_X2 _31137_ (.A(_05935_),
    .Z(_05936_));
 NAND2_X1 _31138_ (.A1(_05934_),
    .A2(_05936_),
    .ZN(_05937_));
 INV_X1 _31139_ (.A(_05844_),
    .ZN(_05938_));
 INV_X2 _31140_ (.A(_05935_),
    .ZN(_05939_));
 OAI21_X1 _31141_ (.A(_05937_),
    .B1(_05938_),
    .B2(_05939_),
    .ZN(_05941_));
 NAND2_X1 _31142_ (.A1(_05855_),
    .A2(_05936_),
    .ZN(_05942_));
 AND2_X2 _31143_ (.A1(_05864_),
    .A2(_05853_),
    .ZN(_05943_));
 INV_X1 _31144_ (.A(_05943_),
    .ZN(_05944_));
 INV_X1 _31145_ (.A(_05876_),
    .ZN(_05945_));
 BUF_X4 _31146_ (.A(_05945_),
    .Z(_05946_));
 OAI21_X1 _31147_ (.A(_05942_),
    .B1(_05944_),
    .B2(_05946_),
    .ZN(_05947_));
 AND2_X1 _31148_ (.A1(_05847_),
    .A2(_05902_),
    .ZN(_05948_));
 BUF_X4 _31149_ (.A(_05948_),
    .Z(_05949_));
 INV_X1 _31150_ (.A(_05949_),
    .ZN(_05950_));
 OAI21_X1 _31151_ (.A(_05854_),
    .B1(_05900_),
    .B2(_05868_),
    .ZN(_05952_));
 NOR2_X1 _31152_ (.A1(_05950_),
    .A2(_05952_),
    .ZN(_05953_));
 INV_X32 _31153_ (.A(_16839_),
    .ZN(_05954_));
 NOR2_X2 _31154_ (.A1(_05954_),
    .A2(_16838_),
    .ZN(_05955_));
 BUF_X4 _31155_ (.A(_05955_),
    .Z(_05956_));
 NAND2_X1 _31156_ (.A1(_05887_),
    .A2(_05956_),
    .ZN(_05957_));
 INV_X1 _31157_ (.A(_05957_),
    .ZN(_05958_));
 AND2_X1 _31158_ (.A1(_05958_),
    .A2(_05949_),
    .ZN(_05959_));
 NOR4_X1 _31159_ (.A1(_05941_),
    .A2(_05947_),
    .A3(_05953_),
    .A4(_05959_),
    .ZN(_05960_));
 AND2_X2 _31160_ (.A1(_05840_),
    .A2(_05858_),
    .ZN(_05961_));
 NAND2_X1 _31161_ (.A1(_05849_),
    .A2(_05961_),
    .ZN(_05963_));
 AND2_X2 _31162_ (.A1(_05955_),
    .A2(_05843_),
    .ZN(_05964_));
 INV_X1 _31163_ (.A(_05964_),
    .ZN(_05965_));
 AND2_X4 _31164_ (.A1(_05955_),
    .A2(_05858_),
    .ZN(_05966_));
 BUF_X4 _31165_ (.A(_05966_),
    .Z(_05967_));
 INV_X4 _31166_ (.A(_05967_),
    .ZN(_05968_));
 NAND2_X2 _31167_ (.A1(_05965_),
    .A2(_05968_),
    .ZN(_05969_));
 AND2_X1 _31168_ (.A1(_05892_),
    .A2(_05902_),
    .ZN(_05970_));
 BUF_X2 _31169_ (.A(_05970_),
    .Z(_05971_));
 BUF_X2 _31170_ (.A(_05971_),
    .Z(_05972_));
 AND2_X1 _31171_ (.A1(_05969_),
    .A2(_05972_),
    .ZN(_05974_));
 INV_X2 _31172_ (.A(_05858_),
    .ZN(_05975_));
 NAND2_X1 _31173_ (.A1(_05975_),
    .A2(_05842_),
    .ZN(_05976_));
 NOR2_X2 _31174_ (.A1(_05976_),
    .A2(_05843_),
    .ZN(_05977_));
 INV_X1 _31175_ (.A(_05977_),
    .ZN(_05978_));
 INV_X1 _31176_ (.A(_05872_),
    .ZN(_05979_));
 AOI21_X1 _31177_ (.A(_05950_),
    .B1(_05978_),
    .B2(_05979_),
    .ZN(_05980_));
 INV_X1 _31178_ (.A(_05976_),
    .ZN(_05981_));
 AND3_X1 _31179_ (.A1(_05981_),
    .A2(_05887_),
    .A3(_05971_),
    .ZN(_05982_));
 AND2_X1 _31180_ (.A1(_05853_),
    .A2(_05871_),
    .ZN(_05983_));
 BUF_X2 _31181_ (.A(_05983_),
    .Z(_05985_));
 AND2_X1 _31182_ (.A1(_05971_),
    .A2(_05985_),
    .ZN(_05986_));
 NOR4_X1 _31183_ (.A1(_05974_),
    .A2(_05980_),
    .A3(_05982_),
    .A4(_05986_),
    .ZN(_05987_));
 AND2_X1 _31184_ (.A1(_05853_),
    .A2(_05843_),
    .ZN(_05988_));
 AND2_X1 _31185_ (.A1(_05920_),
    .A2(_05988_),
    .ZN(_05989_));
 AND2_X1 _31186_ (.A1(_05849_),
    .A2(_05934_),
    .ZN(_05990_));
 AND2_X2 _31187_ (.A1(_05847_),
    .A2(_05878_),
    .ZN(_05991_));
 BUF_X2 _31188_ (.A(_05991_),
    .Z(_05992_));
 AND2_X1 _31189_ (.A1(_05992_),
    .A2(_05844_),
    .ZN(_05993_));
 NOR3_X1 _31190_ (.A1(_05989_),
    .A2(_05990_),
    .A3(_05993_),
    .ZN(_05994_));
 INV_X1 _31191_ (.A(_05925_),
    .ZN(_05996_));
 AND2_X4 _31192_ (.A1(_05889_),
    .A2(_05955_),
    .ZN(_05997_));
 INV_X1 _31193_ (.A(_05997_),
    .ZN(_05998_));
 BUF_X4 _31194_ (.A(_05842_),
    .Z(_05999_));
 NAND2_X1 _31195_ (.A1(_05887_),
    .A2(_05999_),
    .ZN(_06000_));
 AOI21_X1 _31196_ (.A(_05996_),
    .B1(_05998_),
    .B2(_06000_),
    .ZN(_06001_));
 BUF_X4 _31197_ (.A(_05903_),
    .Z(_06002_));
 NAND3_X1 _31198_ (.A1(_06002_),
    .A2(_05999_),
    .A3(_05864_),
    .ZN(_06003_));
 AND2_X2 _31199_ (.A1(_05857_),
    .A2(_05869_),
    .ZN(_06004_));
 INV_X1 _31200_ (.A(_06004_),
    .ZN(_06005_));
 INV_X4 _31201_ (.A(_05903_),
    .ZN(_06007_));
 OAI21_X1 _31202_ (.A(_06003_),
    .B1(_06005_),
    .B2(_06007_),
    .ZN(_06008_));
 AND2_X1 _31203_ (.A1(_05964_),
    .A2(_06002_),
    .ZN(_06009_));
 AND2_X2 _31204_ (.A1(_05869_),
    .A2(_05843_),
    .ZN(_06010_));
 AND3_X1 _31205_ (.A1(_06010_),
    .A2(_05902_),
    .A3(_05847_),
    .ZN(_06011_));
 NOR4_X1 _31206_ (.A1(_06001_),
    .A2(_06008_),
    .A3(_06009_),
    .A4(_06011_),
    .ZN(_06012_));
 AND4_X1 _31207_ (.A1(_05963_),
    .A2(_05987_),
    .A3(_05994_),
    .A4(_06012_),
    .ZN(_06013_));
 NAND4_X1 _31208_ (.A1(_05891_),
    .A2(_05932_),
    .A3(_05960_),
    .A4(_06013_),
    .ZN(_06014_));
 AND2_X2 _31209_ (.A1(_05892_),
    .A2(_05875_),
    .ZN(_06015_));
 AND2_X2 _31210_ (.A1(_05864_),
    .A2(_05955_),
    .ZN(_06016_));
 AND2_X1 _31211_ (.A1(_06015_),
    .A2(_06016_),
    .ZN(_06018_));
 AND2_X4 _31212_ (.A1(_06015_),
    .A2(_05967_),
    .ZN(_06019_));
 NAND2_X1 _31213_ (.A1(_05955_),
    .A2(_05900_),
    .ZN(_06020_));
 INV_X1 _31214_ (.A(_06020_),
    .ZN(_06021_));
 BUF_X2 _31215_ (.A(_06021_),
    .Z(_06022_));
 AOI211_X2 _31216_ (.A(_06018_),
    .B(_06019_),
    .C1(_06015_),
    .C2(_06022_),
    .ZN(_06023_));
 BUF_X4 _31217_ (.A(_06015_),
    .Z(_06024_));
 AND2_X2 _31218_ (.A1(_05842_),
    .A2(_05851_),
    .ZN(_06025_));
 OAI21_X1 _31219_ (.A(_06024_),
    .B1(_06025_),
    .B2(_05943_),
    .ZN(_06026_));
 AND2_X1 _31220_ (.A1(_05851_),
    .A2(_05870_),
    .ZN(_06027_));
 BUF_X4 _31221_ (.A(_06027_),
    .Z(_06029_));
 OAI21_X1 _31222_ (.A(_06024_),
    .B1(_06029_),
    .B2(_05934_),
    .ZN(_06030_));
 NAND3_X1 _31223_ (.A1(_06023_),
    .A2(_06026_),
    .A3(_06030_),
    .ZN(_06031_));
 AND2_X2 _31224_ (.A1(_05847_),
    .A2(_05875_),
    .ZN(_06032_));
 BUF_X2 _31225_ (.A(_06032_),
    .Z(_06033_));
 BUF_X4 _31226_ (.A(_16836_),
    .Z(_06034_));
 AND2_X1 _31227_ (.A1(_05884_),
    .A2(_06034_),
    .ZN(_06035_));
 AOI22_X1 _31228_ (.A1(_06033_),
    .A2(_06035_),
    .B1(_05936_),
    .B2(_05985_),
    .ZN(_06036_));
 INV_X1 _31229_ (.A(_05956_),
    .ZN(_06037_));
 OAI21_X1 _31230_ (.A(_06036_),
    .B1(_06037_),
    .B2(_05939_),
    .ZN(_06038_));
 OAI21_X1 _31231_ (.A(_05954_),
    .B1(_05887_),
    .B2(_16838_),
    .ZN(_06040_));
 AND3_X1 _31232_ (.A1(_05902_),
    .A2(_05837_),
    .A3(_05954_),
    .ZN(_06041_));
 AND2_X1 _31233_ (.A1(_06040_),
    .A2(_06041_),
    .ZN(_06042_));
 BUF_X2 _31234_ (.A(_05876_),
    .Z(_06043_));
 BUF_X2 _31235_ (.A(_05901_),
    .Z(_06044_));
 NAND2_X1 _31236_ (.A1(_06043_),
    .A2(_06044_),
    .ZN(_06045_));
 AND2_X1 _31237_ (.A1(_05956_),
    .A2(_06034_),
    .ZN(_06046_));
 INV_X1 _31238_ (.A(_06046_),
    .ZN(_06047_));
 OAI21_X1 _31239_ (.A(_06045_),
    .B1(_06047_),
    .B2(_05946_),
    .ZN(_06048_));
 NOR4_X1 _31240_ (.A1(_06031_),
    .A2(_06038_),
    .A3(_06042_),
    .A4(_06048_),
    .ZN(_06049_));
 OAI21_X1 _31241_ (.A(_05921_),
    .B1(_06029_),
    .B2(_05934_),
    .ZN(_06051_));
 NAND3_X1 _31242_ (.A1(_05967_),
    .A2(_05836_),
    .A3(_05880_),
    .ZN(_06052_));
 NAND2_X1 _31243_ (.A1(_06051_),
    .A2(_06052_),
    .ZN(_06053_));
 AND2_X2 _31244_ (.A1(_05893_),
    .A2(_05837_),
    .ZN(_06054_));
 BUF_X2 _31245_ (.A(_06054_),
    .Z(_06055_));
 AND2_X1 _31246_ (.A1(_05854_),
    .A2(_05850_),
    .ZN(_06056_));
 OAI21_X1 _31247_ (.A(_06055_),
    .B1(_06046_),
    .B2(_06056_),
    .ZN(_06057_));
 INV_X1 _31248_ (.A(_06054_),
    .ZN(_06058_));
 INV_X1 _31249_ (.A(_05864_),
    .ZN(_06059_));
 NAND2_X1 _31250_ (.A1(_06059_),
    .A2(_05842_),
    .ZN(_06060_));
 OAI21_X1 _31251_ (.A(_06057_),
    .B1(_06058_),
    .B2(_06060_),
    .ZN(_06062_));
 BUF_X2 _31252_ (.A(_05892_),
    .Z(_06063_));
 NAND3_X1 _31253_ (.A1(_06004_),
    .A2(_06063_),
    .A3(_05836_),
    .ZN(_06064_));
 INV_X4 _31254_ (.A(_05906_),
    .ZN(_06065_));
 OAI21_X1 _31255_ (.A(_06064_),
    .B1(_06065_),
    .B2(_06047_),
    .ZN(_06066_));
 NAND2_X1 _31256_ (.A1(_05887_),
    .A2(_05853_),
    .ZN(_06067_));
 NOR2_X1 _31257_ (.A1(_06007_),
    .A2(_06067_),
    .ZN(_06068_));
 NOR4_X1 _31258_ (.A1(_06053_),
    .A2(_06062_),
    .A3(_06066_),
    .A4(_06068_),
    .ZN(_06069_));
 AND2_X4 _31259_ (.A1(_05969_),
    .A2(_05849_),
    .ZN(_06070_));
 NAND2_X1 _31260_ (.A1(_05849_),
    .A2(_05997_),
    .ZN(_06071_));
 OAI21_X1 _31261_ (.A(_05854_),
    .B1(_05900_),
    .B2(_16836_),
    .ZN(_06073_));
 OAI21_X1 _31262_ (.A(_06071_),
    .B1(_06065_),
    .B2(_06073_),
    .ZN(_06074_));
 INV_X1 _31263_ (.A(_05927_),
    .ZN(_06075_));
 AND2_X1 _31264_ (.A1(_06075_),
    .A2(_06054_),
    .ZN(_06076_));
 OR3_X1 _31265_ (.A1(_06070_),
    .A2(_06074_),
    .A3(_06076_),
    .ZN(_06077_));
 OAI21_X1 _31266_ (.A(_05992_),
    .B1(_06004_),
    .B2(_06044_),
    .ZN(_06078_));
 NAND4_X1 _31267_ (.A1(_05889_),
    .A2(_05956_),
    .A3(_05847_),
    .A4(_05893_),
    .ZN(_06079_));
 NAND2_X1 _31268_ (.A1(_06078_),
    .A2(_06079_),
    .ZN(_06080_));
 INV_X1 _31269_ (.A(_05882_),
    .ZN(_06081_));
 NOR2_X1 _31270_ (.A1(_06081_),
    .A2(_06060_),
    .ZN(_06082_));
 OR2_X1 _31271_ (.A1(_06037_),
    .A2(_05889_),
    .ZN(_06084_));
 INV_X2 _31272_ (.A(_06032_),
    .ZN(_06085_));
 NOR2_X1 _31273_ (.A1(_06084_),
    .A2(_06085_),
    .ZN(_06086_));
 NOR4_X2 _31274_ (.A1(_06077_),
    .A2(_06080_),
    .A3(_06082_),
    .A4(_06086_),
    .ZN(_06087_));
 AND2_X1 _31275_ (.A1(_05915_),
    .A2(_06032_),
    .ZN(_06088_));
 BUF_X4 _31276_ (.A(_05838_),
    .Z(_06089_));
 INV_X1 _31277_ (.A(_06089_),
    .ZN(_06090_));
 AOI22_X1 _31278_ (.A1(_05975_),
    .A2(_05884_),
    .B1(_05956_),
    .B2(_06034_),
    .ZN(_06091_));
 NOR2_X1 _31279_ (.A1(_06090_),
    .A2(_06091_),
    .ZN(_06092_));
 INV_X1 _31280_ (.A(_05859_),
    .ZN(_06093_));
 INV_X1 _31281_ (.A(_05988_),
    .ZN(_06095_));
 NAND2_X1 _31282_ (.A1(_06093_),
    .A2(_06095_),
    .ZN(_06096_));
 AOI211_X4 _31283_ (.A(_06088_),
    .B(_06092_),
    .C1(_06096_),
    .C2(_06033_),
    .ZN(_06097_));
 NAND4_X1 _31284_ (.A1(_06049_),
    .A2(_06069_),
    .A3(_06087_),
    .A4(_06097_),
    .ZN(_06098_));
 NOR2_X2 _31285_ (.A1(_06014_),
    .A2(_06098_),
    .ZN(_06099_));
 INV_X1 _31286_ (.A(_06099_),
    .ZN(_06100_));
 INV_X32 _31287_ (.A(_16882_),
    .ZN(_06101_));
 NOR2_X1 _31288_ (.A1(_06101_),
    .A2(_16883_),
    .ZN(_06102_));
 BUF_X2 _31289_ (.A(_06102_),
    .Z(_06103_));
 INV_X32 _31290_ (.A(_16881_),
    .ZN(_06104_));
 NOR2_X4 _31291_ (.A1(_06104_),
    .A2(_16880_),
    .ZN(_06106_));
 BUF_X4 _31292_ (.A(_06106_),
    .Z(_06107_));
 AND2_X2 _31293_ (.A1(_06103_),
    .A2(_06107_),
    .ZN(_06108_));
 INV_X32 _31294_ (.A(_16878_),
    .ZN(_06109_));
 NOR2_X4 _31295_ (.A1(_06109_),
    .A2(_16879_),
    .ZN(_06110_));
 AND2_X4 _31296_ (.A1(_16876_),
    .A2(_16877_),
    .ZN(_06111_));
 AND2_X1 _31297_ (.A1(_06110_),
    .A2(_06111_),
    .ZN(_06112_));
 BUF_X2 _31298_ (.A(_06112_),
    .Z(_06113_));
 AND2_X1 _31299_ (.A1(_06108_),
    .A2(_06113_),
    .ZN(_06114_));
 INV_X1 _31300_ (.A(_06108_),
    .ZN(_06115_));
 INV_X32 _31301_ (.A(_16879_),
    .ZN(_06117_));
 NOR2_X1 _31302_ (.A1(_06117_),
    .A2(_16878_),
    .ZN(_06118_));
 INV_X32 _31303_ (.A(_16876_),
    .ZN(_06119_));
 NOR2_X4 _31304_ (.A1(_06119_),
    .A2(_16877_),
    .ZN(_06120_));
 AND2_X1 _31305_ (.A1(_06118_),
    .A2(_06120_),
    .ZN(_06121_));
 INV_X4 _31306_ (.A(_06121_),
    .ZN(_06122_));
 AND2_X4 _31307_ (.A1(_16879_),
    .A2(_16878_),
    .ZN(_06123_));
 BUF_X16 _31308_ (.A(_06123_),
    .Z(_06124_));
 AND2_X4 _31309_ (.A1(_06124_),
    .A2(_16877_),
    .ZN(_06125_));
 INV_X1 _31310_ (.A(_06125_),
    .ZN(_06126_));
 AOI21_X1 _31311_ (.A(_06115_),
    .B1(_06122_),
    .B2(_06126_),
    .ZN(_06128_));
 NOR2_X4 _31312_ (.A1(_16879_),
    .A2(_16878_),
    .ZN(_06129_));
 INV_X8 _31313_ (.A(_16877_),
    .ZN(_06130_));
 AND2_X1 _31314_ (.A1(_06129_),
    .A2(_06130_),
    .ZN(_06131_));
 AND2_X1 _31315_ (.A1(_06108_),
    .A2(_06131_),
    .ZN(_06132_));
 NAND2_X1 _31316_ (.A1(_06109_),
    .A2(_16877_),
    .ZN(_06133_));
 NOR2_X1 _31317_ (.A1(_06133_),
    .A2(_16879_),
    .ZN(_06134_));
 AND2_X1 _31318_ (.A1(_06108_),
    .A2(_06134_),
    .ZN(_06135_));
 OR4_X4 _31319_ (.A1(_06114_),
    .A2(_06128_),
    .A3(_06132_),
    .A4(_06135_),
    .ZN(_06136_));
 NOR2_X4 _31320_ (.A1(_16876_),
    .A2(_16877_),
    .ZN(_06137_));
 BUF_X4 _31321_ (.A(_06137_),
    .Z(_06139_));
 INV_X4 _31322_ (.A(_06139_),
    .ZN(_06140_));
 NAND2_X4 _31323_ (.A1(_06140_),
    .A2(_06124_),
    .ZN(_06141_));
 INV_X1 _31324_ (.A(_06141_),
    .ZN(_06142_));
 AND2_X4 _31325_ (.A1(_16881_),
    .A2(_16880_),
    .ZN(_06143_));
 AND2_X2 _31326_ (.A1(_06103_),
    .A2(_06143_),
    .ZN(_06144_));
 AND2_X1 _31327_ (.A1(_06142_),
    .A2(_06144_),
    .ZN(_06145_));
 AND2_X1 _31328_ (.A1(_06118_),
    .A2(_06130_),
    .ZN(_06146_));
 BUF_X2 _31329_ (.A(_06146_),
    .Z(_06147_));
 AND2_X1 _31330_ (.A1(_06144_),
    .A2(_06147_),
    .ZN(_06148_));
 BUF_X32 _31331_ (.A(_16876_),
    .Z(_06150_));
 NOR2_X4 _31332_ (.A1(_06130_),
    .A2(_06150_),
    .ZN(_06151_));
 AND2_X1 _31333_ (.A1(_06118_),
    .A2(_06151_),
    .ZN(_06152_));
 BUF_X4 _31334_ (.A(_06152_),
    .Z(_06153_));
 AND2_X1 _31335_ (.A1(_06153_),
    .A2(_06144_),
    .ZN(_06154_));
 OR2_X1 _31336_ (.A1(_06148_),
    .A2(_06154_),
    .ZN(_06155_));
 AND2_X2 _31337_ (.A1(_06110_),
    .A2(_06130_),
    .ZN(_06156_));
 AND2_X1 _31338_ (.A1(_06156_),
    .A2(_06144_),
    .ZN(_06157_));
 AND2_X1 _31339_ (.A1(_06112_),
    .A2(_06144_),
    .ZN(_06158_));
 AND2_X1 _31340_ (.A1(_06129_),
    .A2(_06150_),
    .ZN(_06159_));
 AND2_X1 _31341_ (.A1(_06144_),
    .A2(_06159_),
    .ZN(_06161_));
 OR3_X1 _31342_ (.A1(_06157_),
    .A2(_06158_),
    .A3(_06161_),
    .ZN(_06162_));
 NOR4_X1 _31343_ (.A1(_06136_),
    .A2(_06145_),
    .A3(_06155_),
    .A4(_06162_),
    .ZN(_06163_));
 AND2_X2 _31344_ (.A1(_06110_),
    .A2(_06139_),
    .ZN(_06164_));
 OR2_X1 _31345_ (.A1(_06164_),
    .A2(_06112_),
    .ZN(_06165_));
 AND2_X4 _31346_ (.A1(_06104_),
    .A2(_16880_),
    .ZN(_06166_));
 NOR2_X4 _31347_ (.A1(_16882_),
    .A2(_16883_),
    .ZN(_06167_));
 AND2_X1 _31348_ (.A1(_06166_),
    .A2(_06167_),
    .ZN(_06168_));
 BUF_X2 _31349_ (.A(_06168_),
    .Z(_06169_));
 AND2_X1 _31350_ (.A1(_06165_),
    .A2(_06169_),
    .ZN(_06170_));
 INV_X1 _31351_ (.A(_06170_),
    .ZN(_06172_));
 AND2_X4 _31352_ (.A1(_06151_),
    .A2(_06129_),
    .ZN(_06173_));
 OAI21_X1 _31353_ (.A(_06169_),
    .B1(_06173_),
    .B2(_06131_),
    .ZN(_06174_));
 NOR2_X1 _31354_ (.A1(_06133_),
    .A2(_06117_),
    .ZN(_06175_));
 OAI21_X1 _31355_ (.A(_06169_),
    .B1(_06147_),
    .B2(_06175_),
    .ZN(_06176_));
 AND2_X4 _31356_ (.A1(_06123_),
    .A2(_06111_),
    .ZN(_06177_));
 AND2_X2 _31357_ (.A1(_06124_),
    .A2(_06130_),
    .ZN(_06178_));
 OAI21_X1 _31358_ (.A(_06169_),
    .B1(_06177_),
    .B2(_06178_),
    .ZN(_06179_));
 AND4_X1 _31359_ (.A1(_06172_),
    .A2(_06174_),
    .A3(_06176_),
    .A4(_06179_),
    .ZN(_06180_));
 BUF_X4 _31360_ (.A(_06110_),
    .Z(_06181_));
 INV_X1 _31361_ (.A(_06181_),
    .ZN(_06183_));
 BUF_X4 _31362_ (.A(_06151_),
    .Z(_06184_));
 NOR2_X4 _31363_ (.A1(_06183_),
    .A2(_06184_),
    .ZN(_06185_));
 INV_X1 _31364_ (.A(_06120_),
    .ZN(_06186_));
 NOR2_X1 _31365_ (.A1(_16881_),
    .A2(_16880_),
    .ZN(_06187_));
 AND2_X2 _31366_ (.A1(_06187_),
    .A2(_06167_),
    .ZN(_06188_));
 BUF_X2 _31367_ (.A(_06188_),
    .Z(_06189_));
 NAND3_X1 _31368_ (.A1(_06185_),
    .A2(_06186_),
    .A3(_06189_),
    .ZN(_06190_));
 BUF_X4 _31369_ (.A(_06124_),
    .Z(_06191_));
 BUF_X4 _31370_ (.A(_06119_),
    .Z(_06192_));
 BUF_X4 _31371_ (.A(_06130_),
    .Z(_06194_));
 OAI211_X2 _31372_ (.A(_06188_),
    .B(_06191_),
    .C1(_06192_),
    .C2(_06194_),
    .ZN(_06195_));
 AND3_X1 _31373_ (.A1(_06180_),
    .A2(_06190_),
    .A3(_06195_),
    .ZN(_06196_));
 AND2_X1 _31374_ (.A1(_06166_),
    .A2(_06102_),
    .ZN(_06197_));
 BUF_X4 _31375_ (.A(_06197_),
    .Z(_06198_));
 AND2_X4 _31376_ (.A1(_06120_),
    .A2(_06110_),
    .ZN(_06199_));
 AND2_X1 _31377_ (.A1(_06151_),
    .A2(_06181_),
    .ZN(_06200_));
 BUF_X4 _31378_ (.A(_06200_),
    .Z(_06201_));
 OAI21_X1 _31379_ (.A(_06198_),
    .B1(_06199_),
    .B2(_06201_),
    .ZN(_06202_));
 BUF_X4 _31380_ (.A(_06166_),
    .Z(_06203_));
 BUF_X4 _31381_ (.A(_06150_),
    .Z(_06205_));
 BUF_X4 _31382_ (.A(_06129_),
    .Z(_06206_));
 NAND4_X1 _31383_ (.A1(_06203_),
    .A2(_06103_),
    .A3(_06205_),
    .A4(_06206_),
    .ZN(_06207_));
 AND2_X1 _31384_ (.A1(_06202_),
    .A2(_06207_),
    .ZN(_06208_));
 NOR3_X2 _31385_ (.A1(_06139_),
    .A2(_06117_),
    .A3(_16878_),
    .ZN(_06209_));
 INV_X1 _31386_ (.A(_06111_),
    .ZN(_06210_));
 BUF_X4 _31387_ (.A(_06210_),
    .Z(_06211_));
 AND2_X1 _31388_ (.A1(_06209_),
    .A2(_06211_),
    .ZN(_06212_));
 OAI21_X1 _31389_ (.A(_06198_),
    .B1(_06212_),
    .B2(_06177_),
    .ZN(_06213_));
 AND2_X2 _31390_ (.A1(_06103_),
    .A2(_06187_),
    .ZN(_06214_));
 BUF_X4 _31391_ (.A(_06214_),
    .Z(_06216_));
 AND2_X1 _31392_ (.A1(_06120_),
    .A2(_06129_),
    .ZN(_06217_));
 BUF_X2 _31393_ (.A(_06217_),
    .Z(_06218_));
 OAI21_X1 _31394_ (.A(_06216_),
    .B1(_06113_),
    .B2(_06218_),
    .ZN(_06219_));
 AND2_X2 _31395_ (.A1(_06124_),
    .A2(_06150_),
    .ZN(_06220_));
 OAI21_X1 _31396_ (.A(_06216_),
    .B1(_06220_),
    .B2(_06175_),
    .ZN(_06221_));
 AND4_X1 _31397_ (.A1(_06208_),
    .A2(_06213_),
    .A3(_06219_),
    .A4(_06221_),
    .ZN(_06222_));
 AND2_X1 _31398_ (.A1(_06106_),
    .A2(_06167_),
    .ZN(_06223_));
 INV_X2 _31399_ (.A(_06223_),
    .ZN(_06224_));
 NAND2_X1 _31400_ (.A1(_06210_),
    .A2(_06129_),
    .ZN(_06225_));
 NOR2_X1 _31401_ (.A1(_06224_),
    .A2(_06225_),
    .ZN(_06227_));
 AND2_X2 _31402_ (.A1(_06110_),
    .A2(_16877_),
    .ZN(_06228_));
 AND2_X1 _31403_ (.A1(_06228_),
    .A2(_06223_),
    .ZN(_06229_));
 AND2_X4 _31404_ (.A1(_06120_),
    .A2(_06124_),
    .ZN(_06230_));
 AND2_X4 _31405_ (.A1(_06223_),
    .A2(_06230_),
    .ZN(_06231_));
 AND3_X1 _31406_ (.A1(_06209_),
    .A2(_06167_),
    .A3(_06107_),
    .ZN(_06232_));
 OR4_X4 _31407_ (.A1(_06227_),
    .A2(_06229_),
    .A3(_06231_),
    .A4(_06232_),
    .ZN(_06233_));
 AND2_X2 _31408_ (.A1(_06143_),
    .A2(_06167_),
    .ZN(_06234_));
 BUF_X4 _31409_ (.A(_06234_),
    .Z(_06235_));
 BUF_X4 _31410_ (.A(_06235_),
    .Z(_06236_));
 AND2_X1 _31411_ (.A1(_06236_),
    .A2(_06159_),
    .ZN(_06238_));
 OAI211_X2 _31412_ (.A(_06236_),
    .B(_06191_),
    .C1(_06139_),
    .C2(_06184_),
    .ZN(_06239_));
 INV_X1 _31413_ (.A(_06175_),
    .ZN(_06240_));
 INV_X1 _31414_ (.A(_06235_),
    .ZN(_06241_));
 OAI21_X1 _31415_ (.A(_06239_),
    .B1(_06240_),
    .B2(_06241_),
    .ZN(_06242_));
 AND3_X1 _31416_ (.A1(_06235_),
    .A2(_06150_),
    .A3(_06181_),
    .ZN(_06243_));
 NOR4_X1 _31417_ (.A1(_06233_),
    .A2(_06238_),
    .A3(_06242_),
    .A4(_06243_),
    .ZN(_06244_));
 AND4_X1 _31418_ (.A1(_06163_),
    .A2(_06196_),
    .A3(_06222_),
    .A4(_06244_),
    .ZN(_06245_));
 AND2_X4 _31419_ (.A1(_16882_),
    .A2(_16883_),
    .ZN(_06246_));
 AND2_X2 _31420_ (.A1(_06106_),
    .A2(_06246_),
    .ZN(_06247_));
 BUF_X4 _31421_ (.A(_06247_),
    .Z(_06249_));
 AND2_X1 _31422_ (.A1(_06173_),
    .A2(_06249_),
    .ZN(_06250_));
 AND2_X1 _31423_ (.A1(_06199_),
    .A2(_06249_),
    .ZN(_06251_));
 AND2_X1 _31424_ (.A1(_06228_),
    .A2(_06249_),
    .ZN(_06252_));
 AND2_X1 _31425_ (.A1(_06249_),
    .A2(_06131_),
    .ZN(_06253_));
 OR4_X2 _31426_ (.A1(_06250_),
    .A2(_06251_),
    .A3(_06252_),
    .A4(_06253_),
    .ZN(_06254_));
 AND2_X4 _31427_ (.A1(_06246_),
    .A2(_06143_),
    .ZN(_06255_));
 BUF_X8 _31428_ (.A(_06255_),
    .Z(_06256_));
 BUF_X4 _31429_ (.A(_06256_),
    .Z(_06257_));
 AND2_X1 _31430_ (.A1(_06191_),
    .A2(_06119_),
    .ZN(_06258_));
 NAND2_X1 _31431_ (.A1(_06257_),
    .A2(_06258_),
    .ZN(_06260_));
 INV_X1 _31432_ (.A(_06256_),
    .ZN(_06261_));
 OAI21_X1 _31433_ (.A(_06260_),
    .B1(_06122_),
    .B2(_06261_),
    .ZN(_06262_));
 BUF_X4 _31434_ (.A(_06118_),
    .Z(_06263_));
 AND3_X1 _31435_ (.A1(_06249_),
    .A2(_06263_),
    .A3(_06186_),
    .ZN(_06264_));
 AND2_X4 _31436_ (.A1(_06124_),
    .A2(_06137_),
    .ZN(_06265_));
 AND2_X1 _31437_ (.A1(_06249_),
    .A2(_06265_),
    .ZN(_06266_));
 AND3_X1 _31438_ (.A1(_06177_),
    .A2(_06246_),
    .A3(_06107_),
    .ZN(_06267_));
 OR3_X1 _31439_ (.A1(_06264_),
    .A2(_06266_),
    .A3(_06267_),
    .ZN(_06268_));
 INV_X1 _31440_ (.A(_06156_),
    .ZN(_06269_));
 AOI21_X1 _31441_ (.A(_06261_),
    .B1(_06269_),
    .B2(_06225_),
    .ZN(_06271_));
 NOR4_X1 _31442_ (.A1(_06254_),
    .A2(_06262_),
    .A3(_06268_),
    .A4(_06271_),
    .ZN(_06272_));
 AND2_X2 _31443_ (.A1(_06246_),
    .A2(_06187_),
    .ZN(_06273_));
 BUF_X4 _31444_ (.A(_06273_),
    .Z(_06274_));
 AND2_X1 _31445_ (.A1(_06147_),
    .A2(_06274_),
    .ZN(_06275_));
 INV_X1 _31446_ (.A(_06275_),
    .ZN(_06276_));
 AND2_X1 _31447_ (.A1(_06166_),
    .A2(_06246_),
    .ZN(_06277_));
 BUF_X4 _31448_ (.A(_06277_),
    .Z(_06278_));
 AND2_X1 _31449_ (.A1(_06278_),
    .A2(_06173_),
    .ZN(_06279_));
 INV_X1 _31450_ (.A(_06279_),
    .ZN(_06280_));
 AND2_X1 _31451_ (.A1(_06278_),
    .A2(_06200_),
    .ZN(_06282_));
 INV_X1 _31452_ (.A(_06282_),
    .ZN(_06283_));
 AND2_X1 _31453_ (.A1(_06118_),
    .A2(_06111_),
    .ZN(_06284_));
 AND2_X1 _31454_ (.A1(_06277_),
    .A2(_06284_),
    .ZN(_06285_));
 INV_X1 _31455_ (.A(_06285_),
    .ZN(_06286_));
 OAI211_X2 _31456_ (.A(_06278_),
    .B(_06191_),
    .C1(_06205_),
    .C2(_06194_),
    .ZN(_06287_));
 AND4_X1 _31457_ (.A1(_06280_),
    .A2(_06283_),
    .A3(_06286_),
    .A4(_06287_),
    .ZN(_06288_));
 BUF_X16 _31458_ (.A(_06181_),
    .Z(_06289_));
 AND3_X1 _31459_ (.A1(_06289_),
    .A2(_06246_),
    .A3(_06187_),
    .ZN(_06290_));
 AND2_X2 _31460_ (.A1(_06137_),
    .A2(_06129_),
    .ZN(_06291_));
 AOI22_X1 _31461_ (.A1(_06290_),
    .A2(_06140_),
    .B1(_06291_),
    .B2(_06274_),
    .ZN(_06293_));
 BUF_X4 _31462_ (.A(_16877_),
    .Z(_06294_));
 OAI211_X2 _31463_ (.A(_06274_),
    .B(_06191_),
    .C1(_06205_),
    .C2(_06294_),
    .ZN(_06295_));
 AND4_X1 _31464_ (.A1(_06276_),
    .A2(_06288_),
    .A3(_06293_),
    .A4(_06295_),
    .ZN(_06296_));
 AND2_X4 _31465_ (.A1(_06101_),
    .A2(_16883_),
    .ZN(_06297_));
 BUF_X4 _31466_ (.A(_06297_),
    .Z(_06298_));
 OAI211_X2 _31467_ (.A(_06203_),
    .B(_06298_),
    .C1(_06228_),
    .C2(_06159_),
    .ZN(_06299_));
 AND2_X1 _31468_ (.A1(_06166_),
    .A2(_06297_),
    .ZN(_06300_));
 BUF_X4 _31469_ (.A(_06300_),
    .Z(_06301_));
 INV_X1 _31470_ (.A(_06177_),
    .ZN(_06302_));
 BUF_X4 _31471_ (.A(_06265_),
    .Z(_06304_));
 INV_X4 _31472_ (.A(_06304_),
    .ZN(_06305_));
 NAND2_X1 _31473_ (.A1(_06302_),
    .A2(_06305_),
    .ZN(_06306_));
 OAI21_X1 _31474_ (.A(_06301_),
    .B1(_06306_),
    .B2(_06212_),
    .ZN(_06307_));
 AND2_X1 _31475_ (.A1(_06297_),
    .A2(_06187_),
    .ZN(_06308_));
 BUF_X2 _31476_ (.A(_06308_),
    .Z(_06309_));
 AND2_X4 _31477_ (.A1(_06111_),
    .A2(_06129_),
    .ZN(_06310_));
 INV_X8 _31478_ (.A(_06310_),
    .ZN(_06311_));
 INV_X1 _31479_ (.A(_06291_),
    .ZN(_06312_));
 NAND2_X4 _31480_ (.A1(_06311_),
    .A2(_06312_),
    .ZN(_06313_));
 OAI21_X1 _31481_ (.A(_06309_),
    .B1(_06313_),
    .B2(_06199_),
    .ZN(_06315_));
 AND2_X1 _31482_ (.A1(_06308_),
    .A2(_06147_),
    .ZN(_06316_));
 INV_X1 _31483_ (.A(_06316_),
    .ZN(_06317_));
 AND4_X1 _31484_ (.A1(_06299_),
    .A2(_06307_),
    .A3(_06315_),
    .A4(_06317_),
    .ZN(_06318_));
 AND2_X4 _31485_ (.A1(_06297_),
    .A2(_06143_),
    .ZN(_06319_));
 AND2_X1 _31486_ (.A1(_06151_),
    .A2(_06123_),
    .ZN(_06320_));
 AND2_X1 _31487_ (.A1(_06319_),
    .A2(_06320_),
    .ZN(_06321_));
 AND2_X1 _31488_ (.A1(_06319_),
    .A2(_06175_),
    .ZN(_06322_));
 NOR2_X1 _31489_ (.A1(_06321_),
    .A2(_06322_),
    .ZN(_06323_));
 AND2_X4 _31490_ (.A1(_06297_),
    .A2(_06106_),
    .ZN(_06324_));
 BUF_X2 _31491_ (.A(_06324_),
    .Z(_06326_));
 AND2_X1 _31492_ (.A1(_06326_),
    .A2(_06291_),
    .ZN(_06327_));
 INV_X1 _31493_ (.A(_06327_),
    .ZN(_06328_));
 OAI221_X1 _31494_ (.A(_06326_),
    .B1(_06192_),
    .B2(_06194_),
    .C1(_06191_),
    .C2(_06263_),
    .ZN(_06329_));
 BUF_X4 _31495_ (.A(_06319_),
    .Z(_06330_));
 BUF_X4 _31496_ (.A(_06131_),
    .Z(_06331_));
 OAI21_X1 _31497_ (.A(_06330_),
    .B1(_06185_),
    .B2(_06331_),
    .ZN(_06332_));
 AND4_X1 _31498_ (.A1(_06323_),
    .A2(_06328_),
    .A3(_06329_),
    .A4(_06332_),
    .ZN(_06333_));
 AND4_X2 _31499_ (.A1(_06272_),
    .A2(_06296_),
    .A3(_06318_),
    .A4(_06333_),
    .ZN(_06334_));
 AND2_X2 _31500_ (.A1(_06245_),
    .A2(_06334_),
    .ZN(_06335_));
 BUF_X8 _31501_ (.A(_06335_),
    .Z(_06337_));
 XNOR2_X1 _31502_ (.A(_06100_),
    .B(_06337_),
    .ZN(_06338_));
 XNOR2_X1 _31503_ (.A(_05833_),
    .B(_06338_),
    .ZN(_06339_));
 MUX2_X1 _31504_ (.A(_05207_),
    .B(_06339_),
    .S(_05156_),
    .Z(_00700_));
 MUX2_X1 _31505_ (.A(_17135_),
    .B(_17007_),
    .S(_05205_),
    .Z(_00855_));
 MUX2_X1 _31506_ (.A(_17136_),
    .B(_17008_),
    .S(_05205_),
    .Z(_00856_));
 MUX2_X1 _31507_ (.A(_17137_),
    .B(_17009_),
    .S(_05205_),
    .Z(_00857_));
 MUX2_X1 _31508_ (.A(_17138_),
    .B(_17010_),
    .S(_05205_),
    .Z(_00858_));
 MUX2_X1 _31509_ (.A(_17013_),
    .B(_16885_),
    .S(_05205_),
    .Z(_00733_));
 BUF_X4 _31510_ (.A(_05189_),
    .Z(_06340_));
 MUX2_X1 _31511_ (.A(_17014_),
    .B(_16886_),
    .S(_06340_),
    .Z(_00734_));
 MUX2_X1 _31512_ (.A(_17015_),
    .B(_16887_),
    .S(_06340_),
    .Z(_00735_));
 MUX2_X1 _31513_ (.A(_17016_),
    .B(_16888_),
    .S(_06340_),
    .Z(_00736_));
 MUX2_X1 _31514_ (.A(_17017_),
    .B(_16889_),
    .S(_06340_),
    .Z(_00737_));
 MUX2_X1 _31515_ (.A(_17018_),
    .B(_16890_),
    .S(_06340_),
    .Z(_00738_));
 XOR2_X1 _31516_ (.A(_17187_),
    .B(_17136_),
    .Z(_06342_));
 NAND2_X1 _31517_ (.A1(_05694_),
    .A2(_05587_),
    .ZN(_06343_));
 INV_X1 _31518_ (.A(_06343_),
    .ZN(_06344_));
 OAI21_X1 _31519_ (.A(_05683_),
    .B1(_06344_),
    .B2(_05685_),
    .ZN(_06345_));
 NAND2_X1 _31520_ (.A1(_06344_),
    .A2(_05708_),
    .ZN(_06346_));
 INV_X1 _31521_ (.A(_05661_),
    .ZN(_06348_));
 INV_X1 _31522_ (.A(_05799_),
    .ZN(_06349_));
 AOI21_X1 _31523_ (.A(_05717_),
    .B1(_06348_),
    .B2(_06349_),
    .ZN(_06350_));
 AOI211_X2 _31524_ (.A(_05730_),
    .B(_06350_),
    .C1(_05631_),
    .C2(_05716_),
    .ZN(_06351_));
 NAND4_X1 _31525_ (.A1(_05745_),
    .A2(_05817_),
    .A3(_05675_),
    .A4(_05624_),
    .ZN(_06352_));
 BUF_X4 _31526_ (.A(_05716_),
    .Z(_06353_));
 INV_X1 _31527_ (.A(_05723_),
    .ZN(_06354_));
 OAI21_X1 _31528_ (.A(_06353_),
    .B1(_06354_),
    .B2(_05666_),
    .ZN(_06355_));
 AND4_X1 _31529_ (.A1(_06346_),
    .A2(_06351_),
    .A3(_06352_),
    .A4(_06355_),
    .ZN(_06356_));
 OAI211_X2 _31530_ (.A(_05683_),
    .B(_05579_),
    .C1(_05712_),
    .C2(_05578_),
    .ZN(_06357_));
 AND2_X1 _31531_ (.A1(_05699_),
    .A2(_05646_),
    .ZN(_06359_));
 INV_X1 _31532_ (.A(_05691_),
    .ZN(_06360_));
 INV_X2 _31533_ (.A(_05631_),
    .ZN(_06361_));
 AOI21_X1 _31534_ (.A(_06360_),
    .B1(_06361_),
    .B2(_05680_),
    .ZN(_06362_));
 AND2_X1 _31535_ (.A1(_05589_),
    .A2(_05596_),
    .ZN(_06363_));
 AOI211_X4 _31536_ (.A(_06359_),
    .B(_06362_),
    .C1(_05699_),
    .C2(_06363_),
    .ZN(_06364_));
 AND4_X2 _31537_ (.A1(_06345_),
    .A2(_06356_),
    .A3(_06357_),
    .A4(_06364_),
    .ZN(_06365_));
 INV_X1 _31538_ (.A(_05576_),
    .ZN(_06366_));
 AOI21_X1 _31539_ (.A(_06366_),
    .B1(_06349_),
    .B2(_05680_),
    .ZN(_06367_));
 INV_X1 _31540_ (.A(_05796_),
    .ZN(_06368_));
 AOI21_X1 _31541_ (.A(_06366_),
    .B1(_06361_),
    .B2(_06368_),
    .ZN(_06370_));
 BUF_X4 _31542_ (.A(_05589_),
    .Z(_06371_));
 AND3_X1 _31543_ (.A1(_05576_),
    .A2(_06371_),
    .A3(_05694_),
    .ZN(_06372_));
 CLKBUF_X2 _31544_ (.A(_05573_),
    .Z(_06373_));
 AND4_X1 _31545_ (.A1(_05818_),
    .A2(_06373_),
    .A3(_05817_),
    .A4(_05827_),
    .ZN(_06374_));
 NOR4_X1 _31546_ (.A1(_06367_),
    .A2(_06370_),
    .A3(_06372_),
    .A4(_06374_),
    .ZN(_06375_));
 AOI21_X1 _31547_ (.A(_05626_),
    .B1(_06361_),
    .B2(_05680_),
    .ZN(_06376_));
 INV_X1 _31548_ (.A(_05684_),
    .ZN(_06377_));
 INV_X1 _31549_ (.A(_05763_),
    .ZN(_06378_));
 AOI21_X1 _31550_ (.A(_05626_),
    .B1(_06377_),
    .B2(_06378_),
    .ZN(_06379_));
 BUF_X2 _31551_ (.A(_05608_),
    .Z(_06381_));
 AOI211_X4 _31552_ (.A(_06376_),
    .B(_06379_),
    .C1(_06381_),
    .C2(_06363_),
    .ZN(_06382_));
 BUF_X4 _31553_ (.A(_05637_),
    .Z(_06383_));
 AND2_X2 _31554_ (.A1(_05738_),
    .A2(_05807_),
    .ZN(_06384_));
 NAND2_X1 _31555_ (.A1(_06383_),
    .A2(_06384_),
    .ZN(_06385_));
 AND2_X2 _31556_ (.A1(_05586_),
    .A2(_05620_),
    .ZN(_06386_));
 AND2_X2 _31557_ (.A1(_05581_),
    .A2(_05591_),
    .ZN(_06387_));
 OAI21_X1 _31558_ (.A(_06383_),
    .B1(_06386_),
    .B2(_06387_),
    .ZN(_06388_));
 INV_X1 _31559_ (.A(_05594_),
    .ZN(_06389_));
 NOR2_X2 _31560_ (.A1(_06389_),
    .A2(_05629_),
    .ZN(_06390_));
 BUF_X4 _31561_ (.A(_05636_),
    .Z(_06392_));
 NAND4_X1 _31562_ (.A1(_06390_),
    .A2(_06392_),
    .A3(_05745_),
    .A4(_06373_),
    .ZN(_06393_));
 NAND2_X1 _31563_ (.A1(_06383_),
    .A2(_05800_),
    .ZN(_06394_));
 AND4_X1 _31564_ (.A1(_06385_),
    .A2(_06388_),
    .A3(_06393_),
    .A4(_06394_),
    .ZN(_06395_));
 AND2_X1 _31565_ (.A1(_05767_),
    .A2(_05655_),
    .ZN(_06396_));
 AND2_X1 _31566_ (.A1(_05581_),
    .A2(_05638_),
    .ZN(_06397_));
 NAND2_X1 _31567_ (.A1(_05655_),
    .A2(_06397_),
    .ZN(_06398_));
 NAND4_X1 _31568_ (.A1(_05587_),
    .A2(_05573_),
    .A3(_05726_),
    .A4(_05651_),
    .ZN(_06399_));
 NAND2_X1 _31569_ (.A1(_06398_),
    .A2(_06399_),
    .ZN(_06400_));
 NAND2_X1 _31570_ (.A1(_05592_),
    .A2(_05600_),
    .ZN(_06401_));
 NOR2_X1 _31571_ (.A1(_06401_),
    .A2(_05620_),
    .ZN(_06403_));
 AOI211_X4 _31572_ (.A(_06396_),
    .B(_06400_),
    .C1(_05656_),
    .C2(_06403_),
    .ZN(_06404_));
 AND4_X1 _31573_ (.A1(_06375_),
    .A2(_06382_),
    .A3(_06395_),
    .A4(_06404_),
    .ZN(_06405_));
 AND2_X1 _31574_ (.A1(_05770_),
    .A2(_05684_),
    .ZN(_06406_));
 AND2_X1 _31575_ (.A1(_05771_),
    .A2(_05794_),
    .ZN(_06407_));
 AOI211_X4 _31576_ (.A(_06406_),
    .B(_06407_),
    .C1(_05763_),
    .C2(_05771_),
    .ZN(_06408_));
 AND3_X1 _31577_ (.A1(_05796_),
    .A2(_05651_),
    .A3(_05735_),
    .ZN(_06409_));
 AND3_X1 _31578_ (.A1(_05631_),
    .A2(_05651_),
    .A3(_05735_),
    .ZN(_06410_));
 AOI211_X4 _31579_ (.A(_06409_),
    .B(_06410_),
    .C1(_05639_),
    .C2(_05751_),
    .ZN(_06411_));
 OAI21_X1 _31580_ (.A(_05751_),
    .B1(_05719_),
    .B2(_05760_),
    .ZN(_06412_));
 INV_X1 _31581_ (.A(_05770_),
    .ZN(_06414_));
 OR2_X1 _31582_ (.A1(_06414_),
    .A2(_05627_),
    .ZN(_06415_));
 NAND4_X1 _31583_ (.A1(_06408_),
    .A2(_06411_),
    .A3(_06412_),
    .A4(_06415_),
    .ZN(_06416_));
 INV_X1 _31584_ (.A(_05757_),
    .ZN(_06417_));
 NOR2_X1 _31585_ (.A1(_06417_),
    .A2(_05749_),
    .ZN(_06418_));
 AND4_X1 _31586_ (.A1(_05630_),
    .A2(_05735_),
    .A3(_05722_),
    .A4(_05677_),
    .ZN(_06419_));
 OR2_X1 _31587_ (.A1(_06418_),
    .A2(_06419_),
    .ZN(_06420_));
 INV_X1 _31588_ (.A(_06401_),
    .ZN(_06421_));
 NAND3_X1 _31589_ (.A1(_06421_),
    .A2(_05758_),
    .A3(_05694_),
    .ZN(_06422_));
 INV_X1 _31590_ (.A(_05641_),
    .ZN(_06423_));
 OAI21_X1 _31591_ (.A(_06422_),
    .B1(_06423_),
    .B2(_06417_),
    .ZN(_06425_));
 AND2_X1 _31592_ (.A1(_05755_),
    .A2(_05762_),
    .ZN(_06426_));
 AND2_X1 _31593_ (.A1(_05755_),
    .A2(_05799_),
    .ZN(_06427_));
 AND2_X1 _31594_ (.A1(_05755_),
    .A2(_05672_),
    .ZN(_06428_));
 AND2_X1 _31595_ (.A1(_05755_),
    .A2(_05611_),
    .ZN(_06429_));
 OR4_X2 _31596_ (.A1(_06426_),
    .A2(_06427_),
    .A3(_06428_),
    .A4(_06429_),
    .ZN(_06430_));
 NOR4_X1 _31597_ (.A1(_06416_),
    .A2(_06420_),
    .A3(_06425_),
    .A4(_06430_),
    .ZN(_06431_));
 AND4_X1 _31598_ (.A1(_05636_),
    .A2(_05601_),
    .A3(_05630_),
    .A4(_05789_),
    .ZN(_06432_));
 AND3_X1 _31599_ (.A1(_05711_),
    .A2(_05636_),
    .A3(_05789_),
    .ZN(_06433_));
 AOI211_X4 _31600_ (.A(_06432_),
    .B(_06433_),
    .C1(_05792_),
    .C2(_05641_),
    .ZN(_06434_));
 NAND4_X1 _31601_ (.A1(_06392_),
    .A2(_05818_),
    .A3(_05809_),
    .A4(_05817_),
    .ZN(_06436_));
 BUF_X2 _31602_ (.A(_05792_),
    .Z(_06437_));
 OAI21_X1 _31603_ (.A(_06437_),
    .B1(_05794_),
    .B2(_05613_),
    .ZN(_06438_));
 AND3_X1 _31604_ (.A1(_06434_),
    .A2(_06436_),
    .A3(_06438_),
    .ZN(_06439_));
 AND3_X2 _31605_ (.A1(_06390_),
    .A2(_05779_),
    .A3(_05744_),
    .ZN(_06440_));
 AOI211_X4 _31606_ (.A(_05602_),
    .B(_05780_),
    .C1(_05712_),
    .C2(_05638_),
    .ZN(_06441_));
 BUF_X4 _31607_ (.A(_05779_),
    .Z(_06442_));
 AOI211_X4 _31608_ (.A(_06440_),
    .B(_06441_),
    .C1(_05719_),
    .C2(_06442_),
    .ZN(_06443_));
 OAI21_X1 _31609_ (.A(_05804_),
    .B1(_05623_),
    .B2(_06387_),
    .ZN(_06444_));
 INV_X1 _31610_ (.A(_05666_),
    .ZN(_06445_));
 OAI21_X1 _31611_ (.A(_06444_),
    .B1(_06445_),
    .B2(_05811_),
    .ZN(_06447_));
 NAND2_X1 _31612_ (.A1(_05804_),
    .A2(_05711_),
    .ZN(_06448_));
 INV_X1 _31613_ (.A(_05713_),
    .ZN(_06449_));
 OAI21_X1 _31614_ (.A(_06448_),
    .B1(_06449_),
    .B2(_05811_),
    .ZN(_06450_));
 BUF_X4 _31615_ (.A(_05804_),
    .Z(_06451_));
 AND2_X1 _31616_ (.A1(_05661_),
    .A2(_06451_),
    .ZN(_06452_));
 NOR3_X1 _31617_ (.A1(_06447_),
    .A2(_06450_),
    .A3(_06452_),
    .ZN(_06453_));
 AND2_X1 _31618_ (.A1(_05609_),
    .A2(_05815_),
    .ZN(_06454_));
 BUF_X4 _31619_ (.A(_05815_),
    .Z(_06455_));
 BUF_X2 _31620_ (.A(_05713_),
    .Z(_06456_));
 AND2_X1 _31621_ (.A1(_06455_),
    .A2(_06456_),
    .ZN(_06458_));
 AND4_X1 _31622_ (.A1(_05809_),
    .A2(_05807_),
    .A3(_05589_),
    .A4(_05652_),
    .ZN(_06459_));
 AND4_X1 _31623_ (.A1(_05809_),
    .A2(_05738_),
    .A3(_05620_),
    .A4(_05652_),
    .ZN(_06460_));
 NOR4_X1 _31624_ (.A1(_06454_),
    .A2(_06458_),
    .A3(_06459_),
    .A4(_06460_),
    .ZN(_06461_));
 AND4_X1 _31625_ (.A1(_06439_),
    .A2(_06443_),
    .A3(_06453_),
    .A4(_06461_),
    .ZN(_06462_));
 NAND4_X1 _31626_ (.A1(_06365_),
    .A2(_06405_),
    .A3(_06431_),
    .A4(_06462_),
    .ZN(_06463_));
 NOR2_X2 _31627_ (.A1(_06463_),
    .A2(_05829_),
    .ZN(_06464_));
 AND4_X1 _31628_ (.A1(_05232_),
    .A2(_05441_),
    .A3(_05240_),
    .A4(_05329_),
    .ZN(_06465_));
 NOR2_X1 _31629_ (.A1(_05443_),
    .A2(_06465_),
    .ZN(_06466_));
 NAND2_X1 _31630_ (.A1(_05496_),
    .A2(_05261_),
    .ZN(_06467_));
 AND3_X1 _31631_ (.A1(_05352_),
    .A2(_05417_),
    .A3(_05282_),
    .ZN(_06469_));
 AND2_X1 _31632_ (.A1(_05424_),
    .A2(_05257_),
    .ZN(_06470_));
 AND2_X2 _31633_ (.A1(_05228_),
    .A2(_05254_),
    .ZN(_06471_));
 AOI211_X2 _31634_ (.A(_06469_),
    .B(_06470_),
    .C1(_06471_),
    .C2(_05496_),
    .ZN(_06472_));
 INV_X1 _31635_ (.A(_05319_),
    .ZN(_06473_));
 OAI21_X1 _31636_ (.A(_05498_),
    .B1(_06473_),
    .B2(_05402_),
    .ZN(_06474_));
 OAI21_X1 _31637_ (.A(_05498_),
    .B1(_05473_),
    .B2(_05447_),
    .ZN(_06475_));
 AND4_X1 _31638_ (.A1(_06467_),
    .A2(_06472_),
    .A3(_06474_),
    .A4(_06475_),
    .ZN(_06476_));
 OAI21_X1 _31639_ (.A(_05444_),
    .B1(_05480_),
    .B2(_05211_),
    .ZN(_06477_));
 AND2_X1 _31640_ (.A1(_05419_),
    .A2(_05497_),
    .ZN(_06478_));
 AND2_X1 _31641_ (.A1(_05341_),
    .A2(_05419_),
    .ZN(_06480_));
 AND2_X1 _31642_ (.A1(_05418_),
    .A2(_05252_),
    .ZN(_06481_));
 AND2_X1 _31643_ (.A1(_05419_),
    .A2(_05307_),
    .ZN(_06482_));
 NOR4_X1 _31644_ (.A1(_06478_),
    .A2(_06480_),
    .A3(_06481_),
    .A4(_06482_),
    .ZN(_06483_));
 AND4_X1 _31645_ (.A1(_06466_),
    .A2(_06476_),
    .A3(_06477_),
    .A4(_06483_),
    .ZN(_06484_));
 AND2_X1 _31646_ (.A1(_05314_),
    .A2(_05245_),
    .ZN(_06485_));
 INV_X1 _31647_ (.A(_05244_),
    .ZN(_06486_));
 OAI21_X1 _31648_ (.A(_05259_),
    .B1(_06486_),
    .B2(_05274_),
    .ZN(_06487_));
 BUF_X2 _31649_ (.A(_05245_),
    .Z(_06488_));
 AOI211_X4 _31650_ (.A(_06485_),
    .B(_06487_),
    .C1(_05252_),
    .C2(_06488_),
    .ZN(_06489_));
 INV_X1 _31651_ (.A(_05250_),
    .ZN(_06491_));
 AOI211_X4 _31652_ (.A(_06491_),
    .B(_05235_),
    .C1(_05246_),
    .C2(_05446_),
    .ZN(_06492_));
 NOR2_X1 _31653_ (.A1(_05235_),
    .A2(_05241_),
    .ZN(_06493_));
 INV_X1 _31654_ (.A(_05224_),
    .ZN(_06494_));
 AOI21_X1 _31655_ (.A(_05235_),
    .B1(_05326_),
    .B2(_06494_),
    .ZN(_06495_));
 NOR4_X1 _31656_ (.A1(_06492_),
    .A2(_05506_),
    .A3(_06493_),
    .A4(_06495_),
    .ZN(_06496_));
 AND2_X1 _31657_ (.A1(_05267_),
    .A2(_05383_),
    .ZN(_06497_));
 INV_X1 _31658_ (.A(_05314_),
    .ZN(_06498_));
 AOI21_X1 _31659_ (.A(_05278_),
    .B1(_06498_),
    .B2(_05326_),
    .ZN(_06499_));
 AND2_X1 _31660_ (.A1(_05229_),
    .A2(_05446_),
    .ZN(_06500_));
 AOI211_X4 _31661_ (.A(_06497_),
    .B(_06499_),
    .C1(_06500_),
    .C2(_05270_),
    .ZN(_06502_));
 BUF_X4 _31662_ (.A(_05289_),
    .Z(_06503_));
 INV_X1 _31663_ (.A(_05274_),
    .ZN(_06504_));
 OAI21_X1 _31664_ (.A(_06503_),
    .B1(_06504_),
    .B2(_05435_),
    .ZN(_06505_));
 AND4_X1 _31665_ (.A1(_06489_),
    .A2(_06496_),
    .A3(_06502_),
    .A4(_06505_),
    .ZN(_06506_));
 AND2_X1 _31666_ (.A1(_05394_),
    .A2(_05311_),
    .ZN(_06507_));
 INV_X1 _31667_ (.A(_06507_),
    .ZN(_06508_));
 NAND2_X1 _31668_ (.A1(_05395_),
    .A2(_05521_),
    .ZN(_06509_));
 OAI21_X1 _31669_ (.A(_05395_),
    .B1(_05493_),
    .B2(_05337_),
    .ZN(_06510_));
 OAI21_X1 _31670_ (.A(_05395_),
    .B1(_05211_),
    .B2(_05296_),
    .ZN(_06511_));
 NAND4_X1 _31671_ (.A1(_06508_),
    .A2(_06509_),
    .A3(_06510_),
    .A4(_06511_),
    .ZN(_06513_));
 BUF_X4 _31672_ (.A(_05230_),
    .Z(_06514_));
 NAND4_X1 _31673_ (.A1(_06514_),
    .A2(_05384_),
    .A3(_05275_),
    .A4(_05233_),
    .ZN(_06515_));
 NAND3_X1 _31674_ (.A1(_05375_),
    .A2(_05290_),
    .A3(_05273_),
    .ZN(_06516_));
 NAND4_X1 _31675_ (.A1(_05562_),
    .A2(_05553_),
    .A3(_06515_),
    .A4(_06516_),
    .ZN(_06517_));
 OAI21_X1 _31676_ (.A(_05392_),
    .B1(_05371_),
    .B2(_05318_),
    .ZN(_06518_));
 NAND2_X1 _31677_ (.A1(_06504_),
    .A2(_05392_),
    .ZN(_06519_));
 BUF_X4 _31678_ (.A(_05250_),
    .Z(_06520_));
 NAND3_X1 _31679_ (.A1(_05384_),
    .A2(_06520_),
    .A3(_05329_),
    .ZN(_06521_));
 BUF_X4 _31680_ (.A(_05248_),
    .Z(_06522_));
 NAND4_X1 _31681_ (.A1(_05384_),
    .A2(_06522_),
    .A3(_05240_),
    .A4(_05329_),
    .ZN(_06524_));
 NAND4_X1 _31682_ (.A1(_06518_),
    .A2(_06519_),
    .A3(_06521_),
    .A4(_06524_),
    .ZN(_06525_));
 OAI21_X1 _31683_ (.A(_05413_),
    .B1(_05371_),
    .B2(_05360_),
    .ZN(_06526_));
 OAI21_X1 _31684_ (.A(_05413_),
    .B1(_05353_),
    .B2(_05356_),
    .ZN(_06527_));
 INV_X1 _31685_ (.A(_06500_),
    .ZN(_06528_));
 OAI211_X2 _31686_ (.A(_06526_),
    .B(_06527_),
    .C1(_06528_),
    .C2(_05406_),
    .ZN(_06529_));
 NOR4_X1 _31687_ (.A1(_06513_),
    .A2(_06517_),
    .A3(_06525_),
    .A4(_06529_),
    .ZN(_06530_));
 BUF_X4 _31688_ (.A(_05305_),
    .Z(_06531_));
 NAND3_X1 _31689_ (.A1(_06531_),
    .A2(_05246_),
    .A3(_05230_),
    .ZN(_06532_));
 OAI211_X2 _31690_ (.A(_05306_),
    .B(_06532_),
    .C1(_05408_),
    .C2(_05320_),
    .ZN(_06533_));
 AOI21_X1 _31691_ (.A(_05320_),
    .B1(_05458_),
    .B2(_05459_),
    .ZN(_06535_));
 AND4_X1 _31692_ (.A1(_05265_),
    .A2(_06520_),
    .A3(_05232_),
    .A4(_05303_),
    .ZN(_06536_));
 NOR3_X1 _31693_ (.A1(_06533_),
    .A2(_06535_),
    .A3(_06536_),
    .ZN(_06537_));
 AND4_X1 _31694_ (.A1(_05272_),
    .A2(_05250_),
    .A3(_05212_),
    .A4(_05303_),
    .ZN(_06538_));
 INV_X1 _31695_ (.A(_05473_),
    .ZN(_06539_));
 AOI21_X1 _31696_ (.A(_05364_),
    .B1(_06539_),
    .B2(_05504_),
    .ZN(_06540_));
 BUF_X4 _31697_ (.A(_05297_),
    .Z(_06541_));
 AOI211_X4 _31698_ (.A(_06538_),
    .B(_06540_),
    .C1(_06541_),
    .C2(_05354_),
    .ZN(_06542_));
 OAI21_X1 _31699_ (.A(_05564_),
    .B1(_05339_),
    .B2(_05381_),
    .ZN(_06543_));
 NAND2_X1 _31700_ (.A1(_05373_),
    .A2(_05564_),
    .ZN(_06544_));
 NAND2_X1 _31701_ (.A1(_05296_),
    .A2(_05564_),
    .ZN(_06546_));
 AND4_X1 _31702_ (.A1(_05472_),
    .A2(_06543_),
    .A3(_06544_),
    .A4(_06546_),
    .ZN(_06547_));
 BUF_X4 _31703_ (.A(_05333_),
    .Z(_06548_));
 AND2_X1 _31704_ (.A1(_06548_),
    .A2(_05497_),
    .ZN(_06549_));
 AND3_X1 _31705_ (.A1(_05521_),
    .A2(_05283_),
    .A3(_05303_),
    .ZN(_06550_));
 AND2_X1 _31706_ (.A1(_05473_),
    .A2(_05333_),
    .ZN(_06551_));
 NOR4_X1 _31707_ (.A1(_05461_),
    .A2(_06549_),
    .A3(_06550_),
    .A4(_06551_),
    .ZN(_06552_));
 AND4_X1 _31708_ (.A1(_06537_),
    .A2(_06542_),
    .A3(_06547_),
    .A4(_06552_),
    .ZN(_06553_));
 NAND4_X1 _31709_ (.A1(_06484_),
    .A2(_06506_),
    .A3(_06530_),
    .A4(_06553_),
    .ZN(_06554_));
 NOR2_X4 _31710_ (.A1(_06554_),
    .A2(_05454_),
    .ZN(_06555_));
 XOR2_X2 _31711_ (.A(_06464_),
    .B(_06555_),
    .Z(_06557_));
 XNOR2_X1 _31712_ (.A(_06557_),
    .B(_05571_),
    .ZN(_06558_));
 AND2_X1 _31713_ (.A1(_06278_),
    .A2(_06147_),
    .ZN(_06559_));
 NAND2_X1 _31714_ (.A1(_06278_),
    .A2(_06153_),
    .ZN(_06560_));
 INV_X1 _31715_ (.A(_06284_),
    .ZN(_06561_));
 INV_X8 _31716_ (.A(_06278_),
    .ZN(_06562_));
 OAI21_X1 _31717_ (.A(_06560_),
    .B1(_06561_),
    .B2(_06562_),
    .ZN(_06563_));
 NOR2_X1 _31718_ (.A1(_06141_),
    .A2(_06111_),
    .ZN(_06564_));
 AOI211_X2 _31719_ (.A(_06559_),
    .B(_06563_),
    .C1(_06278_),
    .C2(_06564_),
    .ZN(_06565_));
 AND2_X1 _31720_ (.A1(_06178_),
    .A2(_06273_),
    .ZN(_06566_));
 AND2_X2 _31721_ (.A1(_06263_),
    .A2(_06150_),
    .ZN(_06568_));
 AND2_X1 _31722_ (.A1(_06125_),
    .A2(_06273_),
    .ZN(_06569_));
 AOI221_X1 _31723_ (.A(_06566_),
    .B1(_06568_),
    .B2(_06274_),
    .C1(_06192_),
    .C2(_06569_),
    .ZN(_06570_));
 NAND3_X1 _31724_ (.A1(_06274_),
    .A2(_06184_),
    .A3(_06206_),
    .ZN(_06571_));
 BUF_X4 _31725_ (.A(_06278_),
    .Z(_06572_));
 OAI21_X1 _31726_ (.A(_06572_),
    .B1(_06199_),
    .B2(_06173_),
    .ZN(_06573_));
 NAND4_X1 _31727_ (.A1(_06565_),
    .A2(_06570_),
    .A3(_06571_),
    .A4(_06573_),
    .ZN(_06574_));
 AND2_X1 _31728_ (.A1(_06249_),
    .A2(_06220_),
    .ZN(_06575_));
 AND2_X4 _31729_ (.A1(_06164_),
    .A2(_06256_),
    .ZN(_06576_));
 INV_X2 _31730_ (.A(_06576_),
    .ZN(_06577_));
 OAI211_X2 _31731_ (.A(_06256_),
    .B(_06129_),
    .C1(_06205_),
    .C2(_06294_),
    .ZN(_06579_));
 OAI21_X1 _31732_ (.A(_06256_),
    .B1(_06147_),
    .B2(_06175_),
    .ZN(_06580_));
 NAND3_X1 _31733_ (.A1(_06256_),
    .A2(_06191_),
    .A3(_06184_),
    .ZN(_06581_));
 NAND4_X1 _31734_ (.A1(_06577_),
    .A2(_06579_),
    .A3(_06580_),
    .A4(_06581_),
    .ZN(_06582_));
 INV_X1 _31735_ (.A(_06249_),
    .ZN(_06583_));
 INV_X4 _31736_ (.A(_06313_),
    .ZN(_06584_));
 AOI21_X1 _31737_ (.A(_06583_),
    .B1(_06584_),
    .B2(_06269_),
    .ZN(_06585_));
 OR4_X2 _31738_ (.A1(_06575_),
    .A2(_06582_),
    .A3(_06585_),
    .A4(_06264_),
    .ZN(_06586_));
 AND2_X1 _31739_ (.A1(_06319_),
    .A2(_06265_),
    .ZN(_06587_));
 AND2_X4 _31740_ (.A1(_06185_),
    .A2(_06319_),
    .ZN(_06588_));
 INV_X1 _31741_ (.A(_06129_),
    .ZN(_06590_));
 NOR2_X1 _31742_ (.A1(_06590_),
    .A2(_06120_),
    .ZN(_06591_));
 AOI211_X2 _31743_ (.A(_06587_),
    .B(_06588_),
    .C1(_06319_),
    .C2(_06591_),
    .ZN(_06592_));
 OAI21_X1 _31744_ (.A(_06326_),
    .B1(_06177_),
    .B2(_06178_),
    .ZN(_06593_));
 BUF_X4 _31745_ (.A(_06263_),
    .Z(_06594_));
 NAND4_X1 _31746_ (.A1(_06298_),
    .A2(_06594_),
    .A3(_06120_),
    .A4(_06107_),
    .ZN(_06595_));
 AND2_X1 _31747_ (.A1(_06324_),
    .A2(_06164_),
    .ZN(_06596_));
 INV_X1 _31748_ (.A(_06596_),
    .ZN(_06597_));
 NAND4_X1 _31749_ (.A1(_06592_),
    .A2(_06593_),
    .A3(_06595_),
    .A4(_06597_),
    .ZN(_06598_));
 AND4_X1 _31750_ (.A1(_06192_),
    .A2(_06298_),
    .A3(_06206_),
    .A4(_06187_),
    .ZN(_06599_));
 AOI21_X1 _31751_ (.A(_06599_),
    .B1(_06185_),
    .B2(_06309_),
    .ZN(_06601_));
 OAI21_X1 _31752_ (.A(_06309_),
    .B1(_06142_),
    .B2(_06568_),
    .ZN(_06602_));
 NOR2_X1 _31753_ (.A1(_06590_),
    .A2(_06139_),
    .ZN(_06603_));
 NAND3_X1 _31754_ (.A1(_06301_),
    .A2(_06603_),
    .A3(_06211_),
    .ZN(_06604_));
 BUF_X8 _31755_ (.A(_06125_),
    .Z(_06605_));
 NAND2_X1 _31756_ (.A1(_06301_),
    .A2(_06605_),
    .ZN(_06606_));
 NAND4_X1 _31757_ (.A1(_06601_),
    .A2(_06602_),
    .A3(_06604_),
    .A4(_06606_),
    .ZN(_06607_));
 NOR4_X2 _31758_ (.A1(_06574_),
    .A2(_06586_),
    .A3(_06598_),
    .A4(_06607_),
    .ZN(_06608_));
 AND2_X1 _31759_ (.A1(_06178_),
    .A2(_06235_),
    .ZN(_06609_));
 AND2_X2 _31760_ (.A1(_06263_),
    .A2(_06139_),
    .ZN(_06610_));
 AND2_X4 _31761_ (.A1(_06605_),
    .A2(_06235_),
    .ZN(_06612_));
 AOI221_X1 _31762_ (.A(_06609_),
    .B1(_06610_),
    .B2(_06235_),
    .C1(_06205_),
    .C2(_06612_),
    .ZN(_06613_));
 NAND2_X1 _31763_ (.A1(_06603_),
    .A2(_06235_),
    .ZN(_06614_));
 INV_X1 _31764_ (.A(_06201_),
    .ZN(_06615_));
 OAI211_X2 _31765_ (.A(_06613_),
    .B(_06614_),
    .C1(_06615_),
    .C2(_06241_),
    .ZN(_06616_));
 INV_X1 _31766_ (.A(_06188_),
    .ZN(_06617_));
 NOR3_X1 _31767_ (.A1(_06617_),
    .A2(_06111_),
    .A3(_06141_),
    .ZN(_06618_));
 NAND2_X1 _31768_ (.A1(_06228_),
    .A2(_06188_),
    .ZN(_06619_));
 INV_X1 _31769_ (.A(_06199_),
    .ZN(_06620_));
 OAI21_X1 _31770_ (.A(_06619_),
    .B1(_06620_),
    .B2(_06617_),
    .ZN(_06621_));
 AOI21_X1 _31771_ (.A(_06617_),
    .B1(_06122_),
    .B2(_06240_),
    .ZN(_06623_));
 AND2_X1 _31772_ (.A1(_06188_),
    .A2(_06134_),
    .ZN(_06624_));
 OR4_X1 _31773_ (.A1(_06618_),
    .A2(_06621_),
    .A3(_06623_),
    .A4(_06624_),
    .ZN(_06625_));
 AOI21_X1 _31774_ (.A(_06224_),
    .B1(_06305_),
    .B2(_06126_),
    .ZN(_06626_));
 BUF_X4 _31775_ (.A(_06223_),
    .Z(_06627_));
 AND4_X1 _31776_ (.A1(_06211_),
    .A2(_06627_),
    .A3(_06140_),
    .A4(_06289_),
    .ZN(_06628_));
 OR4_X2 _31777_ (.A1(_06227_),
    .A2(_06626_),
    .A3(_06628_),
    .A4(_06232_),
    .ZN(_06629_));
 AND2_X1 _31778_ (.A1(_06169_),
    .A2(_06610_),
    .ZN(_06630_));
 BUF_X2 _31779_ (.A(_06284_),
    .Z(_06631_));
 AND2_X1 _31780_ (.A1(_06169_),
    .A2(_06631_),
    .ZN(_06632_));
 NOR2_X1 _31781_ (.A1(_06630_),
    .A2(_06632_),
    .ZN(_06634_));
 BUF_X4 _31782_ (.A(_06169_),
    .Z(_06635_));
 OAI21_X1 _31783_ (.A(_06635_),
    .B1(_06199_),
    .B2(_06201_),
    .ZN(_06636_));
 INV_X1 _31784_ (.A(_06168_),
    .ZN(_06637_));
 INV_X1 _31785_ (.A(_06134_),
    .ZN(_06638_));
 OAI211_X2 _31786_ (.A(_06634_),
    .B(_06636_),
    .C1(_06637_),
    .C2(_06638_),
    .ZN(_06639_));
 NOR4_X2 _31787_ (.A1(_06616_),
    .A2(_06625_),
    .A3(_06629_),
    .A4(_06639_),
    .ZN(_06640_));
 BUF_X4 _31788_ (.A(_06198_),
    .Z(_06641_));
 BUF_X4 _31789_ (.A(_06310_),
    .Z(_06642_));
 OAI21_X1 _31790_ (.A(_06641_),
    .B1(_06642_),
    .B2(_06331_),
    .ZN(_06643_));
 AND2_X1 _31791_ (.A1(_06164_),
    .A2(_06216_),
    .ZN(_06645_));
 OAI21_X1 _31792_ (.A(_06214_),
    .B1(_06320_),
    .B2(_06178_),
    .ZN(_06646_));
 NAND4_X1 _31793_ (.A1(_06263_),
    .A2(_06103_),
    .A3(_06150_),
    .A4(_06187_),
    .ZN(_06647_));
 NAND2_X1 _31794_ (.A1(_06646_),
    .A2(_06647_),
    .ZN(_06648_));
 AOI211_X2 _31795_ (.A(_06645_),
    .B(_06648_),
    .C1(_06331_),
    .C2(_06216_),
    .ZN(_06649_));
 OAI21_X1 _31796_ (.A(_06641_),
    .B1(_06568_),
    .B2(_06177_),
    .ZN(_06650_));
 NAND2_X1 _31797_ (.A1(_06641_),
    .A2(_06228_),
    .ZN(_06651_));
 AND4_X1 _31798_ (.A1(_06643_),
    .A2(_06649_),
    .A3(_06650_),
    .A4(_06651_),
    .ZN(_06652_));
 NAND3_X1 _31799_ (.A1(_06142_),
    .A2(_06211_),
    .A3(_06144_),
    .ZN(_06653_));
 NAND2_X1 _31800_ (.A1(_06631_),
    .A2(_06144_),
    .ZN(_06654_));
 AND2_X1 _31801_ (.A1(_06653_),
    .A2(_06654_),
    .ZN(_06656_));
 AND2_X2 _31802_ (.A1(_06181_),
    .A2(_06150_),
    .ZN(_06657_));
 BUF_X2 _31803_ (.A(_06144_),
    .Z(_06658_));
 AND2_X1 _31804_ (.A1(_06657_),
    .A2(_06658_),
    .ZN(_06659_));
 AND2_X1 _31805_ (.A1(_06218_),
    .A2(_06658_),
    .ZN(_06660_));
 AND2_X1 _31806_ (.A1(_06658_),
    .A2(_06642_),
    .ZN(_06661_));
 AND2_X1 _31807_ (.A1(_06144_),
    .A2(_06291_),
    .ZN(_06662_));
 NOR4_X1 _31808_ (.A1(_06659_),
    .A2(_06660_),
    .A3(_06661_),
    .A4(_06662_),
    .ZN(_06663_));
 AOI21_X1 _31809_ (.A(_16879_),
    .B1(_06192_),
    .B2(_06109_),
    .ZN(_06664_));
 NAND3_X1 _31810_ (.A1(_06664_),
    .A2(_06103_),
    .A3(_06107_),
    .ZN(_06665_));
 BUF_X2 _31811_ (.A(_06108_),
    .Z(_06667_));
 NOR3_X1 _31812_ (.A1(_06151_),
    .A2(_06117_),
    .A3(_16878_),
    .ZN(_06668_));
 OAI21_X1 _31813_ (.A(_06667_),
    .B1(_06668_),
    .B2(_06320_),
    .ZN(_06669_));
 AND4_X1 _31814_ (.A1(_06656_),
    .A2(_06663_),
    .A3(_06665_),
    .A4(_06669_),
    .ZN(_06670_));
 NAND4_X1 _31815_ (.A1(_06608_),
    .A2(_06640_),
    .A3(_06652_),
    .A4(_06670_),
    .ZN(_06671_));
 OAI21_X1 _31816_ (.A(_06117_),
    .B1(_06140_),
    .B2(_16878_),
    .ZN(_06672_));
 AND3_X1 _31817_ (.A1(_06187_),
    .A2(_06167_),
    .A3(_06117_),
    .ZN(_06673_));
 AND2_X1 _31818_ (.A1(_06672_),
    .A2(_06673_),
    .ZN(_06674_));
 NOR2_X2 _31819_ (.A1(_06671_),
    .A2(_06674_),
    .ZN(_06675_));
 XOR2_X2 _31820_ (.A(_06675_),
    .B(_06337_),
    .Z(_06676_));
 OAI21_X1 _31821_ (.A(_06089_),
    .B1(_05981_),
    .B2(_05923_),
    .ZN(_06678_));
 AND2_X4 _31822_ (.A1(_05955_),
    .A2(_16837_),
    .ZN(_06679_));
 BUF_X2 _31823_ (.A(_06679_),
    .Z(_06680_));
 OAI21_X1 _31824_ (.A(_05838_),
    .B1(_06022_),
    .B2(_06680_),
    .ZN(_06681_));
 OAI21_X1 _31825_ (.A(_06089_),
    .B1(_06027_),
    .B2(_05934_),
    .ZN(_06682_));
 AND3_X1 _31826_ (.A1(_06678_),
    .A2(_06681_),
    .A3(_06682_),
    .ZN(_06683_));
 INV_X1 _31827_ (.A(_05961_),
    .ZN(_06684_));
 AOI21_X1 _31828_ (.A(_06065_),
    .B1(_06095_),
    .B2(_06684_),
    .ZN(_06685_));
 INV_X1 _31829_ (.A(_06016_),
    .ZN(_06686_));
 AOI21_X1 _31830_ (.A(_06065_),
    .B1(_06020_),
    .B2(_06686_),
    .ZN(_06687_));
 NAND2_X1 _31831_ (.A1(_06059_),
    .A2(_05870_),
    .ZN(_06689_));
 NOR2_X1 _31832_ (.A1(_06689_),
    .A2(_05851_),
    .ZN(_06690_));
 AOI211_X4 _31833_ (.A(_06685_),
    .B(_06687_),
    .C1(_05906_),
    .C2(_06690_),
    .ZN(_06691_));
 INV_X2 _31834_ (.A(_06067_),
    .ZN(_06692_));
 AND2_X1 _31835_ (.A1(_06692_),
    .A2(_05848_),
    .ZN(_06693_));
 NAND2_X1 _31836_ (.A1(_05848_),
    .A2(_05872_),
    .ZN(_06694_));
 INV_X1 _31837_ (.A(_05848_),
    .ZN(_06695_));
 INV_X1 _31838_ (.A(_06679_),
    .ZN(_06696_));
 OAI22_X1 _31839_ (.A1(_06694_),
    .A2(_06034_),
    .B1(_06695_),
    .B2(_06696_),
    .ZN(_06697_));
 AND2_X1 _31840_ (.A1(_05840_),
    .A2(_05850_),
    .ZN(_06698_));
 AOI211_X4 _31841_ (.A(_06693_),
    .B(_06697_),
    .C1(_06698_),
    .C2(_05849_),
    .ZN(_06700_));
 AND2_X1 _31842_ (.A1(_06075_),
    .A2(_05920_),
    .ZN(_06701_));
 NAND2_X1 _31843_ (.A1(_05919_),
    .A2(_05923_),
    .ZN(_06702_));
 INV_X1 _31844_ (.A(_05919_),
    .ZN(_06703_));
 OAI21_X1 _31845_ (.A(_06702_),
    .B1(_06703_),
    .B2(_05938_),
    .ZN(_06704_));
 NOR3_X1 _31846_ (.A1(_05858_),
    .A2(_16838_),
    .A3(_05954_),
    .ZN(_06705_));
 AND2_X2 _31847_ (.A1(_06705_),
    .A2(_05887_),
    .ZN(_06706_));
 AOI211_X4 _31848_ (.A(_06701_),
    .B(_06704_),
    .C1(_05920_),
    .C2(_06706_),
    .ZN(_06707_));
 AND4_X4 _31849_ (.A1(_06683_),
    .A2(_06691_),
    .A3(_06700_),
    .A4(_06707_),
    .ZN(_06708_));
 AND3_X1 _31850_ (.A1(_05925_),
    .A2(_05999_),
    .A3(_05864_),
    .ZN(_06709_));
 NAND3_X1 _31851_ (.A1(_05925_),
    .A2(_05842_),
    .A3(_05843_),
    .ZN(_06711_));
 INV_X1 _31852_ (.A(_06025_),
    .ZN(_06712_));
 OAI21_X1 _31853_ (.A(_06711_),
    .B1(_06712_),
    .B2(_05996_),
    .ZN(_06713_));
 AOI211_X4 _31854_ (.A(_06709_),
    .B(_06713_),
    .C1(_05985_),
    .C2(_05926_),
    .ZN(_06714_));
 AND2_X4 _31855_ (.A1(_05970_),
    .A2(_06680_),
    .ZN(_06715_));
 INV_X1 _31856_ (.A(_05970_),
    .ZN(_06716_));
 INV_X1 _31857_ (.A(_06698_),
    .ZN(_06717_));
 INV_X1 _31858_ (.A(_05911_),
    .ZN(_06718_));
 AOI21_X1 _31859_ (.A(_06716_),
    .B1(_06717_),
    .B2(_06718_),
    .ZN(_06719_));
 AOI211_X4 _31860_ (.A(_06715_),
    .B(_06719_),
    .C1(_05933_),
    .C2(_05970_),
    .ZN(_06720_));
 AND3_X1 _31861_ (.A1(_05926_),
    .A2(_05864_),
    .A3(_05955_),
    .ZN(_06722_));
 AND2_X1 _31862_ (.A1(_05967_),
    .A2(_05926_),
    .ZN(_06723_));
 AND2_X1 _31863_ (.A1(_05901_),
    .A2(_05925_),
    .ZN(_06724_));
 AND2_X1 _31864_ (.A1(_05872_),
    .A2(_05925_),
    .ZN(_06725_));
 NOR4_X1 _31865_ (.A1(_06722_),
    .A2(_06723_),
    .A3(_06724_),
    .A4(_06725_),
    .ZN(_06726_));
 NOR2_X1 _31866_ (.A1(_05888_),
    .A2(_05851_),
    .ZN(_06727_));
 OAI21_X1 _31867_ (.A(_05948_),
    .B1(_05981_),
    .B2(_06727_),
    .ZN(_06728_));
 OAI21_X1 _31868_ (.A(_05903_),
    .B1(_06692_),
    .B2(_05922_),
    .ZN(_06729_));
 OAI211_X2 _31869_ (.A(_05903_),
    .B(_05955_),
    .C1(_05900_),
    .C2(_06034_),
    .ZN(_06730_));
 OAI211_X2 _31870_ (.A(_05903_),
    .B(_05870_),
    .C1(_05900_),
    .C2(_05850_),
    .ZN(_06731_));
 AND4_X1 _31871_ (.A1(_06728_),
    .A2(_06729_),
    .A3(_06730_),
    .A4(_06731_),
    .ZN(_06733_));
 AND4_X1 _31872_ (.A1(_06714_),
    .A2(_06720_),
    .A3(_06726_),
    .A4(_06733_),
    .ZN(_06734_));
 OAI211_X2 _31873_ (.A(_05882_),
    .B(_05884_),
    .C1(_05889_),
    .C2(_05864_),
    .ZN(_06735_));
 OAI21_X1 _31874_ (.A(_05882_),
    .B1(_05865_),
    .B2(_06056_),
    .ZN(_06736_));
 NAND4_X1 _31875_ (.A1(_05956_),
    .A2(_05893_),
    .A3(_06034_),
    .A4(_05880_),
    .ZN(_06737_));
 AND3_X1 _31876_ (.A1(_06735_),
    .A2(_06736_),
    .A3(_06737_),
    .ZN(_06738_));
 AND2_X1 _31877_ (.A1(_06021_),
    .A2(_05991_),
    .ZN(_06739_));
 AND2_X1 _31878_ (.A1(_05991_),
    .A2(_05966_),
    .ZN(_06740_));
 NOR2_X1 _31879_ (.A1(_06739_),
    .A2(_06740_),
    .ZN(_06741_));
 INV_X1 _31880_ (.A(_06741_),
    .ZN(_06742_));
 AND2_X1 _31881_ (.A1(_05992_),
    .A2(_05855_),
    .ZN(_06744_));
 AND2_X1 _31882_ (.A1(_06025_),
    .A2(_05991_),
    .ZN(_06745_));
 AND2_X1 _31883_ (.A1(_05991_),
    .A2(_05985_),
    .ZN(_06746_));
 NOR4_X1 _31884_ (.A1(_06742_),
    .A2(_06744_),
    .A3(_06745_),
    .A4(_06746_),
    .ZN(_06747_));
 INV_X1 _31885_ (.A(_05922_),
    .ZN(_06748_));
 AOI21_X1 _31886_ (.A(_06058_),
    .B1(_06748_),
    .B2(_05944_),
    .ZN(_06749_));
 AND3_X1 _31887_ (.A1(_06054_),
    .A2(_05887_),
    .A3(_06705_),
    .ZN(_06750_));
 AND2_X1 _31888_ (.A1(_05915_),
    .A2(_06054_),
    .ZN(_06751_));
 AND2_X1 _31889_ (.A1(_06054_),
    .A2(_06004_),
    .ZN(_06752_));
 NOR4_X1 _31890_ (.A1(_06749_),
    .A2(_06750_),
    .A3(_06751_),
    .A4(_06752_),
    .ZN(_06753_));
 NAND2_X1 _31891_ (.A1(_05894_),
    .A2(_05943_),
    .ZN(_06755_));
 OAI21_X1 _31892_ (.A(_05894_),
    .B1(_05873_),
    .B2(_05901_),
    .ZN(_06756_));
 NAND2_X1 _31893_ (.A1(_05894_),
    .A2(_05915_),
    .ZN(_06757_));
 NAND2_X1 _31894_ (.A1(_05894_),
    .A2(_06021_),
    .ZN(_06758_));
 AND4_X1 _31895_ (.A1(_06755_),
    .A2(_06756_),
    .A3(_06757_),
    .A4(_06758_),
    .ZN(_06759_));
 AND4_X1 _31896_ (.A1(_06738_),
    .A2(_06747_),
    .A3(_06753_),
    .A4(_06759_),
    .ZN(_06760_));
 INV_X1 _31897_ (.A(_06096_),
    .ZN(_06761_));
 AOI21_X1 _31898_ (.A(_05945_),
    .B1(_06761_),
    .B2(_06748_),
    .ZN(_06762_));
 AND2_X1 _31899_ (.A1(_05967_),
    .A2(_05876_),
    .ZN(_06763_));
 AND2_X1 _31900_ (.A1(_06010_),
    .A2(_05876_),
    .ZN(_06764_));
 NOR4_X1 _31901_ (.A1(_06762_),
    .A2(_05877_),
    .A3(_06763_),
    .A4(_06764_),
    .ZN(_06766_));
 NAND3_X1 _31902_ (.A1(_06010_),
    .A2(_05875_),
    .A3(_05847_),
    .ZN(_06767_));
 OAI21_X1 _31903_ (.A(_06767_),
    .B1(_06085_),
    .B2(_06005_),
    .ZN(_06768_));
 AOI21_X1 _31904_ (.A(_06085_),
    .B1(_06020_),
    .B2(_06686_),
    .ZN(_06769_));
 AND2_X1 _31905_ (.A1(_05909_),
    .A2(_06032_),
    .ZN(_06770_));
 AOI211_X4 _31906_ (.A(_06768_),
    .B(_06769_),
    .C1(_05868_),
    .C2(_06770_),
    .ZN(_06771_));
 INV_X1 _31907_ (.A(_06015_),
    .ZN(_06772_));
 INV_X1 _31908_ (.A(_05923_),
    .ZN(_06773_));
 AOI21_X1 _31909_ (.A(_06772_),
    .B1(_06000_),
    .B2(_06773_),
    .ZN(_06774_));
 AND2_X1 _31910_ (.A1(_06015_),
    .A2(_06004_),
    .ZN(_06775_));
 AND3_X1 _31911_ (.A1(_06010_),
    .A2(_06063_),
    .A3(_05875_),
    .ZN(_06777_));
 NOR4_X1 _31912_ (.A1(_06774_),
    .A2(_06018_),
    .A3(_06775_),
    .A4(_06777_),
    .ZN(_06778_));
 AOI21_X1 _31913_ (.A(_05939_),
    .B1(_05968_),
    .B2(_05979_),
    .ZN(_06779_));
 AND2_X1 _31914_ (.A1(_05844_),
    .A2(_05935_),
    .ZN(_06780_));
 AND2_X1 _31915_ (.A1(_05865_),
    .A2(_05935_),
    .ZN(_06781_));
 AND3_X1 _31916_ (.A1(_05935_),
    .A2(_05999_),
    .A3(_05851_),
    .ZN(_06782_));
 NOR4_X1 _31917_ (.A1(_06779_),
    .A2(_06780_),
    .A3(_06781_),
    .A4(_06782_),
    .ZN(_06783_));
 AND4_X1 _31918_ (.A1(_06766_),
    .A2(_06771_),
    .A3(_06778_),
    .A4(_06783_),
    .ZN(_06784_));
 NAND4_X1 _31919_ (.A1(_06708_),
    .A2(_06734_),
    .A3(_06760_),
    .A4(_06784_),
    .ZN(_06785_));
 NOR2_X2 _31920_ (.A1(_06785_),
    .A2(_06042_),
    .ZN(_06786_));
 XNOR2_X1 _31921_ (.A(_06786_),
    .B(_14401_),
    .ZN(_06788_));
 XNOR2_X1 _31922_ (.A(_06676_),
    .B(_06788_),
    .ZN(_06789_));
 XNOR2_X1 _31923_ (.A(_06558_),
    .B(_06789_),
    .ZN(_06790_));
 MUX2_X1 _31924_ (.A(_06342_),
    .B(_06790_),
    .S(_05156_),
    .Z(_00701_));
 MUX2_X1 _31925_ (.A(_17019_),
    .B(_16891_),
    .S(_06340_),
    .Z(_00739_));
 MUX2_X1 _31926_ (.A(_17020_),
    .B(_16892_),
    .S(_06340_),
    .Z(_00740_));
 MUX2_X1 _31927_ (.A(_17021_),
    .B(_16893_),
    .S(_06340_),
    .Z(_00741_));
 MUX2_X1 _31928_ (.A(_17022_),
    .B(_16894_),
    .S(_06340_),
    .Z(_00742_));
 MUX2_X1 _31929_ (.A(_17024_),
    .B(_16896_),
    .S(_06340_),
    .Z(_00744_));
 BUF_X4 _31930_ (.A(_05189_),
    .Z(_06791_));
 MUX2_X1 _31931_ (.A(_17025_),
    .B(_16897_),
    .S(_06791_),
    .Z(_00745_));
 MUX2_X1 _31932_ (.A(_17026_),
    .B(_16898_),
    .S(_06791_),
    .Z(_00746_));
 MUX2_X1 _31933_ (.A(_17027_),
    .B(_16899_),
    .S(_06791_),
    .Z(_00747_));
 MUX2_X1 _31934_ (.A(_17028_),
    .B(_16900_),
    .S(_06791_),
    .Z(_00748_));
 MUX2_X1 _31935_ (.A(_17029_),
    .B(_16901_),
    .S(_06791_),
    .Z(_00749_));
 XOR2_X1 _31936_ (.A(_17198_),
    .B(_17137_),
    .Z(_06793_));
 AOI211_X4 _31937_ (.A(_05602_),
    .B(_05743_),
    .C1(_05712_),
    .C2(_05818_),
    .ZN(_06794_));
 INV_X1 _31938_ (.A(_05611_),
    .ZN(_06795_));
 AOI21_X1 _31939_ (.A(_05743_),
    .B1(_05721_),
    .B2(_06795_),
    .ZN(_06796_));
 AND4_X1 _31940_ (.A1(_05603_),
    .A2(_05736_),
    .A3(_05672_),
    .A4(_05652_),
    .ZN(_06797_));
 OR4_X2 _31941_ (.A1(_05747_),
    .A2(_06794_),
    .A3(_06796_),
    .A4(_06797_),
    .ZN(_06799_));
 OAI211_X2 _31942_ (.A(_05758_),
    .B(_05579_),
    .C1(_05805_),
    .C2(_05585_),
    .ZN(_06800_));
 OAI21_X1 _31943_ (.A(_05758_),
    .B1(_05611_),
    .B2(_05613_),
    .ZN(_06801_));
 OAI21_X1 _31944_ (.A(_05758_),
    .B1(_05623_),
    .B2(_05646_),
    .ZN(_06802_));
 NAND3_X1 _31945_ (.A1(_06800_),
    .A2(_06801_),
    .A3(_06802_),
    .ZN(_06803_));
 OAI211_X2 _31946_ (.A(_06392_),
    .B(_05736_),
    .C1(_05661_),
    .C2(_05800_),
    .ZN(_06804_));
 NAND3_X1 _31947_ (.A1(_05729_),
    .A2(_06392_),
    .A3(_05736_),
    .ZN(_06805_));
 INV_X1 _31948_ (.A(_05754_),
    .ZN(_06806_));
 OAI211_X2 _31949_ (.A(_06804_),
    .B(_06805_),
    .C1(_06377_),
    .C2(_06806_),
    .ZN(_06807_));
 AND2_X1 _31950_ (.A1(_05771_),
    .A2(_06384_),
    .ZN(_06808_));
 INV_X1 _31951_ (.A(_06808_),
    .ZN(_06810_));
 OAI21_X1 _31952_ (.A(_05771_),
    .B1(_05794_),
    .B2(_05613_),
    .ZN(_06811_));
 OAI211_X2 _31953_ (.A(_06810_),
    .B(_06811_),
    .C1(_05658_),
    .C2(_06414_),
    .ZN(_06812_));
 NOR4_X1 _31954_ (.A1(_06799_),
    .A2(_06803_),
    .A3(_06807_),
    .A4(_06812_),
    .ZN(_06813_));
 AND2_X1 _31955_ (.A1(_05792_),
    .A2(_05713_),
    .ZN(_06814_));
 AOI211_X4 _31956_ (.A(_06433_),
    .B(_06814_),
    .C1(_06437_),
    .C2(_06403_),
    .ZN(_06815_));
 NAND3_X1 _31957_ (.A1(_05613_),
    .A2(_06392_),
    .A3(_05809_),
    .ZN(_06816_));
 OAI21_X1 _31958_ (.A(_06437_),
    .B1(_05763_),
    .B2(_05685_),
    .ZN(_06817_));
 AND3_X1 _31959_ (.A1(_06815_),
    .A2(_06816_),
    .A3(_06817_),
    .ZN(_06818_));
 NAND2_X1 _31960_ (.A1(_06390_),
    .A2(_06442_),
    .ZN(_06819_));
 AND2_X1 _31961_ (.A1(_05784_),
    .A2(_05744_),
    .ZN(_06821_));
 OAI21_X1 _31962_ (.A(_06455_),
    .B1(_06821_),
    .B2(_05611_),
    .ZN(_06822_));
 OAI21_X1 _31963_ (.A(_06442_),
    .B1(_06403_),
    .B2(_05613_),
    .ZN(_06823_));
 BUF_X2 _31964_ (.A(_05679_),
    .Z(_06824_));
 OAI21_X1 _31965_ (.A(_06455_),
    .B1(_06824_),
    .B2(_05788_),
    .ZN(_06825_));
 AND4_X1 _31966_ (.A1(_06819_),
    .A2(_06822_),
    .A3(_06823_),
    .A4(_06825_),
    .ZN(_06826_));
 AND2_X1 _31967_ (.A1(_06451_),
    .A2(_05685_),
    .ZN(_06827_));
 NAND3_X1 _31968_ (.A1(_06451_),
    .A2(_05712_),
    .A3(_06371_),
    .ZN(_06828_));
 OAI21_X1 _31969_ (.A(_06828_),
    .B1(_06795_),
    .B2(_05811_),
    .ZN(_06829_));
 OAI22_X1 _31970_ (.A1(_05582_),
    .A2(_05602_),
    .B1(_05745_),
    .B2(_05598_),
    .ZN(_06830_));
 AOI211_X4 _31971_ (.A(_06827_),
    .B(_06829_),
    .C1(_06451_),
    .C2(_06830_),
    .ZN(_06832_));
 NAND4_X1 _31972_ (.A1(_06813_),
    .A2(_06818_),
    .A3(_06826_),
    .A4(_06832_),
    .ZN(_06833_));
 OAI21_X1 _31973_ (.A(_06381_),
    .B1(_05659_),
    .B2(_05696_),
    .ZN(_06834_));
 AND2_X1 _31974_ (.A1(_05794_),
    .A2(_06381_),
    .ZN(_06835_));
 INV_X1 _31975_ (.A(_06835_),
    .ZN(_06836_));
 NAND2_X1 _31976_ (.A1(_05608_),
    .A2(_06386_),
    .ZN(_06837_));
 AND4_X1 _31977_ (.A1(_05618_),
    .A2(_06834_),
    .A3(_06836_),
    .A4(_06837_),
    .ZN(_06838_));
 OAI21_X1 _31978_ (.A(_05656_),
    .B1(_05796_),
    .B2(_05800_),
    .ZN(_06839_));
 AND4_X1 _31979_ (.A1(_05663_),
    .A2(_06838_),
    .A3(_05667_),
    .A4(_06839_),
    .ZN(_06840_));
 AND2_X1 _31980_ (.A1(_05693_),
    .A2(_05601_),
    .ZN(_06841_));
 OAI21_X1 _31981_ (.A(_05708_),
    .B1(_06841_),
    .B2(_05641_),
    .ZN(_06843_));
 AND2_X4 _31982_ (.A1(_05738_),
    .A2(_05726_),
    .ZN(_06844_));
 OAI21_X1 _31983_ (.A(_06353_),
    .B1(_06844_),
    .B2(_05788_),
    .ZN(_06845_));
 NAND4_X1 _31984_ (.A1(_05652_),
    .A2(_05817_),
    .A3(_05675_),
    .A4(_05805_),
    .ZN(_06846_));
 NAND4_X1 _31985_ (.A1(_06353_),
    .A2(_06371_),
    .A3(_05694_),
    .A4(_05592_),
    .ZN(_06847_));
 AND3_X1 _31986_ (.A1(_06845_),
    .A2(_06846_),
    .A3(_06847_),
    .ZN(_06848_));
 NAND2_X1 _31987_ (.A1(_05708_),
    .A2(_05784_),
    .ZN(_06849_));
 OAI21_X1 _31988_ (.A(_05708_),
    .B1(_05611_),
    .B2(_05613_),
    .ZN(_06850_));
 AND4_X1 _31989_ (.A1(_06843_),
    .A2(_06848_),
    .A3(_06849_),
    .A4(_06850_),
    .ZN(_06851_));
 OAI21_X1 _31990_ (.A(_05576_),
    .B1(_05794_),
    .B2(_05762_),
    .ZN(_06852_));
 OAI21_X1 _31991_ (.A(_06383_),
    .B1(_05794_),
    .B2(_05623_),
    .ZN(_06854_));
 OAI21_X1 _31992_ (.A(_06383_),
    .B1(_06384_),
    .B2(_05788_),
    .ZN(_06855_));
 OAI21_X1 _31993_ (.A(_05576_),
    .B1(_06384_),
    .B2(_06456_),
    .ZN(_06856_));
 AND4_X1 _31994_ (.A1(_06852_),
    .A2(_06854_),
    .A3(_06855_),
    .A4(_06856_),
    .ZN(_06857_));
 OAI21_X1 _31995_ (.A(_05699_),
    .B1(_05719_),
    .B2(_05623_),
    .ZN(_06858_));
 OAI21_X1 _31996_ (.A(_05699_),
    .B1(_05661_),
    .B2(_05800_),
    .ZN(_06859_));
 NAND3_X1 _31997_ (.A1(_05729_),
    .A2(_05636_),
    .A3(_05670_),
    .ZN(_06860_));
 NAND3_X1 _31998_ (.A1(_06858_),
    .A2(_06859_),
    .A3(_06860_),
    .ZN(_06861_));
 OAI21_X1 _31999_ (.A(_05671_),
    .B1(_05641_),
    .B2(_05729_),
    .ZN(_06862_));
 NAND3_X1 _32000_ (.A1(_05683_),
    .A2(_05738_),
    .A3(_05807_),
    .ZN(_06863_));
 NAND2_X1 _32001_ (.A1(_06862_),
    .A2(_06863_),
    .ZN(_06865_));
 NOR3_X1 _32002_ (.A1(_05681_),
    .A2(_05620_),
    .A3(_05723_),
    .ZN(_06866_));
 NOR4_X1 _32003_ (.A1(_06861_),
    .A2(_06865_),
    .A3(_05688_),
    .A4(_06866_),
    .ZN(_06867_));
 NAND4_X1 _32004_ (.A1(_06840_),
    .A2(_06851_),
    .A3(_06857_),
    .A4(_06867_),
    .ZN(_06868_));
 NOR2_X4 _32005_ (.A1(_06833_),
    .A2(_06868_),
    .ZN(_06869_));
 OAI21_X1 _32006_ (.A(_06548_),
    .B1(_05480_),
    .B2(_05399_),
    .ZN(_06870_));
 NAND2_X1 _32007_ (.A1(_05529_),
    .A2(_05333_),
    .ZN(_06871_));
 OAI21_X1 _32008_ (.A(_05354_),
    .B1(_05360_),
    .B2(_05345_),
    .ZN(_06872_));
 OAI21_X1 _32009_ (.A(_05354_),
    .B1(_05339_),
    .B2(_05341_),
    .ZN(_06873_));
 AND4_X1 _32010_ (.A1(_06870_),
    .A2(_06871_),
    .A3(_06872_),
    .A4(_06873_),
    .ZN(_06874_));
 OAI21_X1 _32011_ (.A(_05444_),
    .B1(_05341_),
    .B2(_05399_),
    .ZN(_06876_));
 AND2_X1 _32012_ (.A1(_05314_),
    .A2(_05439_),
    .ZN(_06877_));
 AOI211_X4 _32013_ (.A(_05466_),
    .B(_06877_),
    .C1(_05444_),
    .C2(_05517_),
    .ZN(_06878_));
 AND2_X1 _32014_ (.A1(_05419_),
    .A2(_05517_),
    .ZN(_06879_));
 AND2_X1 _32015_ (.A1(_05418_),
    .A2(_05356_),
    .ZN(_06880_));
 AND2_X1 _32016_ (.A1(_05418_),
    .A2(_05373_),
    .ZN(_06881_));
 NOR4_X1 _32017_ (.A1(_06478_),
    .A2(_06879_),
    .A3(_06880_),
    .A4(_06881_),
    .ZN(_06882_));
 OAI21_X1 _32018_ (.A(_05444_),
    .B1(_05378_),
    .B2(_05383_),
    .ZN(_06883_));
 AND4_X1 _32019_ (.A1(_06876_),
    .A2(_06878_),
    .A3(_06882_),
    .A4(_06883_),
    .ZN(_06884_));
 OAI21_X1 _32020_ (.A(_06531_),
    .B1(_05353_),
    .B2(_05356_),
    .ZN(_06885_));
 NAND3_X1 _32021_ (.A1(_05290_),
    .A2(_06531_),
    .A3(_05273_),
    .ZN(_06887_));
 OAI21_X1 _32022_ (.A(_06531_),
    .B1(_05296_),
    .B2(_06541_),
    .ZN(_06888_));
 NAND4_X1 _32023_ (.A1(_06885_),
    .A2(_06887_),
    .A3(_06888_),
    .A4(_06532_),
    .ZN(_06889_));
 AOI21_X1 _32024_ (.A(_05327_),
    .B1(_05504_),
    .B2(_05483_),
    .ZN(_06890_));
 OAI211_X2 _32025_ (.A(_05564_),
    .B(_06520_),
    .C1(_05246_),
    .C2(_05248_),
    .ZN(_06891_));
 NAND2_X1 _32026_ (.A1(_05318_),
    .A2(_05564_),
    .ZN(_06892_));
 NAND2_X1 _32027_ (.A1(_06891_),
    .A2(_06892_),
    .ZN(_06893_));
 AND2_X1 _32028_ (.A1(_05564_),
    .A2(_05356_),
    .ZN(_06894_));
 NOR4_X1 _32029_ (.A1(_06889_),
    .A2(_06890_),
    .A3(_06893_),
    .A4(_06894_),
    .ZN(_06895_));
 OAI211_X2 _32030_ (.A(_05496_),
    .B(_06514_),
    .C1(_05246_),
    .C2(_06522_),
    .ZN(_06896_));
 OAI211_X2 _32031_ (.A(_05536_),
    .B(_06896_),
    .C1(_05428_),
    .C2(_05319_),
    .ZN(_06898_));
 AOI21_X1 _32032_ (.A(_05431_),
    .B1(_06539_),
    .B2(_05504_),
    .ZN(_06899_));
 NAND4_X1 _32033_ (.A1(_06520_),
    .A2(_05232_),
    .A3(_05441_),
    .A4(_05233_),
    .ZN(_06900_));
 NAND4_X1 _32034_ (.A1(_05441_),
    .A2(_05252_),
    .A3(_05233_),
    .A4(_05446_),
    .ZN(_06901_));
 OAI211_X2 _32035_ (.A(_06900_),
    .B(_06901_),
    .C1(_05431_),
    .C2(_05363_),
    .ZN(_06902_));
 NOR4_X1 _32036_ (.A1(_06898_),
    .A2(_05436_),
    .A3(_06899_),
    .A4(_06902_),
    .ZN(_06903_));
 AND4_X1 _32037_ (.A1(_06874_),
    .A2(_06884_),
    .A3(_06895_),
    .A4(_06903_),
    .ZN(_06904_));
 AND2_X1 _32038_ (.A1(_05382_),
    .A2(_05380_),
    .ZN(_06905_));
 OAI21_X1 _32039_ (.A(_05413_),
    .B1(_06473_),
    .B2(_05263_),
    .ZN(_06906_));
 OAI21_X1 _32040_ (.A(_05375_),
    .B1(_05497_),
    .B2(_05318_),
    .ZN(_06907_));
 NAND2_X1 _32041_ (.A1(_05413_),
    .A2(_06471_),
    .ZN(_06909_));
 NAND2_X1 _32042_ (.A1(_05413_),
    .A2(_05353_),
    .ZN(_06910_));
 AND3_X1 _32043_ (.A1(_05552_),
    .A2(_06909_),
    .A3(_06910_),
    .ZN(_06911_));
 AND4_X1 _32044_ (.A1(_06905_),
    .A2(_06906_),
    .A3(_06907_),
    .A4(_06911_),
    .ZN(_06912_));
 OR2_X1 _32045_ (.A1(_05528_),
    .A2(_06486_),
    .ZN(_06913_));
 NAND4_X1 _32046_ (.A1(_06488_),
    .A2(_05246_),
    .A3(_05446_),
    .A4(_06520_),
    .ZN(_06914_));
 NAND2_X1 _32047_ (.A1(_06913_),
    .A2(_06914_),
    .ZN(_06915_));
 OAI21_X1 _32048_ (.A(_05270_),
    .B1(_05473_),
    .B2(_05378_),
    .ZN(_06916_));
 OAI211_X2 _32049_ (.A(_05270_),
    .B(_06520_),
    .C1(_05310_),
    .C2(_06522_),
    .ZN(_06917_));
 OAI211_X2 _32050_ (.A(_06916_),
    .B(_06917_),
    .C1(_05278_),
    .C2(_06494_),
    .ZN(_06918_));
 AND2_X1 _32051_ (.A1(_05399_),
    .A2(_06488_),
    .ZN(_06920_));
 AND2_X1 _32052_ (.A1(_05421_),
    .A2(_06488_),
    .ZN(_06921_));
 NOR4_X1 _32053_ (.A1(_06915_),
    .A2(_06918_),
    .A3(_06920_),
    .A4(_06921_),
    .ZN(_06922_));
 OAI21_X1 _32054_ (.A(_05392_),
    .B1(_06471_),
    .B2(_05307_),
    .ZN(_06923_));
 OAI21_X1 _32055_ (.A(_05395_),
    .B1(_06471_),
    .B2(_05378_),
    .ZN(_06924_));
 OAI21_X1 _32056_ (.A(_05392_),
    .B1(_05521_),
    .B2(_06541_),
    .ZN(_06925_));
 OAI21_X1 _32057_ (.A(_05395_),
    .B1(_05521_),
    .B2(_05345_),
    .ZN(_06926_));
 AND4_X1 _32058_ (.A1(_06923_),
    .A2(_06924_),
    .A3(_06925_),
    .A4(_06926_),
    .ZN(_06927_));
 BUF_X4 _32059_ (.A(_05216_),
    .Z(_06928_));
 AND2_X1 _32060_ (.A1(_05250_),
    .A2(_05275_),
    .ZN(_06929_));
 OAI21_X1 _32061_ (.A(_06928_),
    .B1(_06929_),
    .B2(_05345_),
    .ZN(_06931_));
 NAND4_X1 _32062_ (.A1(_05233_),
    .A2(_05240_),
    .A3(_05215_),
    .A4(_05310_),
    .ZN(_06932_));
 NAND4_X1 _32063_ (.A1(_06928_),
    .A2(_05273_),
    .A3(_05237_),
    .A4(_05230_),
    .ZN(_06933_));
 AND3_X1 _32064_ (.A1(_06931_),
    .A2(_06932_),
    .A3(_06933_),
    .ZN(_06934_));
 NAND2_X1 _32065_ (.A1(_06503_),
    .A2(_05211_),
    .ZN(_06935_));
 NAND3_X1 _32066_ (.A1(_05521_),
    .A2(_05283_),
    .A3(_05215_),
    .ZN(_06936_));
 NAND3_X1 _32067_ (.A1(_05497_),
    .A2(_05283_),
    .A3(_05215_),
    .ZN(_06937_));
 AND3_X1 _32068_ (.A1(_06935_),
    .A2(_06936_),
    .A3(_06937_),
    .ZN(_06938_));
 NAND2_X1 _32069_ (.A1(_05398_),
    .A2(_06503_),
    .ZN(_06939_));
 OAI21_X1 _32070_ (.A(_06503_),
    .B1(_05341_),
    .B2(_05399_),
    .ZN(_06940_));
 AND4_X1 _32071_ (.A1(_06934_),
    .A2(_06938_),
    .A3(_06939_),
    .A4(_06940_),
    .ZN(_06942_));
 AND4_X1 _32072_ (.A1(_06912_),
    .A2(_06922_),
    .A3(_06927_),
    .A4(_06942_),
    .ZN(_06943_));
 NAND2_X1 _32073_ (.A1(_06904_),
    .A2(_06943_),
    .ZN(_06944_));
 XOR2_X1 _32074_ (.A(_06869_),
    .B(_06944_),
    .Z(_06945_));
 BUF_X4 _32075_ (.A(_05949_),
    .Z(_06946_));
 OAI21_X1 _32076_ (.A(_06946_),
    .B1(_06705_),
    .B2(_06004_),
    .ZN(_06947_));
 AND2_X1 _32077_ (.A1(_06015_),
    .A2(_05855_),
    .ZN(_06948_));
 AND2_X1 _32078_ (.A1(_06016_),
    .A2(_05991_),
    .ZN(_06949_));
 AND2_X2 _32079_ (.A1(_05934_),
    .A2(_05882_),
    .ZN(_06950_));
 NOR3_X1 _32080_ (.A1(_06948_),
    .A2(_06949_),
    .A3(_06950_),
    .ZN(_06951_));
 AOI221_X2 _32081_ (.A(_06777_),
    .B1(_06025_),
    .B2(_05991_),
    .C1(_06027_),
    .C2(_05920_),
    .ZN(_06953_));
 OAI21_X1 _32082_ (.A(_05883_),
    .B1(_05865_),
    .B2(_05964_),
    .ZN(_06954_));
 AOI22_X1 _32083_ (.A1(_05967_),
    .A2(_05894_),
    .B1(_05992_),
    .B2(_05909_),
    .ZN(_06955_));
 AND4_X1 _32084_ (.A1(_06951_),
    .A2(_06953_),
    .A3(_06954_),
    .A4(_06955_),
    .ZN(_06956_));
 INV_X1 _32085_ (.A(_06073_),
    .ZN(_06957_));
 NAND2_X1 _32086_ (.A1(_06946_),
    .A2(_06957_),
    .ZN(_06958_));
 INV_X1 _32087_ (.A(_06035_),
    .ZN(_06959_));
 AOI21_X1 _32088_ (.A(_05939_),
    .B1(_06761_),
    .B2(_06959_),
    .ZN(_06960_));
 NOR2_X1 _32089_ (.A1(_06085_),
    .A2(_06689_),
    .ZN(_06961_));
 NOR2_X1 _32090_ (.A1(_06960_),
    .A2(_06961_),
    .ZN(_06962_));
 AND4_X2 _32091_ (.A1(_06947_),
    .A2(_06956_),
    .A3(_06958_),
    .A4(_06962_),
    .ZN(_06964_));
 NAND2_X1 _32092_ (.A1(_06680_),
    .A2(_05936_),
    .ZN(_06965_));
 NAND2_X1 _32093_ (.A1(_05915_),
    .A2(_05936_),
    .ZN(_06966_));
 AND2_X1 _32094_ (.A1(_05849_),
    .A2(_06029_),
    .ZN(_06967_));
 NOR2_X1 _32095_ (.A1(_05990_),
    .A2(_06967_),
    .ZN(_06968_));
 NAND2_X1 _32096_ (.A1(_05895_),
    .A2(_06044_),
    .ZN(_06969_));
 NAND2_X1 _32097_ (.A1(_05920_),
    .A2(_06022_),
    .ZN(_06970_));
 AND4_X1 _32098_ (.A1(_06966_),
    .A2(_06968_),
    .A3(_06969_),
    .A4(_06970_),
    .ZN(_06971_));
 OAI21_X1 _32099_ (.A(_05915_),
    .B1(_06946_),
    .B2(_05883_),
    .ZN(_06972_));
 AND4_X1 _32100_ (.A1(_06965_),
    .A2(_06971_),
    .A3(_06758_),
    .A4(_06972_),
    .ZN(_06973_));
 NAND2_X1 _32101_ (.A1(_05914_),
    .A2(_06025_),
    .ZN(_06975_));
 NAND2_X1 _32102_ (.A1(_05844_),
    .A2(_06043_),
    .ZN(_06976_));
 AND2_X1 _32103_ (.A1(_06975_),
    .A2(_06976_),
    .ZN(_06977_));
 NAND2_X1 _32104_ (.A1(_05908_),
    .A2(_06016_),
    .ZN(_06978_));
 NAND2_X1 _32105_ (.A1(_05908_),
    .A2(_06025_),
    .ZN(_06979_));
 NAND3_X1 _32106_ (.A1(_05972_),
    .A2(_06698_),
    .A3(_05871_),
    .ZN(_06980_));
 NAND4_X1 _32107_ (.A1(_06977_),
    .A2(_06978_),
    .A3(_06979_),
    .A4(_06980_),
    .ZN(_06981_));
 OAI21_X1 _32108_ (.A(_06043_),
    .B1(_06029_),
    .B2(_06046_),
    .ZN(_06982_));
 NAND2_X1 _32109_ (.A1(_06016_),
    .A2(_06043_),
    .ZN(_06983_));
 NAND2_X1 _32110_ (.A1(_06982_),
    .A2(_06983_),
    .ZN(_06984_));
 NOR2_X1 _32111_ (.A1(_05946_),
    .A2(_06000_),
    .ZN(_06986_));
 AND2_X1 _32112_ (.A1(_06054_),
    .A2(_06957_),
    .ZN(_06987_));
 NOR4_X1 _32113_ (.A1(_06981_),
    .A2(_06984_),
    .A3(_06986_),
    .A4(_06987_),
    .ZN(_06988_));
 NAND3_X1 _32114_ (.A1(_06075_),
    .A2(_05975_),
    .A3(_05992_),
    .ZN(_06989_));
 AOI21_X1 _32115_ (.A(_06007_),
    .B1(_05978_),
    .B2(_06718_),
    .ZN(_06990_));
 AND4_X1 _32116_ (.A1(_06034_),
    .A2(_05884_),
    .A3(_05880_),
    .A4(_05902_),
    .ZN(_06991_));
 NOR3_X1 _32117_ (.A1(_06990_),
    .A2(_06009_),
    .A3(_06991_),
    .ZN(_06992_));
 NOR2_X1 _32118_ (.A1(_05996_),
    .A2(_06689_),
    .ZN(_06993_));
 NOR2_X1 _32119_ (.A1(_06993_),
    .A2(_06722_),
    .ZN(_06994_));
 AND2_X1 _32120_ (.A1(_05894_),
    .A2(_05985_),
    .ZN(_06995_));
 INV_X1 _32121_ (.A(_06995_),
    .ZN(_06997_));
 NAND2_X1 _32122_ (.A1(_06706_),
    .A2(_05883_),
    .ZN(_06998_));
 OAI21_X1 _32123_ (.A(_06089_),
    .B1(_06025_),
    .B2(_05943_),
    .ZN(_06999_));
 OAI21_X1 _32124_ (.A(_06089_),
    .B1(_06016_),
    .B2(_05873_),
    .ZN(_07000_));
 AND4_X1 _32125_ (.A1(_06997_),
    .A2(_06998_),
    .A3(_06999_),
    .A4(_07000_),
    .ZN(_07001_));
 AND4_X1 _32126_ (.A1(_06989_),
    .A2(_06992_),
    .A3(_06994_),
    .A4(_07001_),
    .ZN(_07002_));
 NAND4_X1 _32127_ (.A1(_06964_),
    .A2(_06973_),
    .A3(_06988_),
    .A4(_07002_),
    .ZN(_07003_));
 NAND2_X1 _32128_ (.A1(_05921_),
    .A2(_05860_),
    .ZN(_07004_));
 AND2_X1 _32129_ (.A1(_05909_),
    .A2(_05926_),
    .ZN(_07005_));
 AND2_X1 _32130_ (.A1(_05920_),
    .A2(_05922_),
    .ZN(_07006_));
 NOR4_X1 _32131_ (.A1(_06070_),
    .A2(_07005_),
    .A3(_06751_),
    .A4(_07006_),
    .ZN(_07008_));
 NAND2_X1 _32132_ (.A1(_05890_),
    .A2(_05883_),
    .ZN(_07009_));
 AND2_X1 _32133_ (.A1(_05906_),
    .A2(_05860_),
    .ZN(_07010_));
 AND3_X1 _32134_ (.A1(_05971_),
    .A2(_05839_),
    .A3(_05858_),
    .ZN(_07011_));
 AND2_X1 _32135_ (.A1(_05914_),
    .A2(_05961_),
    .ZN(_07012_));
 NOR4_X1 _32136_ (.A1(_07010_),
    .A2(_07011_),
    .A3(_05856_),
    .A4(_07012_),
    .ZN(_07013_));
 AND4_X1 _32137_ (.A1(_07004_),
    .A2(_07008_),
    .A3(_07009_),
    .A4(_07013_),
    .ZN(_07014_));
 NAND2_X1 _32138_ (.A1(_06043_),
    .A2(_05985_),
    .ZN(_07015_));
 AND2_X1 _32139_ (.A1(_05970_),
    .A2(_05901_),
    .ZN(_07016_));
 AOI221_X4 _32140_ (.A(_07016_),
    .B1(_06022_),
    .B2(_05971_),
    .C1(_05926_),
    .C2(_05898_),
    .ZN(_07017_));
 AND3_X1 _32141_ (.A1(_06032_),
    .A2(_05887_),
    .A3(_06705_),
    .ZN(_07019_));
 AOI211_X4 _32142_ (.A(_06770_),
    .B(_07019_),
    .C1(_05909_),
    .C2(_05949_),
    .ZN(_07020_));
 NAND3_X1 _32143_ (.A1(_06035_),
    .A2(_06063_),
    .A3(_05836_),
    .ZN(_07021_));
 AND4_X1 _32144_ (.A1(_07015_),
    .A2(_07017_),
    .A3(_07020_),
    .A4(_07021_),
    .ZN(_07022_));
 AND2_X1 _32145_ (.A1(_06022_),
    .A2(_06055_),
    .ZN(_07023_));
 AND2_X1 _32146_ (.A1(_05909_),
    .A2(_06055_),
    .ZN(_07024_));
 AND2_X1 _32147_ (.A1(_06680_),
    .A2(_06055_),
    .ZN(_07025_));
 AND2_X1 _32148_ (.A1(_06054_),
    .A2(_05901_),
    .ZN(_07026_));
 NOR4_X1 _32149_ (.A1(_07023_),
    .A2(_07024_),
    .A3(_07025_),
    .A4(_07026_),
    .ZN(_07027_));
 AND2_X1 _32150_ (.A1(_06024_),
    .A2(_05873_),
    .ZN(_07028_));
 AND3_X1 _32151_ (.A1(_06015_),
    .A2(_05871_),
    .A3(_05954_),
    .ZN(_07030_));
 AOI211_X4 _32152_ (.A(_07028_),
    .B(_07030_),
    .C1(_06024_),
    .C2(_06706_),
    .ZN(_07031_));
 NAND4_X1 _32153_ (.A1(_07014_),
    .A2(_07022_),
    .A3(_07027_),
    .A4(_07031_),
    .ZN(_07032_));
 NOR2_X4 _32154_ (.A1(_07003_),
    .A2(_07032_),
    .ZN(_07033_));
 XNOR2_X1 _32155_ (.A(_07033_),
    .B(_00991_),
    .ZN(_07034_));
 XNOR2_X1 _32156_ (.A(_06945_),
    .B(_07034_),
    .ZN(_07035_));
 AND2_X1 _32157_ (.A1(_06188_),
    .A2(_06175_),
    .ZN(_07036_));
 AND3_X1 _32158_ (.A1(_06188_),
    .A2(_06210_),
    .A3(_06289_),
    .ZN(_07037_));
 AND2_X1 _32159_ (.A1(_06188_),
    .A2(_06124_),
    .ZN(_07038_));
 NOR4_X1 _32160_ (.A1(_07036_),
    .A2(_07037_),
    .A3(_06624_),
    .A4(_07038_),
    .ZN(_07039_));
 AND2_X4 _32161_ (.A1(_06169_),
    .A2(_06131_),
    .ZN(_07041_));
 NAND2_X1 _32162_ (.A1(_06168_),
    .A2(_06320_),
    .ZN(_07042_));
 OAI21_X1 _32163_ (.A(_07042_),
    .B1(_06637_),
    .B2(_06240_),
    .ZN(_07043_));
 AND2_X1 _32164_ (.A1(_06181_),
    .A2(_06119_),
    .ZN(_07044_));
 AOI211_X4 _32165_ (.A(_07041_),
    .B(_07043_),
    .C1(_07044_),
    .C2(_06169_),
    .ZN(_07045_));
 NAND2_X1 _32166_ (.A1(_06210_),
    .A2(_06181_),
    .ZN(_07046_));
 NOR2_X1 _32167_ (.A1(_06224_),
    .A2(_07046_),
    .ZN(_07047_));
 INV_X1 _32168_ (.A(_06173_),
    .ZN(_07048_));
 AOI21_X1 _32169_ (.A(_06224_),
    .B1(_07048_),
    .B2(_06311_),
    .ZN(_07049_));
 AOI211_X4 _32170_ (.A(_07047_),
    .B(_07049_),
    .C1(_06627_),
    .C2(_06291_),
    .ZN(_07050_));
 INV_X1 _32171_ (.A(_06243_),
    .ZN(_07052_));
 OAI211_X2 _32172_ (.A(_06235_),
    .B(_06263_),
    .C1(_06150_),
    .C2(_06194_),
    .ZN(_07053_));
 OAI211_X2 _32173_ (.A(_06235_),
    .B(_06124_),
    .C1(_06119_),
    .C2(_06194_),
    .ZN(_07054_));
 AND4_X1 _32174_ (.A1(_07052_),
    .A2(_07053_),
    .A3(_07054_),
    .A4(_06614_),
    .ZN(_07055_));
 AND4_X1 _32175_ (.A1(_07039_),
    .A2(_07045_),
    .A3(_07050_),
    .A4(_07055_),
    .ZN(_07056_));
 INV_X1 _32176_ (.A(_06319_),
    .ZN(_07057_));
 OR2_X1 _32177_ (.A1(_06141_),
    .A2(_06111_),
    .ZN(_07058_));
 INV_X1 _32178_ (.A(_06568_),
    .ZN(_07059_));
 AOI21_X1 _32179_ (.A(_07057_),
    .B1(_07058_),
    .B2(_07059_),
    .ZN(_07060_));
 INV_X1 _32180_ (.A(_06228_),
    .ZN(_07061_));
 AOI211_X2 _32181_ (.A(_06150_),
    .B(_07057_),
    .C1(_06590_),
    .C2(_07061_),
    .ZN(_07063_));
 AND2_X1 _32182_ (.A1(_06324_),
    .A2(_06668_),
    .ZN(_07064_));
 NAND2_X1 _32183_ (.A1(_06324_),
    .A2(_06217_),
    .ZN(_07065_));
 NAND3_X1 _32184_ (.A1(_06199_),
    .A2(_06297_),
    .A3(_06107_),
    .ZN(_07066_));
 INV_X1 _32185_ (.A(_06324_),
    .ZN(_07067_));
 OAI211_X2 _32186_ (.A(_07065_),
    .B(_07066_),
    .C1(_07067_),
    .C2(_06638_),
    .ZN(_07068_));
 OR4_X1 _32187_ (.A1(_07060_),
    .A2(_07063_),
    .A3(_07064_),
    .A4(_07068_),
    .ZN(_07069_));
 NAND4_X1 _32188_ (.A1(_06209_),
    .A2(_06298_),
    .A3(_06211_),
    .A4(_06187_),
    .ZN(_07070_));
 INV_X1 _32189_ (.A(_06308_),
    .ZN(_07071_));
 OAI21_X1 _32190_ (.A(_07070_),
    .B1(_07071_),
    .B2(_06302_),
    .ZN(_07072_));
 NOR2_X1 _32191_ (.A1(_06185_),
    .A2(_06173_),
    .ZN(_07074_));
 NOR2_X1 _32192_ (.A1(_07074_),
    .A2(_07071_),
    .ZN(_07075_));
 AND2_X1 _32193_ (.A1(_06301_),
    .A2(_06124_),
    .ZN(_07076_));
 AND2_X1 _32194_ (.A1(_06300_),
    .A2(_06156_),
    .ZN(_07077_));
 AND2_X1 _32195_ (.A1(_06300_),
    .A2(_06146_),
    .ZN(_07078_));
 AND3_X1 _32196_ (.A1(_06173_),
    .A2(_06203_),
    .A3(_06297_),
    .ZN(_07079_));
 OR4_X4 _32197_ (.A1(_07076_),
    .A2(_07077_),
    .A3(_07078_),
    .A4(_07079_),
    .ZN(_07080_));
 NOR4_X2 _32198_ (.A1(_07069_),
    .A2(_07072_),
    .A3(_07075_),
    .A4(_07080_),
    .ZN(_07081_));
 INV_X1 _32199_ (.A(_06214_),
    .ZN(_07082_));
 NOR2_X1 _32200_ (.A1(_07082_),
    .A2(_07046_),
    .ZN(_07083_));
 INV_X1 _32201_ (.A(_07083_),
    .ZN(_07085_));
 AND2_X1 _32202_ (.A1(_06214_),
    .A2(_06263_),
    .ZN(_07086_));
 INV_X1 _32203_ (.A(_07086_),
    .ZN(_07087_));
 OAI21_X1 _32204_ (.A(_06216_),
    .B1(_06564_),
    .B2(_06159_),
    .ZN(_07088_));
 AND3_X1 _32205_ (.A1(_07085_),
    .A2(_07087_),
    .A3(_07088_),
    .ZN(_07089_));
 AND2_X1 _32206_ (.A1(_06198_),
    .A2(_06147_),
    .ZN(_07090_));
 INV_X1 _32207_ (.A(_07090_),
    .ZN(_07091_));
 NAND2_X1 _32208_ (.A1(_06198_),
    .A2(_06153_),
    .ZN(_07092_));
 OAI21_X1 _32209_ (.A(_06198_),
    .B1(_06113_),
    .B2(_06291_),
    .ZN(_07093_));
 OAI21_X1 _32210_ (.A(_06198_),
    .B1(_06177_),
    .B2(_06265_),
    .ZN(_07094_));
 AND4_X1 _32211_ (.A1(_07091_),
    .A2(_07092_),
    .A3(_07093_),
    .A4(_07094_),
    .ZN(_07096_));
 INV_X1 _32212_ (.A(_06320_),
    .ZN(_07097_));
 AOI21_X1 _32213_ (.A(_06115_),
    .B1(_06240_),
    .B2(_07097_),
    .ZN(_07098_));
 AND2_X1 _32214_ (.A1(_06108_),
    .A2(_06217_),
    .ZN(_07099_));
 AND4_X1 _32215_ (.A1(_06119_),
    .A2(_06181_),
    .A3(_06103_),
    .A4(_06107_),
    .ZN(_07100_));
 NOR4_X1 _32216_ (.A1(_07098_),
    .A2(_06135_),
    .A3(_07099_),
    .A4(_07100_),
    .ZN(_07101_));
 AND4_X1 _32217_ (.A1(_06210_),
    .A2(_06209_),
    .A3(_06103_),
    .A4(_06143_),
    .ZN(_07102_));
 AND4_X1 _32218_ (.A1(_06139_),
    .A2(_06181_),
    .A3(_06103_),
    .A4(_06143_),
    .ZN(_07103_));
 NOR4_X1 _32219_ (.A1(_06145_),
    .A2(_07102_),
    .A3(_06161_),
    .A4(_07103_),
    .ZN(_07104_));
 AND4_X1 _32220_ (.A1(_07089_),
    .A2(_07096_),
    .A3(_07101_),
    .A4(_07104_),
    .ZN(_07105_));
 NAND3_X1 _32221_ (.A1(_06278_),
    .A2(_06140_),
    .A3(_06664_),
    .ZN(_07107_));
 OAI21_X1 _32222_ (.A(_06256_),
    .B1(_06631_),
    .B2(_06125_),
    .ZN(_07108_));
 AND2_X1 _32223_ (.A1(_06152_),
    .A2(_06247_),
    .ZN(_07109_));
 AND2_X1 _32224_ (.A1(_06146_),
    .A2(_06247_),
    .ZN(_07110_));
 NOR4_X2 _32225_ (.A1(_06266_),
    .A2(_07109_),
    .A3(_07110_),
    .A4(_06267_),
    .ZN(_07111_));
 NAND2_X1 _32226_ (.A1(_06200_),
    .A2(_06249_),
    .ZN(_07112_));
 OAI211_X2 _32227_ (.A(_06256_),
    .B(_06181_),
    .C1(_06119_),
    .C2(_06194_),
    .ZN(_07113_));
 AND4_X1 _32228_ (.A1(_07108_),
    .A2(_07111_),
    .A3(_07112_),
    .A4(_07113_),
    .ZN(_07114_));
 INV_X1 _32229_ (.A(_06273_),
    .ZN(_07115_));
 INV_X1 _32230_ (.A(_06657_),
    .ZN(_07116_));
 AOI21_X1 _32231_ (.A(_07115_),
    .B1(_06584_),
    .B2(_07116_),
    .ZN(_07118_));
 AND2_X1 _32232_ (.A1(_06265_),
    .A2(_06273_),
    .ZN(_07119_));
 AND2_X1 _32233_ (.A1(_06284_),
    .A2(_06273_),
    .ZN(_07120_));
 NOR4_X1 _32234_ (.A1(_07118_),
    .A2(_06569_),
    .A3(_07119_),
    .A4(_07120_),
    .ZN(_07121_));
 OAI21_X1 _32235_ (.A(_06278_),
    .B1(_06306_),
    .B2(_06153_),
    .ZN(_07122_));
 AND4_X1 _32236_ (.A1(_07107_),
    .A2(_07114_),
    .A3(_07121_),
    .A4(_07122_),
    .ZN(_07123_));
 AND4_X2 _32237_ (.A1(_07056_),
    .A2(_07081_),
    .A3(_07105_),
    .A4(_07123_),
    .ZN(_07124_));
 INV_X1 _32238_ (.A(_06674_),
    .ZN(_07125_));
 NAND2_X2 _32239_ (.A1(_07124_),
    .A2(_07125_),
    .ZN(_07126_));
 XNOR2_X1 _32240_ (.A(_07126_),
    .B(_06555_),
    .ZN(_07127_));
 XNOR2_X1 _32241_ (.A(_07035_),
    .B(_07127_),
    .ZN(_07129_));
 MUX2_X1 _32242_ (.A(_06793_),
    .B(_07129_),
    .S(_05156_),
    .Z(_00702_));
 MUX2_X1 _32243_ (.A(_17030_),
    .B(_16902_),
    .S(_06791_),
    .Z(_00750_));
 MUX2_X1 _32244_ (.A(_17031_),
    .B(_16903_),
    .S(_06791_),
    .Z(_00751_));
 MUX2_X1 _32245_ (.A(_17032_),
    .B(_16904_),
    .S(_06791_),
    .Z(_00752_));
 MUX2_X1 _32246_ (.A(_17033_),
    .B(_16905_),
    .S(_06791_),
    .Z(_00753_));
 MUX2_X1 _32247_ (.A(_17035_),
    .B(_16907_),
    .S(_06791_),
    .Z(_00755_));
 MUX2_X1 _32248_ (.A(_17036_),
    .B(_16908_),
    .S(_03836_),
    .Z(_00756_));
 MUX2_X1 _32249_ (.A(_17037_),
    .B(_16909_),
    .S(_03836_),
    .Z(_00757_));
 MUX2_X1 _32250_ (.A(_17038_),
    .B(_16910_),
    .S(_03836_),
    .Z(_00758_));
 MUX2_X1 _32251_ (.A(_17039_),
    .B(_16911_),
    .S(_03836_),
    .Z(_00759_));
 MUX2_X1 _32252_ (.A(_17040_),
    .B(_16912_),
    .S(_03836_),
    .Z(_00760_));
 XOR2_X1 _32253_ (.A(_17201_),
    .B(_17138_),
    .Z(_07131_));
 NOR2_X1 _32254_ (.A1(_05945_),
    .A2(_06020_),
    .ZN(_07132_));
 NOR2_X1 _32255_ (.A1(_06060_),
    .A2(_05889_),
    .ZN(_07133_));
 AOI221_X4 _32256_ (.A(_07132_),
    .B1(_05912_),
    .B2(_06043_),
    .C1(_06002_),
    .C2(_07133_),
    .ZN(_07134_));
 AND2_X1 _32257_ (.A1(_05908_),
    .A2(_06022_),
    .ZN(_07135_));
 INV_X1 _32258_ (.A(_07135_),
    .ZN(_07136_));
 AND2_X1 _32259_ (.A1(_05906_),
    .A2(_05933_),
    .ZN(_07137_));
 INV_X1 _32260_ (.A(_07137_),
    .ZN(_07138_));
 NAND4_X1 _32261_ (.A1(_06063_),
    .A2(_05836_),
    .A3(_05900_),
    .A4(_05884_),
    .ZN(_07140_));
 AND3_X1 _32262_ (.A1(_07138_),
    .A2(_06064_),
    .A3(_07140_),
    .ZN(_07141_));
 AND2_X1 _32263_ (.A1(_06706_),
    .A2(_05894_),
    .ZN(_07142_));
 INV_X1 _32264_ (.A(_07142_),
    .ZN(_07143_));
 NAND3_X1 _32265_ (.A1(_05922_),
    .A2(_06063_),
    .A3(_05893_),
    .ZN(_07144_));
 AND4_X1 _32266_ (.A1(_07136_),
    .A2(_07141_),
    .A3(_07143_),
    .A4(_07144_),
    .ZN(_07145_));
 AND2_X1 _32267_ (.A1(_05908_),
    .A2(_05922_),
    .ZN(_07146_));
 AOI221_X4 _32268_ (.A(_07146_),
    .B1(_06680_),
    .B2(_05908_),
    .C1(_05972_),
    .C2(_05915_),
    .ZN(_07147_));
 OAI21_X1 _32269_ (.A(_06089_),
    .B1(_05997_),
    .B2(_06727_),
    .ZN(_07148_));
 NOR3_X1 _32270_ (.A1(_06772_),
    .A2(_05889_),
    .A3(_06060_),
    .ZN(_07149_));
 INV_X1 _32271_ (.A(_07149_),
    .ZN(_07151_));
 AND2_X1 _32272_ (.A1(_05992_),
    .A2(_05961_),
    .ZN(_07152_));
 NOR2_X1 _32273_ (.A1(_05993_),
    .A2(_07152_),
    .ZN(_07153_));
 NAND2_X1 _32274_ (.A1(_05949_),
    .A2(_05922_),
    .ZN(_07154_));
 AND4_X1 _32275_ (.A1(_07148_),
    .A2(_07151_),
    .A3(_07153_),
    .A4(_07154_),
    .ZN(_07155_));
 AND4_X1 _32276_ (.A1(_07134_),
    .A2(_07145_),
    .A3(_07147_),
    .A4(_07155_),
    .ZN(_07156_));
 AOI21_X1 _32277_ (.A(_06693_),
    .B1(_05981_),
    .B2(_06089_),
    .ZN(_07157_));
 AND2_X1 _32278_ (.A1(_05844_),
    .A2(_06043_),
    .ZN(_07158_));
 AND3_X1 _32279_ (.A1(_05901_),
    .A2(_05925_),
    .A3(_05868_),
    .ZN(_07159_));
 NOR4_X1 _32280_ (.A1(_06948_),
    .A2(_06949_),
    .A3(_07158_),
    .A4(_07159_),
    .ZN(_07160_));
 INV_X1 _32281_ (.A(_05992_),
    .ZN(_07162_));
 OAI22_X1 _32282_ (.A1(_07162_),
    .A2(_06005_),
    .B1(_05968_),
    .B2(_05946_),
    .ZN(_07163_));
 AND2_X1 _32283_ (.A1(_05844_),
    .A2(_06055_),
    .ZN(_07164_));
 AND3_X1 _32284_ (.A1(_06033_),
    .A2(_05868_),
    .A3(_06044_),
    .ZN(_07165_));
 NOR4_X1 _32285_ (.A1(_07163_),
    .A2(_07164_),
    .A3(_07165_),
    .A4(_06780_),
    .ZN(_07166_));
 AOI21_X1 _32286_ (.A(_05939_),
    .B1(_06684_),
    .B2(_06095_),
    .ZN(_07167_));
 AND2_X1 _32287_ (.A1(_05967_),
    .A2(_06033_),
    .ZN(_07168_));
 AND2_X1 _32288_ (.A1(_05997_),
    .A2(_05936_),
    .ZN(_07169_));
 AND3_X1 _32289_ (.A1(_06010_),
    .A2(_06063_),
    .A3(_05902_),
    .ZN(_07170_));
 NOR4_X1 _32290_ (.A1(_07167_),
    .A2(_07168_),
    .A3(_07169_),
    .A4(_07170_),
    .ZN(_07171_));
 AND4_X1 _32291_ (.A1(_07157_),
    .A2(_07160_),
    .A3(_07166_),
    .A4(_07171_),
    .ZN(_07173_));
 NAND4_X1 _32292_ (.A1(_05893_),
    .A2(_06034_),
    .A3(_05880_),
    .A4(_05854_),
    .ZN(_07174_));
 AND4_X1 _32293_ (.A1(_05871_),
    .A2(_05893_),
    .A3(_05884_),
    .A4(_05880_),
    .ZN(_07175_));
 AND2_X1 _32294_ (.A1(_06027_),
    .A2(_05882_),
    .ZN(_07176_));
 AOI211_X4 _32295_ (.A(_07175_),
    .B(_07176_),
    .C1(_05969_),
    .C2(_05883_),
    .ZN(_07177_));
 AOI21_X1 _32296_ (.A(_05996_),
    .B1(_05978_),
    .B2(_06773_),
    .ZN(_07178_));
 AOI211_X4 _32297_ (.A(_06987_),
    .B(_07178_),
    .C1(_05884_),
    .C2(_05895_),
    .ZN(_07179_));
 OAI211_X2 _32298_ (.A(_05883_),
    .B(_05999_),
    .C1(_05871_),
    .C2(_05868_),
    .ZN(_07180_));
 AND4_X1 _32299_ (.A1(_07174_),
    .A2(_07177_),
    .A3(_07179_),
    .A4(_07180_),
    .ZN(_07181_));
 OAI21_X1 _32300_ (.A(_06033_),
    .B1(_05855_),
    .B2(_05873_),
    .ZN(_07182_));
 NOR2_X1 _32301_ (.A1(_06019_),
    .A2(_07028_),
    .ZN(_07184_));
 AND2_X1 _32302_ (.A1(_05956_),
    .A2(_05868_),
    .ZN(_07185_));
 OAI21_X1 _32303_ (.A(_05921_),
    .B1(_05977_),
    .B2(_07185_),
    .ZN(_07186_));
 AND2_X1 _32304_ (.A1(_05971_),
    .A2(_06727_),
    .ZN(_07187_));
 INV_X1 _32305_ (.A(_07187_),
    .ZN(_07188_));
 AND4_X1 _32306_ (.A1(_07182_),
    .A2(_07184_),
    .A3(_07186_),
    .A4(_07188_),
    .ZN(_07189_));
 NAND4_X1 _32307_ (.A1(_07156_),
    .A2(_07173_),
    .A3(_07181_),
    .A4(_07189_),
    .ZN(_07190_));
 NAND2_X1 _32308_ (.A1(_05928_),
    .A2(_06055_),
    .ZN(_07191_));
 AOI221_X4 _32309_ (.A(_07010_),
    .B1(_05949_),
    .B2(_05855_),
    .C1(_05972_),
    .C2(_05969_),
    .ZN(_07192_));
 AND2_X1 _32310_ (.A1(_05870_),
    .A2(_05850_),
    .ZN(_07193_));
 AOI221_X4 _32311_ (.A(_06723_),
    .B1(_05860_),
    .B2(_05920_),
    .C1(_06089_),
    .C2(_07193_),
    .ZN(_07195_));
 AOI221_X4 _32312_ (.A(_06088_),
    .B1(_05985_),
    .B2(_05935_),
    .C1(_06044_),
    .C2(_06043_),
    .ZN(_07196_));
 AND4_X1 _32313_ (.A1(_07191_),
    .A2(_07192_),
    .A3(_07195_),
    .A4(_07196_),
    .ZN(_07197_));
 AOI22_X1 _32314_ (.A1(_05914_),
    .A2(_05873_),
    .B1(_05895_),
    .B2(_05985_),
    .ZN(_07198_));
 OR2_X1 _32315_ (.A1(_06746_),
    .A2(_05877_),
    .ZN(_07199_));
 AND2_X1 _32316_ (.A1(_05914_),
    .A2(_06046_),
    .ZN(_07200_));
 OAI21_X1 _32317_ (.A(_06965_),
    .B1(_06085_),
    .B2(_06020_),
    .ZN(_07201_));
 NOR4_X1 _32318_ (.A1(_07199_),
    .A2(_07200_),
    .A3(_07025_),
    .A4(_07201_),
    .ZN(_07202_));
 AND2_X1 _32319_ (.A1(_05933_),
    .A2(_05925_),
    .ZN(_07203_));
 INV_X1 _32320_ (.A(_07203_),
    .ZN(_07204_));
 INV_X1 _32321_ (.A(_06029_),
    .ZN(_07206_));
 OAI211_X2 _32322_ (.A(_07204_),
    .B(_05937_),
    .C1(_07206_),
    .C2(_06703_),
    .ZN(_07207_));
 NAND2_X1 _32323_ (.A1(_05949_),
    .A2(_06029_),
    .ZN(_07208_));
 NAND3_X1 _32324_ (.A1(_06044_),
    .A2(_06002_),
    .A3(_05868_),
    .ZN(_07209_));
 OAI211_X2 _32325_ (.A(_07208_),
    .B(_07209_),
    .C1(_05944_),
    .C2(_06085_),
    .ZN(_07210_));
 OAI21_X1 _32326_ (.A(_06975_),
    .B1(_06695_),
    .B2(_07206_),
    .ZN(_07211_));
 NAND2_X1 _32327_ (.A1(_05865_),
    .A2(_06033_),
    .ZN(_07212_));
 OAI21_X1 _32328_ (.A(_07212_),
    .B1(_06093_),
    .B2(_05946_),
    .ZN(_07213_));
 NOR4_X1 _32329_ (.A1(_07207_),
    .A2(_07210_),
    .A3(_07211_),
    .A4(_07213_),
    .ZN(_07214_));
 NAND4_X1 _32330_ (.A1(_07197_),
    .A2(_07198_),
    .A3(_07202_),
    .A4(_07214_),
    .ZN(_07215_));
 NOR2_X4 _32331_ (.A1(_07190_),
    .A2(_07215_),
    .ZN(_07217_));
 XNOR2_X1 _32332_ (.A(_07217_),
    .B(_14561_),
    .ZN(_07218_));
 XOR2_X1 _32333_ (.A(_05570_),
    .B(_06944_),
    .Z(_07219_));
 XOR2_X1 _32334_ (.A(_07218_),
    .B(_07219_),
    .Z(_07220_));
 INV_X1 _32335_ (.A(_06252_),
    .ZN(_07221_));
 BUF_X4 _32336_ (.A(_06249_),
    .Z(_07222_));
 AND3_X1 _32337_ (.A1(_07222_),
    .A2(_06211_),
    .A3(_06209_),
    .ZN(_07223_));
 NOR3_X1 _32338_ (.A1(_07223_),
    .A2(_06266_),
    .A3(_06575_),
    .ZN(_07224_));
 OAI21_X1 _32339_ (.A(_06257_),
    .B1(_06220_),
    .B2(_06175_),
    .ZN(_07225_));
 OAI21_X1 _32340_ (.A(_06257_),
    .B1(_06313_),
    .B2(_06156_),
    .ZN(_07226_));
 AND4_X1 _32341_ (.A1(_07221_),
    .A2(_07224_),
    .A3(_07225_),
    .A4(_07226_),
    .ZN(_07228_));
 NAND2_X1 _32342_ (.A1(_06330_),
    .A2(_06591_),
    .ZN(_07229_));
 AND4_X1 _32343_ (.A1(_06298_),
    .A2(_06263_),
    .A3(_06184_),
    .A4(_06143_),
    .ZN(_07230_));
 AOI21_X1 _32344_ (.A(_07057_),
    .B1(_06305_),
    .B2(_07097_),
    .ZN(_07231_));
 AOI211_X4 _32345_ (.A(_07230_),
    .B(_07231_),
    .C1(_06330_),
    .C2(_06147_),
    .ZN(_07232_));
 AND2_X2 _32346_ (.A1(_06324_),
    .A2(_06153_),
    .ZN(_07233_));
 OAI21_X1 _32347_ (.A(_07066_),
    .B1(_07067_),
    .B2(_07061_),
    .ZN(_07234_));
 AOI211_X4 _32348_ (.A(_07233_),
    .B(_07234_),
    .C1(_06326_),
    .C2(_06564_),
    .ZN(_07235_));
 OAI21_X1 _32349_ (.A(_06330_),
    .B1(_06201_),
    .B2(_06156_),
    .ZN(_07236_));
 AND4_X1 _32350_ (.A1(_07229_),
    .A2(_07232_),
    .A3(_07235_),
    .A4(_07236_),
    .ZN(_07237_));
 OAI21_X1 _32351_ (.A(_06572_),
    .B1(_06121_),
    .B2(_06153_),
    .ZN(_07239_));
 OAI21_X1 _32352_ (.A(_06572_),
    .B1(_06218_),
    .B2(_06134_),
    .ZN(_07240_));
 OAI21_X1 _32353_ (.A(_06572_),
    .B1(_06304_),
    .B2(_06605_),
    .ZN(_07241_));
 NAND3_X1 _32354_ (.A1(_06228_),
    .A2(_06203_),
    .A3(_06246_),
    .ZN(_07242_));
 NAND4_X1 _32355_ (.A1(_07239_),
    .A2(_07240_),
    .A3(_07241_),
    .A4(_07242_),
    .ZN(_07243_));
 OAI21_X1 _32356_ (.A(_06273_),
    .B1(_06568_),
    .B2(_06230_),
    .ZN(_07244_));
 NAND2_X1 _32357_ (.A1(_06153_),
    .A2(_06273_),
    .ZN(_07245_));
 NAND2_X1 _32358_ (.A1(_07244_),
    .A2(_07245_),
    .ZN(_07246_));
 AND2_X1 _32359_ (.A1(_06274_),
    .A2(_06134_),
    .ZN(_07247_));
 NOR4_X1 _32360_ (.A1(_07243_),
    .A2(_07246_),
    .A3(_06290_),
    .A4(_07247_),
    .ZN(_07248_));
 AND2_X1 _32361_ (.A1(_06301_),
    .A2(_06134_),
    .ZN(_07250_));
 INV_X1 _32362_ (.A(_07250_),
    .ZN(_07251_));
 INV_X1 _32363_ (.A(_07078_),
    .ZN(_07252_));
 NAND2_X1 _32364_ (.A1(_06301_),
    .A2(_06178_),
    .ZN(_07253_));
 NAND3_X1 _32365_ (.A1(_06631_),
    .A2(_06203_),
    .A3(_06298_),
    .ZN(_07254_));
 NAND4_X1 _32366_ (.A1(_07251_),
    .A2(_07252_),
    .A3(_07253_),
    .A4(_07254_),
    .ZN(_07255_));
 AOI211_X4 _32367_ (.A(_06117_),
    .B(_07071_),
    .C1(_06294_),
    .C2(_16878_),
    .ZN(_07256_));
 AND2_X1 _32368_ (.A1(_06309_),
    .A2(_06289_),
    .ZN(_07257_));
 INV_X1 _32369_ (.A(_06184_),
    .ZN(_07258_));
 NAND2_X1 _32370_ (.A1(_07258_),
    .A2(_06206_),
    .ZN(_07259_));
 NOR2_X1 _32371_ (.A1(_07071_),
    .A2(_07259_),
    .ZN(_07261_));
 NOR4_X1 _32372_ (.A1(_07255_),
    .A2(_07256_),
    .A3(_07257_),
    .A4(_07261_),
    .ZN(_07262_));
 AND4_X1 _32373_ (.A1(_07228_),
    .A2(_07237_),
    .A3(_07248_),
    .A4(_07262_),
    .ZN(_07263_));
 NAND2_X1 _32374_ (.A1(_06635_),
    .A2(_06201_),
    .ZN(_07264_));
 NAND2_X1 _32375_ (.A1(_06635_),
    .A2(_06642_),
    .ZN(_07265_));
 NAND2_X1 _32376_ (.A1(_07264_),
    .A2(_07265_),
    .ZN(_07266_));
 INV_X1 _32377_ (.A(_06147_),
    .ZN(_07267_));
 AOI21_X1 _32378_ (.A(_06637_),
    .B1(_06561_),
    .B2(_07267_),
    .ZN(_07268_));
 AOI211_X4 _32379_ (.A(_07266_),
    .B(_07268_),
    .C1(_06178_),
    .C2(_06635_),
    .ZN(_07269_));
 AND2_X1 _32380_ (.A1(_07038_),
    .A2(_07258_),
    .ZN(_07270_));
 AND3_X1 _32381_ (.A1(_06189_),
    .A2(_06594_),
    .A3(_06184_),
    .ZN(_07272_));
 NOR2_X1 _32382_ (.A1(_07270_),
    .A2(_07272_),
    .ZN(_07273_));
 NAND3_X1 _32383_ (.A1(_06603_),
    .A2(_06211_),
    .A3(_06189_),
    .ZN(_07274_));
 NAND4_X1 _32384_ (.A1(_07269_),
    .A2(_06619_),
    .A3(_07273_),
    .A4(_07274_),
    .ZN(_07275_));
 AND2_X1 _32385_ (.A1(_06658_),
    .A2(_06230_),
    .ZN(_07276_));
 NOR4_X1 _32386_ (.A1(_07276_),
    .A2(_06148_),
    .A3(_06659_),
    .A4(_06661_),
    .ZN(_07277_));
 AND3_X1 _32387_ (.A1(_06668_),
    .A2(_06667_),
    .A3(_06186_),
    .ZN(_07278_));
 AND2_X1 _32388_ (.A1(_06667_),
    .A2(_06320_),
    .ZN(_07279_));
 AND2_X1 _32389_ (.A1(_06667_),
    .A2(_06230_),
    .ZN(_07280_));
 NOR3_X1 _32390_ (.A1(_07278_),
    .A2(_07279_),
    .A3(_07280_),
    .ZN(_07281_));
 AND2_X1 _32391_ (.A1(_06199_),
    .A2(_06667_),
    .ZN(_07283_));
 NOR3_X1 _32392_ (.A1(_06114_),
    .A2(_07283_),
    .A3(_07099_),
    .ZN(_07284_));
 OAI21_X1 _32393_ (.A(_06216_),
    .B1(_06199_),
    .B2(_06173_),
    .ZN(_07285_));
 OAI21_X1 _32394_ (.A(_06641_),
    .B1(_06199_),
    .B2(_06642_),
    .ZN(_07286_));
 OAI21_X1 _32395_ (.A(_06641_),
    .B1(_06153_),
    .B2(_06220_),
    .ZN(_07287_));
 OAI21_X1 _32396_ (.A(_06216_),
    .B1(_06153_),
    .B2(_06605_),
    .ZN(_07288_));
 AND4_X1 _32397_ (.A1(_07285_),
    .A2(_07286_),
    .A3(_07287_),
    .A4(_07288_),
    .ZN(_07289_));
 NAND4_X1 _32398_ (.A1(_07277_),
    .A2(_07281_),
    .A3(_07284_),
    .A4(_07289_),
    .ZN(_07290_));
 NAND4_X1 _32399_ (.A1(_06594_),
    .A2(_06184_),
    .A3(_06107_),
    .A4(_06167_),
    .ZN(_07291_));
 NAND4_X1 _32400_ (.A1(_06107_),
    .A2(_06191_),
    .A3(_06111_),
    .A4(_06167_),
    .ZN(_07292_));
 OAI211_X2 _32401_ (.A(_07291_),
    .B(_07292_),
    .C1(_06224_),
    .C2(_07267_),
    .ZN(_07294_));
 AND2_X1 _32402_ (.A1(_06156_),
    .A2(_06627_),
    .ZN(_07295_));
 NOR2_X1 _32403_ (.A1(_06224_),
    .A2(_07259_),
    .ZN(_07296_));
 OR4_X1 _32404_ (.A1(_06229_),
    .A2(_07294_),
    .A3(_07295_),
    .A4(_07296_),
    .ZN(_07297_));
 NOR2_X1 _32405_ (.A1(_07046_),
    .A2(_06139_),
    .ZN(_07298_));
 OAI21_X1 _32406_ (.A(_06236_),
    .B1(_07298_),
    .B2(_06331_),
    .ZN(_07299_));
 OAI21_X1 _32407_ (.A(_06236_),
    .B1(_06610_),
    .B2(_06220_),
    .ZN(_07300_));
 NAND2_X1 _32408_ (.A1(_07299_),
    .A2(_07300_),
    .ZN(_07301_));
 NOR4_X1 _32409_ (.A1(_07275_),
    .A2(_07290_),
    .A3(_07297_),
    .A4(_07301_),
    .ZN(_07302_));
 NAND2_X1 _32410_ (.A1(_07263_),
    .A2(_07302_),
    .ZN(_07303_));
 XNOR2_X1 _32411_ (.A(_06337_),
    .B(_07303_),
    .ZN(_07305_));
 AND4_X1 _32412_ (.A1(_05818_),
    .A2(_05735_),
    .A3(_05722_),
    .A4(_05651_),
    .ZN(_07306_));
 AND4_X1 _32413_ (.A1(_05589_),
    .A2(_05735_),
    .A3(_05726_),
    .A4(_05651_),
    .ZN(_07307_));
 AOI211_X4 _32414_ (.A(_07306_),
    .B(_07307_),
    .C1(_05751_),
    .C2(_05613_),
    .ZN(_07308_));
 AND4_X1 _32415_ (.A1(_05738_),
    .A2(_05741_),
    .A3(_05748_),
    .A4(_05745_),
    .ZN(_07309_));
 AOI211_X2 _32416_ (.A(_06409_),
    .B(_07309_),
    .C1(_06456_),
    .C2(_05751_),
    .ZN(_07310_));
 AND2_X1 _32417_ (.A1(_05770_),
    .A2(_06386_),
    .ZN(_07311_));
 NOR3_X1 _32418_ (.A1(_05773_),
    .A2(_06406_),
    .A3(_07311_),
    .ZN(_07312_));
 OAI21_X1 _32419_ (.A(_05771_),
    .B1(_06384_),
    .B2(_05641_),
    .ZN(_07313_));
 AND4_X1 _32420_ (.A1(_07308_),
    .A2(_07310_),
    .A3(_07312_),
    .A4(_07313_),
    .ZN(_07314_));
 AND2_X4 _32421_ (.A1(_05601_),
    .A2(_05673_),
    .ZN(_07316_));
 NAND2_X1 _32422_ (.A1(_07316_),
    .A2(_05815_),
    .ZN(_07317_));
 NAND2_X1 _32423_ (.A1(_06824_),
    .A2(_06455_),
    .ZN(_07318_));
 AND3_X1 _32424_ (.A1(_07317_),
    .A2(_07318_),
    .A3(_05822_),
    .ZN(_07319_));
 OAI211_X2 _32425_ (.A(_06442_),
    .B(_05817_),
    .C1(_05807_),
    .C2(_05673_),
    .ZN(_07320_));
 OAI211_X2 _32426_ (.A(_05779_),
    .B(_06371_),
    .C1(_05805_),
    .C2(_05603_),
    .ZN(_07321_));
 OAI21_X1 _32427_ (.A(_06442_),
    .B1(_05661_),
    .B2(_05800_),
    .ZN(_07322_));
 OAI21_X1 _32428_ (.A(_06442_),
    .B1(_05711_),
    .B2(_06456_),
    .ZN(_07323_));
 AND4_X1 _32429_ (.A1(_07320_),
    .A2(_07321_),
    .A3(_07322_),
    .A4(_07323_),
    .ZN(_07324_));
 OAI21_X1 _32430_ (.A(_06455_),
    .B1(_06387_),
    .B2(_05685_),
    .ZN(_07325_));
 OAI211_X2 _32431_ (.A(_06455_),
    .B(_06371_),
    .C1(_05620_),
    .C2(_05726_),
    .ZN(_07327_));
 AND4_X1 _32432_ (.A1(_07319_),
    .A2(_07324_),
    .A3(_07325_),
    .A4(_07327_),
    .ZN(_07328_));
 AND4_X1 _32433_ (.A1(_05809_),
    .A2(_05587_),
    .A3(_05726_),
    .A4(_05677_),
    .ZN(_07329_));
 AND2_X2 _32434_ (.A1(_05623_),
    .A2(_05804_),
    .ZN(_07330_));
 AOI211_X2 _32435_ (.A(_07329_),
    .B(_07330_),
    .C1(_06451_),
    .C2(_05646_),
    .ZN(_07331_));
 AND4_X1 _32436_ (.A1(_06437_),
    .A2(_05748_),
    .A3(_06371_),
    .A4(_05745_),
    .ZN(_07332_));
 AND3_X1 _32437_ (.A1(_05763_),
    .A2(_06392_),
    .A3(_05809_),
    .ZN(_07333_));
 AND2_X1 _32438_ (.A1(_05792_),
    .A2(_05660_),
    .ZN(_07334_));
 NOR4_X1 _32439_ (.A1(_07332_),
    .A2(_07333_),
    .A3(_07334_),
    .A4(_06814_),
    .ZN(_07335_));
 OAI21_X1 _32440_ (.A(_06451_),
    .B1(_06456_),
    .B2(_05729_),
    .ZN(_07336_));
 OAI211_X2 _32441_ (.A(_06451_),
    .B(_05738_),
    .C1(_05805_),
    .C2(_05818_),
    .ZN(_07338_));
 AND4_X1 _32442_ (.A1(_07331_),
    .A2(_07335_),
    .A3(_07336_),
    .A4(_07338_),
    .ZN(_07339_));
 OAI21_X1 _32443_ (.A(_05758_),
    .B1(_05659_),
    .B2(_06824_),
    .ZN(_07340_));
 NAND4_X1 _32444_ (.A1(_05736_),
    .A2(_06371_),
    .A3(_05726_),
    .A4(_05827_),
    .ZN(_07341_));
 NAND3_X1 _32445_ (.A1(_07340_),
    .A2(_06802_),
    .A3(_07341_),
    .ZN(_07342_));
 AND2_X1 _32446_ (.A1(_06403_),
    .A2(_05754_),
    .ZN(_07343_));
 AOI21_X1 _32447_ (.A(_06806_),
    .B1(_06445_),
    .B2(_06377_),
    .ZN(_07344_));
 NOR4_X1 _32448_ (.A1(_07342_),
    .A2(_07343_),
    .A3(_06428_),
    .A4(_07344_),
    .ZN(_07345_));
 NAND4_X1 _32449_ (.A1(_07314_),
    .A2(_07328_),
    .A3(_07339_),
    .A4(_07345_),
    .ZN(_07346_));
 AND3_X1 _32450_ (.A1(_05683_),
    .A2(_05630_),
    .A3(_05587_),
    .ZN(_07347_));
 AOI211_X4 _32451_ (.A(_05689_),
    .B(_07347_),
    .C1(_05683_),
    .C2(_06397_),
    .ZN(_07349_));
 INV_X1 _32452_ (.A(_05711_),
    .ZN(_07350_));
 AOI21_X1 _32453_ (.A(_05681_),
    .B1(_06361_),
    .B2(_07350_),
    .ZN(_07351_));
 AOI21_X1 _32454_ (.A(_07351_),
    .B1(_05683_),
    .B2(_05661_),
    .ZN(_07352_));
 OAI21_X1 _32455_ (.A(_05699_),
    .B1(_06387_),
    .B2(_05685_),
    .ZN(_07353_));
 NAND2_X1 _32456_ (.A1(_05691_),
    .A2(_05609_),
    .ZN(_07354_));
 AND2_X1 _32457_ (.A1(_07353_),
    .A2(_07354_),
    .ZN(_07355_));
 OAI21_X1 _32458_ (.A(_05699_),
    .B1(_05696_),
    .B2(_05711_),
    .ZN(_07356_));
 AND4_X1 _32459_ (.A1(_07349_),
    .A2(_07352_),
    .A3(_07355_),
    .A4(_07356_),
    .ZN(_07357_));
 NOR2_X1 _32460_ (.A1(_05638_),
    .A2(_05578_),
    .ZN(_07358_));
 AND2_X1 _32461_ (.A1(_07358_),
    .A2(_05579_),
    .ZN(_07360_));
 OAI21_X1 _32462_ (.A(_05656_),
    .B1(_05796_),
    .B2(_07360_),
    .ZN(_07361_));
 NOR2_X1 _32463_ (.A1(_06379_),
    .A2(_06835_),
    .ZN(_07362_));
 NAND3_X1 _32464_ (.A1(_05692_),
    .A2(_05656_),
    .A3(_05694_),
    .ZN(_07363_));
 AND2_X1 _32465_ (.A1(_07363_),
    .A2(_05663_),
    .ZN(_07364_));
 OAI21_X1 _32466_ (.A(_06381_),
    .B1(_05767_),
    .B2(_05639_),
    .ZN(_07365_));
 AND4_X1 _32467_ (.A1(_07361_),
    .A2(_07362_),
    .A3(_07364_),
    .A4(_07365_),
    .ZN(_07366_));
 AOI211_X4 _32468_ (.A(_05783_),
    .B(_06366_),
    .C1(_05805_),
    .C2(_05818_),
    .ZN(_07367_));
 OAI21_X1 _32469_ (.A(_06383_),
    .B1(_05666_),
    .B2(_05623_),
    .ZN(_07368_));
 NAND2_X1 _32470_ (.A1(_06383_),
    .A2(_05679_),
    .ZN(_07369_));
 NAND2_X1 _32471_ (.A1(_05637_),
    .A2(_05672_),
    .ZN(_07371_));
 NAND4_X1 _32472_ (.A1(_07368_),
    .A2(_06394_),
    .A3(_07369_),
    .A4(_07371_),
    .ZN(_07372_));
 NAND4_X1 _32473_ (.A1(_05738_),
    .A2(_05673_),
    .A3(_06373_),
    .A4(_05827_),
    .ZN(_07373_));
 AND2_X1 _32474_ (.A1(_05595_),
    .A2(_05596_),
    .ZN(_07374_));
 INV_X1 _32475_ (.A(_07374_),
    .ZN(_07375_));
 OAI21_X1 _32476_ (.A(_07373_),
    .B1(_06366_),
    .B2(_07375_),
    .ZN(_07376_));
 NOR4_X1 _32477_ (.A1(_07367_),
    .A2(_07372_),
    .A3(_06372_),
    .A4(_07376_),
    .ZN(_07377_));
 OAI21_X1 _32478_ (.A(_06353_),
    .B1(_05772_),
    .B2(_06386_),
    .ZN(_07378_));
 OAI211_X2 _32479_ (.A(_05708_),
    .B(_05664_),
    .C1(_05805_),
    .C2(_05578_),
    .ZN(_07379_));
 NAND2_X1 _32480_ (.A1(_05711_),
    .A2(_06353_),
    .ZN(_07380_));
 NAND2_X1 _32481_ (.A1(_05705_),
    .A2(_05657_),
    .ZN(_07382_));
 AND4_X1 _32482_ (.A1(_07378_),
    .A2(_07379_),
    .A3(_07380_),
    .A4(_07382_),
    .ZN(_07383_));
 NAND4_X1 _32483_ (.A1(_07357_),
    .A2(_07366_),
    .A3(_07377_),
    .A4(_07383_),
    .ZN(_07384_));
 NOR2_X2 _32484_ (.A1(_07346_),
    .A2(_07384_),
    .ZN(_07385_));
 AOI21_X1 _32485_ (.A(_06877_),
    .B1(_06473_),
    .B2(_05444_),
    .ZN(_07386_));
 NAND4_X1 _32486_ (.A1(_06514_),
    .A2(_05275_),
    .A3(_05441_),
    .A4(_05329_),
    .ZN(_07387_));
 AND3_X1 _32487_ (.A1(_07386_),
    .A2(_06883_),
    .A3(_07387_),
    .ZN(_07388_));
 AND3_X1 _32488_ (.A1(_05419_),
    .A2(_06522_),
    .A3(_05230_),
    .ZN(_07389_));
 NOR4_X1 _32489_ (.A1(_05481_),
    .A2(_06481_),
    .A3(_06880_),
    .A4(_07389_),
    .ZN(_07390_));
 NAND4_X1 _32490_ (.A1(_05441_),
    .A2(_06522_),
    .A3(_05233_),
    .A4(_05240_),
    .ZN(_07391_));
 NAND4_X1 _32491_ (.A1(_06514_),
    .A2(_05275_),
    .A3(_05441_),
    .A4(_05233_),
    .ZN(_07393_));
 OAI211_X2 _32492_ (.A(_07391_),
    .B(_07393_),
    .C1(_05483_),
    .C2(_05431_),
    .ZN(_07394_));
 INV_X1 _32493_ (.A(_05297_),
    .ZN(_07395_));
 AOI21_X1 _32494_ (.A(_05431_),
    .B1(_07395_),
    .B2(_05550_),
    .ZN(_07396_));
 AND3_X1 _32495_ (.A1(_05261_),
    .A2(_05498_),
    .A3(_05262_),
    .ZN(_07397_));
 NOR3_X1 _32496_ (.A1(_07394_),
    .A2(_07396_),
    .A3(_07397_),
    .ZN(_07398_));
 NAND2_X1 _32497_ (.A1(_05493_),
    .A2(_05496_),
    .ZN(_07399_));
 OAI21_X1 _32498_ (.A(_07399_),
    .B1(_05427_),
    .B2(_05428_),
    .ZN(_07400_));
 AND2_X1 _32499_ (.A1(_05496_),
    .A2(_05211_),
    .ZN(_07401_));
 NOR4_X1 _32500_ (.A1(_07400_),
    .A2(_05535_),
    .A3(_07401_),
    .A4(_06470_),
    .ZN(_07402_));
 NAND4_X1 _32501_ (.A1(_07388_),
    .A2(_07390_),
    .A3(_07398_),
    .A4(_07402_),
    .ZN(_07404_));
 OAI211_X2 _32502_ (.A(_05564_),
    .B(_06520_),
    .C1(_05310_),
    .C2(_06522_),
    .ZN(_07405_));
 AND3_X1 _32503_ (.A1(_05472_),
    .A2(_05325_),
    .A3(_07405_),
    .ZN(_07406_));
 OAI21_X1 _32504_ (.A(_05564_),
    .B1(_05398_),
    .B2(_05349_),
    .ZN(_07407_));
 OAI21_X1 _32505_ (.A(_06531_),
    .B1(_05502_),
    .B2(_05353_),
    .ZN(_07408_));
 OAI21_X1 _32506_ (.A(_06531_),
    .B1(_05373_),
    .B2(_06541_),
    .ZN(_07409_));
 NAND4_X1 _32507_ (.A1(_07406_),
    .A2(_07407_),
    .A3(_07408_),
    .A4(_07409_),
    .ZN(_07410_));
 OAI211_X2 _32508_ (.A(_05354_),
    .B(_06520_),
    .C1(_05246_),
    .C2(_06522_),
    .ZN(_07411_));
 OAI211_X2 _32509_ (.A(_05354_),
    .B(_06514_),
    .C1(_05272_),
    .C2(_05275_),
    .ZN(_07412_));
 OAI21_X1 _32510_ (.A(_05354_),
    .B1(_05337_),
    .B2(_05356_),
    .ZN(_07413_));
 NAND4_X1 _32511_ (.A1(_07411_),
    .A2(_07412_),
    .A3(_05362_),
    .A4(_07413_),
    .ZN(_07415_));
 OAI211_X2 _32512_ (.A(_06548_),
    .B(_06514_),
    .C1(_05310_),
    .C2(_05446_),
    .ZN(_07416_));
 OAI21_X1 _32513_ (.A(_06548_),
    .B1(_05353_),
    .B2(_05307_),
    .ZN(_07417_));
 OAI21_X1 _32514_ (.A(_06548_),
    .B1(_05497_),
    .B2(_05373_),
    .ZN(_07418_));
 OAI21_X1 _32515_ (.A(_06548_),
    .B1(_05296_),
    .B2(_06541_),
    .ZN(_07419_));
 NAND4_X1 _32516_ (.A1(_07416_),
    .A2(_07417_),
    .A3(_07418_),
    .A4(_07419_),
    .ZN(_07420_));
 NOR4_X1 _32517_ (.A1(_07404_),
    .A2(_07410_),
    .A3(_07415_),
    .A4(_07420_),
    .ZN(_07421_));
 OAI211_X2 _32518_ (.A(_05384_),
    .B(_05283_),
    .C1(_05318_),
    .C2(_06541_),
    .ZN(_07422_));
 NAND2_X1 _32519_ (.A1(_05405_),
    .A2(_05402_),
    .ZN(_07423_));
 NAND4_X1 _32520_ (.A1(_06527_),
    .A2(_07422_),
    .A3(_06909_),
    .A4(_07423_),
    .ZN(_07424_));
 AND2_X1 _32521_ (.A1(_05219_),
    .A2(_05446_),
    .ZN(_07426_));
 INV_X1 _32522_ (.A(_07426_),
    .ZN(_07427_));
 AOI21_X1 _32523_ (.A(_05556_),
    .B1(_07427_),
    .B2(_05550_),
    .ZN(_07428_));
 AOI21_X1 _32524_ (.A(_05556_),
    .B1(_05277_),
    .B2(_05336_),
    .ZN(_07429_));
 NOR3_X1 _32525_ (.A1(_07424_),
    .A2(_07428_),
    .A3(_07429_),
    .ZN(_07430_));
 OAI21_X1 _32526_ (.A(_05270_),
    .B1(_05263_),
    .B2(_05296_),
    .ZN(_07431_));
 OAI21_X1 _32527_ (.A(_05270_),
    .B1(_05337_),
    .B2(_05356_),
    .ZN(_07432_));
 OAI211_X2 _32528_ (.A(_07431_),
    .B(_07432_),
    .C1(_05504_),
    .C2(_05278_),
    .ZN(_07433_));
 OAI21_X1 _32529_ (.A(_06928_),
    .B1(_05349_),
    .B2(_05493_),
    .ZN(_07434_));
 OAI21_X1 _32530_ (.A(_06503_),
    .B1(_05381_),
    .B2(_05353_),
    .ZN(_07435_));
 NAND2_X1 _32531_ (.A1(_05296_),
    .A2(_06928_),
    .ZN(_07437_));
 NAND4_X1 _32532_ (.A1(_07434_),
    .A2(_07435_),
    .A3(_07437_),
    .A4(_05547_),
    .ZN(_07438_));
 NAND3_X1 _32533_ (.A1(_06488_),
    .A2(_05255_),
    .A3(_06514_),
    .ZN(_07439_));
 NAND3_X1 _32534_ (.A1(_06488_),
    .A2(_05232_),
    .A3(_06514_),
    .ZN(_07440_));
 OAI211_X2 _32535_ (.A(_07439_),
    .B(_07440_),
    .C1(_05408_),
    .C2(_06486_),
    .ZN(_07441_));
 NAND2_X1 _32536_ (.A1(_05296_),
    .A2(_05244_),
    .ZN(_07442_));
 NAND4_X1 _32537_ (.A1(_06520_),
    .A2(_05272_),
    .A3(_05329_),
    .A4(_05215_),
    .ZN(_07443_));
 OAI211_X2 _32538_ (.A(_07442_),
    .B(_07443_),
    .C1(_05326_),
    .C2(_06486_),
    .ZN(_07444_));
 NOR4_X1 _32539_ (.A1(_07433_),
    .A2(_07438_),
    .A3(_07441_),
    .A4(_07444_),
    .ZN(_07445_));
 OAI21_X1 _32540_ (.A(_05392_),
    .B1(_05541_),
    .B2(_05507_),
    .ZN(_07446_));
 OAI211_X2 _32541_ (.A(_05384_),
    .B(_05329_),
    .C1(_05337_),
    .C2(_05356_),
    .ZN(_07448_));
 AND3_X1 _32542_ (.A1(_07446_),
    .A2(_06519_),
    .A3(_07448_),
    .ZN(_07449_));
 INV_X1 _32543_ (.A(_05394_),
    .ZN(_07450_));
 AOI21_X1 _32544_ (.A(_07450_),
    .B1(_06498_),
    .B2(_05363_),
    .ZN(_07451_));
 AND2_X1 _32545_ (.A1(_05381_),
    .A2(_05395_),
    .ZN(_07452_));
 AND2_X1 _32546_ (.A1(_05395_),
    .A2(_05378_),
    .ZN(_07453_));
 AND3_X1 _32547_ (.A1(_05369_),
    .A2(_05265_),
    .A3(_05252_),
    .ZN(_07454_));
 NOR4_X1 _32548_ (.A1(_07451_),
    .A2(_07452_),
    .A3(_07453_),
    .A4(_07454_),
    .ZN(_07455_));
 AND4_X1 _32549_ (.A1(_07430_),
    .A2(_07445_),
    .A3(_07449_),
    .A4(_07455_),
    .ZN(_07456_));
 NAND2_X1 _32550_ (.A1(_07421_),
    .A2(_07456_),
    .ZN(_07457_));
 XOR2_X1 _32551_ (.A(_07385_),
    .B(_07457_),
    .Z(_07459_));
 XNOR2_X2 _32552_ (.A(_07305_),
    .B(_07459_),
    .ZN(_07460_));
 XNOR2_X1 _32553_ (.A(_07220_),
    .B(_07460_),
    .ZN(_07461_));
 MUX2_X1 _32554_ (.A(_07131_),
    .B(_07461_),
    .S(_05156_),
    .Z(_00703_));
 MUX2_X1 _32555_ (.A(_17041_),
    .B(_16913_),
    .S(_03836_),
    .Z(_00761_));
 MUX2_X1 _32556_ (.A(_17042_),
    .B(_16914_),
    .S(_03836_),
    .Z(_00762_));
 XOR2_X1 _32557_ (.A(_17202_),
    .B(_17013_),
    .Z(_07462_));
 NAND2_X1 _32558_ (.A1(_06326_),
    .A2(_06113_),
    .ZN(_07463_));
 NAND2_X1 _32559_ (.A1(_06597_),
    .A2(_07463_),
    .ZN(_07464_));
 INV_X1 _32560_ (.A(_07233_),
    .ZN(_07465_));
 OAI21_X1 _32561_ (.A(_07465_),
    .B1(_06302_),
    .B2(_07067_),
    .ZN(_07467_));
 AOI211_X4 _32562_ (.A(_07464_),
    .B(_07467_),
    .C1(_06326_),
    .C2(_06134_),
    .ZN(_07468_));
 AND2_X1 _32563_ (.A1(_06319_),
    .A2(_06230_),
    .ZN(_07469_));
 AND3_X1 _32564_ (.A1(_06319_),
    .A2(_06186_),
    .A3(_06668_),
    .ZN(_07470_));
 AOI211_X4 _32565_ (.A(_07469_),
    .B(_07470_),
    .C1(_06605_),
    .C2(_06319_),
    .ZN(_07471_));
 NAND4_X1 _32566_ (.A1(_06298_),
    .A2(_06205_),
    .A3(_06143_),
    .A4(_06206_),
    .ZN(_07472_));
 OAI211_X2 _32567_ (.A(_06330_),
    .B(_06289_),
    .C1(_06192_),
    .C2(_06294_),
    .ZN(_07473_));
 AND3_X4 _32568_ (.A1(_07471_),
    .A2(_07472_),
    .A3(_07473_),
    .ZN(_07474_));
 NOR2_X1 _32569_ (.A1(_07058_),
    .A2(_07071_),
    .ZN(_07475_));
 AND2_X1 _32570_ (.A1(_06309_),
    .A2(_06164_),
    .ZN(_07476_));
 AND2_X1 _32571_ (.A1(_06309_),
    .A2(_06175_),
    .ZN(_07478_));
 NOR4_X1 _32572_ (.A1(_07475_),
    .A2(_07261_),
    .A3(_07476_),
    .A4(_07478_),
    .ZN(_07479_));
 AND2_X1 _32573_ (.A1(_06212_),
    .A2(_06301_),
    .ZN(_07480_));
 AND3_X1 _32574_ (.A1(_06657_),
    .A2(_06203_),
    .A3(_06298_),
    .ZN(_07481_));
 NOR4_X1 _32575_ (.A1(_07480_),
    .A2(_07076_),
    .A3(_07250_),
    .A4(_07481_),
    .ZN(_07482_));
 NAND4_X1 _32576_ (.A1(_07468_),
    .A2(_07474_),
    .A3(_07479_),
    .A4(_07482_),
    .ZN(_07483_));
 OAI211_X2 _32577_ (.A(_06257_),
    .B(_06594_),
    .C1(_06205_),
    .C2(_06294_),
    .ZN(_07484_));
 OAI211_X2 _32578_ (.A(_06257_),
    .B(_06289_),
    .C1(_06111_),
    .C2(_06139_),
    .ZN(_07485_));
 OAI21_X1 _32579_ (.A(_06257_),
    .B1(_06291_),
    .B2(_06134_),
    .ZN(_07486_));
 NAND4_X1 _32580_ (.A1(_07484_),
    .A2(_07485_),
    .A3(_06581_),
    .A4(_07486_),
    .ZN(_07487_));
 OAI211_X2 _32581_ (.A(_07222_),
    .B(_06289_),
    .C1(_06192_),
    .C2(_06194_),
    .ZN(_07489_));
 OAI211_X2 _32582_ (.A(_07222_),
    .B(_06206_),
    .C1(_06120_),
    .C2(_06184_),
    .ZN(_07490_));
 OAI211_X2 _32583_ (.A(_07222_),
    .B(_06594_),
    .C1(_06205_),
    .C2(_06194_),
    .ZN(_07491_));
 OAI21_X1 _32584_ (.A(_07222_),
    .B1(_06304_),
    .B2(_06605_),
    .ZN(_07492_));
 NAND4_X1 _32585_ (.A1(_07489_),
    .A2(_07490_),
    .A3(_07491_),
    .A4(_07492_),
    .ZN(_07493_));
 AND2_X1 _32586_ (.A1(_06273_),
    .A2(_06331_),
    .ZN(_07494_));
 INV_X1 _32587_ (.A(_07494_),
    .ZN(_07495_));
 NAND3_X1 _32588_ (.A1(_06274_),
    .A2(_06139_),
    .A3(_06289_),
    .ZN(_07496_));
 OAI211_X2 _32589_ (.A(_07495_),
    .B(_07496_),
    .C1(_07115_),
    .C2(_06311_),
    .ZN(_07497_));
 AOI21_X1 _32590_ (.A(_07115_),
    .B1(_06561_),
    .B2(_07267_),
    .ZN(_07498_));
 NOR4_X1 _32591_ (.A1(_07497_),
    .A2(_06569_),
    .A3(_06566_),
    .A4(_07498_),
    .ZN(_07500_));
 OAI21_X1 _32592_ (.A(_06572_),
    .B1(_06164_),
    .B2(_06113_),
    .ZN(_07501_));
 NAND2_X1 _32593_ (.A1(_06572_),
    .A2(_06605_),
    .ZN(_07502_));
 NAND3_X1 _32594_ (.A1(_06218_),
    .A2(_06203_),
    .A3(_06246_),
    .ZN(_07503_));
 AND4_X1 _32595_ (.A1(_06286_),
    .A2(_07501_),
    .A3(_07502_),
    .A4(_07503_),
    .ZN(_07504_));
 NAND2_X1 _32596_ (.A1(_07500_),
    .A2(_07504_),
    .ZN(_07505_));
 NOR4_X2 _32597_ (.A1(_07483_),
    .A2(_07487_),
    .A3(_07493_),
    .A4(_07505_),
    .ZN(_07506_));
 AOI211_X4 _32598_ (.A(_06630_),
    .B(_06632_),
    .C1(_06304_),
    .C2(_06635_),
    .ZN(_07507_));
 OAI21_X1 _32599_ (.A(_06189_),
    .B1(_07298_),
    .B2(_06159_),
    .ZN(_07508_));
 AND2_X1 _32600_ (.A1(_06304_),
    .A2(_06188_),
    .ZN(_07509_));
 AOI221_X4 _32601_ (.A(_07509_),
    .B1(_06631_),
    .B2(_06189_),
    .C1(_06184_),
    .C2(_07038_),
    .ZN(_07511_));
 OAI21_X1 _32602_ (.A(_06635_),
    .B1(_06156_),
    .B2(_06591_),
    .ZN(_07512_));
 NAND4_X1 _32603_ (.A1(_07507_),
    .A2(_07508_),
    .A3(_07511_),
    .A4(_07512_),
    .ZN(_07513_));
 AND2_X1 _32604_ (.A1(_06108_),
    .A2(_06568_),
    .ZN(_07514_));
 AND3_X1 _32605_ (.A1(_06220_),
    .A2(_06103_),
    .A3(_06107_),
    .ZN(_07515_));
 AOI221_X4 _32606_ (.A(_07514_),
    .B1(_06605_),
    .B2(_06108_),
    .C1(_06194_),
    .C2(_07515_),
    .ZN(_07516_));
 AND2_X1 _32607_ (.A1(_06594_),
    .A2(_06192_),
    .ZN(_07517_));
 OAI21_X1 _32608_ (.A(_06658_),
    .B1(_06230_),
    .B2(_07517_),
    .ZN(_07518_));
 OAI21_X1 _32609_ (.A(_06658_),
    .B1(_07298_),
    .B2(_06642_),
    .ZN(_07519_));
 NOR3_X1 _32610_ (.A1(_06135_),
    .A2(_07283_),
    .A3(_07099_),
    .ZN(_07520_));
 NAND4_X1 _32611_ (.A1(_07516_),
    .A2(_07518_),
    .A3(_07519_),
    .A4(_07520_),
    .ZN(_07522_));
 NAND2_X1 _32612_ (.A1(_06641_),
    .A2(_06175_),
    .ZN(_07523_));
 NAND2_X1 _32613_ (.A1(_06641_),
    .A2(_06191_),
    .ZN(_07524_));
 OAI21_X1 _32614_ (.A(_06198_),
    .B1(_06657_),
    .B2(_06642_),
    .ZN(_07525_));
 AND4_X1 _32615_ (.A1(_07091_),
    .A2(_07523_),
    .A3(_07524_),
    .A4(_07525_),
    .ZN(_07526_));
 OAI211_X2 _32616_ (.A(_06216_),
    .B(_06206_),
    .C1(_06192_),
    .C2(_06294_),
    .ZN(_07527_));
 OAI21_X1 _32617_ (.A(_06216_),
    .B1(_06121_),
    .B2(_06258_),
    .ZN(_07528_));
 NAND4_X1 _32618_ (.A1(_07526_),
    .A2(_07085_),
    .A3(_07527_),
    .A4(_07528_),
    .ZN(_07529_));
 INV_X1 _32619_ (.A(_06231_),
    .ZN(_07530_));
 NAND2_X1 _32620_ (.A1(_06304_),
    .A2(_06236_),
    .ZN(_07531_));
 NAND3_X1 _32621_ (.A1(_06185_),
    .A2(_06186_),
    .A3(_06236_),
    .ZN(_07533_));
 OAI21_X1 _32622_ (.A(_06627_),
    .B1(_06218_),
    .B2(_06657_),
    .ZN(_07534_));
 NAND4_X1 _32623_ (.A1(_07530_),
    .A2(_07531_),
    .A3(_07533_),
    .A4(_07534_),
    .ZN(_07535_));
 NOR4_X1 _32624_ (.A1(_07513_),
    .A2(_07522_),
    .A3(_07529_),
    .A4(_07535_),
    .ZN(_07536_));
 AND2_X2 _32625_ (.A1(_07506_),
    .A2(_07536_),
    .ZN(_07537_));
 XOR2_X2 _32626_ (.A(_07537_),
    .B(_06337_),
    .Z(_07538_));
 OAI21_X1 _32627_ (.A(_06946_),
    .B1(_05964_),
    .B2(_05967_),
    .ZN(_07539_));
 AND4_X1 _32628_ (.A1(_05999_),
    .A2(_05858_),
    .A3(_05902_),
    .A4(_05880_),
    .ZN(_07540_));
 AOI21_X1 _32629_ (.A(_06007_),
    .B1(_05998_),
    .B2(_05979_),
    .ZN(_07541_));
 AOI211_X2 _32630_ (.A(_07540_),
    .B(_07541_),
    .C1(_05915_),
    .C2(_06002_),
    .ZN(_07542_));
 OAI211_X2 _32631_ (.A(_06946_),
    .B(_05975_),
    .C1(_05999_),
    .C2(_05854_),
    .ZN(_07544_));
 OAI21_X1 _32632_ (.A(_06946_),
    .B1(_05873_),
    .B2(_06044_),
    .ZN(_07545_));
 AND4_X1 _32633_ (.A1(_07539_),
    .A2(_07542_),
    .A3(_07544_),
    .A4(_07545_),
    .ZN(_07546_));
 INV_X1 _32634_ (.A(_05866_),
    .ZN(_07547_));
 NAND2_X1 _32635_ (.A1(_05914_),
    .A2(_06046_),
    .ZN(_07548_));
 NAND3_X1 _32636_ (.A1(_05914_),
    .A2(_06059_),
    .A3(_06727_),
    .ZN(_07549_));
 OAI211_X2 _32637_ (.A(_05914_),
    .B(_05884_),
    .C1(_05900_),
    .C2(_05868_),
    .ZN(_07550_));
 NAND4_X1 _32638_ (.A1(_07547_),
    .A2(_07548_),
    .A3(_07549_),
    .A4(_07550_),
    .ZN(_07551_));
 AND2_X1 _32639_ (.A1(_05920_),
    .A2(_05999_),
    .ZN(_07552_));
 OAI21_X1 _32640_ (.A(_05921_),
    .B1(_05873_),
    .B2(_06044_),
    .ZN(_07553_));
 NAND2_X1 _32641_ (.A1(_05921_),
    .A2(_06016_),
    .ZN(_07555_));
 NAND3_X1 _32642_ (.A1(_07553_),
    .A2(_06970_),
    .A3(_07555_),
    .ZN(_07556_));
 NOR4_X1 _32643_ (.A1(_07551_),
    .A2(_05989_),
    .A3(_07552_),
    .A4(_07556_),
    .ZN(_07557_));
 AND3_X1 _32644_ (.A1(_05860_),
    .A2(_05837_),
    .A3(_05836_),
    .ZN(_07558_));
 AOI211_X4 _32645_ (.A(_07558_),
    .B(_05845_),
    .C1(_05865_),
    .C2(_06089_),
    .ZN(_07559_));
 OAI21_X1 _32646_ (.A(_05908_),
    .B1(_06025_),
    .B2(_05909_),
    .ZN(_07560_));
 NAND2_X1 _32647_ (.A1(_05908_),
    .A2(_05912_),
    .ZN(_07561_));
 AND2_X1 _32648_ (.A1(_07560_),
    .A2(_07561_),
    .ZN(_07562_));
 OAI21_X1 _32649_ (.A(_05908_),
    .B1(_05934_),
    .B2(_06680_),
    .ZN(_07563_));
 AND4_X1 _32650_ (.A1(_06681_),
    .A2(_07559_),
    .A3(_07562_),
    .A4(_07563_),
    .ZN(_07564_));
 NAND2_X1 _32651_ (.A1(_06692_),
    .A2(_05926_),
    .ZN(_07566_));
 NAND2_X1 _32652_ (.A1(_05972_),
    .A2(_05860_),
    .ZN(_07567_));
 OR2_X1 _32653_ (.A1(_06716_),
    .A2(_06060_),
    .ZN(_07568_));
 NAND2_X1 _32654_ (.A1(_05972_),
    .A2(_05997_),
    .ZN(_07569_));
 OAI21_X1 _32655_ (.A(_05972_),
    .B1(_05934_),
    .B2(_06010_),
    .ZN(_07570_));
 AND4_X1 _32656_ (.A1(_07567_),
    .A2(_07568_),
    .A3(_07569_),
    .A4(_07570_),
    .ZN(_07571_));
 AOI21_X1 _32657_ (.A(_06993_),
    .B1(_05964_),
    .B2(_05926_),
    .ZN(_07572_));
 AND4_X1 _32658_ (.A1(_07566_),
    .A2(_07571_),
    .A3(_06711_),
    .A4(_07572_),
    .ZN(_07573_));
 NAND4_X1 _32659_ (.A1(_07546_),
    .A2(_07557_),
    .A3(_07564_),
    .A4(_07573_),
    .ZN(_07574_));
 OAI21_X1 _32660_ (.A(_05895_),
    .B1(_05865_),
    .B2(_05860_),
    .ZN(_07575_));
 NOR4_X1 _32661_ (.A1(_06749_),
    .A2(_06076_),
    .A3(_06751_),
    .A4(_07025_),
    .ZN(_07577_));
 NAND4_X1 _32662_ (.A1(_06063_),
    .A2(_05956_),
    .A3(_05893_),
    .A4(_05871_),
    .ZN(_07578_));
 OAI21_X1 _32663_ (.A(_05895_),
    .B1(_06004_),
    .B2(_06044_),
    .ZN(_07579_));
 AND4_X1 _32664_ (.A1(_07575_),
    .A2(_07577_),
    .A3(_07578_),
    .A4(_07579_),
    .ZN(_07580_));
 AOI21_X1 _32665_ (.A(_06085_),
    .B1(_06748_),
    .B2(_06067_),
    .ZN(_07581_));
 AOI21_X1 _32666_ (.A(_06085_),
    .B1(_06959_),
    .B2(_06020_),
    .ZN(_07582_));
 AOI21_X1 _32667_ (.A(_05939_),
    .B1(_05998_),
    .B2(_05886_),
    .ZN(_07583_));
 NOR4_X1 _32668_ (.A1(_07581_),
    .A2(_07582_),
    .A3(_07583_),
    .A4(_06780_),
    .ZN(_07584_));
 OAI211_X2 _32669_ (.A(_06024_),
    .B(_05956_),
    .C1(_05871_),
    .C2(_06034_),
    .ZN(_07585_));
 OAI21_X1 _32670_ (.A(_07585_),
    .B1(_06772_),
    .B2(_05979_),
    .ZN(_07586_));
 OAI21_X1 _32671_ (.A(_06024_),
    .B1(_05943_),
    .B2(_05912_),
    .ZN(_07588_));
 NAND2_X1 _32672_ (.A1(_06024_),
    .A2(_05865_),
    .ZN(_07589_));
 NAND2_X1 _32673_ (.A1(_07588_),
    .A2(_07589_),
    .ZN(_07590_));
 AOI21_X1 _32674_ (.A(_05946_),
    .B1(_06717_),
    .B2(_06718_),
    .ZN(_07591_));
 NOR4_X1 _32675_ (.A1(_07586_),
    .A2(_06984_),
    .A3(_07590_),
    .A4(_07591_),
    .ZN(_07592_));
 INV_X1 _32676_ (.A(_06706_),
    .ZN(_07593_));
 AOI21_X1 _32677_ (.A(_06081_),
    .B1(_07593_),
    .B2(_07206_),
    .ZN(_07594_));
 AOI21_X1 _32678_ (.A(_06081_),
    .B1(_06712_),
    .B2(_05944_),
    .ZN(_07595_));
 AOI21_X1 _32679_ (.A(_07162_),
    .B1(_06684_),
    .B2(_05897_),
    .ZN(_07596_));
 NOR4_X1 _32680_ (.A1(_07594_),
    .A2(_06080_),
    .A3(_07595_),
    .A4(_07596_),
    .ZN(_07597_));
 NAND4_X1 _32681_ (.A1(_07580_),
    .A2(_07584_),
    .A3(_07592_),
    .A4(_07597_),
    .ZN(_07599_));
 NOR2_X2 _32682_ (.A1(_07574_),
    .A2(_07599_),
    .ZN(_07600_));
 XOR2_X1 _32683_ (.A(_07538_),
    .B(_07600_),
    .Z(_07601_));
 OAI21_X1 _32684_ (.A(_06353_),
    .B1(_07316_),
    .B2(_05713_),
    .ZN(_07602_));
 OAI211_X2 _32685_ (.A(_06353_),
    .B(_05589_),
    .C1(_05805_),
    .C2(_05818_),
    .ZN(_07603_));
 AND2_X1 _32686_ (.A1(_07602_),
    .A2(_07603_),
    .ZN(_07604_));
 AOI21_X1 _32687_ (.A(_06360_),
    .B1(_06361_),
    .B2(_07350_),
    .ZN(_07605_));
 INV_X1 _32688_ (.A(_06386_),
    .ZN(_07606_));
 OAI21_X1 _32689_ (.A(_07354_),
    .B1(_06360_),
    .B2(_07606_),
    .ZN(_07607_));
 AND3_X1 _32690_ (.A1(_05622_),
    .A2(_06392_),
    .A3(_05675_),
    .ZN(_07608_));
 AND3_X1 _32691_ (.A1(_07316_),
    .A2(_06392_),
    .A3(_05675_),
    .ZN(_07610_));
 NOR4_X1 _32692_ (.A1(_07605_),
    .A2(_07607_),
    .A3(_07608_),
    .A4(_07610_),
    .ZN(_07611_));
 NAND2_X1 _32693_ (.A1(_06354_),
    .A2(_05671_),
    .ZN(_07612_));
 AND3_X1 _32694_ (.A1(_05671_),
    .A2(_05601_),
    .A3(_05591_),
    .ZN(_07613_));
 INV_X1 _32695_ (.A(_07613_),
    .ZN(_07614_));
 NAND3_X1 _32696_ (.A1(_05683_),
    .A2(_05589_),
    .A3(_05726_),
    .ZN(_07615_));
 AND4_X1 _32697_ (.A1(_07612_),
    .A2(_07614_),
    .A3(_06862_),
    .A4(_07615_),
    .ZN(_07616_));
 OAI21_X1 _32698_ (.A(_05708_),
    .B1(_05696_),
    .B2(_05672_),
    .ZN(_07617_));
 AND3_X1 _32699_ (.A1(_07617_),
    .A2(_05704_),
    .A3(_06346_),
    .ZN(_07618_));
 AND4_X1 _32700_ (.A1(_07604_),
    .A2(_07611_),
    .A3(_07616_),
    .A4(_07618_),
    .ZN(_07619_));
 NAND2_X1 _32701_ (.A1(_05656_),
    .A2(_05613_),
    .ZN(_07621_));
 INV_X1 _32702_ (.A(_05655_),
    .ZN(_07622_));
 OAI21_X1 _32703_ (.A(_07621_),
    .B1(_07622_),
    .B2(_06795_),
    .ZN(_07623_));
 NAND4_X1 _32704_ (.A1(_06373_),
    .A2(_05672_),
    .A3(_05652_),
    .A4(_05805_),
    .ZN(_07624_));
 OAI21_X1 _32705_ (.A(_07624_),
    .B1(_07622_),
    .B2(_06449_),
    .ZN(_07625_));
 AND2_X1 _32706_ (.A1(_06841_),
    .A2(_05655_),
    .ZN(_07626_));
 AND4_X1 _32707_ (.A1(_05817_),
    .A2(_06373_),
    .A3(_05726_),
    .A4(_05652_),
    .ZN(_07627_));
 NOR4_X1 _32708_ (.A1(_07623_),
    .A2(_07625_),
    .A3(_07626_),
    .A4(_07627_),
    .ZN(_07628_));
 AOI211_X4 _32709_ (.A(_06389_),
    .B(_05626_),
    .C1(_05712_),
    .C2(_05818_),
    .ZN(_07629_));
 AND2_X1 _32710_ (.A1(_06381_),
    .A2(_05639_),
    .ZN(_07630_));
 AND2_X1 _32711_ (.A1(_06821_),
    .A2(_06381_),
    .ZN(_07632_));
 AND2_X1 _32712_ (.A1(_05719_),
    .A2(_06381_),
    .ZN(_07633_));
 NOR4_X1 _32713_ (.A1(_07629_),
    .A2(_07630_),
    .A3(_07632_),
    .A4(_07633_),
    .ZN(_07634_));
 AND2_X1 _32714_ (.A1(_05637_),
    .A2(_05794_),
    .ZN(_07635_));
 INV_X1 _32715_ (.A(_07635_),
    .ZN(_07636_));
 NAND3_X1 _32716_ (.A1(_07636_),
    .A2(_05645_),
    .A3(_05647_),
    .ZN(_07637_));
 NAND2_X1 _32717_ (.A1(_05772_),
    .A2(_05576_),
    .ZN(_07638_));
 NAND4_X1 _32718_ (.A1(_05573_),
    .A2(_05722_),
    .A3(_05620_),
    .A4(_05677_),
    .ZN(_07639_));
 OAI211_X2 _32719_ (.A(_07638_),
    .B(_07639_),
    .C1(_05721_),
    .C2(_06366_),
    .ZN(_07640_));
 OAI21_X1 _32720_ (.A(_07369_),
    .B1(_07371_),
    .B2(_05748_),
    .ZN(_07641_));
 NOR4_X1 _32721_ (.A1(_07637_),
    .A2(_06367_),
    .A3(_07640_),
    .A4(_07641_),
    .ZN(_07643_));
 NAND4_X1 _32722_ (.A1(_07619_),
    .A2(_07628_),
    .A3(_07634_),
    .A4(_07643_),
    .ZN(_07644_));
 AOI221_X1 _32723_ (.A(_07311_),
    .B1(_05616_),
    .B2(_05770_),
    .C1(_05596_),
    .C2(_06406_),
    .ZN(_07645_));
 OAI21_X1 _32724_ (.A(_05751_),
    .B1(_05794_),
    .B2(_05762_),
    .ZN(_07646_));
 OAI21_X1 _32725_ (.A(_05751_),
    .B1(_06403_),
    .B2(_05796_),
    .ZN(_07647_));
 AND4_X1 _32726_ (.A1(_05740_),
    .A2(_07645_),
    .A3(_07646_),
    .A4(_07647_),
    .ZN(_07648_));
 NAND3_X1 _32727_ (.A1(_05719_),
    .A2(_05636_),
    .A3(_05789_),
    .ZN(_07649_));
 AND4_X1 _32728_ (.A1(_05596_),
    .A2(_05587_),
    .A3(_05789_),
    .A4(_05677_),
    .ZN(_07650_));
 AND2_X1 _32729_ (.A1(_05803_),
    .A2(_05583_),
    .ZN(_07651_));
 AOI211_X2 _32730_ (.A(_07650_),
    .B(_07651_),
    .C1(_05804_),
    .C2(_06830_),
    .ZN(_07652_));
 OAI21_X1 _32731_ (.A(_06437_),
    .B1(_05762_),
    .B2(_05646_),
    .ZN(_07654_));
 OAI21_X1 _32732_ (.A(_06437_),
    .B1(_06421_),
    .B2(_06456_),
    .ZN(_07655_));
 AND4_X1 _32733_ (.A1(_07649_),
    .A2(_07652_),
    .A3(_07654_),
    .A4(_07655_),
    .ZN(_07656_));
 OAI211_X2 _32734_ (.A(_06455_),
    .B(_05579_),
    .C1(_05578_),
    .C2(_05673_),
    .ZN(_07657_));
 OAI21_X1 _32735_ (.A(_05779_),
    .B1(_05664_),
    .B2(_05685_),
    .ZN(_07658_));
 OAI21_X1 _32736_ (.A(_05779_),
    .B1(_05788_),
    .B2(_05800_),
    .ZN(_07659_));
 AND4_X1 _32737_ (.A1(_05821_),
    .A2(_07657_),
    .A3(_07658_),
    .A4(_07659_),
    .ZN(_07660_));
 INV_X1 _32738_ (.A(_06420_),
    .ZN(_07661_));
 OAI21_X1 _32739_ (.A(_05755_),
    .B1(_05719_),
    .B2(_05623_),
    .ZN(_07662_));
 OAI21_X1 _32740_ (.A(_05758_),
    .B1(_05767_),
    .B2(_06824_),
    .ZN(_07663_));
 OAI21_X1 _32741_ (.A(_05755_),
    .B1(_06390_),
    .B2(_06824_),
    .ZN(_07665_));
 AND4_X1 _32742_ (.A1(_07661_),
    .A2(_07662_),
    .A3(_07663_),
    .A4(_07665_),
    .ZN(_07666_));
 NAND4_X1 _32743_ (.A1(_07648_),
    .A2(_07656_),
    .A3(_07660_),
    .A4(_07666_),
    .ZN(_07667_));
 NOR2_X2 _32744_ (.A1(_07644_),
    .A2(_07667_),
    .ZN(_07668_));
 OAI21_X1 _32745_ (.A(_05375_),
    .B1(_05521_),
    .B2(_05497_),
    .ZN(_07669_));
 AND4_X1 _32746_ (.A1(_05369_),
    .A2(_05275_),
    .A3(_05239_),
    .A4(_05212_),
    .ZN(_07670_));
 AND2_X1 _32747_ (.A1(_05399_),
    .A2(_05370_),
    .ZN(_07671_));
 AOI211_X2 _32748_ (.A(_07670_),
    .B(_07671_),
    .C1(_05341_),
    .C2(_05375_),
    .ZN(_07672_));
 OAI21_X1 _32749_ (.A(_05375_),
    .B1(_06541_),
    .B2(_05517_),
    .ZN(_07673_));
 OAI21_X1 _32750_ (.A(_05405_),
    .B1(_05339_),
    .B2(_05473_),
    .ZN(_07674_));
 OAI211_X2 _32751_ (.A(_05384_),
    .B(_05283_),
    .C1(_05371_),
    .C2(_05517_),
    .ZN(_07676_));
 AND3_X1 _32752_ (.A1(_07674_),
    .A2(_07423_),
    .A3(_07676_),
    .ZN(_07677_));
 AND4_X1 _32753_ (.A1(_07669_),
    .A2(_07672_),
    .A3(_07673_),
    .A4(_07677_),
    .ZN(_07678_));
 INV_X1 _32754_ (.A(_06471_),
    .ZN(_07679_));
 AOI21_X1 _32755_ (.A(_07450_),
    .B1(_07679_),
    .B2(_05483_),
    .ZN(_07680_));
 AOI21_X1 _32756_ (.A(_07450_),
    .B1(_06498_),
    .B2(_05326_),
    .ZN(_07681_));
 OAI21_X2 _32757_ (.A(_05392_),
    .B1(_06500_),
    .B2(_05378_),
    .ZN(_07682_));
 NAND2_X1 _32758_ (.A1(_07682_),
    .A2(_06521_),
    .ZN(_07683_));
 AND2_X1 _32759_ (.A1(_05395_),
    .A2(_05383_),
    .ZN(_07684_));
 NOR4_X2 _32760_ (.A1(_07680_),
    .A2(_07681_),
    .A3(_07683_),
    .A4(_07684_),
    .ZN(_07685_));
 INV_X1 _32761_ (.A(_05241_),
    .ZN(_07687_));
 NAND2_X1 _32762_ (.A1(_07687_),
    .A2(_06488_),
    .ZN(_07688_));
 NAND2_X1 _32763_ (.A1(_05267_),
    .A2(_05334_),
    .ZN(_07689_));
 OAI211_X2 _32764_ (.A(_05267_),
    .B(_05229_),
    .C1(_05310_),
    .C2(_05248_),
    .ZN(_07690_));
 OAI21_X1 _32765_ (.A(_05267_),
    .B1(_05371_),
    .B2(_05296_),
    .ZN(_07691_));
 NAND2_X1 _32766_ (.A1(_05541_),
    .A2(_05267_),
    .ZN(_07692_));
 AND4_X1 _32767_ (.A1(_07689_),
    .A2(_07690_),
    .A3(_07691_),
    .A4(_07692_),
    .ZN(_07693_));
 NAND3_X1 _32768_ (.A1(_06488_),
    .A2(_05275_),
    .A3(_05230_),
    .ZN(_07694_));
 AND2_X4 _32769_ (.A1(_06929_),
    .A2(_05245_),
    .ZN(_07695_));
 AOI21_X1 _32770_ (.A(_07695_),
    .B1(_05529_),
    .B2(_05245_),
    .ZN(_07696_));
 AND4_X1 _32771_ (.A1(_07688_),
    .A2(_07693_),
    .A3(_07694_),
    .A4(_07696_),
    .ZN(_07698_));
 OAI211_X2 _32772_ (.A(_06928_),
    .B(_05230_),
    .C1(_05310_),
    .C2(_06522_),
    .ZN(_07699_));
 OAI21_X1 _32773_ (.A(_06503_),
    .B1(_05263_),
    .B2(_05252_),
    .ZN(_07700_));
 OAI21_X1 _32774_ (.A(_06928_),
    .B1(_05541_),
    .B2(_05297_),
    .ZN(_07701_));
 OAI211_X2 _32775_ (.A(_05289_),
    .B(_05273_),
    .C1(_05240_),
    .C2(_05230_),
    .ZN(_07702_));
 AND4_X1 _32776_ (.A1(_07699_),
    .A2(_07700_),
    .A3(_07701_),
    .A4(_07702_),
    .ZN(_07703_));
 NAND4_X1 _32777_ (.A1(_07678_),
    .A2(_07685_),
    .A3(_07698_),
    .A4(_07703_),
    .ZN(_07704_));
 OAI21_X1 _32778_ (.A(_05350_),
    .B1(_05297_),
    .B2(_05517_),
    .ZN(_07705_));
 AND3_X1 _32779_ (.A1(_05543_),
    .A2(_05351_),
    .A3(_07705_),
    .ZN(_07706_));
 OAI21_X1 _32780_ (.A(_06548_),
    .B1(_05353_),
    .B2(_05356_),
    .ZN(_07707_));
 OAI21_X1 _32781_ (.A(_05333_),
    .B1(_05497_),
    .B2(_05345_),
    .ZN(_07709_));
 AND4_X1 _32782_ (.A1(_05462_),
    .A2(_07706_),
    .A3(_07707_),
    .A4(_07709_),
    .ZN(_07710_));
 OAI211_X2 _32783_ (.A(_06531_),
    .B(_06520_),
    .C1(_05246_),
    .C2(_06522_),
    .ZN(_07711_));
 OAI21_X1 _32784_ (.A(_07711_),
    .B1(_07395_),
    .B2(_05320_),
    .ZN(_07712_));
 NAND2_X4 _32785_ (.A1(_06531_),
    .A2(_05383_),
    .ZN(_07713_));
 NAND3_X1 _32786_ (.A1(_05474_),
    .A2(_05308_),
    .A3(_07713_),
    .ZN(_07714_));
 AOI21_X1 _32787_ (.A(_05327_),
    .B1(_06528_),
    .B2(_05463_),
    .ZN(_07715_));
 NOR4_X1 _32788_ (.A1(_07712_),
    .A2(_07714_),
    .A3(_07715_),
    .A4(_06893_),
    .ZN(_07716_));
 AOI22_X1 _32789_ (.A1(_06481_),
    .A2(_05396_),
    .B1(_05360_),
    .B2(_05419_),
    .ZN(_07717_));
 OAI21_X1 _32790_ (.A(_05444_),
    .B1(_05450_),
    .B2(_05360_),
    .ZN(_07718_));
 OAI21_X1 _32791_ (.A(_05419_),
    .B1(_05473_),
    .B2(_05378_),
    .ZN(_07720_));
 AND4_X1 _32792_ (.A1(_06466_),
    .A2(_07717_),
    .A3(_07718_),
    .A4(_07720_),
    .ZN(_07721_));
 OAI21_X1 _32793_ (.A(_05496_),
    .B1(_05353_),
    .B2(_05307_),
    .ZN(_07722_));
 NAND4_X1 _32794_ (.A1(_07722_),
    .A2(_05425_),
    .A3(_05426_),
    .A4(_07399_),
    .ZN(_07723_));
 AOI21_X1 _32795_ (.A(_05431_),
    .B1(_07679_),
    .B2(_05514_),
    .ZN(_07724_));
 AND2_X1 _32796_ (.A1(_05498_),
    .A2(_05318_),
    .ZN(_07725_));
 AND3_X1 _32797_ (.A1(_05290_),
    .A2(_05273_),
    .A3(_05498_),
    .ZN(_07726_));
 NOR4_X1 _32798_ (.A1(_07723_),
    .A2(_07724_),
    .A3(_07725_),
    .A4(_07726_),
    .ZN(_07727_));
 NAND4_X1 _32799_ (.A1(_07710_),
    .A2(_07716_),
    .A3(_07721_),
    .A4(_07727_),
    .ZN(_07728_));
 NOR2_X4 _32800_ (.A1(_07704_),
    .A2(_07728_),
    .ZN(_07729_));
 XOR2_X2 _32801_ (.A(_07668_),
    .B(_07729_),
    .Z(_07731_));
 XNOR2_X1 _32802_ (.A(_07731_),
    .B(_00993_),
    .ZN(_07732_));
 XOR2_X1 _32803_ (.A(_05570_),
    .B(_07457_),
    .Z(_07733_));
 XNOR2_X1 _32804_ (.A(_07732_),
    .B(_07733_),
    .ZN(_07734_));
 XNOR2_X1 _32805_ (.A(_07601_),
    .B(_07734_),
    .ZN(_07735_));
 MUX2_X1 _32806_ (.A(_07462_),
    .B(_07735_),
    .S(_05156_),
    .Z(_00704_));
 XOR2_X1 _32807_ (.A(_17203_),
    .B(_17014_),
    .Z(_07736_));
 AND3_X1 _32808_ (.A1(_05683_),
    .A2(_05805_),
    .A3(_05589_),
    .ZN(_07737_));
 NAND2_X1 _32809_ (.A1(_06361_),
    .A2(_06348_),
    .ZN(_07738_));
 OAI21_X1 _32810_ (.A(_05656_),
    .B1(_07738_),
    .B2(_05796_),
    .ZN(_07739_));
 OAI211_X2 _32811_ (.A(_07739_),
    .B(_07612_),
    .C1(_07350_),
    .C2(_05681_),
    .ZN(_07741_));
 OAI211_X2 _32812_ (.A(_06346_),
    .B(_06849_),
    .C1(_05626_),
    .C2(_05723_),
    .ZN(_07742_));
 OR4_X1 _32813_ (.A1(_07737_),
    .A2(_07741_),
    .A3(_07347_),
    .A4(_07742_),
    .ZN(_07743_));
 AND2_X1 _32814_ (.A1(_06824_),
    .A2(_05683_),
    .ZN(_07744_));
 AOI22_X1 _32815_ (.A1(_05751_),
    .A2(_06844_),
    .B1(_06437_),
    .B2(_05661_),
    .ZN(_07745_));
 OAI221_X1 _32816_ (.A(_07745_),
    .B1(_06449_),
    .B2(_05681_),
    .C1(_07606_),
    .C2(_05743_),
    .ZN(_07746_));
 OAI22_X1 _32817_ (.A1(_06806_),
    .A2(_06795_),
    .B1(_07622_),
    .B2(_06349_),
    .ZN(_07747_));
 OR4_X1 _32818_ (.A1(_07744_),
    .A2(_07746_),
    .A3(_07630_),
    .A4(_07747_),
    .ZN(_07748_));
 NAND2_X1 _32819_ (.A1(_06437_),
    .A2(_05646_),
    .ZN(_07749_));
 NAND3_X1 _32820_ (.A1(_05729_),
    .A2(_05652_),
    .A3(_05736_),
    .ZN(_07750_));
 NOR2_X1 _32821_ (.A1(_05749_),
    .A2(_05673_),
    .ZN(_07752_));
 INV_X1 _32822_ (.A(_07752_),
    .ZN(_07753_));
 OAI211_X2 _32823_ (.A(_07749_),
    .B(_07750_),
    .C1(_07753_),
    .C2(_06360_),
    .ZN(_07754_));
 AND2_X1 _32824_ (.A1(_05656_),
    .A2(_05763_),
    .ZN(_07755_));
 AOI221_X1 _32825_ (.A(_07755_),
    .B1(_05719_),
    .B2(_06381_),
    .C1(_05763_),
    .C2(_06455_),
    .ZN(_07756_));
 NAND2_X1 _32826_ (.A1(_05815_),
    .A2(_07374_),
    .ZN(_07757_));
 AOI22_X1 _32827_ (.A1(_06403_),
    .A2(_05755_),
    .B1(_05788_),
    .B2(_06381_),
    .ZN(_07758_));
 NAND4_X1 _32828_ (.A1(_07756_),
    .A2(_07621_),
    .A3(_07757_),
    .A4(_07758_),
    .ZN(_07759_));
 NOR4_X1 _32829_ (.A1(_07743_),
    .A2(_07748_),
    .A3(_07754_),
    .A4(_07759_),
    .ZN(_07760_));
 NAND4_X1 _32830_ (.A1(_06390_),
    .A2(_05745_),
    .A3(_05677_),
    .A4(_05735_),
    .ZN(_07761_));
 NAND4_X1 _32831_ (.A1(_05736_),
    .A2(_05738_),
    .A3(_05673_),
    .A4(_05677_),
    .ZN(_07763_));
 OAI211_X2 _32832_ (.A(_07761_),
    .B(_07763_),
    .C1(_05680_),
    .C2(_06417_),
    .ZN(_07764_));
 AOI221_X4 _32833_ (.A(_07764_),
    .B1(_05623_),
    .B2(_05758_),
    .C1(_05576_),
    .C2(_05604_),
    .ZN(_07765_));
 OAI21_X1 _32834_ (.A(_06442_),
    .B1(_07738_),
    .B2(_05593_),
    .ZN(_07766_));
 OAI21_X1 _32835_ (.A(_06383_),
    .B1(_05719_),
    .B2(_05611_),
    .ZN(_07767_));
 OAI21_X1 _32836_ (.A(_06383_),
    .B1(_06844_),
    .B2(_06824_),
    .ZN(_07768_));
 AND3_X1 _32837_ (.A1(_07767_),
    .A2(_07768_),
    .A3(_05648_),
    .ZN(_07769_));
 OR2_X1 _32838_ (.A1(_05796_),
    .A2(_06844_),
    .ZN(_07770_));
 NAND2_X2 _32839_ (.A1(_06361_),
    .A2(_05680_),
    .ZN(_07771_));
 OAI21_X1 _32840_ (.A(_05699_),
    .B1(_07770_),
    .B2(_07771_),
    .ZN(_07772_));
 NAND4_X1 _32841_ (.A1(_07765_),
    .A2(_07766_),
    .A3(_07769_),
    .A4(_07772_),
    .ZN(_07774_));
 AND2_X1 _32842_ (.A1(_07771_),
    .A2(_05741_),
    .ZN(_07775_));
 AND4_X1 _32843_ (.A1(_05818_),
    .A2(_06371_),
    .A3(_06373_),
    .A4(_05827_),
    .ZN(_07776_));
 AND4_X1 _32844_ (.A1(_05807_),
    .A2(_06373_),
    .A3(_05817_),
    .A4(_05827_),
    .ZN(_07777_));
 NOR3_X1 _32845_ (.A1(_07775_),
    .A2(_07776_),
    .A3(_07777_),
    .ZN(_07778_));
 OAI21_X1 _32846_ (.A(_06451_),
    .B1(_05796_),
    .B2(_07360_),
    .ZN(_07779_));
 OAI21_X1 _32847_ (.A(_06451_),
    .B1(_05685_),
    .B2(_05646_),
    .ZN(_07780_));
 NAND4_X1 _32848_ (.A1(_06451_),
    .A2(_06371_),
    .A3(_05694_),
    .A4(_05592_),
    .ZN(_07781_));
 AND3_X1 _32849_ (.A1(_07779_),
    .A2(_07780_),
    .A3(_07781_),
    .ZN(_07782_));
 AND2_X1 _32850_ (.A1(_05661_),
    .A2(_06353_),
    .ZN(_07783_));
 INV_X1 _32851_ (.A(_07783_),
    .ZN(_07785_));
 OAI21_X1 _32852_ (.A(_06353_),
    .B1(_06456_),
    .B2(_05729_),
    .ZN(_07786_));
 NAND4_X1 _32853_ (.A1(_05807_),
    .A2(_05817_),
    .A3(_05652_),
    .A4(_05675_),
    .ZN(_07787_));
 AND3_X1 _32854_ (.A1(_07785_),
    .A2(_07786_),
    .A3(_07787_),
    .ZN(_07788_));
 AND2_X1 _32855_ (.A1(_06824_),
    .A2(_05708_),
    .ZN(_07789_));
 AND3_X1 _32856_ (.A1(_05800_),
    .A2(_05675_),
    .A3(_05624_),
    .ZN(_07790_));
 AND4_X1 _32857_ (.A1(_05603_),
    .A2(_05624_),
    .A3(_05672_),
    .A4(_05675_),
    .ZN(_07791_));
 NOR4_X1 _32858_ (.A1(_05829_),
    .A2(_07789_),
    .A3(_07790_),
    .A4(_07791_),
    .ZN(_07792_));
 NAND4_X1 _32859_ (.A1(_07778_),
    .A2(_07782_),
    .A3(_07788_),
    .A4(_07792_),
    .ZN(_07793_));
 AND2_X1 _32860_ (.A1(_05755_),
    .A2(_06387_),
    .ZN(_07794_));
 OR4_X1 _32861_ (.A1(_05747_),
    .A2(_07794_),
    .A3(_07613_),
    .A4(_07608_),
    .ZN(_07796_));
 AND4_X1 _32862_ (.A1(_05807_),
    .A2(_05735_),
    .A3(_05589_),
    .A4(_05624_),
    .ZN(_07797_));
 AOI221_X4 _32863_ (.A(_07797_),
    .B1(_05771_),
    .B2(_05646_),
    .C1(_06406_),
    .C2(_05603_),
    .ZN(_07798_));
 OAI22_X1 _32864_ (.A1(_05748_),
    .A2(_05590_),
    .B1(_05578_),
    .B2(_05728_),
    .ZN(_07799_));
 OAI21_X1 _32865_ (.A(_06437_),
    .B1(_07799_),
    .B2(_05685_),
    .ZN(_07800_));
 OAI21_X1 _32866_ (.A(_06455_),
    .B1(_05759_),
    .B2(_06384_),
    .ZN(_07801_));
 OAI21_X1 _32867_ (.A(_05771_),
    .B1(_06824_),
    .B2(_06456_),
    .ZN(_07802_));
 NAND4_X1 _32868_ (.A1(_07798_),
    .A2(_07800_),
    .A3(_07801_),
    .A4(_07802_),
    .ZN(_07803_));
 NOR4_X1 _32869_ (.A1(_07774_),
    .A2(_07793_),
    .A3(_07796_),
    .A4(_07803_),
    .ZN(_07804_));
 AND2_X2 _32870_ (.A1(_07760_),
    .A2(_07804_),
    .ZN(_07805_));
 NAND3_X1 _32871_ (.A1(_05277_),
    .A2(_07427_),
    .A3(_05550_),
    .ZN(_07807_));
 OAI21_X1 _32872_ (.A(_05564_),
    .B1(_07807_),
    .B2(_05240_),
    .ZN(_07808_));
 AOI211_X4 _32873_ (.A(_06491_),
    .B(_07450_),
    .C1(_05310_),
    .C2(_06522_),
    .ZN(_07809_));
 AOI21_X1 _32874_ (.A(_07450_),
    .B1(_05504_),
    .B2(_06539_),
    .ZN(_07810_));
 NOR3_X1 _32875_ (.A1(_07809_),
    .A2(_07453_),
    .A3(_07810_),
    .ZN(_07811_));
 OAI21_X1 _32876_ (.A(_05444_),
    .B1(_05460_),
    .B2(_05290_),
    .ZN(_07812_));
 OAI21_X1 _32877_ (.A(_06548_),
    .B1(_05349_),
    .B2(_05383_),
    .ZN(_07813_));
 OAI21_X1 _32878_ (.A(_06548_),
    .B1(_05371_),
    .B2(_05373_),
    .ZN(_07814_));
 AND2_X1 _32879_ (.A1(_07813_),
    .A2(_07814_),
    .ZN(_07815_));
 AND4_X1 _32880_ (.A1(_07808_),
    .A2(_07811_),
    .A3(_07812_),
    .A4(_07815_),
    .ZN(_07816_));
 OAI21_X1 _32881_ (.A(_05270_),
    .B1(_06473_),
    .B2(_05360_),
    .ZN(_07818_));
 NAND2_X1 _32882_ (.A1(_05493_),
    .A2(_05498_),
    .ZN(_07819_));
 NAND2_X1 _32883_ (.A1(_05375_),
    .A2(_05353_),
    .ZN(_07820_));
 NAND2_X1 _32884_ (.A1(_06929_),
    .A2(_05270_),
    .ZN(_07821_));
 AND4_X1 _32885_ (.A1(_07819_),
    .A2(_05474_),
    .A3(_07820_),
    .A4(_07821_),
    .ZN(_07822_));
 OAI21_X1 _32886_ (.A(_05496_),
    .B1(_05307_),
    .B2(_05383_),
    .ZN(_07823_));
 OAI21_X1 _32887_ (.A(_05496_),
    .B1(_05360_),
    .B2(_06541_),
    .ZN(_07824_));
 NAND4_X1 _32888_ (.A1(_06514_),
    .A2(_05283_),
    .A3(_05232_),
    .A4(_05441_),
    .ZN(_07825_));
 AND3_X1 _32889_ (.A1(_07823_),
    .A2(_07824_),
    .A3(_07825_),
    .ZN(_07826_));
 AND4_X1 _32890_ (.A1(_05377_),
    .A2(_07818_),
    .A3(_07822_),
    .A4(_07826_),
    .ZN(_07827_));
 NOR2_X1 _32891_ (.A1(_06480_),
    .A2(_06485_),
    .ZN(_07829_));
 OAI21_X1 _32892_ (.A(_05354_),
    .B1(_05341_),
    .B2(_05507_),
    .ZN(_07830_));
 AND4_X1 _32893_ (.A1(_05538_),
    .A2(_05455_),
    .A3(_07830_),
    .A4(_05355_),
    .ZN(_07831_));
 NAND3_X1 _32894_ (.A1(_05413_),
    .A2(_05237_),
    .A3(_05240_),
    .ZN(_07832_));
 NAND3_X1 _32895_ (.A1(_05356_),
    .A2(_05265_),
    .A3(_05303_),
    .ZN(_07833_));
 AND3_X1 _32896_ (.A1(_07832_),
    .A2(_06937_),
    .A3(_07833_),
    .ZN(_07834_));
 AND4_X1 _32897_ (.A1(_07829_),
    .A2(_07831_),
    .A3(_06939_),
    .A4(_07834_),
    .ZN(_07835_));
 OAI21_X1 _32898_ (.A(_07442_),
    .B1(_05482_),
    .B2(_05338_),
    .ZN(_07836_));
 AOI221_X1 _32899_ (.A(_07836_),
    .B1(_05307_),
    .B2(_06928_),
    .C1(_05493_),
    .C2(_05354_),
    .ZN(_07837_));
 AOI22_X1 _32900_ (.A1(_05521_),
    .A2(_05354_),
    .B1(_06541_),
    .B2(_06488_),
    .ZN(_07838_));
 AND4_X1 _32901_ (.A1(_07688_),
    .A2(_07837_),
    .A3(_07689_),
    .A4(_07838_),
    .ZN(_07840_));
 NAND4_X1 _32902_ (.A1(_07816_),
    .A2(_07827_),
    .A3(_07835_),
    .A4(_07840_),
    .ZN(_07841_));
 AND2_X1 _32903_ (.A1(_05498_),
    .A2(_05517_),
    .ZN(_07842_));
 OR4_X2 _32904_ (.A1(_05531_),
    .A2(_07671_),
    .A3(_05436_),
    .A4(_07842_),
    .ZN(_07843_));
 OAI21_X1 _32905_ (.A(_06503_),
    .B1(_05360_),
    .B2(_05507_),
    .ZN(_07844_));
 NAND3_X1 _32906_ (.A1(_07844_),
    .A2(_07713_),
    .A3(_07423_),
    .ZN(_07845_));
 OAI221_X1 _32907_ (.A(_05312_),
    .B1(_07395_),
    .B2(_05235_),
    .C1(_05406_),
    .C2(_05347_),
    .ZN(_07846_));
 NOR4_X1 _32908_ (.A1(_07843_),
    .A2(_05503_),
    .A3(_07845_),
    .A4(_07846_),
    .ZN(_07847_));
 OAI21_X1 _32909_ (.A(_06928_),
    .B1(_05373_),
    .B2(_05517_),
    .ZN(_07848_));
 AND2_X1 _32910_ (.A1(_05444_),
    .A2(_05378_),
    .ZN(_07849_));
 AOI21_X1 _32911_ (.A(_07849_),
    .B1(_05498_),
    .B2(_06929_),
    .ZN(_07851_));
 AOI21_X1 _32912_ (.A(_07695_),
    .B1(_05473_),
    .B2(_05413_),
    .ZN(_07852_));
 OAI21_X1 _32913_ (.A(_05392_),
    .B1(_05381_),
    .B2(_05307_),
    .ZN(_07853_));
 AND4_X1 _32914_ (.A1(_07848_),
    .A2(_07851_),
    .A3(_07852_),
    .A4(_07853_),
    .ZN(_07854_));
 AOI21_X1 _32915_ (.A(_05527_),
    .B1(_05480_),
    .B2(_05419_),
    .ZN(_07855_));
 OAI21_X1 _32916_ (.A(_06504_),
    .B1(_06503_),
    .B2(_06488_),
    .ZN(_07856_));
 AND3_X1 _32917_ (.A1(_07856_),
    .A2(_05389_),
    .A3(_05388_),
    .ZN(_07857_));
 NAND4_X1 _32918_ (.A1(_07847_),
    .A2(_07854_),
    .A3(_07855_),
    .A4(_07857_),
    .ZN(_07858_));
 NOR2_X2 _32919_ (.A1(_07841_),
    .A2(_07858_),
    .ZN(_07859_));
 XNOR2_X1 _32920_ (.A(_07805_),
    .B(_07859_),
    .ZN(_07860_));
 AND2_X1 _32921_ (.A1(_05991_),
    .A2(_05988_),
    .ZN(_07862_));
 AND3_X1 _32922_ (.A1(_05988_),
    .A2(_06063_),
    .A3(_05893_),
    .ZN(_07863_));
 NOR2_X1 _32923_ (.A1(_07862_),
    .A2(_07863_),
    .ZN(_07864_));
 OAI21_X1 _32924_ (.A(_07589_),
    .B1(_05965_),
    .B2(_06081_),
    .ZN(_07865_));
 AND2_X1 _32925_ (.A1(_05961_),
    .A2(_05936_),
    .ZN(_07866_));
 NOR4_X1 _32926_ (.A1(_07865_),
    .A2(_06019_),
    .A3(_07176_),
    .A4(_07866_),
    .ZN(_07867_));
 OAI21_X1 _32927_ (.A(_05942_),
    .B1(_06686_),
    .B2(_05939_),
    .ZN(_07868_));
 AND2_X1 _32928_ (.A1(_05865_),
    .A2(_05992_),
    .ZN(_07869_));
 AND2_X1 _32929_ (.A1(_05967_),
    .A2(_06002_),
    .ZN(_07870_));
 NOR4_X1 _32930_ (.A1(_07868_),
    .A2(_06740_),
    .A3(_07869_),
    .A4(_07870_),
    .ZN(_07871_));
 AOI221_X4 _32931_ (.A(_07159_),
    .B1(_06016_),
    .B2(_05992_),
    .C1(_05860_),
    .C2(_06054_),
    .ZN(_07873_));
 AND4_X1 _32932_ (.A1(_07864_),
    .A2(_07867_),
    .A3(_07871_),
    .A4(_07873_),
    .ZN(_07874_));
 INV_X1 _32933_ (.A(_05855_),
    .ZN(_07875_));
 OAI22_X1 _32934_ (.A1(_06703_),
    .A2(_07875_),
    .B1(_05944_),
    .B2(_06007_),
    .ZN(_07876_));
 AOI221_X1 _32935_ (.A(_07876_),
    .B1(_05964_),
    .B2(_05971_),
    .C1(_05961_),
    .C2(_05882_),
    .ZN(_07877_));
 NAND2_X1 _32936_ (.A1(_06029_),
    .A2(_06043_),
    .ZN(_07878_));
 AND2_X1 _32937_ (.A1(_05972_),
    .A2(_05860_),
    .ZN(_07879_));
 NOR4_X1 _32938_ (.A1(_07879_),
    .A2(_05866_),
    .A3(_06715_),
    .A4(_06725_),
    .ZN(_07880_));
 AND4_X1 _32939_ (.A1(_05905_),
    .A2(_07877_),
    .A3(_07878_),
    .A4(_07880_),
    .ZN(_07881_));
 OAI21_X1 _32940_ (.A(_05972_),
    .B1(_07133_),
    .B2(_05928_),
    .ZN(_07882_));
 OAI221_X1 _32941_ (.A(_07882_),
    .B1(_06959_),
    .B2(_06695_),
    .C1(_05979_),
    .C2(_07162_),
    .ZN(_07884_));
 NAND2_X1 _32942_ (.A1(_06024_),
    .A2(_05985_),
    .ZN(_07885_));
 OAI211_X2 _32943_ (.A(_07548_),
    .B(_07885_),
    .C1(_06718_),
    .C2(_05946_),
    .ZN(_07886_));
 NAND4_X1 _32944_ (.A1(_06970_),
    .A2(_06757_),
    .A3(_06966_),
    .A4(_07015_),
    .ZN(_07887_));
 NOR4_X1 _32945_ (.A1(_07884_),
    .A2(_07142_),
    .A3(_07886_),
    .A4(_07887_),
    .ZN(_07888_));
 AOI22_X1 _32946_ (.A1(_07552_),
    .A2(_05871_),
    .B1(_05992_),
    .B2(_05898_),
    .ZN(_07889_));
 NAND2_X1 _32947_ (.A1(_05844_),
    .A2(_06033_),
    .ZN(_07890_));
 AOI22_X1 _32948_ (.A1(_06024_),
    .A2(_05912_),
    .B1(_05873_),
    .B2(_06002_),
    .ZN(_07891_));
 AND4_X1 _32949_ (.A1(_07009_),
    .A2(_07889_),
    .A3(_07890_),
    .A4(_07891_),
    .ZN(_07892_));
 AND4_X1 _32950_ (.A1(_07874_),
    .A2(_07881_),
    .A3(_07888_),
    .A4(_07892_),
    .ZN(_07893_));
 AND2_X1 _32951_ (.A1(_06680_),
    .A2(_05882_),
    .ZN(_07895_));
 OR2_X1 _32952_ (.A1(_06950_),
    .A2(_07895_),
    .ZN(_07896_));
 INV_X1 _32953_ (.A(_07185_),
    .ZN(_07897_));
 AOI21_X1 _32954_ (.A(_05946_),
    .B1(_05978_),
    .B2(_07897_),
    .ZN(_07898_));
 AOI21_X1 _32955_ (.A(_06090_),
    .B1(_06748_),
    .B2(_05944_),
    .ZN(_07899_));
 NOR3_X1 _32956_ (.A1(_07896_),
    .A2(_07898_),
    .A3(_07899_),
    .ZN(_07900_));
 INV_X1 _32957_ (.A(_06053_),
    .ZN(_07901_));
 OAI21_X1 _32958_ (.A(_05976_),
    .B1(_05889_),
    .B2(_06037_),
    .ZN(_07902_));
 NAND2_X1 _32959_ (.A1(_07902_),
    .A2(_05926_),
    .ZN(_07903_));
 NAND4_X1 _32960_ (.A1(_07900_),
    .A2(_07566_),
    .A3(_07901_),
    .A4(_07903_),
    .ZN(_07904_));
 AOI22_X1 _32961_ (.A1(_05981_),
    .A2(_06946_),
    .B1(_06692_),
    .B2(_05914_),
    .ZN(_07906_));
 OAI21_X1 _32962_ (.A(_06946_),
    .B1(_07193_),
    .B2(_05956_),
    .ZN(_07907_));
 NAND3_X1 _32963_ (.A1(_07906_),
    .A2(_06958_),
    .A3(_07907_),
    .ZN(_07908_));
 AOI22_X1 _32964_ (.A1(_06024_),
    .A2(_06022_),
    .B1(_06033_),
    .B2(_05912_),
    .ZN(_07909_));
 OAI21_X1 _32965_ (.A(_06033_),
    .B1(_05934_),
    .B2(_05967_),
    .ZN(_07910_));
 OAI211_X2 _32966_ (.A(_07909_),
    .B(_07910_),
    .C1(_06090_),
    .C2(_06091_),
    .ZN(_07911_));
 OAI21_X1 _32967_ (.A(_06055_),
    .B1(_06690_),
    .B2(_05958_),
    .ZN(_07912_));
 OAI21_X1 _32968_ (.A(_05908_),
    .B1(_07902_),
    .B2(_05860_),
    .ZN(_07913_));
 INV_X1 _32969_ (.A(_06042_),
    .ZN(_07914_));
 AND2_X1 _32970_ (.A1(_05936_),
    .A2(_07193_),
    .ZN(_07915_));
 INV_X1 _32971_ (.A(_07915_),
    .ZN(_07917_));
 NAND4_X1 _32972_ (.A1(_07912_),
    .A2(_07913_),
    .A3(_07914_),
    .A4(_07917_),
    .ZN(_07918_));
 NOR4_X1 _32973_ (.A1(_07904_),
    .A2(_07908_),
    .A3(_07911_),
    .A4(_07918_),
    .ZN(_07919_));
 NAND2_X2 _32974_ (.A1(_07893_),
    .A2(_07919_),
    .ZN(_07920_));
 XNOR2_X1 _32975_ (.A(_07920_),
    .B(_00994_),
    .ZN(_07921_));
 XOR2_X1 _32976_ (.A(_07860_),
    .B(_07921_),
    .Z(_07922_));
 NAND2_X1 _32977_ (.A1(_07076_),
    .A2(_07258_),
    .ZN(_07923_));
 AOI211_X4 _32978_ (.A(_07478_),
    .B(_07075_),
    .C1(_06142_),
    .C2(_06309_),
    .ZN(_07924_));
 OAI21_X1 _32979_ (.A(_06301_),
    .B1(_06201_),
    .B2(_06642_),
    .ZN(_07925_));
 NAND4_X1 _32980_ (.A1(_06203_),
    .A2(_06298_),
    .A3(_06594_),
    .A4(_06294_),
    .ZN(_07926_));
 AND4_X1 _32981_ (.A1(_07923_),
    .A2(_07924_),
    .A3(_07925_),
    .A4(_07926_),
    .ZN(_07928_));
 AOI211_X4 _32982_ (.A(_07494_),
    .B(_07246_),
    .C1(_07044_),
    .C2(_06274_),
    .ZN(_07929_));
 AND2_X1 _32983_ (.A1(_06572_),
    .A2(_06331_),
    .ZN(_07930_));
 NOR3_X1 _32984_ (.A1(_06282_),
    .A2(_06279_),
    .A3(_07930_),
    .ZN(_07931_));
 OAI211_X2 _32985_ (.A(_06572_),
    .B(_06594_),
    .C1(_06205_),
    .C2(_06294_),
    .ZN(_07932_));
 AND4_X1 _32986_ (.A1(_07502_),
    .A2(_07929_),
    .A3(_07931_),
    .A4(_07932_),
    .ZN(_07933_));
 OAI21_X1 _32987_ (.A(_07222_),
    .B1(_06657_),
    .B2(_06603_),
    .ZN(_07934_));
 OAI211_X2 _32988_ (.A(_06257_),
    .B(_16879_),
    .C1(_16878_),
    .C2(_06120_),
    .ZN(_07935_));
 OAI21_X1 _32989_ (.A(_07222_),
    .B1(_06147_),
    .B2(_06220_),
    .ZN(_07936_));
 AND4_X1 _32990_ (.A1(_06577_),
    .A2(_07934_),
    .A3(_07935_),
    .A4(_07936_),
    .ZN(_07937_));
 OAI21_X1 _32991_ (.A(_06326_),
    .B1(_06173_),
    .B2(_06218_),
    .ZN(_07939_));
 NAND4_X1 _32992_ (.A1(_07939_),
    .A2(_06593_),
    .A3(_06595_),
    .A4(_07463_),
    .ZN(_07940_));
 AOI21_X1 _32993_ (.A(_07057_),
    .B1(_06620_),
    .B2(_07048_),
    .ZN(_07941_));
 AND2_X1 _32994_ (.A1(_06212_),
    .A2(_06330_),
    .ZN(_07942_));
 NOR4_X1 _32995_ (.A1(_07940_),
    .A2(_07941_),
    .A3(_07942_),
    .A4(_07469_),
    .ZN(_07943_));
 NAND4_X1 _32996_ (.A1(_07928_),
    .A2(_07933_),
    .A3(_07937_),
    .A4(_07943_),
    .ZN(_07944_));
 OAI21_X1 _32997_ (.A(_06635_),
    .B1(_06121_),
    .B2(_06258_),
    .ZN(_07945_));
 AND2_X1 _32998_ (.A1(_06169_),
    .A2(_06310_),
    .ZN(_07946_));
 AND3_X1 _32999_ (.A1(_06113_),
    .A2(_06203_),
    .A3(_06167_),
    .ZN(_07947_));
 AOI211_X4 _33000_ (.A(_07946_),
    .B(_07947_),
    .C1(_06156_),
    .C2(_06635_),
    .ZN(_07948_));
 OAI21_X1 _33001_ (.A(_06189_),
    .B1(_06164_),
    .B2(_06603_),
    .ZN(_07950_));
 AOI22_X1 _33002_ (.A1(_07038_),
    .A2(_07258_),
    .B1(_06189_),
    .B2(_06610_),
    .ZN(_07951_));
 AND4_X1 _33003_ (.A1(_07945_),
    .A2(_07948_),
    .A3(_07950_),
    .A4(_07951_),
    .ZN(_07952_));
 OAI211_X2 _33004_ (.A(_06658_),
    .B(_16879_),
    .C1(_16878_),
    .C2(_06211_),
    .ZN(_07953_));
 NAND2_X1 _33005_ (.A1(_06667_),
    .A2(_06304_),
    .ZN(_07954_));
 INV_X1 _33006_ (.A(_06230_),
    .ZN(_07955_));
 OAI21_X1 _33007_ (.A(_07954_),
    .B1(_06115_),
    .B2(_07955_),
    .ZN(_07956_));
 NOR3_X1 _33008_ (.A1(_07956_),
    .A2(_07514_),
    .A3(_07279_),
    .ZN(_07957_));
 AND2_X1 _33009_ (.A1(_06228_),
    .A2(_06658_),
    .ZN(_07958_));
 NOR3_X1 _33010_ (.A1(_06157_),
    .A2(_07958_),
    .A3(_06662_),
    .ZN(_07959_));
 OAI21_X1 _33011_ (.A(_06667_),
    .B1(_06313_),
    .B2(_06201_),
    .ZN(_07961_));
 AND4_X1 _33012_ (.A1(_07953_),
    .A2(_07957_),
    .A3(_07959_),
    .A4(_07961_),
    .ZN(_07962_));
 NAND2_X1 _33013_ (.A1(_06641_),
    .A2(_06331_),
    .ZN(_07963_));
 INV_X1 _33014_ (.A(_06198_),
    .ZN(_07964_));
 OAI211_X2 _33015_ (.A(_07963_),
    .B(_06651_),
    .C1(_07964_),
    .C2(_06620_),
    .ZN(_07965_));
 OAI21_X1 _33016_ (.A(_07523_),
    .B1(_07964_),
    .B2(_07097_),
    .ZN(_07966_));
 INV_X1 _33017_ (.A(_07044_),
    .ZN(_07967_));
 AOI21_X1 _33018_ (.A(_07082_),
    .B1(_07967_),
    .B2(_06311_),
    .ZN(_07968_));
 NOR4_X1 _33019_ (.A1(_07965_),
    .A2(_07966_),
    .A3(_07968_),
    .A4(_07086_),
    .ZN(_07969_));
 AND2_X4 _33020_ (.A1(_06627_),
    .A2(_06304_),
    .ZN(_07970_));
 AOI211_X4 _33021_ (.A(_07970_),
    .B(_06231_),
    .C1(_06605_),
    .C2(_06627_),
    .ZN(_07972_));
 AND2_X1 _33022_ (.A1(_06121_),
    .A2(_06235_),
    .ZN(_07973_));
 AOI211_X4 _33023_ (.A(_06612_),
    .B(_07973_),
    .C1(_06185_),
    .C2(_06236_),
    .ZN(_07974_));
 NAND3_X1 _33024_ (.A1(_06668_),
    .A2(_06627_),
    .A3(_06186_),
    .ZN(_07975_));
 OAI211_X2 _33025_ (.A(_06627_),
    .B(_06211_),
    .C1(_06206_),
    .C2(_06289_),
    .ZN(_07976_));
 AND4_X4 _33026_ (.A1(_07972_),
    .A2(_07974_),
    .A3(_07975_),
    .A4(_07976_),
    .ZN(_07977_));
 NAND4_X1 _33027_ (.A1(_07952_),
    .A2(_07962_),
    .A3(_07969_),
    .A4(_07977_),
    .ZN(_07978_));
 NOR2_X2 _33028_ (.A1(_07944_),
    .A2(_07978_),
    .ZN(_07979_));
 XOR2_X1 _33029_ (.A(_07979_),
    .B(_07729_),
    .Z(_07980_));
 XNOR2_X1 _33030_ (.A(_07922_),
    .B(_07980_),
    .ZN(_07981_));
 MUX2_X1 _33031_ (.A(_07736_),
    .B(_07981_),
    .S(_05156_),
    .Z(_00705_));
 XOR2_X1 _33032_ (.A(_17204_),
    .B(_17015_),
    .Z(_07983_));
 OAI21_X1 _33033_ (.A(_05270_),
    .B1(_05341_),
    .B2(_05399_),
    .ZN(_07984_));
 OAI21_X1 _33034_ (.A(_05270_),
    .B1(_05541_),
    .B2(_06541_),
    .ZN(_07985_));
 NAND3_X1 _33035_ (.A1(_07984_),
    .A2(_07432_),
    .A3(_07985_),
    .ZN(_07986_));
 AOI22_X1 _33036_ (.A1(_05211_),
    .A2(_05439_),
    .B1(_05373_),
    .B2(_06928_),
    .ZN(_07987_));
 OAI211_X2 _33037_ (.A(_07987_),
    .B(_06546_),
    .C1(_05556_),
    .C2(_05449_),
    .ZN(_07988_));
 AOI21_X1 _33038_ (.A(_05364_),
    .B1(_07679_),
    .B2(_05483_),
    .ZN(_07989_));
 AOI211_X2 _33039_ (.A(_05208_),
    .B(_05364_),
    .C1(_07427_),
    .C2(_05347_),
    .ZN(_07990_));
 NOR3_X4 _33040_ (.A1(_05493_),
    .A2(_05521_),
    .A3(_05352_),
    .ZN(_07991_));
 NOR2_X1 _33041_ (.A1(_07991_),
    .A2(_05327_),
    .ZN(_07993_));
 OAI211_X2 _33042_ (.A(_05439_),
    .B(_05446_),
    .C1(_05219_),
    .C2(_05228_),
    .ZN(_07994_));
 NAND4_X1 _33043_ (.A1(_05265_),
    .A2(_05417_),
    .A3(_05272_),
    .A4(_05252_),
    .ZN(_07995_));
 OAI211_X2 _33044_ (.A(_07994_),
    .B(_07995_),
    .C1(_06494_),
    .C2(_05482_),
    .ZN(_07996_));
 OR4_X4 _33045_ (.A1(_07989_),
    .A2(_07990_),
    .A3(_07993_),
    .A4(_07996_),
    .ZN(_07997_));
 NOR2_X1 _33046_ (.A1(_06507_),
    .A2(_07454_),
    .ZN(_07998_));
 NAND4_X1 _33047_ (.A1(_07998_),
    .A2(_06871_),
    .A3(_05411_),
    .A4(_06467_),
    .ZN(_07999_));
 AOI22_X1 _33048_ (.A1(_05352_),
    .A2(_05289_),
    .B1(_05333_),
    .B2(_05373_),
    .ZN(_08000_));
 AOI22_X1 _33049_ (.A1(_05337_),
    .A2(_05418_),
    .B1(_05296_),
    .B2(_05216_),
    .ZN(_08001_));
 OAI211_X2 _33050_ (.A(_08000_),
    .B(_08001_),
    .C1(_07450_),
    .C2(_05397_),
    .ZN(_08002_));
 OR4_X4 _33051_ (.A1(_07988_),
    .A2(_07997_),
    .A3(_07999_),
    .A4(_08002_),
    .ZN(_08004_));
 NAND2_X1 _33052_ (.A1(_07807_),
    .A2(_05392_),
    .ZN(_08005_));
 OAI211_X2 _33053_ (.A(_05459_),
    .B(_05463_),
    .C1(_05246_),
    .C2(_05409_),
    .ZN(_08006_));
 OAI21_X1 _33054_ (.A(_05413_),
    .B1(_08006_),
    .B2(_05378_),
    .ZN(_08007_));
 NOR4_X1 _33055_ (.A1(_05276_),
    .A2(_05383_),
    .A3(_05378_),
    .A4(_05497_),
    .ZN(_08008_));
 OAI211_X2 _33056_ (.A(_08005_),
    .B(_08007_),
    .C1(_05431_),
    .C2(_08008_),
    .ZN(_08009_));
 INV_X1 _33057_ (.A(_05217_),
    .ZN(_08010_));
 OAI21_X1 _33058_ (.A(_06503_),
    .B1(_05399_),
    .B2(_05360_),
    .ZN(_08011_));
 AND3_X1 _33059_ (.A1(_05524_),
    .A2(_08010_),
    .A3(_08011_),
    .ZN(_08012_));
 AND2_X1 _33060_ (.A1(_05314_),
    .A2(_05498_),
    .ZN(_08013_));
 AOI221_X4 _33061_ (.A(_08013_),
    .B1(_05341_),
    .B2(_05333_),
    .C1(_05439_),
    .C2(_05517_),
    .ZN(_08015_));
 NAND2_X1 _33062_ (.A1(_05419_),
    .A2(_05497_),
    .ZN(_08016_));
 NAND4_X1 _33063_ (.A1(_08012_),
    .A2(_08015_),
    .A3(_05470_),
    .A4(_08016_),
    .ZN(_08017_));
 OR4_X4 _33064_ (.A1(_07986_),
    .A2(_08004_),
    .A3(_08009_),
    .A4(_08017_),
    .ZN(_08018_));
 AOI21_X1 _33065_ (.A(_06486_),
    .B1(_05409_),
    .B2(_05241_),
    .ZN(_08019_));
 AND3_X1 _33066_ (.A1(_05447_),
    .A2(_05384_),
    .A3(_05233_),
    .ZN(_08020_));
 NAND2_X1 _33067_ (.A1(_06503_),
    .A2(_05517_),
    .ZN(_08021_));
 OAI21_X1 _33068_ (.A(_08021_),
    .B1(_05428_),
    .B2(_07395_),
    .ZN(_08022_));
 NOR4_X1 _33069_ (.A1(_06915_),
    .A2(_08019_),
    .A3(_08020_),
    .A4(_08022_),
    .ZN(_08023_));
 AND2_X1 _33070_ (.A1(_05502_),
    .A2(_05496_),
    .ZN(_08024_));
 NOR4_X1 _33071_ (.A1(_08024_),
    .A2(_07842_),
    .A3(_06880_),
    .A4(_07452_),
    .ZN(_08026_));
 OAI22_X1 _33072_ (.A1(_05554_),
    .A2(_05556_),
    .B1(_05428_),
    .B2(_05338_),
    .ZN(_08027_));
 AND2_X1 _33073_ (.A1(_06928_),
    .A2(_05407_),
    .ZN(_08028_));
 AND2_X1 _33074_ (.A1(_06548_),
    .A2(_05383_),
    .ZN(_08029_));
 NOR4_X1 _33075_ (.A1(_08027_),
    .A2(_08028_),
    .A3(_08029_),
    .A4(_05465_),
    .ZN(_08030_));
 OAI21_X1 _33076_ (.A(_06531_),
    .B1(_07426_),
    .B2(_05318_),
    .ZN(_08031_));
 NAND3_X1 _33077_ (.A1(_06531_),
    .A2(_05435_),
    .A3(_05396_),
    .ZN(_08032_));
 NAND4_X1 _33078_ (.A1(_06514_),
    .A2(_05446_),
    .A3(_05265_),
    .A4(_05303_),
    .ZN(_08033_));
 AND4_X1 _33079_ (.A1(_05455_),
    .A2(_08031_),
    .A3(_08032_),
    .A4(_08033_),
    .ZN(_08034_));
 NAND4_X1 _33080_ (.A1(_08023_),
    .A2(_08026_),
    .A3(_08030_),
    .A4(_08034_),
    .ZN(_08035_));
 NOR2_X4 _33081_ (.A1(_08018_),
    .A2(_08035_),
    .ZN(_08037_));
 AND4_X1 _33082_ (.A1(_05722_),
    .A2(_05734_),
    .A3(_05620_),
    .A4(_05651_),
    .ZN(_08038_));
 AND2_X1 _33083_ (.A1(_05741_),
    .A2(_05583_),
    .ZN(_08039_));
 AND2_X1 _33084_ (.A1(_05692_),
    .A2(_05694_),
    .ZN(_08040_));
 AOI211_X2 _33085_ (.A(_08038_),
    .B(_08039_),
    .C1(_08040_),
    .C2(_05751_),
    .ZN(_08041_));
 OAI21_X1 _33086_ (.A(_05751_),
    .B1(_06824_),
    .B2(_05800_),
    .ZN(_08042_));
 AND3_X1 _33087_ (.A1(_08041_),
    .A2(_07750_),
    .A3(_08042_),
    .ZN(_08043_));
 AOI211_X4 _33088_ (.A(_05783_),
    .B(_06806_),
    .C1(_05582_),
    .C2(_05638_),
    .ZN(_08044_));
 AOI211_X4 _33089_ (.A(_06427_),
    .B(_08044_),
    .C1(_05748_),
    .C2(_06428_),
    .ZN(_08045_));
 AOI211_X4 _33090_ (.A(_06389_),
    .B(_06417_),
    .C1(_05712_),
    .C2(_05603_),
    .ZN(_08046_));
 AND3_X1 _33091_ (.A1(_05758_),
    .A2(_05745_),
    .A3(_05784_),
    .ZN(_08048_));
 AND4_X1 _33092_ (.A1(_05603_),
    .A2(_05736_),
    .A3(_05589_),
    .A4(_05827_),
    .ZN(_08049_));
 AND4_X1 _33093_ (.A1(_05579_),
    .A2(_05736_),
    .A3(_05827_),
    .A4(_07358_),
    .ZN(_08050_));
 NOR4_X1 _33094_ (.A1(_08046_),
    .A2(_08048_),
    .A3(_08049_),
    .A4(_08050_),
    .ZN(_08051_));
 NAND2_X1 _33095_ (.A1(_05771_),
    .A2(_06456_),
    .ZN(_08052_));
 NOR2_X1 _33096_ (.A1(_05773_),
    .A2(_07311_),
    .ZN(_08053_));
 NAND2_X1 _33097_ (.A1(_05771_),
    .A2(_06387_),
    .ZN(_08054_));
 AND4_X1 _33098_ (.A1(_08052_),
    .A2(_08053_),
    .A3(_06415_),
    .A4(_08054_),
    .ZN(_08055_));
 AND4_X2 _33099_ (.A1(_08043_),
    .A2(_08045_),
    .A3(_08051_),
    .A4(_08055_),
    .ZN(_08056_));
 OAI21_X1 _33100_ (.A(_05699_),
    .B1(_05611_),
    .B2(_05613_),
    .ZN(_08057_));
 OAI21_X1 _33101_ (.A(_05699_),
    .B1(_07316_),
    .B2(_06456_),
    .ZN(_08059_));
 AND3_X1 _33102_ (.A1(_08057_),
    .A2(_08059_),
    .A3(_07353_),
    .ZN(_08060_));
 INV_X1 _33103_ (.A(_07612_),
    .ZN(_08061_));
 NOR4_X1 _33104_ (.A1(_06865_),
    .A2(_08061_),
    .A3(_07737_),
    .A4(_05688_),
    .ZN(_08062_));
 NAND2_X1 _33105_ (.A1(_05705_),
    .A2(_05612_),
    .ZN(_08063_));
 NAND2_X1 _33106_ (.A1(_05763_),
    .A2(_05708_),
    .ZN(_08064_));
 NAND2_X1 _33107_ (.A1(_08063_),
    .A2(_08064_),
    .ZN(_08065_));
 AND3_X1 _33108_ (.A1(_05729_),
    .A2(_05675_),
    .A3(_05624_),
    .ZN(_08066_));
 NOR3_X1 _33109_ (.A1(_08065_),
    .A2(_07789_),
    .A3(_08066_),
    .ZN(_08067_));
 AND2_X1 _33110_ (.A1(_05711_),
    .A2(_06353_),
    .ZN(_08068_));
 AND2_X1 _33111_ (.A1(_05716_),
    .A2(_06397_),
    .ZN(_08070_));
 NOR4_X1 _33112_ (.A1(_07783_),
    .A2(_05725_),
    .A3(_08068_),
    .A4(_08070_),
    .ZN(_08071_));
 AND4_X1 _33113_ (.A1(_08060_),
    .A2(_08062_),
    .A3(_08067_),
    .A4(_08071_),
    .ZN(_08072_));
 NAND4_X1 _33114_ (.A1(_06373_),
    .A2(_05579_),
    .A3(_05827_),
    .A4(_07358_),
    .ZN(_08073_));
 OAI21_X1 _33115_ (.A(_08073_),
    .B1(_06368_),
    .B2(_06366_),
    .ZN(_08074_));
 AOI21_X1 _33116_ (.A(_08074_),
    .B1(_08040_),
    .B2(_05576_),
    .ZN(_08075_));
 OAI21_X1 _33117_ (.A(_05625_),
    .B1(_05626_),
    .B2(_05584_),
    .ZN(_08076_));
 AND2_X1 _33118_ (.A1(_06381_),
    .A2(_05611_),
    .ZN(_08077_));
 AND4_X1 _33119_ (.A1(_05672_),
    .A2(_05624_),
    .A3(_06373_),
    .A4(_05726_),
    .ZN(_08078_));
 NOR4_X1 _33120_ (.A1(_08076_),
    .A2(_05628_),
    .A3(_08077_),
    .A4(_08078_),
    .ZN(_08079_));
 AND2_X1 _33121_ (.A1(_06384_),
    .A2(_05656_),
    .ZN(_08081_));
 AND2_X1 _33122_ (.A1(_05656_),
    .A2(_06386_),
    .ZN(_08082_));
 AND4_X1 _33123_ (.A1(_05603_),
    .A2(_06373_),
    .A3(_05817_),
    .A4(_05652_),
    .ZN(_08083_));
 NOR4_X1 _33124_ (.A1(_06396_),
    .A2(_08081_),
    .A3(_08082_),
    .A4(_08083_),
    .ZN(_08084_));
 OAI21_X1 _33125_ (.A(_06383_),
    .B1(_05666_),
    .B2(_05784_),
    .ZN(_08085_));
 AND3_X1 _33126_ (.A1(_08085_),
    .A2(_06394_),
    .A3(_07371_),
    .ZN(_08086_));
 AND4_X1 _33127_ (.A1(_08075_),
    .A2(_08079_),
    .A3(_08084_),
    .A4(_08086_),
    .ZN(_08087_));
 OAI21_X1 _33128_ (.A(_06455_),
    .B1(_07770_),
    .B2(_05692_),
    .ZN(_08088_));
 OAI21_X1 _33129_ (.A(_05804_),
    .B1(_06386_),
    .B2(_05763_),
    .ZN(_08089_));
 NAND2_X1 _33130_ (.A1(_05804_),
    .A2(_05799_),
    .ZN(_08090_));
 NAND4_X1 _33131_ (.A1(_05738_),
    .A2(_05807_),
    .A3(_05809_),
    .A4(_05827_),
    .ZN(_08092_));
 AND4_X1 _33132_ (.A1(_06448_),
    .A2(_08089_),
    .A3(_08090_),
    .A4(_08092_),
    .ZN(_08093_));
 OAI21_X1 _33133_ (.A(_06437_),
    .B1(_05796_),
    .B2(_07360_),
    .ZN(_08094_));
 NAND4_X1 _33134_ (.A1(_05784_),
    .A2(_06392_),
    .A3(_05809_),
    .A4(_05745_),
    .ZN(_08095_));
 NAND4_X1 _33135_ (.A1(_06392_),
    .A2(_06371_),
    .A3(_05603_),
    .A4(_05809_),
    .ZN(_08096_));
 AND3_X1 _33136_ (.A1(_08094_),
    .A2(_08095_),
    .A3(_08096_),
    .ZN(_08097_));
 NAND2_X1 _33137_ (.A1(_05611_),
    .A2(_06442_),
    .ZN(_08098_));
 NAND2_X1 _33138_ (.A1(_05661_),
    .A2(_06442_),
    .ZN(_08099_));
 NAND2_X1 _33139_ (.A1(_06442_),
    .A2(_05646_),
    .ZN(_08100_));
 AND4_X1 _33140_ (.A1(_08098_),
    .A2(_06819_),
    .A3(_08099_),
    .A4(_08100_),
    .ZN(_08101_));
 AND4_X1 _33141_ (.A1(_08088_),
    .A2(_08093_),
    .A3(_08097_),
    .A4(_08101_),
    .ZN(_08103_));
 NAND4_X1 _33142_ (.A1(_08056_),
    .A2(_08072_),
    .A3(_08087_),
    .A4(_08103_),
    .ZN(_08104_));
 NOR2_X1 _33143_ (.A1(_08104_),
    .A2(_05829_),
    .ZN(_08105_));
 XOR2_X2 _33144_ (.A(_08037_),
    .B(_08105_),
    .Z(_08106_));
 AND4_X1 _33145_ (.A1(_05854_),
    .A2(_05893_),
    .A3(_05858_),
    .A4(_05880_),
    .ZN(_08107_));
 AND2_X1 _33146_ (.A1(_05882_),
    .A2(_05912_),
    .ZN(_08108_));
 AOI211_X4 _33147_ (.A(_08107_),
    .B(_08108_),
    .C1(_05977_),
    .C2(_05883_),
    .ZN(_08109_));
 OAI21_X1 _33148_ (.A(_05883_),
    .B1(_06029_),
    .B2(_06010_),
    .ZN(_08110_));
 OAI21_X1 _33149_ (.A(_05883_),
    .B1(_06022_),
    .B2(_06680_),
    .ZN(_08111_));
 AND3_X1 _33150_ (.A1(_08109_),
    .A2(_08110_),
    .A3(_08111_),
    .ZN(_08112_));
 AND2_X1 _33151_ (.A1(_05971_),
    .A2(_06004_),
    .ZN(_08114_));
 INV_X1 _33152_ (.A(_08114_),
    .ZN(_08115_));
 NAND2_X1 _33153_ (.A1(_07864_),
    .A2(_08115_),
    .ZN(_08116_));
 AND3_X1 _33154_ (.A1(_05920_),
    .A2(_05999_),
    .A3(_05858_),
    .ZN(_08117_));
 NOR4_X1 _33155_ (.A1(_08116_),
    .A2(_06070_),
    .A3(_06074_),
    .A4(_08117_),
    .ZN(_08118_));
 NOR4_X1 _33156_ (.A1(_06742_),
    .A2(_06701_),
    .A3(_06961_),
    .A4(_07187_),
    .ZN(_08119_));
 AND2_X1 _33157_ (.A1(_05914_),
    .A2(_06010_),
    .ZN(_08120_));
 AND2_X1 _33158_ (.A1(_05921_),
    .A2(_06016_),
    .ZN(_08121_));
 NOR4_X1 _33159_ (.A1(_08120_),
    .A2(_08121_),
    .A3(_07168_),
    .A4(_07866_),
    .ZN(_08122_));
 OAI21_X1 _33160_ (.A(_06055_),
    .B1(_07185_),
    .B2(_06698_),
    .ZN(_08123_));
 NAND3_X1 _33161_ (.A1(_05895_),
    .A2(_06059_),
    .A3(_05884_),
    .ZN(_08125_));
 AND3_X1 _33162_ (.A1(_07568_),
    .A2(_08123_),
    .A3(_08125_),
    .ZN(_08126_));
 AND4_X1 _33163_ (.A1(_08118_),
    .A2(_08119_),
    .A3(_08122_),
    .A4(_08126_),
    .ZN(_08127_));
 NAND3_X1 _33164_ (.A1(_07141_),
    .A2(_07136_),
    .A3(_06994_),
    .ZN(_08128_));
 AOI21_X1 _33165_ (.A(_06772_),
    .B1(_06761_),
    .B2(_06717_),
    .ZN(_08129_));
 AOI21_X1 _33166_ (.A(_06772_),
    .B1(_07206_),
    .B2(_07897_),
    .ZN(_08130_));
 NOR4_X1 _33167_ (.A1(_08128_),
    .A2(_06042_),
    .A3(_08129_),
    .A4(_08130_),
    .ZN(_08131_));
 AND2_X1 _33168_ (.A1(_05895_),
    .A2(_06022_),
    .ZN(_08132_));
 AND2_X1 _33169_ (.A1(_05909_),
    .A2(_05949_),
    .ZN(_08133_));
 OR4_X1 _33170_ (.A1(_06995_),
    .A2(_08132_),
    .A3(_08133_),
    .A4(_07026_),
    .ZN(_08134_));
 OAI221_X1 _33171_ (.A(_05916_),
    .B1(_06773_),
    .B2(_06007_),
    .C1(_05978_),
    .C2(_06090_),
    .ZN(_08136_));
 NOR3_X1 _33172_ (.A1(_08134_),
    .A2(_06088_),
    .A3(_08136_),
    .ZN(_08137_));
 AND4_X1 _33173_ (.A1(_08112_),
    .A2(_08127_),
    .A3(_08131_),
    .A4(_08137_),
    .ZN(_08138_));
 AOI221_X4 _33174_ (.A(_07870_),
    .B1(_05934_),
    .B2(_05972_),
    .C1(_05977_),
    .C2(_05936_),
    .ZN(_08139_));
 OR4_X1 _33175_ (.A1(_05993_),
    .A2(_07146_),
    .A3(_07152_),
    .A4(_07132_),
    .ZN(_08140_));
 AND2_X1 _33176_ (.A1(_06946_),
    .A2(_06044_),
    .ZN(_08141_));
 OAI22_X1 _33177_ (.A1(_06695_),
    .A2(_06718_),
    .B1(_07162_),
    .B2(_05979_),
    .ZN(_08142_));
 OAI22_X1 _33178_ (.A1(_06090_),
    .A2(_07897_),
    .B1(_06085_),
    .B2(_06718_),
    .ZN(_08143_));
 NOR4_X1 _33179_ (.A1(_08140_),
    .A2(_08141_),
    .A3(_08142_),
    .A4(_08143_),
    .ZN(_08144_));
 AND4_X1 _33180_ (.A1(_06983_),
    .A2(_06980_),
    .A3(_07569_),
    .A4(_07209_),
    .ZN(_08145_));
 NOR3_X1 _33181_ (.A1(_05861_),
    .A2(_06752_),
    .A3(_06764_),
    .ZN(_08147_));
 AOI22_X1 _33182_ (.A1(_06680_),
    .A2(_06946_),
    .B1(_06004_),
    .B2(_06002_),
    .ZN(_08148_));
 AOI22_X1 _33183_ (.A1(_06029_),
    .A2(_06089_),
    .B1(_05949_),
    .B2(_05855_),
    .ZN(_08149_));
 AND4_X1 _33184_ (.A1(_08145_),
    .A2(_08147_),
    .A3(_08148_),
    .A4(_08149_),
    .ZN(_08150_));
 OAI21_X1 _33185_ (.A(_06043_),
    .B1(_05855_),
    .B2(_05961_),
    .ZN(_08151_));
 OAI21_X1 _33186_ (.A(_08151_),
    .B1(_06761_),
    .B2(_06058_),
    .ZN(_08152_));
 NOR2_X1 _33187_ (.A1(_05996_),
    .A2(_06040_),
    .ZN(_08153_));
 AND2_X1 _33188_ (.A1(_05921_),
    .A2(_06056_),
    .ZN(_08154_));
 AOI21_X1 _33189_ (.A(_05939_),
    .B1(_07206_),
    .B2(_05965_),
    .ZN(_08155_));
 NOR4_X1 _33190_ (.A1(_08152_),
    .A2(_08153_),
    .A3(_08154_),
    .A4(_08155_),
    .ZN(_08156_));
 AND4_X1 _33191_ (.A1(_08139_),
    .A2(_08144_),
    .A3(_08150_),
    .A4(_08156_),
    .ZN(_08158_));
 NAND2_X1 _33192_ (.A1(_08138_),
    .A2(_08158_),
    .ZN(_08159_));
 XNOR2_X1 _33193_ (.A(_08159_),
    .B(_00995_),
    .ZN(_08160_));
 XNOR2_X1 _33194_ (.A(_08106_),
    .B(_08160_),
    .ZN(_08161_));
 OAI22_X1 _33195_ (.A1(_06615_),
    .A2(_07067_),
    .B1(_07071_),
    .B2(_06311_),
    .ZN(_08162_));
 AOI221_X4 _33196_ (.A(_08162_),
    .B1(_06631_),
    .B2(_06326_),
    .C1(_06330_),
    .C2(_06610_),
    .ZN(_08163_));
 NAND2_X1 _33197_ (.A1(_06603_),
    .A2(_06189_),
    .ZN(_08164_));
 NAND3_X1 _33198_ (.A1(_06189_),
    .A2(_06594_),
    .A3(_06186_),
    .ZN(_08165_));
 AND4_X1 _33199_ (.A1(_06323_),
    .A2(_06656_),
    .A3(_08164_),
    .A4(_08165_),
    .ZN(_08166_));
 NOR4_X1 _33200_ (.A1(_07047_),
    .A2(_06135_),
    .A3(_07099_),
    .A4(_07037_),
    .ZN(_08167_));
 AND4_X1 _33201_ (.A1(_07229_),
    .A2(_08163_),
    .A3(_08166_),
    .A4(_08167_),
    .ZN(_08169_));
 INV_X1 _33202_ (.A(_07298_),
    .ZN(_08170_));
 INV_X1 _33203_ (.A(_07517_),
    .ZN(_08171_));
 AOI21_X1 _33204_ (.A(_07115_),
    .B1(_08170_),
    .B2(_08171_),
    .ZN(_08172_));
 AOI21_X1 _33205_ (.A(_07082_),
    .B1(_07116_),
    .B2(_07048_),
    .ZN(_08173_));
 AND3_X1 _33206_ (.A1(_06326_),
    .A2(_06211_),
    .A3(_06206_),
    .ZN(_08174_));
 NOR4_X1 _33207_ (.A1(_08172_),
    .A2(_08173_),
    .A3(_07296_),
    .A4(_08174_),
    .ZN(_08175_));
 NAND2_X1 _33208_ (.A1(_06304_),
    .A2(_06189_),
    .ZN(_08176_));
 AND2_X1 _33209_ (.A1(_06113_),
    .A2(_06256_),
    .ZN(_08177_));
 AOI221_X4 _33210_ (.A(_08177_),
    .B1(_06301_),
    .B2(_06291_),
    .C1(_06201_),
    .C2(_06667_),
    .ZN(_08178_));
 AOI22_X1 _33211_ (.A1(_06164_),
    .A2(_07222_),
    .B1(_06631_),
    .B2(_06236_),
    .ZN(_08180_));
 NAND2_X1 _33212_ (.A1(_06330_),
    .A2(_06113_),
    .ZN(_08181_));
 AND3_X1 _33213_ (.A1(_08180_),
    .A2(_08181_),
    .A3(_07265_),
    .ZN(_08182_));
 NAND2_X1 _33214_ (.A1(_06173_),
    .A2(_06236_),
    .ZN(_08183_));
 OAI21_X1 _33215_ (.A(_06257_),
    .B1(_06153_),
    .B2(_06218_),
    .ZN(_08184_));
 AND3_X1 _33216_ (.A1(_07465_),
    .A2(_08183_),
    .A3(_08184_),
    .ZN(_08185_));
 AND4_X1 _33217_ (.A1(_08176_),
    .A2(_08178_),
    .A3(_08182_),
    .A4(_08185_),
    .ZN(_08186_));
 NAND2_X1 _33218_ (.A1(_06186_),
    .A2(_06263_),
    .ZN(_08187_));
 AOI21_X1 _33219_ (.A(_07964_),
    .B1(_07046_),
    .B2(_08187_),
    .ZN(_08188_));
 AOI21_X1 _33220_ (.A(_08188_),
    .B1(_06641_),
    .B2(_06642_),
    .ZN(_08189_));
 OAI21_X1 _33221_ (.A(_06309_),
    .B1(_06306_),
    .B2(_06209_),
    .ZN(_08191_));
 OAI21_X1 _33222_ (.A(_06627_),
    .B1(_06258_),
    .B2(_06594_),
    .ZN(_08192_));
 AND4_X1 _33223_ (.A1(_07125_),
    .A2(_08189_),
    .A3(_08191_),
    .A4(_08192_),
    .ZN(_08193_));
 AND4_X1 _33224_ (.A1(_08169_),
    .A2(_08175_),
    .A3(_08186_),
    .A4(_08193_),
    .ZN(_08194_));
 AND2_X1 _33225_ (.A1(_06326_),
    .A2(_06605_),
    .ZN(_08195_));
 AND2_X1 _33226_ (.A1(_06330_),
    .A2(_06178_),
    .ZN(_08196_));
 OR2_X1 _33227_ (.A1(_08195_),
    .A2(_08196_),
    .ZN(_08197_));
 AOI21_X1 _33228_ (.A(_06637_),
    .B1(_07058_),
    .B2(_08187_),
    .ZN(_08198_));
 AOI21_X1 _33229_ (.A(_06583_),
    .B1(_06561_),
    .B2(_07097_),
    .ZN(_08199_));
 NOR4_X1 _33230_ (.A1(_08197_),
    .A2(_06648_),
    .A3(_08198_),
    .A4(_08199_),
    .ZN(_08200_));
 OR4_X1 _33231_ (.A1(_06609_),
    .A2(_07077_),
    .A3(_06559_),
    .A4(_07247_),
    .ZN(_08202_));
 OAI22_X1 _33232_ (.A1(_06562_),
    .A2(_06638_),
    .B1(_06115_),
    .B2(_07059_),
    .ZN(_08203_));
 NOR4_X1 _33233_ (.A1(_08202_),
    .A2(_07494_),
    .A3(_07958_),
    .A4(_08203_),
    .ZN(_08204_));
 OAI21_X1 _33234_ (.A(_06260_),
    .B1(_06269_),
    .B2(_06261_),
    .ZN(_08205_));
 AND3_X1 _33235_ (.A1(_06188_),
    .A2(_06294_),
    .A3(_06191_),
    .ZN(_08206_));
 NOR4_X1 _33236_ (.A1(_08205_),
    .A2(_06148_),
    .A3(_06253_),
    .A4(_08206_),
    .ZN(_08207_));
 AOI22_X1 _33237_ (.A1(_06572_),
    .A2(_06201_),
    .B1(_06230_),
    .B2(_06274_),
    .ZN(_08208_));
 AOI22_X1 _33238_ (.A1(_06631_),
    .A2(_06572_),
    .B1(_06218_),
    .B2(_06658_),
    .ZN(_08209_));
 AND4_X1 _33239_ (.A1(_06172_),
    .A2(_08207_),
    .A3(_08208_),
    .A4(_08209_),
    .ZN(_08210_));
 NOR4_X1 _33240_ (.A1(_07480_),
    .A2(_07930_),
    .A3(_06612_),
    .A4(_07515_),
    .ZN(_08211_));
 AND4_X1 _33241_ (.A1(_08200_),
    .A2(_08204_),
    .A3(_08210_),
    .A4(_08211_),
    .ZN(_08213_));
 NAND2_X1 _33242_ (.A1(_08194_),
    .A2(_08213_),
    .ZN(_08214_));
 XNOR2_X1 _33243_ (.A(_08214_),
    .B(_07859_),
    .ZN(_08215_));
 XNOR2_X1 _33244_ (.A(_08161_),
    .B(_08215_),
    .ZN(_08216_));
 MUX2_X2 _33245_ (.A(_07983_),
    .B(_08216_),
    .S(_05156_),
    .Z(_00706_));
 XOR2_X1 _33246_ (.A(_17205_),
    .B(_17016_),
    .Z(_08217_));
 AOI211_X2 _33247_ (.A(_05783_),
    .B(_05780_),
    .C1(_16797_),
    .C2(_05638_),
    .ZN(_08218_));
 AND2_X2 _33248_ (.A1(_05692_),
    .A2(_05779_),
    .ZN(_08219_));
 OR4_X4 _33249_ (.A1(_05782_),
    .A2(_08218_),
    .A3(_06440_),
    .A4(_08219_),
    .ZN(_08220_));
 AND3_X1 _33250_ (.A1(_05815_),
    .A2(_05722_),
    .A3(_05694_),
    .ZN(_08221_));
 NAND2_X1 _33251_ (.A1(_07317_),
    .A2(_07757_),
    .ZN(_08223_));
 NOR4_X4 _33252_ (.A1(_08220_),
    .A2(_06454_),
    .A3(_08221_),
    .A4(_08223_),
    .ZN(_08224_));
 AOI221_X4 _33253_ (.A(_06414_),
    .B1(_05712_),
    .B2(_05748_),
    .C1(_05602_),
    .C2(_06389_),
    .ZN(_08225_));
 AND2_X1 _33254_ (.A1(_05770_),
    .A2(_06387_),
    .ZN(_08226_));
 AOI21_X1 _33255_ (.A(_05743_),
    .B1(_05749_),
    .B2(_05584_),
    .ZN(_08227_));
 NOR4_X1 _33256_ (.A1(_08225_),
    .A2(_07775_),
    .A3(_08226_),
    .A4(_08227_),
    .ZN(_08228_));
 NAND3_X1 _33257_ (.A1(_05762_),
    .A2(_05636_),
    .A3(_05789_),
    .ZN(_08229_));
 NAND2_X1 _33258_ (.A1(_08229_),
    .A2(_07649_),
    .ZN(_08230_));
 AND3_X1 _33259_ (.A1(_06390_),
    .A2(_05636_),
    .A3(_05789_),
    .ZN(_08231_));
 NOR3_X1 _33260_ (.A1(_08230_),
    .A2(_07334_),
    .A3(_08231_),
    .ZN(_08232_));
 OAI21_X1 _33261_ (.A(_05804_),
    .B1(_05692_),
    .B2(_06387_),
    .ZN(_08234_));
 OAI211_X2 _33262_ (.A(_05803_),
    .B(_05595_),
    .C1(_05712_),
    .C2(_05638_),
    .ZN(_08235_));
 AND4_X1 _33263_ (.A1(_08090_),
    .A2(_08232_),
    .A3(_08234_),
    .A4(_08235_),
    .ZN(_08236_));
 NAND3_X1 _33264_ (.A1(_05799_),
    .A2(_05677_),
    .A3(_05735_),
    .ZN(_08237_));
 AND3_X1 _33265_ (.A1(_05754_),
    .A2(_05744_),
    .A3(_06390_),
    .ZN(_08238_));
 NOR2_X1 _33266_ (.A1(_07343_),
    .A2(_08238_),
    .ZN(_08239_));
 OAI21_X1 _33267_ (.A(_05757_),
    .B1(_06821_),
    .B2(_05794_),
    .ZN(_08240_));
 OAI211_X2 _33268_ (.A(_05636_),
    .B(_05735_),
    .C1(_05612_),
    .C2(_06397_),
    .ZN(_08241_));
 AND4_X1 _33269_ (.A1(_08237_),
    .A2(_08239_),
    .A3(_08240_),
    .A4(_08241_),
    .ZN(_08242_));
 AND4_X4 _33270_ (.A1(_08224_),
    .A2(_08228_),
    .A3(_08236_),
    .A4(_08242_),
    .ZN(_08243_));
 OAI21_X1 _33271_ (.A(_05637_),
    .B1(_06403_),
    .B2(_05641_),
    .ZN(_08245_));
 NAND4_X1 _33272_ (.A1(_05636_),
    .A2(_05573_),
    .A3(_05638_),
    .A4(_05722_),
    .ZN(_08246_));
 OAI21_X1 _33273_ (.A(_05637_),
    .B1(_05793_),
    .B2(_05719_),
    .ZN(_08247_));
 NAND3_X1 _33274_ (.A1(_08245_),
    .A2(_08246_),
    .A3(_08247_),
    .ZN(_08248_));
 INV_X1 _33275_ (.A(_08248_),
    .ZN(_08249_));
 OAI21_X1 _33276_ (.A(_05576_),
    .B1(_06386_),
    .B2(_05763_),
    .ZN(_08250_));
 OAI21_X1 _33277_ (.A(_05576_),
    .B1(_05679_),
    .B2(_05788_),
    .ZN(_08251_));
 AND3_X1 _33278_ (.A1(_08249_),
    .A2(_08250_),
    .A3(_08251_),
    .ZN(_08252_));
 NAND4_X1 _33279_ (.A1(_05707_),
    .A2(_05704_),
    .A3(_08063_),
    .A4(_07382_),
    .ZN(_08253_));
 AND2_X1 _33280_ (.A1(_05666_),
    .A2(_05716_),
    .ZN(_08254_));
 AOI21_X1 _33281_ (.A(_05717_),
    .B1(_05680_),
    .B2(_07375_),
    .ZN(_08256_));
 NOR4_X1 _33282_ (.A1(_08253_),
    .A2(_08254_),
    .A3(_08070_),
    .A4(_08256_),
    .ZN(_08257_));
 OAI21_X1 _33283_ (.A(_05608_),
    .B1(_07316_),
    .B2(_05713_),
    .ZN(_08258_));
 OAI21_X1 _33284_ (.A(_05608_),
    .B1(_05684_),
    .B2(_05583_),
    .ZN(_08259_));
 NAND3_X1 _33285_ (.A1(_08258_),
    .A2(_08259_),
    .A3(_06837_),
    .ZN(_08260_));
 OAI21_X1 _33286_ (.A(_06398_),
    .B1(_07622_),
    .B2(_05749_),
    .ZN(_08261_));
 NOR4_X1 _33287_ (.A1(_08260_),
    .A2(_08261_),
    .A3(_07626_),
    .A4(_06396_),
    .ZN(_08262_));
 OAI21_X1 _33288_ (.A(_05691_),
    .B1(_05762_),
    .B2(_05583_),
    .ZN(_08263_));
 OAI21_X1 _33289_ (.A(_08263_),
    .B1(_07753_),
    .B2(_06360_),
    .ZN(_08264_));
 AOI21_X1 _33290_ (.A(_05681_),
    .B1(_07753_),
    .B2(_05597_),
    .ZN(_08265_));
 OAI21_X1 _33291_ (.A(_05691_),
    .B1(_05679_),
    .B2(_05799_),
    .ZN(_08267_));
 OAI211_X2 _33292_ (.A(_08267_),
    .B(_06860_),
    .C1(_06360_),
    .C2(_06423_),
    .ZN(_08268_));
 NOR3_X1 _33293_ (.A1(_08264_),
    .A2(_08265_),
    .A3(_08268_),
    .ZN(_08269_));
 AND4_X1 _33294_ (.A1(_08252_),
    .A2(_08257_),
    .A3(_08262_),
    .A4(_08269_),
    .ZN(_08270_));
 AND2_X4 _33295_ (.A1(_08243_),
    .A2(_08270_),
    .ZN(_08271_));
 BUF_X8 _33296_ (.A(_08271_),
    .Z(_08272_));
 XNOR2_X2 _33297_ (.A(_08272_),
    .B(_05570_),
    .ZN(_08273_));
 AND2_X1 _33298_ (.A1(_06025_),
    .A2(_06033_),
    .ZN(_08274_));
 AND2_X1 _33299_ (.A1(_05943_),
    .A2(_06032_),
    .ZN(_08275_));
 AND2_X1 _33300_ (.A1(_06032_),
    .A2(_05912_),
    .ZN(_08276_));
 OR4_X1 _33301_ (.A1(_08274_),
    .A2(_06770_),
    .A3(_08275_),
    .A4(_08276_),
    .ZN(_08278_));
 NOR2_X1 _33302_ (.A1(_06780_),
    .A2(_06782_),
    .ZN(_08279_));
 OAI21_X1 _33303_ (.A(_05936_),
    .B1(_05997_),
    .B2(_07193_),
    .ZN(_08280_));
 OAI211_X2 _33304_ (.A(_08279_),
    .B(_08280_),
    .C1(_05939_),
    .C2(_05952_),
    .ZN(_08281_));
 NOR4_X1 _33305_ (.A1(_08278_),
    .A2(_08281_),
    .A3(_06086_),
    .A4(_06768_),
    .ZN(_08282_));
 AND2_X1 _33306_ (.A1(_07030_),
    .A2(_05868_),
    .ZN(_08283_));
 AND2_X1 _33307_ (.A1(_06015_),
    .A2(_05901_),
    .ZN(_08284_));
 OR4_X1 _33308_ (.A1(_06019_),
    .A2(_08283_),
    .A3(_08284_),
    .A4(_06775_),
    .ZN(_08285_));
 AOI21_X1 _33309_ (.A(_05946_),
    .B1(_06000_),
    .B2(_06095_),
    .ZN(_08286_));
 AOI21_X1 _33310_ (.A(_05946_),
    .B1(_07206_),
    .B2(_05979_),
    .ZN(_08287_));
 NOR4_X2 _33311_ (.A1(_08285_),
    .A2(_07132_),
    .A3(_08286_),
    .A4(_08287_),
    .ZN(_08289_));
 NAND2_X1 _33312_ (.A1(_06022_),
    .A2(_06055_),
    .ZN(_08290_));
 OAI21_X1 _33313_ (.A(_05895_),
    .B1(_06690_),
    .B2(_06706_),
    .ZN(_08291_));
 OAI21_X1 _33314_ (.A(_05895_),
    .B1(_05909_),
    .B2(_05923_),
    .ZN(_08292_));
 OAI21_X1 _33315_ (.A(_06055_),
    .B1(_06096_),
    .B2(_06025_),
    .ZN(_08293_));
 AND4_X1 _33316_ (.A1(_08290_),
    .A2(_08291_),
    .A3(_08292_),
    .A4(_08293_),
    .ZN(_08294_));
 AND3_X1 _33317_ (.A1(_05991_),
    .A2(_05975_),
    .A3(_05870_),
    .ZN(_08295_));
 OR4_X1 _33318_ (.A1(_06739_),
    .A2(_08295_),
    .A3(_06949_),
    .A4(_07862_),
    .ZN(_08296_));
 NOR4_X1 _33319_ (.A1(_08296_),
    .A2(_06082_),
    .A3(_07896_),
    .A4(_08108_),
    .ZN(_08297_));
 AND4_X1 _33320_ (.A1(_08282_),
    .A2(_08289_),
    .A3(_08294_),
    .A4(_08297_),
    .ZN(_08298_));
 OAI211_X2 _33321_ (.A(_05847_),
    .B(_05836_),
    .C1(_05985_),
    .C2(_05912_),
    .ZN(_08300_));
 AND4_X1 _33322_ (.A1(_06071_),
    .A2(_08300_),
    .A3(_06694_),
    .A4(_05963_),
    .ZN(_08301_));
 OAI21_X1 _33323_ (.A(_05921_),
    .B1(_06075_),
    .B2(_06705_),
    .ZN(_08302_));
 OAI21_X1 _33324_ (.A(_05921_),
    .B1(_05915_),
    .B2(_05961_),
    .ZN(_08303_));
 AND4_X1 _33325_ (.A1(_06702_),
    .A2(_08301_),
    .A3(_08302_),
    .A4(_08303_),
    .ZN(_08304_));
 AND3_X1 _33326_ (.A1(_05943_),
    .A2(_06063_),
    .A3(_05902_),
    .ZN(_08305_));
 NOR3_X1 _33327_ (.A1(_06716_),
    .A2(_05889_),
    .A3(_06060_),
    .ZN(_08306_));
 AOI211_X4 _33328_ (.A(_08305_),
    .B(_08306_),
    .C1(_05971_),
    .C2(_05912_),
    .ZN(_08307_));
 AOI211_X4 _33329_ (.A(_06724_),
    .B(_07203_),
    .C1(_05926_),
    .C2(_07133_),
    .ZN(_08308_));
 OAI21_X1 _33330_ (.A(_05971_),
    .B1(_05997_),
    .B2(_05964_),
    .ZN(_08309_));
 INV_X1 _33331_ (.A(_08309_),
    .ZN(_08311_));
 NOR4_X1 _33332_ (.A1(_08311_),
    .A2(_06715_),
    .A3(_07016_),
    .A4(_08114_),
    .ZN(_08312_));
 AND3_X1 _33333_ (.A1(_08307_),
    .A2(_08308_),
    .A3(_08312_),
    .ZN(_08313_));
 AOI21_X1 _33334_ (.A(_06065_),
    .B1(_07593_),
    .B2(_06005_),
    .ZN(_08314_));
 NAND3_X1 _33335_ (.A1(_05865_),
    .A2(_06063_),
    .A3(_05836_),
    .ZN(_08315_));
 OAI211_X2 _33336_ (.A(_06979_),
    .B(_08315_),
    .C1(_06065_),
    .C2(_06773_),
    .ZN(_08316_));
 AOI21_X1 _33337_ (.A(_06090_),
    .B1(_07875_),
    .B2(_06684_),
    .ZN(_08317_));
 AOI21_X1 _33338_ (.A(_06090_),
    .B1(_06959_),
    .B2(_06696_),
    .ZN(_08318_));
 NOR4_X1 _33339_ (.A1(_08314_),
    .A2(_08316_),
    .A3(_08317_),
    .A4(_08318_),
    .ZN(_08319_));
 OAI21_X1 _33340_ (.A(_06002_),
    .B1(_06680_),
    .B2(_07193_),
    .ZN(_08320_));
 NOR2_X1 _33341_ (.A1(_05953_),
    .A2(_08133_),
    .ZN(_08322_));
 OAI21_X1 _33342_ (.A(_05949_),
    .B1(_05958_),
    .B2(_06029_),
    .ZN(_08323_));
 OAI211_X2 _33343_ (.A(_06002_),
    .B(_06034_),
    .C1(_05999_),
    .C2(_05854_),
    .ZN(_08324_));
 AND4_X1 _33344_ (.A1(_08320_),
    .A2(_08322_),
    .A3(_08323_),
    .A4(_08324_),
    .ZN(_08325_));
 AND4_X1 _33345_ (.A1(_08304_),
    .A2(_08313_),
    .A3(_08319_),
    .A4(_08325_),
    .ZN(_08326_));
 AND2_X2 _33346_ (.A1(_08298_),
    .A2(_08326_),
    .ZN(_08327_));
 BUF_X8 _33347_ (.A(_08327_),
    .Z(_08328_));
 XNOR2_X1 _33348_ (.A(_08328_),
    .B(_00996_),
    .ZN(_08329_));
 XNOR2_X1 _33349_ (.A(_08273_),
    .B(_08329_),
    .ZN(_08330_));
 INV_X1 _33350_ (.A(_07970_),
    .ZN(_08331_));
 OAI211_X2 _33351_ (.A(_07530_),
    .B(_08331_),
    .C1(_06240_),
    .C2(_06224_),
    .ZN(_08333_));
 NAND2_X1 _33352_ (.A1(_06218_),
    .A2(_06627_),
    .ZN(_08334_));
 OAI21_X1 _33353_ (.A(_08334_),
    .B1(_07061_),
    .B2(_06224_),
    .ZN(_08335_));
 NAND2_X1 _33354_ (.A1(_06631_),
    .A2(_06236_),
    .ZN(_08336_));
 OAI211_X2 _33355_ (.A(_08336_),
    .B(_07531_),
    .C1(_06302_),
    .C2(_06241_),
    .ZN(_08337_));
 OR4_X4 _33356_ (.A1(_06238_),
    .A2(_08333_),
    .A3(_08335_),
    .A4(_08337_),
    .ZN(_08338_));
 OAI21_X1 _33357_ (.A(_07273_),
    .B1(_06617_),
    .B2(_06672_),
    .ZN(_08339_));
 OAI21_X1 _33358_ (.A(_06635_),
    .B1(_06201_),
    .B2(_06113_),
    .ZN(_08340_));
 NAND3_X1 _33359_ (.A1(_06591_),
    .A2(_06203_),
    .A3(_06167_),
    .ZN(_08341_));
 OAI211_X2 _33360_ (.A(_08340_),
    .B(_08341_),
    .C1(_06269_),
    .C2(_06637_),
    .ZN(_08342_));
 NAND2_X1 _33361_ (.A1(_06635_),
    .A2(_06177_),
    .ZN(_08344_));
 OAI211_X2 _33362_ (.A(_08344_),
    .B(_07042_),
    .C1(_06637_),
    .C2(_06122_),
    .ZN(_08345_));
 NOR4_X2 _33363_ (.A1(_08338_),
    .A2(_08339_),
    .A3(_08342_),
    .A4(_08345_),
    .ZN(_08346_));
 AND3_X1 _33364_ (.A1(_06658_),
    .A2(_06192_),
    .A3(_06206_),
    .ZN(_08347_));
 OR4_X1 _33365_ (.A1(_06145_),
    .A2(_08347_),
    .A3(_06154_),
    .A4(_06158_),
    .ZN(_08348_));
 NAND2_X1 _33366_ (.A1(_06641_),
    .A2(_06657_),
    .ZN(_08349_));
 NAND4_X1 _33367_ (.A1(_07091_),
    .A2(_08349_),
    .A3(_06643_),
    .A4(_07524_),
    .ZN(_08350_));
 OAI21_X1 _33368_ (.A(_06216_),
    .B1(_06230_),
    .B2(_07517_),
    .ZN(_08351_));
 OAI21_X1 _33369_ (.A(_08351_),
    .B1(_08170_),
    .B2(_07082_),
    .ZN(_08352_));
 OAI21_X1 _33370_ (.A(_06667_),
    .B1(_06668_),
    .B2(_06304_),
    .ZN(_08353_));
 OAI21_X1 _33371_ (.A(_06667_),
    .B1(_06642_),
    .B2(_06331_),
    .ZN(_08355_));
 OAI211_X2 _33372_ (.A(_08353_),
    .B(_08355_),
    .C1(_06269_),
    .C2(_06115_),
    .ZN(_08356_));
 NOR4_X1 _33373_ (.A1(_08348_),
    .A2(_08350_),
    .A3(_08352_),
    .A4(_08356_),
    .ZN(_08357_));
 OR4_X1 _33374_ (.A1(_06327_),
    .A2(_07464_),
    .A3(_08195_),
    .A4(_07064_),
    .ZN(_08358_));
 OAI21_X1 _33375_ (.A(_06309_),
    .B1(_06313_),
    .B2(_07044_),
    .ZN(_08359_));
 OAI21_X1 _33376_ (.A(_06309_),
    .B1(_06177_),
    .B2(_06178_),
    .ZN(_08360_));
 OAI211_X2 _33377_ (.A(_08359_),
    .B(_08360_),
    .C1(_07071_),
    .C2(_08171_),
    .ZN(_08361_));
 NAND2_X1 _33378_ (.A1(_06301_),
    .A2(_06291_),
    .ZN(_08362_));
 NAND4_X1 _33379_ (.A1(_07923_),
    .A2(_07251_),
    .A3(_07252_),
    .A4(_08362_),
    .ZN(_08363_));
 OAI211_X2 _33380_ (.A(_06330_),
    .B(_16879_),
    .C1(_06194_),
    .C2(_06109_),
    .ZN(_08364_));
 OAI211_X2 _33381_ (.A(_06298_),
    .B(_06143_),
    .C1(_06642_),
    .C2(_06331_),
    .ZN(_08366_));
 OAI211_X2 _33382_ (.A(_08364_),
    .B(_08366_),
    .C1(_08170_),
    .C2(_07057_),
    .ZN(_08367_));
 NOR4_X1 _33383_ (.A1(_08358_),
    .A2(_08361_),
    .A3(_08363_),
    .A4(_08367_),
    .ZN(_08368_));
 AOI211_X4 _33384_ (.A(_06266_),
    .B(_06575_),
    .C1(_06631_),
    .C2(_07222_),
    .ZN(_08369_));
 OAI21_X1 _33385_ (.A(_06257_),
    .B1(_06230_),
    .B2(_06610_),
    .ZN(_08370_));
 OAI21_X1 _33386_ (.A(_07222_),
    .B1(_06156_),
    .B2(_06331_),
    .ZN(_08371_));
 OAI211_X2 _33387_ (.A(_06257_),
    .B(_06289_),
    .C1(_06205_),
    .C2(_06294_),
    .ZN(_08372_));
 NAND4_X1 _33388_ (.A1(_08369_),
    .A2(_08370_),
    .A3(_08371_),
    .A4(_08372_),
    .ZN(_08373_));
 AOI21_X1 _33389_ (.A(_06562_),
    .B1(_06584_),
    .B2(_07967_),
    .ZN(_08374_));
 AOI21_X1 _33390_ (.A(_06562_),
    .B1(_07955_),
    .B2(_08171_),
    .ZN(_08375_));
 INV_X1 _33391_ (.A(_07119_),
    .ZN(_08377_));
 OAI21_X1 _33392_ (.A(_06274_),
    .B1(_06113_),
    .B2(_06218_),
    .ZN(_08378_));
 NAND4_X1 _33393_ (.A1(_06276_),
    .A2(_08377_),
    .A3(_07245_),
    .A4(_08378_),
    .ZN(_08379_));
 NOR4_X1 _33394_ (.A1(_08373_),
    .A2(_08374_),
    .A3(_08375_),
    .A4(_08379_),
    .ZN(_08380_));
 NAND4_X1 _33395_ (.A1(_08346_),
    .A2(_08357_),
    .A3(_08368_),
    .A4(_08380_),
    .ZN(_08381_));
 NOR2_X2 _33396_ (.A1(_08381_),
    .A2(_06674_),
    .ZN(_08382_));
 XOR2_X1 _33397_ (.A(_08037_),
    .B(_08382_),
    .Z(_08383_));
 XNOR2_X1 _33398_ (.A(_08330_),
    .B(_08383_),
    .ZN(_08384_));
 BUF_X4 _33399_ (.A(_09098_),
    .Z(_08385_));
 MUX2_X1 _33400_ (.A(_08217_),
    .B(_08384_),
    .S(_08385_),
    .Z(_00707_));
 XOR2_X1 _33401_ (.A(_17206_),
    .B(_17017_),
    .Z(_08387_));
 XNOR2_X1 _33402_ (.A(_06676_),
    .B(_00997_),
    .ZN(_08388_));
 XNOR2_X1 _33403_ (.A(_05457_),
    .B(_05831_),
    .ZN(_08389_));
 XNOR2_X1 _33404_ (.A(_08389_),
    .B(_08328_),
    .ZN(_08390_));
 XNOR2_X1 _33405_ (.A(_08388_),
    .B(_08390_),
    .ZN(_08391_));
 MUX2_X1 _33406_ (.A(_08387_),
    .B(_08391_),
    .S(_08385_),
    .Z(_00668_));
 XOR2_X1 _33407_ (.A(_17207_),
    .B(_17018_),
    .Z(_08392_));
 XNOR2_X1 _33408_ (.A(_07126_),
    .B(_00998_),
    .ZN(_08393_));
 XOR2_X1 _33409_ (.A(_06676_),
    .B(_08393_),
    .Z(_08394_));
 XNOR2_X2 _33410_ (.A(_08328_),
    .B(_06100_),
    .ZN(_08395_));
 XNOR2_X1 _33411_ (.A(_06557_),
    .B(_08395_),
    .ZN(_08397_));
 XNOR2_X1 _33412_ (.A(_08394_),
    .B(_08397_),
    .ZN(_08398_));
 MUX2_X1 _33413_ (.A(_08392_),
    .B(_08398_),
    .S(_08385_),
    .Z(_00669_));
 XOR2_X1 _33414_ (.A(_17177_),
    .B(_17019_),
    .Z(_08399_));
 XOR2_X2 _33415_ (.A(_07126_),
    .B(_06786_),
    .Z(_08400_));
 XNOR2_X1 _33416_ (.A(_08400_),
    .B(_06945_),
    .ZN(_08401_));
 XNOR2_X1 _33417_ (.A(_07303_),
    .B(_00999_),
    .ZN(_08402_));
 XNOR2_X1 _33418_ (.A(_08401_),
    .B(_08402_),
    .ZN(_08403_));
 MUX2_X1 _33419_ (.A(_08399_),
    .B(_08403_),
    .S(_08385_),
    .Z(_00670_));
 XOR2_X1 _33420_ (.A(_17178_),
    .B(_17020_),
    .Z(_08404_));
 XOR2_X2 _33421_ (.A(_08328_),
    .B(_07033_),
    .Z(_08406_));
 XNOR2_X1 _33422_ (.A(_07537_),
    .B(_01000_),
    .ZN(_08407_));
 XNOR2_X1 _33423_ (.A(_08406_),
    .B(_08407_),
    .ZN(_08408_));
 XOR2_X1 _33424_ (.A(_08408_),
    .B(_07460_),
    .Z(_08409_));
 MUX2_X1 _33425_ (.A(_08404_),
    .B(_08409_),
    .S(_08385_),
    .Z(_00671_));
 XOR2_X1 _33426_ (.A(_17179_),
    .B(_17021_),
    .Z(_08410_));
 XNOR2_X1 _33427_ (.A(_07731_),
    .B(_01001_),
    .ZN(_08411_));
 XNOR2_X1 _33428_ (.A(_08328_),
    .B(_07217_),
    .ZN(_08412_));
 XOR2_X1 _33429_ (.A(_08411_),
    .B(_08412_),
    .Z(_08413_));
 XNOR2_X1 _33430_ (.A(_07538_),
    .B(_07979_),
    .ZN(_08414_));
 XNOR2_X1 _33431_ (.A(_08413_),
    .B(_08414_),
    .ZN(_08416_));
 MUX2_X1 _33432_ (.A(_08410_),
    .B(_08416_),
    .S(_08385_),
    .Z(_00672_));
 XOR2_X1 _33433_ (.A(_17180_),
    .B(_17022_),
    .Z(_08417_));
 XNOR2_X1 _33434_ (.A(_07805_),
    .B(_01002_),
    .ZN(_08418_));
 XNOR2_X1 _33435_ (.A(_07979_),
    .B(_07600_),
    .ZN(_08419_));
 XNOR2_X1 _33436_ (.A(_08418_),
    .B(_08419_),
    .ZN(_08420_));
 XNOR2_X1 _33437_ (.A(_08420_),
    .B(_08215_),
    .ZN(_08421_));
 MUX2_X1 _33438_ (.A(_08417_),
    .B(_08421_),
    .S(_08385_),
    .Z(_00673_));
 XOR2_X1 _33439_ (.A(_17181_),
    .B(_17024_),
    .Z(_08422_));
 XNOR2_X1 _33440_ (.A(_08382_),
    .B(_15485_),
    .ZN(_08423_));
 XNOR2_X1 _33441_ (.A(_08106_),
    .B(_08423_),
    .ZN(_08425_));
 XOR2_X1 _33442_ (.A(_08214_),
    .B(_07920_),
    .Z(_08426_));
 XNOR2_X1 _33443_ (.A(_08425_),
    .B(_08426_),
    .ZN(_08427_));
 MUX2_X1 _33444_ (.A(_08422_),
    .B(_08427_),
    .S(_08385_),
    .Z(_00674_));
 XOR2_X1 _33445_ (.A(_17182_),
    .B(_17025_),
    .Z(_08428_));
 XNOR2_X1 _33446_ (.A(_08159_),
    .B(_01004_),
    .ZN(_08429_));
 XNOR2_X1 _33447_ (.A(_08273_),
    .B(_08429_),
    .ZN(_08430_));
 XNOR2_X1 _33448_ (.A(_08382_),
    .B(_06337_),
    .ZN(_08431_));
 XNOR2_X1 _33449_ (.A(_08430_),
    .B(_08431_),
    .ZN(_08432_));
 MUX2_X1 _33450_ (.A(_08428_),
    .B(_08432_),
    .S(_08385_),
    .Z(_00675_));
 XOR2_X1 _33451_ (.A(_17183_),
    .B(_17026_),
    .Z(_08434_));
 XNOR2_X1 _33452_ (.A(_06675_),
    .B(_05457_),
    .ZN(_08435_));
 XOR2_X1 _33453_ (.A(_08435_),
    .B(_08272_),
    .Z(_08436_));
 XNOR2_X1 _33454_ (.A(_08395_),
    .B(_01005_),
    .ZN(_08437_));
 XNOR2_X1 _33455_ (.A(_08436_),
    .B(_08437_),
    .ZN(_08438_));
 MUX2_X1 _33456_ (.A(_08434_),
    .B(_08438_),
    .S(_08385_),
    .Z(_00636_));
 XOR2_X1 _33457_ (.A(_17184_),
    .B(_17027_),
    .Z(_08439_));
 XOR2_X1 _33458_ (.A(_08400_),
    .B(_08395_),
    .Z(_08440_));
 XOR2_X1 _33459_ (.A(_08272_),
    .B(_05831_),
    .Z(_08441_));
 XNOR2_X1 _33460_ (.A(_06555_),
    .B(_15887_),
    .ZN(_08442_));
 XNOR2_X1 _33461_ (.A(_08441_),
    .B(_08442_),
    .ZN(_08444_));
 XNOR2_X1 _33462_ (.A(_08440_),
    .B(_08444_),
    .ZN(_08445_));
 BUF_X4 _33463_ (.A(_09098_),
    .Z(_08446_));
 MUX2_X1 _33464_ (.A(_08439_),
    .B(_08445_),
    .S(_08446_),
    .Z(_00637_));
 XOR2_X1 _33465_ (.A(_17185_),
    .B(_17028_),
    .Z(_08447_));
 XOR2_X1 _33466_ (.A(_07033_),
    .B(_07303_),
    .Z(_08448_));
 XNOR2_X1 _33467_ (.A(_08448_),
    .B(_06464_),
    .ZN(_08449_));
 XNOR2_X1 _33468_ (.A(_06944_),
    .B(_01007_),
    .ZN(_08450_));
 XNOR2_X1 _33469_ (.A(_08450_),
    .B(_06786_),
    .ZN(_08451_));
 XNOR2_X1 _33470_ (.A(_08449_),
    .B(_08451_),
    .ZN(_08452_));
 MUX2_X1 _33471_ (.A(_08447_),
    .B(_08452_),
    .S(_08446_),
    .Z(_00638_));
 XOR2_X1 _33472_ (.A(_17186_),
    .B(_17029_),
    .Z(_08454_));
 XNOR2_X1 _33473_ (.A(_08272_),
    .B(_06869_),
    .ZN(_08455_));
 XNOR2_X1 _33474_ (.A(_07457_),
    .B(_01008_),
    .ZN(_08456_));
 XOR2_X1 _33475_ (.A(_08455_),
    .B(_08456_),
    .Z(_08457_));
 XNOR2_X1 _33476_ (.A(_07537_),
    .B(_07217_),
    .ZN(_08458_));
 XNOR2_X1 _33477_ (.A(_08406_),
    .B(_08458_),
    .ZN(_08459_));
 XNOR2_X1 _33478_ (.A(_08457_),
    .B(_08459_),
    .ZN(_08460_));
 MUX2_X1 _33479_ (.A(_08454_),
    .B(_08460_),
    .S(_08446_),
    .Z(_00639_));
 XOR2_X1 _33480_ (.A(_08272_),
    .B(_07385_),
    .Z(_08461_));
 XNOR2_X1 _33481_ (.A(_08461_),
    .B(_08419_),
    .ZN(_08463_));
 XNOR2_X1 _33482_ (.A(_07729_),
    .B(_01009_),
    .ZN(_08464_));
 XNOR2_X1 _33483_ (.A(_08412_),
    .B(_08464_),
    .ZN(_08465_));
 OR2_X1 _33484_ (.A1(_08463_),
    .A2(_08465_),
    .ZN(_08466_));
 AOI21_X1 _33485_ (.A(_01331_),
    .B1(_08463_),
    .B2(_08465_),
    .ZN(_08467_));
 XNOR2_X1 _33486_ (.A(_17188_),
    .B(_17030_),
    .ZN(_08468_));
 AOI22_X1 _33487_ (.A1(_08466_),
    .A2(_08467_),
    .B1(_01331_),
    .B2(_08468_),
    .ZN(_00640_));
 XOR2_X1 _33488_ (.A(_17189_),
    .B(_17031_),
    .Z(_08469_));
 XNOR2_X1 _33489_ (.A(_08426_),
    .B(_07668_),
    .ZN(_08470_));
 XNOR2_X1 _33490_ (.A(_07600_),
    .B(_01010_),
    .ZN(_08471_));
 XNOR2_X1 _33491_ (.A(_08471_),
    .B(_07859_),
    .ZN(_08473_));
 XNOR2_X1 _33492_ (.A(_08470_),
    .B(_08473_),
    .ZN(_08474_));
 MUX2_X1 _33493_ (.A(_08469_),
    .B(_08474_),
    .S(_08446_),
    .Z(_00641_));
 XOR2_X1 _33494_ (.A(_17190_),
    .B(_17032_),
    .Z(_08475_));
 XNOR2_X1 _33495_ (.A(_07920_),
    .B(_01011_),
    .ZN(_08476_));
 XOR2_X1 _33496_ (.A(_08037_),
    .B(_08476_),
    .Z(_08477_));
 XNOR2_X1 _33497_ (.A(_07805_),
    .B(_08159_),
    .ZN(_08478_));
 XNOR2_X1 _33498_ (.A(_08478_),
    .B(_08382_),
    .ZN(_08479_));
 XNOR2_X1 _33499_ (.A(_08477_),
    .B(_08479_),
    .ZN(_08480_));
 MUX2_X1 _33500_ (.A(_08475_),
    .B(_08480_),
    .S(_08446_),
    .Z(_00642_));
 XOR2_X1 _33501_ (.A(_17191_),
    .B(_17033_),
    .Z(_08482_));
 XNOR2_X1 _33502_ (.A(_06337_),
    .B(_01012_),
    .ZN(_08483_));
 XNOR2_X1 _33503_ (.A(_08483_),
    .B(_08105_),
    .ZN(_08484_));
 XNOR2_X1 _33504_ (.A(_08159_),
    .B(_05570_),
    .ZN(_08485_));
 XNOR2_X1 _33505_ (.A(_08485_),
    .B(_08328_),
    .ZN(_08486_));
 XNOR2_X1 _33506_ (.A(_08484_),
    .B(_08486_),
    .ZN(_08487_));
 MUX2_X1 _33507_ (.A(_08482_),
    .B(_08487_),
    .S(_08446_),
    .Z(_00643_));
 XOR2_X1 _33508_ (.A(_17192_),
    .B(_17035_),
    .Z(_08488_));
 XNOR2_X2 _33509_ (.A(_08273_),
    .B(_05831_),
    .ZN(_08489_));
 XNOR2_X2 _33510_ (.A(_08489_),
    .B(_06099_),
    .ZN(_08490_));
 XNOR2_X2 _33511_ (.A(_08490_),
    .B(_06675_),
    .ZN(_08492_));
 XNOR2_X1 _33512_ (.A(_08492_),
    .B(_01014_),
    .ZN(_08493_));
 MUX2_X1 _33513_ (.A(_08488_),
    .B(_08493_),
    .S(_08446_),
    .Z(_00604_));
 XOR2_X1 _33514_ (.A(_17193_),
    .B(_17036_),
    .Z(_08494_));
 XOR2_X1 _33515_ (.A(_08441_),
    .B(_05571_),
    .Z(_08495_));
 XOR2_X1 _33516_ (.A(_08400_),
    .B(_06464_),
    .Z(_08496_));
 XNOR2_X1 _33517_ (.A(_08495_),
    .B(_08496_),
    .ZN(_08497_));
 INV_X1 _33518_ (.A(_01016_),
    .ZN(_08498_));
 XNOR2_X1 _33519_ (.A(_08497_),
    .B(_08498_),
    .ZN(_08499_));
 MUX2_X1 _33520_ (.A(_08494_),
    .B(_08499_),
    .S(_08446_),
    .Z(_00605_));
 XOR2_X1 _33521_ (.A(_17194_),
    .B(_17037_),
    .Z(_08501_));
 XNOR2_X1 _33522_ (.A(_06557_),
    .B(_01018_),
    .ZN(_08502_));
 XNOR2_X1 _33523_ (.A(_08448_),
    .B(_06869_),
    .ZN(_08503_));
 XNOR2_X1 _33524_ (.A(_08502_),
    .B(_08503_),
    .ZN(_08504_));
 MUX2_X1 _33525_ (.A(_08501_),
    .B(_08504_),
    .S(_08446_),
    .Z(_00606_));
 XOR2_X1 _33526_ (.A(_17195_),
    .B(_17038_),
    .Z(_08505_));
 XNOR2_X1 _33527_ (.A(_08455_),
    .B(_08458_),
    .ZN(_08506_));
 XNOR2_X1 _33528_ (.A(_07385_),
    .B(_01020_),
    .ZN(_08507_));
 XOR2_X1 _33529_ (.A(_07219_),
    .B(_08507_),
    .Z(_08508_));
 XNOR2_X1 _33530_ (.A(_08506_),
    .B(_08508_),
    .ZN(_08509_));
 MUX2_X1 _33531_ (.A(_08505_),
    .B(_08509_),
    .S(_08446_),
    .Z(_00607_));
 XOR2_X1 _33532_ (.A(_17196_),
    .B(_17039_),
    .Z(_08511_));
 XOR2_X1 _33533_ (.A(_07668_),
    .B(_01022_),
    .Z(_08512_));
 XOR2_X1 _33534_ (.A(_07733_),
    .B(_08512_),
    .Z(_08513_));
 XNOR2_X1 _33535_ (.A(_08463_),
    .B(_08513_),
    .ZN(_08514_));
 MUX2_X1 _33536_ (.A(_08511_),
    .B(_08514_),
    .S(_09099_),
    .Z(_00608_));
 XOR2_X1 _33537_ (.A(_17197_),
    .B(_17040_),
    .Z(_08515_));
 XNOR2_X1 _33538_ (.A(_07920_),
    .B(_01024_),
    .ZN(_08516_));
 XNOR2_X1 _33539_ (.A(_08516_),
    .B(_07805_),
    .ZN(_08517_));
 XNOR2_X1 _33540_ (.A(_07731_),
    .B(_08214_),
    .ZN(_08518_));
 XNOR2_X1 _33541_ (.A(_08517_),
    .B(_08518_),
    .ZN(_08520_));
 MUX2_X1 _33542_ (.A(_08515_),
    .B(_08520_),
    .S(_09099_),
    .Z(_00609_));
 XOR2_X1 _33543_ (.A(_17199_),
    .B(_17041_),
    .Z(_08521_));
 XNOR2_X1 _33544_ (.A(_08382_),
    .B(_01026_),
    .ZN(_08522_));
 XNOR2_X1 _33545_ (.A(_08522_),
    .B(_07860_),
    .ZN(_08523_));
 XNOR2_X1 _33546_ (.A(_08105_),
    .B(_08159_),
    .ZN(_08524_));
 XNOR2_X1 _33547_ (.A(_08523_),
    .B(_08524_),
    .ZN(_08525_));
 MUX2_X1 _33548_ (.A(_08521_),
    .B(_08525_),
    .S(_09099_),
    .Z(_00610_));
 XOR2_X1 _33549_ (.A(_17200_),
    .B(_17042_),
    .Z(_08526_));
 XOR2_X1 _33550_ (.A(_08272_),
    .B(_01028_),
    .Z(_08527_));
 XNOR2_X1 _33551_ (.A(_08106_),
    .B(_08527_),
    .ZN(_08529_));
 XOR2_X1 _33552_ (.A(_08328_),
    .B(_06337_),
    .Z(_08530_));
 XNOR2_X1 _33553_ (.A(_08529_),
    .B(_08530_),
    .ZN(_08531_));
 MUX2_X2 _33554_ (.A(_08526_),
    .B(_08531_),
    .S(_09099_),
    .Z(_00611_));
 AND3_X1 _33555_ (.A1(_05158_),
    .A2(_05159_),
    .A3(_01198_),
    .ZN(_00603_));
 XNOR2_X1 _33556_ (.A(_05457_),
    .B(_01014_),
    .ZN(_00884_));
 XNOR2_X1 _33557_ (.A(_06555_),
    .B(_08498_),
    .ZN(_00885_));
 XNOR2_X1 _33558_ (.A(_06944_),
    .B(_03694_),
    .ZN(_00886_));
 XOR2_X1 _33559_ (.A(_07457_),
    .B(_17195_),
    .Z(_00887_));
 XNOR2_X1 _33560_ (.A(_07729_),
    .B(_17196_),
    .ZN(_00888_));
 XOR2_X1 _33561_ (.A(_07859_),
    .B(_01024_),
    .Z(_00889_));
 XOR2_X1 _33562_ (.A(_08037_),
    .B(_01026_),
    .Z(_00890_));
 XNOR2_X1 _33563_ (.A(_05570_),
    .B(_17200_),
    .ZN(_00891_));
 XOR2_X1 _33564_ (.A(_02677_),
    .B(_01042_),
    .Z(_00980_));
 XNOR2_X1 _33565_ (.A(_03015_),
    .B(_05129_),
    .ZN(_00981_));
 XNOR2_X1 _33566_ (.A(_03503_),
    .B(_17226_),
    .ZN(_00982_));
 XNOR2_X1 _33567_ (.A(_03971_),
    .B(_01713_),
    .ZN(_00983_));
 XNOR2_X1 _33568_ (.A(_04246_),
    .B(_01717_),
    .ZN(_00984_));
 XOR2_X1 _33569_ (.A(_04380_),
    .B(_01044_),
    .Z(_00985_));
 XOR2_X1 _33570_ (.A(_04701_),
    .B(_01048_),
    .Z(_00986_));
 XNOR2_X1 _33571_ (.A(_02580_),
    .B(_17232_),
    .ZN(_00987_));
 XOR2_X1 _33572_ (.A(_11857_),
    .B(_01033_),
    .Z(_00940_));
 XNOR2_X1 _33573_ (.A(_12256_),
    .B(_01843_),
    .ZN(_00941_));
 XNOR2_X1 _33574_ (.A(_12661_),
    .B(_17258_),
    .ZN(_00942_));
 XNOR2_X1 _33575_ (.A(_13129_),
    .B(_17259_),
    .ZN(_00943_));
 XNOR2_X1 _33576_ (.A(_13332_),
    .B(_17260_),
    .ZN(_00944_));
 XNOR2_X1 _33577_ (.A(_13508_),
    .B(_01867_),
    .ZN(_00945_));
 XNOR2_X1 _33578_ (.A(_13846_),
    .B(_01036_),
    .ZN(_00946_));
 XNOR2_X1 _33579_ (.A(_11958_),
    .B(_17264_),
    .ZN(_00947_));
 XOR2_X1 _33580_ (.A(_08787_),
    .B(_01054_),
    .Z(_00908_));
 XOR2_X1 _33581_ (.A(_09287_),
    .B(_01055_),
    .Z(_00909_));
 XNOR2_X1 _33582_ (.A(_09684_),
    .B(_17162_),
    .ZN(_00910_));
 XNOR2_X1 _33583_ (.A(_09986_),
    .B(_17163_),
    .ZN(_00911_));
 XNOR2_X1 _33584_ (.A(_10270_),
    .B(_17164_),
    .ZN(_00912_));
 XOR2_X1 _33585_ (.A(_10564_),
    .B(_01056_),
    .Z(_00913_));
 XOR2_X1 _33586_ (.A(_10669_),
    .B(_01057_),
    .Z(_00914_));
 XNOR2_X1 _33587_ (.A(_08887_),
    .B(_17168_),
    .ZN(_00915_));
 XNOR2_X1 _33588_ (.A(_05831_),
    .B(_01005_),
    .ZN(_00876_));
 XNOR2_X1 _33589_ (.A(_06464_),
    .B(_15887_),
    .ZN(_00877_));
 XNOR2_X1 _33590_ (.A(_06869_),
    .B(_17185_),
    .ZN(_00878_));
 XNOR2_X1 _33591_ (.A(_07385_),
    .B(_17186_),
    .ZN(_00879_));
 XNOR2_X1 _33592_ (.A(_07668_),
    .B(_17188_),
    .ZN(_00880_));
 XOR2_X1 _33593_ (.A(_07805_),
    .B(_01010_),
    .Z(_00881_));
 XNOR2_X1 _33594_ (.A(_08105_),
    .B(_16245_),
    .ZN(_00882_));
 XNOR2_X1 _33595_ (.A(_08272_),
    .B(_17191_),
    .ZN(_00883_));
 XNOR2_X1 _33596_ (.A(_02361_),
    .B(_01038_),
    .ZN(_00972_));
 XNOR2_X1 _33597_ (.A(_03116_),
    .B(_05071_),
    .ZN(_00973_));
 XNOR2_X1 _33598_ (.A(_03427_),
    .B(_17217_),
    .ZN(_00974_));
 XNOR2_X1 _33599_ (.A(_03892_),
    .B(_01820_),
    .ZN(_00975_));
 XNOR2_X1 _33600_ (.A(_04178_),
    .B(_17220_),
    .ZN(_00976_));
 XNOR2_X1 _33601_ (.A(_04442_),
    .B(_05102_),
    .ZN(_00977_));
 XOR2_X1 _33602_ (.A(_04635_),
    .B(_01041_),
    .Z(_00978_));
 XNOR2_X1 _33603_ (.A(_05005_),
    .B(_17223_),
    .ZN(_00979_));
 XOR2_X1 _33604_ (.A(_11387_),
    .B(_01029_),
    .Z(_00932_));
 XOR2_X1 _33605_ (.A(_12357_),
    .B(_01030_),
    .Z(_00933_));
 XNOR2_X1 _33606_ (.A(_12736_),
    .B(_17249_),
    .ZN(_00934_));
 XNOR2_X1 _33607_ (.A(_13058_),
    .B(_17250_),
    .ZN(_00935_));
 XNOR2_X1 _33608_ (.A(_13389_),
    .B(_17252_),
    .ZN(_00936_));
 XOR2_X1 _33609_ (.A(_13568_),
    .B(_01031_),
    .Z(_00937_));
 XOR2_X1 _33610_ (.A(_13797_),
    .B(_01032_),
    .Z(_00938_));
 XNOR2_X1 _33611_ (.A(_13960_),
    .B(_17255_),
    .ZN(_00939_));
 XOR2_X1 _33612_ (.A(_08560_),
    .B(_01050_),
    .Z(_00900_));
 XOR2_X1 _33613_ (.A(_09213_),
    .B(_01051_),
    .Z(_00901_));
 XNOR2_X1 _33614_ (.A(_09616_),
    .B(_11068_),
    .ZN(_00902_));
 XNOR2_X1 _33615_ (.A(_10065_),
    .B(_17154_),
    .ZN(_00903_));
 XNOR2_X1 _33616_ (.A(_10327_),
    .B(_17156_),
    .ZN(_00904_));
 XOR2_X1 _33617_ (.A(_10514_),
    .B(_01052_),
    .Z(_00905_));
 XOR2_X1 _33618_ (.A(_10717_),
    .B(_01053_),
    .Z(_00906_));
 XNOR2_X1 _33619_ (.A(_10886_),
    .B(_17159_),
    .ZN(_00907_));
 XNOR2_X1 _33620_ (.A(_06099_),
    .B(_17206_),
    .ZN(_00868_));
 XNOR2_X1 _33621_ (.A(_06786_),
    .B(_17207_),
    .ZN(_00869_));
 XNOR2_X1 _33622_ (.A(_07033_),
    .B(_17177_),
    .ZN(_00870_));
 XNOR2_X1 _33623_ (.A(_07217_),
    .B(_17178_),
    .ZN(_00871_));
 XNOR2_X1 _33624_ (.A(_07600_),
    .B(_17179_),
    .ZN(_00872_));
 XOR2_X1 _33625_ (.A(_07920_),
    .B(_17180_),
    .Z(_00873_));
 XOR2_X1 _33626_ (.A(_08159_),
    .B(_17181_),
    .Z(_00874_));
 XNOR2_X1 _33627_ (.A(_08328_),
    .B(_17182_),
    .ZN(_00875_));
 XNOR2_X1 _33628_ (.A(_02128_),
    .B(_17238_),
    .ZN(_00956_));
 XNOR2_X1 _33629_ (.A(_03212_),
    .B(_17239_),
    .ZN(_00957_));
 XNOR2_X1 _33630_ (.A(_03577_),
    .B(_05030_),
    .ZN(_00958_));
 XNOR2_X1 _33631_ (.A(_03805_),
    .B(_17210_),
    .ZN(_00959_));
 XNOR2_X1 _33632_ (.A(_04108_),
    .B(_17211_),
    .ZN(_00960_));
 XNOR2_X1 _33633_ (.A(_04513_),
    .B(_05048_),
    .ZN(_00961_));
 XNOR2_X1 _33634_ (.A(_04771_),
    .B(_17213_),
    .ZN(_00962_));
 XNOR2_X1 _33635_ (.A(_04950_),
    .B(_17214_),
    .ZN(_00963_));
 XNOR2_X1 _33636_ (.A(_11624_),
    .B(_17270_),
    .ZN(_00924_));
 XNOR2_X1 _33637_ (.A(_12472_),
    .B(_17271_),
    .ZN(_00925_));
 XNOR2_X1 _33638_ (.A(_12823_),
    .B(_17241_),
    .ZN(_00926_));
 XNOR2_X1 _33639_ (.A(_12982_),
    .B(_17242_),
    .ZN(_00927_));
 XNOR2_X1 _33640_ (.A(_13444_),
    .B(_01806_),
    .ZN(_00928_));
 XNOR2_X1 _33641_ (.A(_13685_),
    .B(_17244_),
    .ZN(_00929_));
 XNOR2_X1 _33642_ (.A(_13743_),
    .B(_17245_),
    .ZN(_00930_));
 XNOR2_X1 _33643_ (.A(_14014_),
    .B(_17246_),
    .ZN(_00931_));
 XNOR2_X1 _33644_ (.A(_06567_),
    .B(_10997_),
    .ZN(_00892_));
 XNOR2_X1 _33645_ (.A(_09528_),
    .B(_11004_),
    .ZN(_00893_));
 XNOR2_X1 _33646_ (.A(_09763_),
    .B(_17145_),
    .ZN(_00894_));
 XNOR2_X1 _33647_ (.A(_10148_),
    .B(_17146_),
    .ZN(_00895_));
 XNOR2_X1 _33648_ (.A(_10212_),
    .B(_17147_),
    .ZN(_00896_));
 XNOR2_X1 _33649_ (.A(_10465_),
    .B(_17148_),
    .ZN(_00897_));
 XNOR2_X1 _33650_ (.A(_10777_),
    .B(_17149_),
    .ZN(_00898_));
 XNOR2_X1 _33651_ (.A(_10934_),
    .B(_17150_),
    .ZN(_00899_));
 XNOR2_X1 _33652_ (.A(_06675_),
    .B(_17176_),
    .ZN(_00860_));
 XOR2_X1 _33653_ (.A(_07126_),
    .B(_17187_),
    .Z(_00861_));
 XOR2_X1 _33654_ (.A(_07303_),
    .B(_17198_),
    .Z(_00862_));
 XNOR2_X1 _33655_ (.A(_07537_),
    .B(_17201_),
    .ZN(_00863_));
 XNOR2_X1 _33656_ (.A(_07979_),
    .B(_17202_),
    .ZN(_00864_));
 XOR2_X1 _33657_ (.A(_08214_),
    .B(_17203_),
    .Z(_00865_));
 XNOR2_X1 _33658_ (.A(_08382_),
    .B(_17204_),
    .ZN(_00866_));
 XNOR2_X1 _33659_ (.A(_06337_),
    .B(_17205_),
    .ZN(_00867_));
 XNOR2_X1 _33660_ (.A(_03316_),
    .B(_02909_),
    .ZN(_00948_));
 XOR2_X1 _33661_ (.A(_03671_),
    .B(_17219_),
    .Z(_00949_));
 XOR2_X1 _33662_ (.A(_04045_),
    .B(_17230_),
    .Z(_00950_));
 XNOR2_X1 _33663_ (.A(_04318_),
    .B(_17233_),
    .ZN(_00951_));
 XNOR2_X1 _33664_ (.A(_04574_),
    .B(_17234_),
    .ZN(_00952_));
 XOR2_X1 _33665_ (.A(_04830_),
    .B(_17235_),
    .Z(_00953_));
 XNOR2_X1 _33666_ (.A(_04893_),
    .B(_17236_),
    .ZN(_00954_));
 XOR2_X1 _33667_ (.A(_02907_),
    .B(_17237_),
    .Z(_00955_));
 XNOR2_X1 _33668_ (.A(_12583_),
    .B(_17240_),
    .ZN(_00916_));
 XNOR2_X1 _33669_ (.A(_12904_),
    .B(_01782_),
    .ZN(_00917_));
 XNOR2_X1 _33670_ (.A(_13199_),
    .B(_01785_),
    .ZN(_00918_));
 XNOR2_X1 _33671_ (.A(_13275_),
    .B(_17265_),
    .ZN(_00919_));
 XNOR2_X1 _33672_ (.A(_13621_),
    .B(_17266_),
    .ZN(_00920_));
 XNOR2_X1 _33673_ (.A(_13903_),
    .B(_17267_),
    .ZN(_00921_));
 XNOR2_X1 _33674_ (.A(_14064_),
    .B(_13905_),
    .ZN(_00922_));
 XNOR2_X1 _33675_ (.A(_12175_),
    .B(_17269_),
    .ZN(_00923_));
 XNOR2_X1 _33676_ (.A(_09412_),
    .B(_04132_),
    .ZN(_00964_));
 XNOR2_X1 _33677_ (.A(_09837_),
    .B(_09101_),
    .ZN(_00965_));
 XNOR2_X1 _33678_ (.A(_09914_),
    .B(_17166_),
    .ZN(_00966_));
 XNOR2_X1 _33679_ (.A(_10401_),
    .B(_17169_),
    .ZN(_00967_));
 XNOR2_X1 _33680_ (.A(_10616_),
    .B(_17170_),
    .ZN(_00968_));
 XNOR2_X1 _33681_ (.A(_10837_),
    .B(_14851_),
    .ZN(_00969_));
 XNOR2_X1 _33682_ (.A(_10989_),
    .B(_17172_),
    .ZN(_00970_));
 XNOR2_X1 _33683_ (.A(_09093_),
    .B(_17173_),
    .ZN(_00971_));
 BUF_X1 _33684_ (.A(ld),
    .Z(_01330_));
 BUF_X1 _33685_ (.A(\u0.r0.rcnt[0] ),
    .Z(_17140_));
 BUF_X1 _33686_ (.A(\u0.r0.rcnt[1] ),
    .Z(_17141_));
 BUF_X1 _33687_ (.A(\u0.r0.rcnt[2] ),
    .Z(_17142_));
 BUF_X1 _33688_ (.A(\u0.r0.rcnt[3] ),
    .Z(_17143_));
 BUF_X1 _33689_ (.A(_01186_),
    .Z(_00587_));
 BUF_X1 _33690_ (.A(_01187_),
    .Z(_00588_));
 BUF_X1 _33691_ (.A(_01188_),
    .Z(_00589_));
 BUF_X1 _33692_ (.A(_01189_),
    .Z(_00590_));
 BUF_X1 _33693_ (.A(_01190_),
    .Z(_00591_));
 BUF_X1 _33694_ (.A(_01191_),
    .Z(_00592_));
 BUF_X1 _33695_ (.A(_01192_),
    .Z(_00593_));
 BUF_X1 _33696_ (.A(_01193_),
    .Z(_00594_));
 BUF_X1 _33697_ (.A(_01194_),
    .Z(_00595_));
 BUF_X1 _33698_ (.A(_01195_),
    .Z(_00596_));
 BUF_X1 _33699_ (.A(_01196_),
    .Z(_00597_));
 BUF_X1 _33700_ (.A(_01197_),
    .Z(_00598_));
 BUF_X1 _33701_ (.A(\sa03[0] ),
    .Z(_16780_));
 BUF_X1 _33702_ (.A(\sa03[1] ),
    .Z(_16781_));
 BUF_X1 _33703_ (.A(\sa03[3] ),
    .Z(_16783_));
 BUF_X1 _33704_ (.A(\sa03[2] ),
    .Z(_16782_));
 BUF_X1 _33705_ (.A(\sa03[5] ),
    .Z(_16785_));
 BUF_X1 _33706_ (.A(\sa03[4] ),
    .Z(_16784_));
 BUF_X1 _33707_ (.A(\sa03[7] ),
    .Z(_16787_));
 BUF_X1 _33708_ (.A(\sa03[6] ),
    .Z(_16786_));
 BUF_X1 _33709_ (.A(\sa10[5] ),
    .Z(_16793_));
 BUF_X1 _33710_ (.A(\sa10[4] ),
    .Z(_16792_));
 BUF_X1 _33711_ (.A(\sa10[7] ),
    .Z(_16795_));
 BUF_X1 _33712_ (.A(\sa10[6] ),
    .Z(_16794_));
 BUF_X1 _33713_ (.A(\sa10[1] ),
    .Z(_16789_));
 BUF_X1 _33714_ (.A(\sa10[0] ),
    .Z(_16788_));
 BUF_X1 _33715_ (.A(\sa10[2] ),
    .Z(_16790_));
 BUF_X1 _33716_ (.A(\sa10[3] ),
    .Z(_16791_));
 BUF_X1 _33717_ (.A(\sa21[5] ),
    .Z(_16833_));
 BUF_X1 _33718_ (.A(\sa21[4] ),
    .Z(_16832_));
 BUF_X1 _33719_ (.A(\sa21[7] ),
    .Z(_16835_));
 BUF_X1 _33720_ (.A(\sa21[6] ),
    .Z(_16834_));
 BUF_X1 _33721_ (.A(\sa21[1] ),
    .Z(_16829_));
 BUF_X1 _33722_ (.A(\sa21[0] ),
    .Z(_16828_));
 BUF_X1 _33723_ (.A(\sa21[2] ),
    .Z(_16830_));
 BUF_X1 _33724_ (.A(\sa21[3] ),
    .Z(_16831_));
 BUF_X1 _33725_ (.A(\sa32[0] ),
    .Z(_16868_));
 BUF_X1 _33726_ (.A(\sa32[1] ),
    .Z(_16869_));
 BUF_X1 _33727_ (.A(\sa32[3] ),
    .Z(_16871_));
 BUF_X1 _33728_ (.A(\sa32[2] ),
    .Z(_16870_));
 BUF_X1 _33729_ (.A(\sa32[5] ),
    .Z(_16873_));
 BUF_X1 _33730_ (.A(\sa32[4] ),
    .Z(_16872_));
 BUF_X1 _33731_ (.A(\sa32[7] ),
    .Z(_16875_));
 BUF_X1 _33732_ (.A(\sa32[6] ),
    .Z(_16874_));
 BUF_X1 _33733_ (.A(\u0.tmp_w[0] ),
    .Z(_17144_));
 BUF_X1 _33734_ (.A(\text_in_r[0] ),
    .Z(_17012_));
 BUF_X1 _33735_ (.A(ld_r),
    .Z(_01331_));
 BUF_X1 _33736_ (.A(_00724_),
    .Z(_00125_));
 BUF_X1 _33737_ (.A(\u0.tmp_w[1] ),
    .Z(_17155_));
 BUF_X1 _33738_ (.A(\text_in_r[1] ),
    .Z(_17051_));
 BUF_X1 _33739_ (.A(_00725_),
    .Z(_00126_));
 BUF_X1 _33740_ (.A(\u0.tmp_w[2] ),
    .Z(_17166_));
 BUF_X1 _33741_ (.A(\text_in_r[2] ),
    .Z(_17062_));
 BUF_X1 _33742_ (.A(_00726_),
    .Z(_00127_));
 BUF_X1 _33743_ (.A(\u0.tmp_w[3] ),
    .Z(_17169_));
 BUF_X1 _33744_ (.A(\text_in_r[3] ),
    .Z(_17073_));
 BUF_X1 _33745_ (.A(_00727_),
    .Z(_00128_));
 BUF_X1 _33746_ (.A(\u0.tmp_w[4] ),
    .Z(_17170_));
 BUF_X1 _33747_ (.A(\text_in_r[4] ),
    .Z(_17084_));
 BUF_X1 _33748_ (.A(_00728_),
    .Z(_00129_));
 BUF_X1 _33749_ (.A(\u0.tmp_w[5] ),
    .Z(_17171_));
 BUF_X1 _33750_ (.A(\text_in_r[5] ),
    .Z(_17095_));
 BUF_X1 _33751_ (.A(_00729_),
    .Z(_00130_));
 BUF_X1 _33752_ (.A(\u0.tmp_w[6] ),
    .Z(_17172_));
 BUF_X1 _33753_ (.A(\text_in_r[6] ),
    .Z(_17106_));
 BUF_X1 _33754_ (.A(_00730_),
    .Z(_00131_));
 BUF_X1 _33755_ (.A(\u0.tmp_w[7] ),
    .Z(_17173_));
 BUF_X1 _33756_ (.A(\text_in_r[7] ),
    .Z(_17117_));
 BUF_X1 _33757_ (.A(_00731_),
    .Z(_00132_));
 BUF_X1 _33758_ (.A(_00450_),
    .Z(_01049_));
 BUF_X1 _33759_ (.A(\text_in_r[8] ),
    .Z(_17128_));
 BUF_X1 _33760_ (.A(\u0.tmp_w[8] ),
    .Z(_17174_));
 BUF_X1 _33761_ (.A(_00692_),
    .Z(_00093_));
 BUF_X1 _33762_ (.A(\u0.tmp_w[9] ),
    .Z(_17175_));
 BUF_X1 _33763_ (.A(\text_in_r[9] ),
    .Z(_17139_));
 BUF_X1 _33764_ (.A(_00693_),
    .Z(_00094_));
 BUF_X1 _33765_ (.A(\u0.tmp_w[10] ),
    .Z(_17145_));
 BUF_X1 _33766_ (.A(\text_in_r[10] ),
    .Z(_17023_));
 BUF_X1 _33767_ (.A(_00694_),
    .Z(_00095_));
 BUF_X1 _33768_ (.A(\u0.tmp_w[11] ),
    .Z(_17146_));
 BUF_X1 _33769_ (.A(\text_in_r[11] ),
    .Z(_17034_));
 BUF_X1 _33770_ (.A(_00695_),
    .Z(_00096_));
 BUF_X1 _33771_ (.A(\u0.tmp_w[12] ),
    .Z(_17147_));
 BUF_X1 _33772_ (.A(\text_in_r[12] ),
    .Z(_17043_));
 BUF_X1 _33773_ (.A(_00696_),
    .Z(_00097_));
 BUF_X1 _33774_ (.A(\u0.tmp_w[13] ),
    .Z(_17148_));
 BUF_X1 _33775_ (.A(\text_in_r[13] ),
    .Z(_17044_));
 BUF_X1 _33776_ (.A(_00697_),
    .Z(_00098_));
 BUF_X1 _33777_ (.A(\u0.tmp_w[14] ),
    .Z(_17149_));
 BUF_X1 _33778_ (.A(\text_in_r[14] ),
    .Z(_17045_));
 BUF_X1 _33779_ (.A(_00698_),
    .Z(_00099_));
 BUF_X1 _33780_ (.A(\u0.tmp_w[15] ),
    .Z(_17150_));
 BUF_X1 _33781_ (.A(\text_in_r[15] ),
    .Z(_17046_));
 BUF_X1 _33782_ (.A(_00699_),
    .Z(_00100_));
 BUF_X1 _33783_ (.A(_00451_),
    .Z(_01050_));
 BUF_X1 _33784_ (.A(\text_in_r[16] ),
    .Z(_17047_));
 BUF_X1 _33785_ (.A(\u0.tmp_w[16] ),
    .Z(_17151_));
 BUF_X1 _33786_ (.A(_00660_),
    .Z(_00061_));
 BUF_X1 _33787_ (.A(_00452_),
    .Z(_01051_));
 BUF_X1 _33788_ (.A(\text_in_r[17] ),
    .Z(_17048_));
 BUF_X1 _33789_ (.A(\u0.tmp_w[17] ),
    .Z(_17152_));
 BUF_X1 _33790_ (.A(_00661_),
    .Z(_00062_));
 BUF_X1 _33791_ (.A(\u0.tmp_w[18] ),
    .Z(_17153_));
 BUF_X1 _33792_ (.A(\text_in_r[18] ),
    .Z(_17049_));
 BUF_X1 _33793_ (.A(_00662_),
    .Z(_00063_));
 BUF_X1 _33794_ (.A(\u0.tmp_w[19] ),
    .Z(_17154_));
 BUF_X1 _33795_ (.A(\text_in_r[19] ),
    .Z(_17050_));
 BUF_X1 _33796_ (.A(_00663_),
    .Z(_00064_));
 BUF_X1 _33797_ (.A(\u0.tmp_w[20] ),
    .Z(_17156_));
 BUF_X1 _33798_ (.A(\text_in_r[20] ),
    .Z(_17052_));
 BUF_X1 _33799_ (.A(_00664_),
    .Z(_00065_));
 BUF_X1 _33800_ (.A(_00453_),
    .Z(_01052_));
 BUF_X1 _33801_ (.A(\text_in_r[21] ),
    .Z(_17053_));
 BUF_X1 _33802_ (.A(\u0.tmp_w[21] ),
    .Z(_17157_));
 BUF_X1 _33803_ (.A(_00665_),
    .Z(_00066_));
 BUF_X1 _33804_ (.A(_00454_),
    .Z(_01053_));
 BUF_X1 _33805_ (.A(\text_in_r[22] ),
    .Z(_17054_));
 BUF_X1 _33806_ (.A(\u0.tmp_w[22] ),
    .Z(_17158_));
 BUF_X1 _33807_ (.A(_00666_),
    .Z(_00067_));
 BUF_X1 _33808_ (.A(\u0.tmp_w[23] ),
    .Z(_17159_));
 BUF_X1 _33809_ (.A(\text_in_r[23] ),
    .Z(_17055_));
 BUF_X1 _33810_ (.A(_00667_),
    .Z(_00068_));
 BUF_X1 _33811_ (.A(_00455_),
    .Z(_01054_));
 BUF_X1 _33812_ (.A(\text_in_r[24] ),
    .Z(_17056_));
 BUF_X1 _33813_ (.A(\u0.tmp_w[24] ),
    .Z(_17160_));
 BUF_X1 _33814_ (.A(_00628_),
    .Z(_00029_));
 BUF_X1 _33815_ (.A(_00456_),
    .Z(_01055_));
 BUF_X1 _33816_ (.A(\text_in_r[25] ),
    .Z(_17057_));
 BUF_X1 _33817_ (.A(\u0.tmp_w[25] ),
    .Z(_17161_));
 BUF_X1 _33818_ (.A(_00629_),
    .Z(_00030_));
 BUF_X1 _33819_ (.A(\u0.tmp_w[26] ),
    .Z(_17162_));
 BUF_X1 _33820_ (.A(\text_in_r[26] ),
    .Z(_17058_));
 BUF_X1 _33821_ (.A(_00630_),
    .Z(_00031_));
 BUF_X1 _33822_ (.A(\u0.tmp_w[27] ),
    .Z(_17163_));
 BUF_X1 _33823_ (.A(\text_in_r[27] ),
    .Z(_17059_));
 BUF_X1 _33824_ (.A(_00631_),
    .Z(_00032_));
 BUF_X1 _33825_ (.A(\u0.tmp_w[28] ),
    .Z(_17164_));
 BUF_X1 _33826_ (.A(\text_in_r[28] ),
    .Z(_17060_));
 BUF_X1 _33827_ (.A(_00632_),
    .Z(_00033_));
 BUF_X1 _33828_ (.A(_00457_),
    .Z(_01056_));
 BUF_X1 _33829_ (.A(\text_in_r[29] ),
    .Z(_17061_));
 BUF_X1 _33830_ (.A(\u0.tmp_w[29] ),
    .Z(_17165_));
 BUF_X1 _33831_ (.A(_00633_),
    .Z(_00034_));
 BUF_X1 _33832_ (.A(_00458_),
    .Z(_01057_));
 BUF_X1 _33833_ (.A(\text_in_r[30] ),
    .Z(_17063_));
 BUF_X1 _33834_ (.A(\u0.tmp_w[30] ),
    .Z(_17167_));
 BUF_X1 _33835_ (.A(_00634_),
    .Z(_00035_));
 BUF_X1 _33836_ (.A(\u0.tmp_w[31] ),
    .Z(_17168_));
 BUF_X1 _33837_ (.A(\text_in_r[31] ),
    .Z(_17064_));
 BUF_X1 _33838_ (.A(_00635_),
    .Z(_00036_));
 BUF_X1 _33839_ (.A(\sa02[0] ),
    .Z(_16772_));
 BUF_X1 _33840_ (.A(\sa02[1] ),
    .Z(_16773_));
 BUF_X1 _33841_ (.A(\sa02[3] ),
    .Z(_16775_));
 BUF_X1 _33842_ (.A(\sa02[2] ),
    .Z(_16774_));
 BUF_X1 _33843_ (.A(\sa02[5] ),
    .Z(_16777_));
 BUF_X1 _33844_ (.A(\sa02[4] ),
    .Z(_16776_));
 BUF_X1 _33845_ (.A(\sa02[7] ),
    .Z(_16779_));
 BUF_X1 _33846_ (.A(\sa02[6] ),
    .Z(_16778_));
 BUF_X1 _33847_ (.A(\sa13[5] ),
    .Z(_16817_));
 BUF_X1 _33848_ (.A(\sa13[4] ),
    .Z(_16816_));
 BUF_X1 _33849_ (.A(\sa13[7] ),
    .Z(_16819_));
 BUF_X1 _33850_ (.A(\sa13[6] ),
    .Z(_16818_));
 BUF_X1 _33851_ (.A(\sa13[1] ),
    .Z(_16813_));
 BUF_X1 _33852_ (.A(\sa13[0] ),
    .Z(_16812_));
 BUF_X1 _33853_ (.A(\sa13[2] ),
    .Z(_16814_));
 BUF_X1 _33854_ (.A(\sa13[3] ),
    .Z(_16815_));
 BUF_X1 _33855_ (.A(\sa20[5] ),
    .Z(_16825_));
 BUF_X1 _33856_ (.A(\sa20[4] ),
    .Z(_16824_));
 BUF_X1 _33857_ (.A(\sa20[7] ),
    .Z(_16827_));
 BUF_X1 _33858_ (.A(\sa20[6] ),
    .Z(_16826_));
 BUF_X1 _33859_ (.A(\sa20[1] ),
    .Z(_16821_));
 BUF_X1 _33860_ (.A(\sa20[0] ),
    .Z(_16820_));
 BUF_X1 _33861_ (.A(\sa20[2] ),
    .Z(_16822_));
 BUF_X1 _33862_ (.A(\sa20[3] ),
    .Z(_16823_));
 BUF_X1 _33863_ (.A(\sa31[0] ),
    .Z(_16860_));
 BUF_X1 _33864_ (.A(\sa31[1] ),
    .Z(_16861_));
 BUF_X1 _33865_ (.A(\sa31[3] ),
    .Z(_16863_));
 BUF_X1 _33866_ (.A(\sa31[2] ),
    .Z(_16862_));
 BUF_X1 _33867_ (.A(\sa31[5] ),
    .Z(_16865_));
 BUF_X1 _33868_ (.A(\sa31[4] ),
    .Z(_16864_));
 BUF_X1 _33869_ (.A(\sa31[7] ),
    .Z(_16867_));
 BUF_X1 _33870_ (.A(\sa31[6] ),
    .Z(_16866_));
 BUF_X1 _33871_ (.A(\u0.w[2][0] ),
    .Z(_17240_));
 BUF_X1 _33872_ (.A(\text_in_r[32] ),
    .Z(_17065_));
 BUF_X1 _33873_ (.A(_00716_),
    .Z(_00117_));
 BUF_X1 _33874_ (.A(\u0.w[2][1] ),
    .Z(_17251_));
 BUF_X1 _33875_ (.A(\text_in_r[33] ),
    .Z(_17066_));
 BUF_X1 _33876_ (.A(_00717_),
    .Z(_00118_));
 BUF_X1 _33877_ (.A(\u0.w[2][2] ),
    .Z(_17262_));
 BUF_X1 _33878_ (.A(\text_in_r[34] ),
    .Z(_17067_));
 BUF_X1 _33879_ (.A(_00718_),
    .Z(_00119_));
 BUF_X1 _33880_ (.A(\u0.w[2][3] ),
    .Z(_17265_));
 BUF_X1 _33881_ (.A(\text_in_r[35] ),
    .Z(_17068_));
 BUF_X1 _33882_ (.A(_00719_),
    .Z(_00120_));
 BUF_X1 _33883_ (.A(\u0.w[2][4] ),
    .Z(_17266_));
 BUF_X1 _33884_ (.A(\text_in_r[36] ),
    .Z(_17069_));
 BUF_X1 _33885_ (.A(_00720_),
    .Z(_00121_));
 BUF_X1 _33886_ (.A(\u0.w[2][5] ),
    .Z(_17267_));
 BUF_X1 _33887_ (.A(\text_in_r[37] ),
    .Z(_17070_));
 BUF_X1 _33888_ (.A(_00721_),
    .Z(_00122_));
 BUF_X1 _33889_ (.A(\u0.w[2][6] ),
    .Z(_17268_));
 BUF_X1 _33890_ (.A(\text_in_r[38] ),
    .Z(_17071_));
 BUF_X1 _33891_ (.A(_00722_),
    .Z(_00123_));
 BUF_X1 _33892_ (.A(\u0.w[2][7] ),
    .Z(_17269_));
 BUF_X1 _33893_ (.A(\text_in_r[39] ),
    .Z(_17072_));
 BUF_X1 _33894_ (.A(_00723_),
    .Z(_00124_));
 BUF_X1 _33895_ (.A(_00389_),
    .Z(_00988_));
 BUF_X1 _33896_ (.A(key[96]),
    .Z(_01325_));
 BUF_X1 _33897_ (.A(_01058_),
    .Z(_00459_));
 BUF_X1 _33898_ (.A(_00390_),
    .Z(_00989_));
 BUF_X1 _33899_ (.A(key[97]),
    .Z(_01326_));
 BUF_X1 _33900_ (.A(_01069_),
    .Z(_00470_));
 BUF_X1 _33901_ (.A(_00391_),
    .Z(_00990_));
 BUF_X1 _33902_ (.A(\u0.w[2][8] ),
    .Z(_17270_));
 BUF_X1 _33903_ (.A(\text_in_r[40] ),
    .Z(_17074_));
 BUF_X1 _33904_ (.A(_00684_),
    .Z(_00085_));
 BUF_X1 _33905_ (.A(_00392_),
    .Z(_00991_));
 BUF_X1 _33906_ (.A(key[98]),
    .Z(_01327_));
 BUF_X1 _33907_ (.A(_01080_),
    .Z(_00481_));
 BUF_X1 _33908_ (.A(_00393_),
    .Z(_00992_));
 BUF_X1 _33909_ (.A(key[99]),
    .Z(_01328_));
 BUF_X1 _33910_ (.A(_01083_),
    .Z(_00484_));
 BUF_X1 _33911_ (.A(_00394_),
    .Z(_00993_));
 BUF_X1 _33912_ (.A(key[100]),
    .Z(_01203_));
 BUF_X1 _33913_ (.A(_01084_),
    .Z(_00485_));
 BUF_X1 _33914_ (.A(_00395_),
    .Z(_00994_));
 BUF_X1 _33915_ (.A(key[101]),
    .Z(_01204_));
 BUF_X1 _33916_ (.A(_01085_),
    .Z(_00486_));
 BUF_X1 _33917_ (.A(_00396_),
    .Z(_00995_));
 BUF_X1 _33918_ (.A(key[102]),
    .Z(_01205_));
 BUF_X1 _33919_ (.A(_01086_),
    .Z(_00487_));
 BUF_X1 _33920_ (.A(_00397_),
    .Z(_00996_));
 BUF_X1 _33921_ (.A(key[103]),
    .Z(_01206_));
 BUF_X1 _33922_ (.A(_01087_),
    .Z(_00488_));
 BUF_X1 _33923_ (.A(_00398_),
    .Z(_00997_));
 BUF_X1 _33924_ (.A(key[104]),
    .Z(_01207_));
 BUF_X1 _33925_ (.A(_01088_),
    .Z(_00489_));
 BUF_X1 _33926_ (.A(_00399_),
    .Z(_00998_));
 BUF_X1 _33927_ (.A(key[105]),
    .Z(_01208_));
 BUF_X1 _33928_ (.A(_01089_),
    .Z(_00490_));
 BUF_X1 _33929_ (.A(_00400_),
    .Z(_00999_));
 BUF_X1 _33930_ (.A(key[106]),
    .Z(_01209_));
 BUF_X1 _33931_ (.A(_01059_),
    .Z(_00460_));
 BUF_X1 _33932_ (.A(_00401_),
    .Z(_01000_));
 BUF_X1 _33933_ (.A(key[107]),
    .Z(_01210_));
 BUF_X1 _33934_ (.A(_01060_),
    .Z(_00461_));
 BUF_X1 _33935_ (.A(\u0.w[2][9] ),
    .Z(_17271_));
 BUF_X1 _33936_ (.A(\text_in_r[41] ),
    .Z(_17075_));
 BUF_X1 _33937_ (.A(_00685_),
    .Z(_00086_));
 BUF_X1 _33938_ (.A(_00402_),
    .Z(_01001_));
 BUF_X1 _33939_ (.A(key[108]),
    .Z(_01211_));
 BUF_X1 _33940_ (.A(_01061_),
    .Z(_00462_));
 BUF_X1 _33941_ (.A(_00403_),
    .Z(_01002_));
 BUF_X1 _33942_ (.A(key[109]),
    .Z(_01212_));
 BUF_X1 _33943_ (.A(_01062_),
    .Z(_00463_));
 BUF_X1 _33944_ (.A(_00404_),
    .Z(_01003_));
 BUF_X1 _33945_ (.A(key[110]),
    .Z(_01214_));
 BUF_X1 _33946_ (.A(_01063_),
    .Z(_00464_));
 BUF_X1 _33947_ (.A(_00405_),
    .Z(_01004_));
 BUF_X1 _33948_ (.A(key[111]),
    .Z(_01215_));
 BUF_X1 _33949_ (.A(_01064_),
    .Z(_00465_));
 BUF_X1 _33950_ (.A(_00406_),
    .Z(_01005_));
 BUF_X1 _33951_ (.A(key[112]),
    .Z(_01216_));
 BUF_X1 _33952_ (.A(_01065_),
    .Z(_00466_));
 BUF_X1 _33953_ (.A(_00407_),
    .Z(_01006_));
 BUF_X1 _33954_ (.A(key[113]),
    .Z(_01217_));
 BUF_X1 _33955_ (.A(_01066_),
    .Z(_00467_));
 BUF_X1 _33956_ (.A(_00408_),
    .Z(_01007_));
 BUF_X1 _33957_ (.A(key[114]),
    .Z(_01218_));
 BUF_X1 _33958_ (.A(_01067_),
    .Z(_00468_));
 BUF_X1 _33959_ (.A(_00409_),
    .Z(_01008_));
 BUF_X1 _33960_ (.A(key[115]),
    .Z(_01219_));
 BUF_X1 _33961_ (.A(_01068_),
    .Z(_00469_));
 BUF_X1 _33962_ (.A(_00410_),
    .Z(_01009_));
 BUF_X1 _33963_ (.A(key[116]),
    .Z(_01220_));
 BUF_X1 _33964_ (.A(_01070_),
    .Z(_00471_));
 BUF_X1 _33965_ (.A(_00411_),
    .Z(_01010_));
 BUF_X1 _33966_ (.A(key[117]),
    .Z(_01221_));
 BUF_X1 _33967_ (.A(_01071_),
    .Z(_00472_));
 BUF_X1 _33968_ (.A(\u0.w[2][10] ),
    .Z(_17241_));
 BUF_X1 _33969_ (.A(\text_in_r[42] ),
    .Z(_17076_));
 BUF_X1 _33970_ (.A(_00686_),
    .Z(_00087_));
 BUF_X1 _33971_ (.A(_00412_),
    .Z(_01011_));
 BUF_X1 _33972_ (.A(key[118]),
    .Z(_01222_));
 BUF_X1 _33973_ (.A(_01072_),
    .Z(_00473_));
 BUF_X1 _33974_ (.A(_00413_),
    .Z(_01012_));
 BUF_X1 _33975_ (.A(key[119]),
    .Z(_01223_));
 BUF_X1 _33976_ (.A(_01073_),
    .Z(_00474_));
 BUF_X1 _33977_ (.A(_00415_),
    .Z(_01014_));
 BUF_X1 _33978_ (.A(_00414_),
    .Z(_01013_));
 BUF_X1 _33979_ (.A(key[120]),
    .Z(_01225_));
 BUF_X1 _33980_ (.A(_01074_),
    .Z(_00475_));
 BUF_X1 _33981_ (.A(_00417_),
    .Z(_01016_));
 BUF_X1 _33982_ (.A(_00416_),
    .Z(_01015_));
 BUF_X1 _33983_ (.A(key[121]),
    .Z(_01226_));
 BUF_X1 _33984_ (.A(_01075_),
    .Z(_00476_));
 BUF_X1 _33985_ (.A(_00419_),
    .Z(_01018_));
 BUF_X1 _33986_ (.A(_00418_),
    .Z(_01017_));
 BUF_X1 _33987_ (.A(key[122]),
    .Z(_01227_));
 BUF_X1 _33988_ (.A(_01076_),
    .Z(_00477_));
 BUF_X1 _33989_ (.A(_00421_),
    .Z(_01020_));
 BUF_X1 _33990_ (.A(_00420_),
    .Z(_01019_));
 BUF_X1 _33991_ (.A(key[123]),
    .Z(_01228_));
 BUF_X1 _33992_ (.A(_01077_),
    .Z(_00478_));
 BUF_X1 _33993_ (.A(_00423_),
    .Z(_01022_));
 BUF_X1 _33994_ (.A(_00422_),
    .Z(_01021_));
 BUF_X1 _33995_ (.A(key[124]),
    .Z(_01229_));
 BUF_X1 _33996_ (.A(_01078_),
    .Z(_00479_));
 BUF_X1 _33997_ (.A(_00425_),
    .Z(_01024_));
 BUF_X1 _33998_ (.A(_00424_),
    .Z(_01023_));
 BUF_X1 _33999_ (.A(key[125]),
    .Z(_01230_));
 BUF_X1 _34000_ (.A(_01079_),
    .Z(_00480_));
 BUF_X1 _34001_ (.A(_00427_),
    .Z(_01026_));
 BUF_X1 _34002_ (.A(_00426_),
    .Z(_01025_));
 BUF_X1 _34003_ (.A(key[126]),
    .Z(_01231_));
 BUF_X1 _34004_ (.A(_01081_),
    .Z(_00482_));
 BUF_X1 _34005_ (.A(_00429_),
    .Z(_01028_));
 BUF_X1 _34006_ (.A(_00428_),
    .Z(_01027_));
 BUF_X1 _34007_ (.A(key[127]),
    .Z(_01232_));
 BUF_X1 _34008_ (.A(_01082_),
    .Z(_00483_));
 BUF_X1 _34009_ (.A(\u0.w[2][11] ),
    .Z(_17242_));
 BUF_X1 _34010_ (.A(\text_in_r[43] ),
    .Z(_17077_));
 BUF_X1 _34011_ (.A(_00687_),
    .Z(_00088_));
 BUF_X1 _34012_ (.A(\u0.w[2][12] ),
    .Z(_17243_));
 BUF_X1 _34013_ (.A(\text_in_r[44] ),
    .Z(_17078_));
 BUF_X1 _34014_ (.A(_00688_),
    .Z(_00089_));
 BUF_X1 _34015_ (.A(\u0.w[2][13] ),
    .Z(_17244_));
 BUF_X1 _34016_ (.A(\text_in_r[45] ),
    .Z(_17079_));
 BUF_X1 _34017_ (.A(_00689_),
    .Z(_00090_));
 BUF_X1 _34018_ (.A(\u0.w[2][14] ),
    .Z(_17245_));
 BUF_X1 _34019_ (.A(\text_in_r[46] ),
    .Z(_17080_));
 BUF_X1 _34020_ (.A(_00690_),
    .Z(_00091_));
 BUF_X1 _34021_ (.A(\u0.w[2][15] ),
    .Z(_17246_));
 BUF_X1 _34022_ (.A(\text_in_r[47] ),
    .Z(_17081_));
 BUF_X1 _34023_ (.A(_00691_),
    .Z(_00092_));
 BUF_X1 _34024_ (.A(\u0.w[1][0] ),
    .Z(_17208_));
 BUF_X1 _34025_ (.A(\u0.w[0][0] ),
    .Z(_17176_));
 BUF_X1 _34026_ (.A(key[64]),
    .Z(_01290_));
 BUF_X1 _34027_ (.A(_01090_),
    .Z(_00491_));
 BUF_X1 _34028_ (.A(\u0.w[1][1] ),
    .Z(_17219_));
 BUF_X1 _34029_ (.A(\u0.w[0][1] ),
    .Z(_17187_));
 BUF_X1 _34030_ (.A(key[65]),
    .Z(_01291_));
 BUF_X1 _34031_ (.A(_01101_),
    .Z(_00502_));
 BUF_X1 _34032_ (.A(\u0.w[1][2] ),
    .Z(_17230_));
 BUF_X1 _34033_ (.A(\u0.w[0][2] ),
    .Z(_17198_));
 BUF_X1 _34034_ (.A(key[66]),
    .Z(_01292_));
 BUF_X1 _34035_ (.A(_01112_),
    .Z(_00513_));
 BUF_X1 _34036_ (.A(\u0.w[1][3] ),
    .Z(_17233_));
 BUF_X1 _34037_ (.A(\u0.w[0][3] ),
    .Z(_17201_));
 BUF_X1 _34038_ (.A(key[67]),
    .Z(_01293_));
 BUF_X1 _34039_ (.A(_01115_),
    .Z(_00516_));
 BUF_X1 _34040_ (.A(\u0.w[1][4] ),
    .Z(_17234_));
 BUF_X1 _34041_ (.A(\u0.w[0][4] ),
    .Z(_17202_));
 BUF_X1 _34042_ (.A(key[68]),
    .Z(_01294_));
 BUF_X1 _34043_ (.A(_01116_),
    .Z(_00517_));
 BUF_X1 _34044_ (.A(\u0.w[1][5] ),
    .Z(_17235_));
 BUF_X1 _34045_ (.A(\u0.w[0][5] ),
    .Z(_17203_));
 BUF_X1 _34046_ (.A(key[69]),
    .Z(_01295_));
 BUF_X1 _34047_ (.A(_01117_),
    .Z(_00518_));
 BUF_X1 _34048_ (.A(\u0.w[1][6] ),
    .Z(_17236_));
 BUF_X1 _34049_ (.A(\u0.w[0][6] ),
    .Z(_17204_));
 BUF_X1 _34050_ (.A(key[70]),
    .Z(_01297_));
 BUF_X1 _34051_ (.A(_01118_),
    .Z(_00519_));
 BUF_X1 _34052_ (.A(\u0.w[1][7] ),
    .Z(_17237_));
 BUF_X1 _34053_ (.A(\u0.w[0][7] ),
    .Z(_17205_));
 BUF_X1 _34054_ (.A(key[71]),
    .Z(_01298_));
 BUF_X1 _34055_ (.A(_01119_),
    .Z(_00520_));
 BUF_X1 _34056_ (.A(\u0.w[1][8] ),
    .Z(_17238_));
 BUF_X1 _34057_ (.A(\u0.w[0][8] ),
    .Z(_17206_));
 BUF_X1 _34058_ (.A(key[72]),
    .Z(_01299_));
 BUF_X1 _34059_ (.A(_01120_),
    .Z(_00521_));
 BUF_X1 _34060_ (.A(\u0.w[1][9] ),
    .Z(_17239_));
 BUF_X1 _34061_ (.A(\u0.w[0][9] ),
    .Z(_17207_));
 BUF_X1 _34062_ (.A(key[73]),
    .Z(_01300_));
 BUF_X1 _34063_ (.A(_01121_),
    .Z(_00522_));
 BUF_X1 _34064_ (.A(\u0.w[1][10] ),
    .Z(_17209_));
 BUF_X1 _34065_ (.A(\u0.w[0][10] ),
    .Z(_17177_));
 BUF_X1 _34066_ (.A(key[74]),
    .Z(_01301_));
 BUF_X1 _34067_ (.A(_01091_),
    .Z(_00492_));
 BUF_X1 _34068_ (.A(\u0.w[1][11] ),
    .Z(_17210_));
 BUF_X1 _34069_ (.A(\u0.w[0][11] ),
    .Z(_17178_));
 BUF_X1 _34070_ (.A(key[75]),
    .Z(_01302_));
 BUF_X1 _34071_ (.A(_01092_),
    .Z(_00493_));
 BUF_X1 _34072_ (.A(\u0.w[1][12] ),
    .Z(_17211_));
 BUF_X1 _34073_ (.A(\u0.w[0][12] ),
    .Z(_17179_));
 BUF_X1 _34074_ (.A(key[76]),
    .Z(_01303_));
 BUF_X1 _34075_ (.A(_01093_),
    .Z(_00494_));
 BUF_X1 _34076_ (.A(\u0.w[1][13] ),
    .Z(_17212_));
 BUF_X1 _34077_ (.A(\u0.w[0][13] ),
    .Z(_17180_));
 BUF_X1 _34078_ (.A(key[77]),
    .Z(_01304_));
 BUF_X1 _34079_ (.A(_01094_),
    .Z(_00495_));
 BUF_X1 _34080_ (.A(\u0.w[1][14] ),
    .Z(_17213_));
 BUF_X1 _34081_ (.A(\u0.w[0][14] ),
    .Z(_17181_));
 BUF_X1 _34082_ (.A(key[78]),
    .Z(_01305_));
 BUF_X1 _34083_ (.A(_01095_),
    .Z(_00496_));
 BUF_X1 _34084_ (.A(\u0.w[1][15] ),
    .Z(_17214_));
 BUF_X1 _34085_ (.A(\u0.w[0][15] ),
    .Z(_17182_));
 BUF_X1 _34086_ (.A(key[79]),
    .Z(_01306_));
 BUF_X1 _34087_ (.A(_01096_),
    .Z(_00497_));
 BUF_X1 _34088_ (.A(\u0.w[1][16] ),
    .Z(_17215_));
 BUF_X1 _34089_ (.A(\u0.w[0][16] ),
    .Z(_17183_));
 BUF_X1 _34090_ (.A(key[80]),
    .Z(_01308_));
 BUF_X1 _34091_ (.A(_01097_),
    .Z(_00498_));
 BUF_X1 _34092_ (.A(\u0.w[1][17] ),
    .Z(_17216_));
 BUF_X1 _34093_ (.A(\u0.w[0][17] ),
    .Z(_17184_));
 BUF_X1 _34094_ (.A(key[81]),
    .Z(_01309_));
 BUF_X1 _34095_ (.A(_01098_),
    .Z(_00499_));
 BUF_X1 _34096_ (.A(\u0.w[1][18] ),
    .Z(_17217_));
 BUF_X1 _34097_ (.A(\u0.w[0][18] ),
    .Z(_17185_));
 BUF_X1 _34098_ (.A(key[82]),
    .Z(_01310_));
 BUF_X1 _34099_ (.A(_01099_),
    .Z(_00500_));
 BUF_X1 _34100_ (.A(\u0.w[1][19] ),
    .Z(_17218_));
 BUF_X1 _34101_ (.A(\u0.w[0][19] ),
    .Z(_17186_));
 BUF_X1 _34102_ (.A(key[83]),
    .Z(_01311_));
 BUF_X1 _34103_ (.A(_01100_),
    .Z(_00501_));
 BUF_X1 _34104_ (.A(\u0.w[1][20] ),
    .Z(_17220_));
 BUF_X1 _34105_ (.A(\u0.w[0][20] ),
    .Z(_17188_));
 BUF_X1 _34106_ (.A(key[84]),
    .Z(_01312_));
 BUF_X1 _34107_ (.A(_01102_),
    .Z(_00503_));
 BUF_X1 _34108_ (.A(\u0.w[1][21] ),
    .Z(_17221_));
 BUF_X1 _34109_ (.A(\u0.w[0][21] ),
    .Z(_17189_));
 BUF_X1 _34110_ (.A(key[85]),
    .Z(_01313_));
 BUF_X1 _34111_ (.A(_01103_),
    .Z(_00504_));
 BUF_X1 _34112_ (.A(\u0.w[1][22] ),
    .Z(_17222_));
 BUF_X1 _34113_ (.A(\u0.w[0][22] ),
    .Z(_17190_));
 BUF_X1 _34114_ (.A(key[86]),
    .Z(_01314_));
 BUF_X1 _34115_ (.A(_01104_),
    .Z(_00505_));
 BUF_X1 _34116_ (.A(\u0.w[1][23] ),
    .Z(_17223_));
 BUF_X1 _34117_ (.A(\u0.w[0][23] ),
    .Z(_17191_));
 BUF_X1 _34118_ (.A(key[87]),
    .Z(_01315_));
 BUF_X1 _34119_ (.A(_01105_),
    .Z(_00506_));
 BUF_X1 _34120_ (.A(\u0.w[0][24] ),
    .Z(_17192_));
 BUF_X1 _34121_ (.A(\u0.w[1][24] ),
    .Z(_17224_));
 BUF_X1 _34122_ (.A(key[88]),
    .Z(_01316_));
 BUF_X1 _34123_ (.A(_01106_),
    .Z(_00507_));
 BUF_X1 _34124_ (.A(\u0.w[0][25] ),
    .Z(_17193_));
 BUF_X1 _34125_ (.A(\u0.w[1][25] ),
    .Z(_17225_));
 BUF_X1 _34126_ (.A(key[89]),
    .Z(_01317_));
 BUF_X1 _34127_ (.A(_01107_),
    .Z(_00508_));
 BUF_X1 _34128_ (.A(\u0.w[0][26] ),
    .Z(_17194_));
 BUF_X1 _34129_ (.A(\u0.w[1][26] ),
    .Z(_17226_));
 BUF_X1 _34130_ (.A(key[90]),
    .Z(_01319_));
 BUF_X1 _34131_ (.A(_01108_),
    .Z(_00509_));
 BUF_X1 _34132_ (.A(\u0.w[0][27] ),
    .Z(_17195_));
 BUF_X1 _34133_ (.A(\u0.w[1][27] ),
    .Z(_17227_));
 BUF_X1 _34134_ (.A(key[91]),
    .Z(_01320_));
 BUF_X1 _34135_ (.A(_01109_),
    .Z(_00510_));
 BUF_X1 _34136_ (.A(\u0.w[0][28] ),
    .Z(_17196_));
 BUF_X1 _34137_ (.A(\u0.w[1][28] ),
    .Z(_17228_));
 BUF_X1 _34138_ (.A(key[92]),
    .Z(_01321_));
 BUF_X1 _34139_ (.A(_01110_),
    .Z(_00511_));
 BUF_X1 _34140_ (.A(\u0.w[0][29] ),
    .Z(_17197_));
 BUF_X1 _34141_ (.A(\u0.w[1][29] ),
    .Z(_17229_));
 BUF_X1 _34142_ (.A(key[93]),
    .Z(_01322_));
 BUF_X1 _34143_ (.A(_01111_),
    .Z(_00512_));
 BUF_X1 _34144_ (.A(\u0.w[0][30] ),
    .Z(_17199_));
 BUF_X1 _34145_ (.A(\u0.w[1][30] ),
    .Z(_17231_));
 BUF_X1 _34146_ (.A(key[94]),
    .Z(_01323_));
 BUF_X1 _34147_ (.A(_01113_),
    .Z(_00514_));
 BUF_X1 _34148_ (.A(\u0.w[0][31] ),
    .Z(_17200_));
 BUF_X1 _34149_ (.A(\u0.w[1][31] ),
    .Z(_17232_));
 BUF_X1 _34150_ (.A(key[95]),
    .Z(_01324_));
 BUF_X1 _34151_ (.A(_01114_),
    .Z(_00515_));
 BUF_X1 _34152_ (.A(_00430_),
    .Z(_01029_));
 BUF_X1 _34153_ (.A(\u0.w[2][16] ),
    .Z(_17247_));
 BUF_X1 _34154_ (.A(\text_in_r[48] ),
    .Z(_17082_));
 BUF_X1 _34155_ (.A(_00652_),
    .Z(_00053_));
 BUF_X1 _34156_ (.A(_00431_),
    .Z(_01030_));
 BUF_X1 _34157_ (.A(\u0.w[2][17] ),
    .Z(_17248_));
 BUF_X1 _34158_ (.A(\text_in_r[49] ),
    .Z(_17083_));
 BUF_X1 _34159_ (.A(_00653_),
    .Z(_00054_));
 BUF_X1 _34160_ (.A(\u0.w[2][18] ),
    .Z(_17249_));
 BUF_X1 _34161_ (.A(\text_in_r[50] ),
    .Z(_17085_));
 BUF_X1 _34162_ (.A(_00654_),
    .Z(_00055_));
 BUF_X1 _34163_ (.A(\u0.w[2][19] ),
    .Z(_17250_));
 BUF_X1 _34164_ (.A(\text_in_r[51] ),
    .Z(_17086_));
 BUF_X1 _34165_ (.A(_00655_),
    .Z(_00056_));
 BUF_X1 _34166_ (.A(\u0.w[2][20] ),
    .Z(_17252_));
 BUF_X1 _34167_ (.A(\text_in_r[52] ),
    .Z(_17087_));
 BUF_X1 _34168_ (.A(_00656_),
    .Z(_00057_));
 BUF_X1 _34169_ (.A(_00432_),
    .Z(_01031_));
 BUF_X1 _34170_ (.A(\u0.w[2][21] ),
    .Z(_17253_));
 BUF_X1 _34171_ (.A(\text_in_r[53] ),
    .Z(_17088_));
 BUF_X1 _34172_ (.A(_00657_),
    .Z(_00058_));
 BUF_X1 _34173_ (.A(_00433_),
    .Z(_01032_));
 BUF_X1 _34174_ (.A(\u0.w[2][22] ),
    .Z(_17254_));
 BUF_X1 _34175_ (.A(\text_in_r[54] ),
    .Z(_17089_));
 BUF_X1 _34176_ (.A(_00658_),
    .Z(_00059_));
 BUF_X1 _34177_ (.A(\u0.w[2][23] ),
    .Z(_17255_));
 BUF_X1 _34178_ (.A(\text_in_r[55] ),
    .Z(_17090_));
 BUF_X1 _34179_ (.A(_00659_),
    .Z(_00060_));
 BUF_X1 _34180_ (.A(key[32]),
    .Z(_01255_));
 BUF_X1 _34181_ (.A(_01122_),
    .Z(_00523_));
 BUF_X1 _34182_ (.A(key[33]),
    .Z(_01256_));
 BUF_X1 _34183_ (.A(_01133_),
    .Z(_00534_));
 BUF_X1 _34184_ (.A(key[34]),
    .Z(_01257_));
 BUF_X1 _34185_ (.A(_01144_),
    .Z(_00545_));
 BUF_X1 _34186_ (.A(key[35]),
    .Z(_01258_));
 BUF_X1 _34187_ (.A(_01147_),
    .Z(_00548_));
 BUF_X1 _34188_ (.A(key[36]),
    .Z(_01259_));
 BUF_X1 _34189_ (.A(_01148_),
    .Z(_00549_));
 BUF_X1 _34190_ (.A(key[37]),
    .Z(_01260_));
 BUF_X1 _34191_ (.A(_01149_),
    .Z(_00550_));
 BUF_X1 _34192_ (.A(key[38]),
    .Z(_01261_));
 BUF_X1 _34193_ (.A(_01150_),
    .Z(_00551_));
 BUF_X1 _34194_ (.A(key[39]),
    .Z(_01262_));
 BUF_X1 _34195_ (.A(_01151_),
    .Z(_00552_));
 BUF_X1 _34196_ (.A(key[40]),
    .Z(_01264_));
 BUF_X1 _34197_ (.A(_01152_),
    .Z(_00553_));
 BUF_X1 _34198_ (.A(key[41]),
    .Z(_01265_));
 BUF_X1 _34199_ (.A(_01153_),
    .Z(_00554_));
 BUF_X1 _34200_ (.A(key[42]),
    .Z(_01266_));
 BUF_X1 _34201_ (.A(_01123_),
    .Z(_00524_));
 BUF_X1 _34202_ (.A(key[43]),
    .Z(_01267_));
 BUF_X1 _34203_ (.A(_01124_),
    .Z(_00525_));
 BUF_X1 _34204_ (.A(key[44]),
    .Z(_01268_));
 BUF_X1 _34205_ (.A(_01125_),
    .Z(_00526_));
 BUF_X1 _34206_ (.A(key[45]),
    .Z(_01269_));
 BUF_X1 _34207_ (.A(_01126_),
    .Z(_00527_));
 BUF_X1 _34208_ (.A(key[46]),
    .Z(_01270_));
 BUF_X1 _34209_ (.A(_01127_),
    .Z(_00528_));
 BUF_X1 _34210_ (.A(key[47]),
    .Z(_01271_));
 BUF_X1 _34211_ (.A(_01128_),
    .Z(_00529_));
 BUF_X1 _34212_ (.A(key[48]),
    .Z(_01272_));
 BUF_X1 _34213_ (.A(_01129_),
    .Z(_00530_));
 BUF_X1 _34214_ (.A(key[49]),
    .Z(_01273_));
 BUF_X1 _34215_ (.A(_01130_),
    .Z(_00531_));
 BUF_X1 _34216_ (.A(key[50]),
    .Z(_01275_));
 BUF_X1 _34217_ (.A(_01131_),
    .Z(_00532_));
 BUF_X1 _34218_ (.A(key[51]),
    .Z(_01276_));
 BUF_X1 _34219_ (.A(_01132_),
    .Z(_00533_));
 BUF_X1 _34220_ (.A(key[52]),
    .Z(_01277_));
 BUF_X1 _34221_ (.A(_01134_),
    .Z(_00535_));
 BUF_X1 _34222_ (.A(key[53]),
    .Z(_01278_));
 BUF_X1 _34223_ (.A(_01135_),
    .Z(_00536_));
 BUF_X1 _34224_ (.A(key[54]),
    .Z(_01279_));
 BUF_X1 _34225_ (.A(_01136_),
    .Z(_00537_));
 BUF_X1 _34226_ (.A(key[55]),
    .Z(_01280_));
 BUF_X1 _34227_ (.A(_01137_),
    .Z(_00538_));
 BUF_X1 _34228_ (.A(\u0.w[2][24] ),
    .Z(_17256_));
 BUF_X1 _34229_ (.A(key[56]),
    .Z(_01281_));
 BUF_X1 _34230_ (.A(_01138_),
    .Z(_00539_));
 BUF_X1 _34231_ (.A(\u0.w[2][25] ),
    .Z(_17257_));
 BUF_X1 _34232_ (.A(key[57]),
    .Z(_01282_));
 BUF_X1 _34233_ (.A(_01139_),
    .Z(_00540_));
 BUF_X1 _34234_ (.A(\u0.w[2][26] ),
    .Z(_17258_));
 BUF_X1 _34235_ (.A(key[58]),
    .Z(_01283_));
 BUF_X1 _34236_ (.A(_01140_),
    .Z(_00541_));
 BUF_X1 _34237_ (.A(\u0.w[2][27] ),
    .Z(_17259_));
 BUF_X1 _34238_ (.A(key[59]),
    .Z(_01284_));
 BUF_X1 _34239_ (.A(_01141_),
    .Z(_00542_));
 BUF_X1 _34240_ (.A(\u0.w[2][28] ),
    .Z(_17260_));
 BUF_X1 _34241_ (.A(key[60]),
    .Z(_01286_));
 BUF_X1 _34242_ (.A(_01142_),
    .Z(_00543_));
 BUF_X1 _34243_ (.A(\u0.w[2][29] ),
    .Z(_17261_));
 BUF_X1 _34244_ (.A(key[61]),
    .Z(_01287_));
 BUF_X1 _34245_ (.A(_01143_),
    .Z(_00544_));
 BUF_X1 _34246_ (.A(\u0.w[2][30] ),
    .Z(_17263_));
 BUF_X1 _34247_ (.A(key[62]),
    .Z(_01288_));
 BUF_X1 _34248_ (.A(_01145_),
    .Z(_00546_));
 BUF_X1 _34249_ (.A(\u0.w[2][31] ),
    .Z(_17264_));
 BUF_X1 _34250_ (.A(key[63]),
    .Z(_01289_));
 BUF_X1 _34251_ (.A(_01146_),
    .Z(_00547_));
 BUF_X1 _34252_ (.A(_00434_),
    .Z(_01033_));
 BUF_X1 _34253_ (.A(\text_in_r[56] ),
    .Z(_17091_));
 BUF_X1 _34254_ (.A(_00620_),
    .Z(_00021_));
 BUF_X1 _34255_ (.A(_00435_),
    .Z(_01034_));
 BUF_X1 _34256_ (.A(\text_in_r[57] ),
    .Z(_17092_));
 BUF_X1 _34257_ (.A(_00621_),
    .Z(_00022_));
 BUF_X1 _34258_ (.A(\text_in_r[58] ),
    .Z(_17093_));
 BUF_X1 _34259_ (.A(_00622_),
    .Z(_00023_));
 BUF_X1 _34260_ (.A(\text_in_r[59] ),
    .Z(_17094_));
 BUF_X1 _34261_ (.A(_00623_),
    .Z(_00024_));
 BUF_X1 _34262_ (.A(\text_in_r[60] ),
    .Z(_17096_));
 BUF_X1 _34263_ (.A(_00624_),
    .Z(_00025_));
 BUF_X1 _34264_ (.A(_00436_),
    .Z(_01035_));
 BUF_X1 _34265_ (.A(\text_in_r[61] ),
    .Z(_17097_));
 BUF_X1 _34266_ (.A(_00625_),
    .Z(_00026_));
 BUF_X1 _34267_ (.A(_00437_),
    .Z(_01036_));
 BUF_X1 _34268_ (.A(\text_in_r[62] ),
    .Z(_17098_));
 BUF_X1 _34269_ (.A(_00626_),
    .Z(_00027_));
 BUF_X1 _34270_ (.A(\text_in_r[63] ),
    .Z(_17099_));
 BUF_X1 _34271_ (.A(_00627_),
    .Z(_00028_));
 BUF_X1 _34272_ (.A(key[0]),
    .Z(_01202_));
 BUF_X1 _34273_ (.A(_01154_),
    .Z(_00555_));
 BUF_X1 _34274_ (.A(key[1]),
    .Z(_01241_));
 BUF_X1 _34275_ (.A(_01165_),
    .Z(_00566_));
 BUF_X1 _34276_ (.A(\sa01[5] ),
    .Z(_16769_));
 BUF_X1 _34277_ (.A(\sa01[4] ),
    .Z(_16768_));
 BUF_X1 _34278_ (.A(\sa01[7] ),
    .Z(_16771_));
 BUF_X1 _34279_ (.A(\sa01[6] ),
    .Z(_16770_));
 BUF_X1 _34280_ (.A(\sa01[1] ),
    .Z(_16765_));
 BUF_X1 _34281_ (.A(\sa01[0] ),
    .Z(_16764_));
 BUF_X1 _34282_ (.A(\sa01[2] ),
    .Z(_16766_));
 BUF_X1 _34283_ (.A(\sa01[3] ),
    .Z(_16767_));
 BUF_X1 _34284_ (.A(\sa12[5] ),
    .Z(_16809_));
 BUF_X1 _34285_ (.A(\sa12[4] ),
    .Z(_16808_));
 BUF_X1 _34286_ (.A(\sa12[7] ),
    .Z(_16811_));
 BUF_X1 _34287_ (.A(\sa12[6] ),
    .Z(_16810_));
 BUF_X1 _34288_ (.A(\sa12[1] ),
    .Z(_16805_));
 BUF_X1 _34289_ (.A(\sa12[0] ),
    .Z(_16804_));
 BUF_X1 _34290_ (.A(\sa12[2] ),
    .Z(_16806_));
 BUF_X1 _34291_ (.A(\sa12[3] ),
    .Z(_16807_));
 BUF_X1 _34292_ (.A(\sa23[5] ),
    .Z(_16849_));
 BUF_X1 _34293_ (.A(\sa23[4] ),
    .Z(_16848_));
 BUF_X1 _34294_ (.A(\sa23[7] ),
    .Z(_16851_));
 BUF_X1 _34295_ (.A(\sa23[6] ),
    .Z(_16850_));
 BUF_X1 _34296_ (.A(\sa23[1] ),
    .Z(_16845_));
 BUF_X1 _34297_ (.A(\sa23[0] ),
    .Z(_16844_));
 BUF_X1 _34298_ (.A(\sa23[2] ),
    .Z(_16846_));
 BUF_X1 _34299_ (.A(\sa23[3] ),
    .Z(_16847_));
 BUF_X1 _34300_ (.A(\sa30[0] ),
    .Z(_16852_));
 BUF_X1 _34301_ (.A(\sa30[1] ),
    .Z(_16853_));
 BUF_X1 _34302_ (.A(\sa30[2] ),
    .Z(_16854_));
 BUF_X1 _34303_ (.A(\sa30[3] ),
    .Z(_16855_));
 BUF_X1 _34304_ (.A(\sa30[5] ),
    .Z(_16857_));
 BUF_X1 _34305_ (.A(\sa30[4] ),
    .Z(_16856_));
 BUF_X1 _34306_ (.A(\sa30[7] ),
    .Z(_16859_));
 BUF_X1 _34307_ (.A(\sa30[6] ),
    .Z(_16858_));
 BUF_X1 _34308_ (.A(\text_in_r[64] ),
    .Z(_17100_));
 BUF_X1 _34309_ (.A(_00708_),
    .Z(_00109_));
 BUF_X1 _34310_ (.A(key[2]),
    .Z(_01252_));
 BUF_X1 _34311_ (.A(_01176_),
    .Z(_00577_));
 BUF_X1 _34312_ (.A(key[3]),
    .Z(_01263_));
 BUF_X1 _34313_ (.A(_01179_),
    .Z(_00580_));
 BUF_X1 _34314_ (.A(key[4]),
    .Z(_01274_));
 BUF_X1 _34315_ (.A(_01180_),
    .Z(_00581_));
 BUF_X1 _34316_ (.A(key[5]),
    .Z(_01285_));
 BUF_X1 _34317_ (.A(_01181_),
    .Z(_00582_));
 BUF_X1 _34318_ (.A(key[6]),
    .Z(_01296_));
 BUF_X1 _34319_ (.A(_01182_),
    .Z(_00583_));
 BUF_X1 _34320_ (.A(key[7]),
    .Z(_01307_));
 BUF_X1 _34321_ (.A(_01183_),
    .Z(_00584_));
 BUF_X1 _34322_ (.A(key[8]),
    .Z(_01318_));
 BUF_X1 _34323_ (.A(_01184_),
    .Z(_00585_));
 BUF_X1 _34324_ (.A(key[9]),
    .Z(_01329_));
 BUF_X1 _34325_ (.A(_01185_),
    .Z(_00586_));
 BUF_X1 _34326_ (.A(key[10]),
    .Z(_01213_));
 BUF_X1 _34327_ (.A(_01155_),
    .Z(_00556_));
 BUF_X1 _34328_ (.A(key[11]),
    .Z(_01224_));
 BUF_X1 _34329_ (.A(_01156_),
    .Z(_00557_));
 BUF_X1 _34330_ (.A(\text_in_r[65] ),
    .Z(_17101_));
 BUF_X1 _34331_ (.A(_00709_),
    .Z(_00110_));
 BUF_X1 _34332_ (.A(key[12]),
    .Z(_01233_));
 BUF_X1 _34333_ (.A(_01157_),
    .Z(_00558_));
 BUF_X1 _34334_ (.A(key[13]),
    .Z(_01234_));
 BUF_X1 _34335_ (.A(_01158_),
    .Z(_00559_));
 BUF_X1 _34336_ (.A(key[14]),
    .Z(_01235_));
 BUF_X1 _34337_ (.A(_01159_),
    .Z(_00560_));
 BUF_X1 _34338_ (.A(key[15]),
    .Z(_01236_));
 BUF_X1 _34339_ (.A(_01160_),
    .Z(_00561_));
 BUF_X1 _34340_ (.A(key[16]),
    .Z(_01237_));
 BUF_X1 _34341_ (.A(_01161_),
    .Z(_00562_));
 BUF_X1 _34342_ (.A(key[17]),
    .Z(_01238_));
 BUF_X1 _34343_ (.A(_01162_),
    .Z(_00563_));
 BUF_X1 _34344_ (.A(key[18]),
    .Z(_01239_));
 BUF_X1 _34345_ (.A(_01163_),
    .Z(_00564_));
 BUF_X1 _34346_ (.A(key[19]),
    .Z(_01240_));
 BUF_X1 _34347_ (.A(_01164_),
    .Z(_00565_));
 BUF_X1 _34348_ (.A(key[20]),
    .Z(_01242_));
 BUF_X1 _34349_ (.A(_01166_),
    .Z(_00567_));
 BUF_X1 _34350_ (.A(key[21]),
    .Z(_01243_));
 BUF_X1 _34351_ (.A(_01167_),
    .Z(_00568_));
 BUF_X1 _34352_ (.A(\text_in_r[66] ),
    .Z(_17102_));
 BUF_X1 _34353_ (.A(_00710_),
    .Z(_00111_));
 BUF_X1 _34354_ (.A(key[22]),
    .Z(_01244_));
 BUF_X1 _34355_ (.A(_01168_),
    .Z(_00569_));
 BUF_X1 _34356_ (.A(key[23]),
    .Z(_01245_));
 BUF_X1 _34357_ (.A(_01169_),
    .Z(_00570_));
 BUF_X1 _34358_ (.A(key[24]),
    .Z(_01246_));
 BUF_X1 _34359_ (.A(_01170_),
    .Z(_00571_));
 BUF_X1 _34360_ (.A(key[25]),
    .Z(_01247_));
 BUF_X1 _34361_ (.A(_01171_),
    .Z(_00572_));
 BUF_X1 _34362_ (.A(key[26]),
    .Z(_01248_));
 BUF_X1 _34363_ (.A(_01172_),
    .Z(_00573_));
 BUF_X1 _34364_ (.A(key[27]),
    .Z(_01249_));
 BUF_X1 _34365_ (.A(_01173_),
    .Z(_00574_));
 BUF_X1 _34366_ (.A(key[28]),
    .Z(_01250_));
 BUF_X1 _34367_ (.A(_01174_),
    .Z(_00575_));
 BUF_X1 _34368_ (.A(key[29]),
    .Z(_01251_));
 BUF_X1 _34369_ (.A(_01175_),
    .Z(_00576_));
 BUF_X1 _34370_ (.A(key[30]),
    .Z(_01253_));
 BUF_X1 _34371_ (.A(_01177_),
    .Z(_00578_));
 BUF_X1 _34372_ (.A(key[31]),
    .Z(_01254_));
 BUF_X1 _34373_ (.A(_01178_),
    .Z(_00579_));
 BUF_X1 _34374_ (.A(\text_in_r[67] ),
    .Z(_17103_));
 BUF_X1 _34375_ (.A(_00711_),
    .Z(_00112_));
 BUF_X1 _34376_ (.A(\text_in_r[68] ),
    .Z(_17104_));
 BUF_X1 _34377_ (.A(_00712_),
    .Z(_00113_));
 BUF_X1 _34378_ (.A(\text_in_r[69] ),
    .Z(_17105_));
 BUF_X1 _34379_ (.A(_00713_),
    .Z(_00114_));
 BUF_X1 _34380_ (.A(\text_in_r[70] ),
    .Z(_17107_));
 BUF_X1 _34381_ (.A(_00714_),
    .Z(_00115_));
 BUF_X1 _34382_ (.A(\text_in_r[71] ),
    .Z(_17108_));
 BUF_X1 _34383_ (.A(_00715_),
    .Z(_00116_));
 BUF_X1 _34384_ (.A(_00438_),
    .Z(_01037_));
 BUF_X1 _34385_ (.A(\text_in_r[72] ),
    .Z(_17109_));
 BUF_X1 _34386_ (.A(_00676_),
    .Z(_00077_));
 BUF_X1 _34387_ (.A(\text_in_r[73] ),
    .Z(_17110_));
 BUF_X1 _34388_ (.A(_00677_),
    .Z(_00078_));
 BUF_X1 _34389_ (.A(\text_in_r[74] ),
    .Z(_17111_));
 BUF_X1 _34390_ (.A(_00678_),
    .Z(_00079_));
 BUF_X1 _34391_ (.A(\text_in_r[75] ),
    .Z(_17112_));
 BUF_X1 _34392_ (.A(_00679_),
    .Z(_00080_));
 BUF_X1 _34393_ (.A(\text_in_r[76] ),
    .Z(_17113_));
 BUF_X1 _34394_ (.A(_00680_),
    .Z(_00081_));
 BUF_X1 _34395_ (.A(\text_in_r[77] ),
    .Z(_17114_));
 BUF_X1 _34396_ (.A(_00681_),
    .Z(_00082_));
 BUF_X1 _34397_ (.A(\text_in_r[78] ),
    .Z(_17115_));
 BUF_X1 _34398_ (.A(_00682_),
    .Z(_00083_));
 BUF_X1 _34399_ (.A(\text_in_r[79] ),
    .Z(_17116_));
 BUF_X1 _34400_ (.A(_00683_),
    .Z(_00084_));
 BUF_X1 _34401_ (.A(_00439_),
    .Z(_01038_));
 BUF_X1 _34402_ (.A(\text_in_r[80] ),
    .Z(_17118_));
 BUF_X1 _34403_ (.A(_00644_),
    .Z(_00045_));
 BUF_X1 _34404_ (.A(_00440_),
    .Z(_01039_));
 BUF_X1 _34405_ (.A(\text_in_r[81] ),
    .Z(_17119_));
 BUF_X1 _34406_ (.A(_00645_),
    .Z(_00046_));
 BUF_X1 _34407_ (.A(\text_in_r[82] ),
    .Z(_17120_));
 BUF_X1 _34408_ (.A(_00646_),
    .Z(_00047_));
 BUF_X1 _34409_ (.A(\text_in_r[83] ),
    .Z(_17121_));
 BUF_X1 _34410_ (.A(_00647_),
    .Z(_00048_));
 BUF_X1 _34411_ (.A(\text_in_r[84] ),
    .Z(_17122_));
 BUF_X1 _34412_ (.A(_00648_),
    .Z(_00049_));
 BUF_X1 _34413_ (.A(_00441_),
    .Z(_01040_));
 BUF_X1 _34414_ (.A(\text_in_r[85] ),
    .Z(_17123_));
 BUF_X1 _34415_ (.A(_00649_),
    .Z(_00050_));
 BUF_X1 _34416_ (.A(_00442_),
    .Z(_01041_));
 BUF_X1 _34417_ (.A(\text_in_r[86] ),
    .Z(_17124_));
 BUF_X1 _34418_ (.A(_00650_),
    .Z(_00051_));
 BUF_X1 _34419_ (.A(\text_in_r[87] ),
    .Z(_17125_));
 BUF_X1 _34420_ (.A(_00651_),
    .Z(_00052_));
 BUF_X1 _34421_ (.A(_00443_),
    .Z(_01042_));
 BUF_X1 _34422_ (.A(\text_in_r[88] ),
    .Z(_17126_));
 BUF_X1 _34423_ (.A(_00612_),
    .Z(_00013_));
 BUF_X1 _34424_ (.A(_00444_),
    .Z(_01043_));
 BUF_X1 _34425_ (.A(\text_in_r[89] ),
    .Z(_17127_));
 BUF_X1 _34426_ (.A(_00613_),
    .Z(_00014_));
 BUF_X1 _34427_ (.A(\text_in_r[90] ),
    .Z(_17129_));
 BUF_X1 _34428_ (.A(_00614_),
    .Z(_00015_));
 BUF_X1 _34429_ (.A(\text_in_r[91] ),
    .Z(_17130_));
 BUF_X1 _34430_ (.A(_00615_),
    .Z(_00016_));
 BUF_X1 _34431_ (.A(\text_in_r[92] ),
    .Z(_17131_));
 BUF_X1 _34432_ (.A(_00616_),
    .Z(_00017_));
 BUF_X1 _34433_ (.A(_00445_),
    .Z(_01044_));
 BUF_X1 _34434_ (.A(\text_in_r[93] ),
    .Z(_17132_));
 BUF_X1 _34435_ (.A(_00617_),
    .Z(_00018_));
 BUF_X1 _34436_ (.A(rst),
    .Z(_16755_));
 BUF_X1 _34437_ (.A(\dcnt[2] ),
    .Z(_01200_));
 BUF_X1 _34438_ (.A(\dcnt[3] ),
    .Z(_01201_));
 BUF_X1 _34439_ (.A(\dcnt[0] ),
    .Z(_01198_));
 BUF_X1 _34440_ (.A(\dcnt[1] ),
    .Z(_01199_));
 BUF_X1 _34441_ (.A(_00599_),
    .Z(_00000_));
 BUF_X1 _34442_ (.A(_00446_),
    .Z(_01045_));
 BUF_X1 _34443_ (.A(_00600_),
    .Z(_00001_));
 BUF_X1 _34444_ (.A(_00447_),
    .Z(_01046_));
 BUF_X1 _34445_ (.A(_00601_),
    .Z(_00002_));
 BUF_X1 _34446_ (.A(_00448_),
    .Z(_01047_));
 BUF_X1 _34447_ (.A(_00602_),
    .Z(_00003_));
 BUF_X1 _34448_ (.A(_00449_),
    .Z(_01048_));
 BUF_X1 _34449_ (.A(\text_in_r[94] ),
    .Z(_17133_));
 BUF_X1 _34450_ (.A(_00618_),
    .Z(_00019_));
 BUF_X1 _34451_ (.A(text_in[0]),
    .Z(_16884_));
 BUF_X1 _34452_ (.A(_00732_),
    .Z(_00133_));
 BUF_X1 _34453_ (.A(text_in[1]),
    .Z(_16923_));
 BUF_X1 _34454_ (.A(_00771_),
    .Z(_00172_));
 BUF_X1 _34455_ (.A(text_in[2]),
    .Z(_16934_));
 BUF_X1 _34456_ (.A(_00782_),
    .Z(_00183_));
 BUF_X1 _34457_ (.A(text_in[3]),
    .Z(_16945_));
 BUF_X1 _34458_ (.A(_00793_),
    .Z(_00194_));
 BUF_X1 _34459_ (.A(text_in[4]),
    .Z(_16956_));
 BUF_X1 _34460_ (.A(_00804_),
    .Z(_00205_));
 BUF_X1 _34461_ (.A(text_in[5]),
    .Z(_16967_));
 BUF_X1 _34462_ (.A(_00815_),
    .Z(_00216_));
 BUF_X1 _34463_ (.A(\text_in_r[95] ),
    .Z(_17134_));
 BUF_X1 _34464_ (.A(_00619_),
    .Z(_00020_));
 BUF_X1 _34465_ (.A(text_in[6]),
    .Z(_16978_));
 BUF_X1 _34466_ (.A(_00826_),
    .Z(_00227_));
 BUF_X1 _34467_ (.A(text_in[7]),
    .Z(_16989_));
 BUF_X1 _34468_ (.A(_00837_),
    .Z(_00238_));
 BUF_X1 _34469_ (.A(text_in[8]),
    .Z(_17000_));
 BUF_X1 _34470_ (.A(_00848_),
    .Z(_00249_));
 BUF_X1 _34471_ (.A(text_in[9]),
    .Z(_17011_));
 BUF_X1 _34472_ (.A(_00859_),
    .Z(_00260_));
 BUF_X1 _34473_ (.A(text_in[10]),
    .Z(_16895_));
 BUF_X1 _34474_ (.A(_00743_),
    .Z(_00144_));
 BUF_X1 _34475_ (.A(text_in[11]),
    .Z(_16906_));
 BUF_X1 _34476_ (.A(_00754_),
    .Z(_00155_));
 BUF_X1 _34477_ (.A(text_in[12]),
    .Z(_16915_));
 BUF_X1 _34478_ (.A(_00763_),
    .Z(_00164_));
 BUF_X1 _34479_ (.A(text_in[13]),
    .Z(_16916_));
 BUF_X1 _34480_ (.A(_00764_),
    .Z(_00165_));
 BUF_X1 _34481_ (.A(text_in[14]),
    .Z(_16917_));
 BUF_X1 _34482_ (.A(_00765_),
    .Z(_00166_));
 BUF_X1 _34483_ (.A(text_in[15]),
    .Z(_16918_));
 BUF_X1 _34484_ (.A(_00766_),
    .Z(_00167_));
 BUF_X1 _34485_ (.A(text_in[16]),
    .Z(_16919_));
 BUF_X1 _34486_ (.A(_00767_),
    .Z(_00168_));
 BUF_X1 _34487_ (.A(text_in[17]),
    .Z(_16920_));
 BUF_X1 _34488_ (.A(_00768_),
    .Z(_00169_));
 BUF_X1 _34489_ (.A(text_in[18]),
    .Z(_16921_));
 BUF_X1 _34490_ (.A(_00769_),
    .Z(_00170_));
 BUF_X1 _34491_ (.A(text_in[19]),
    .Z(_16922_));
 BUF_X1 _34492_ (.A(_00770_),
    .Z(_00171_));
 BUF_X1 _34493_ (.A(text_in[20]),
    .Z(_16924_));
 BUF_X1 _34494_ (.A(_00772_),
    .Z(_00173_));
 BUF_X1 _34495_ (.A(text_in[21]),
    .Z(_16925_));
 BUF_X1 _34496_ (.A(_00773_),
    .Z(_00174_));
 BUF_X1 _34497_ (.A(text_in[22]),
    .Z(_16926_));
 BUF_X1 _34498_ (.A(_00774_),
    .Z(_00175_));
 BUF_X1 _34499_ (.A(text_in[23]),
    .Z(_16927_));
 BUF_X1 _34500_ (.A(_00775_),
    .Z(_00176_));
 BUF_X1 _34501_ (.A(text_in[24]),
    .Z(_16928_));
 BUF_X1 _34502_ (.A(_00776_),
    .Z(_00177_));
 BUF_X1 _34503_ (.A(text_in[25]),
    .Z(_16929_));
 BUF_X1 _34504_ (.A(_00777_),
    .Z(_00178_));
 BUF_X1 _34505_ (.A(text_in[26]),
    .Z(_16930_));
 BUF_X1 _34506_ (.A(_00778_),
    .Z(_00179_));
 BUF_X1 _34507_ (.A(text_in[27]),
    .Z(_16931_));
 BUF_X1 _34508_ (.A(_00779_),
    .Z(_00180_));
 BUF_X1 _34509_ (.A(text_in[28]),
    .Z(_16932_));
 BUF_X1 _34510_ (.A(_00780_),
    .Z(_00181_));
 BUF_X1 _34511_ (.A(text_in[29]),
    .Z(_16933_));
 BUF_X1 _34512_ (.A(_00781_),
    .Z(_00182_));
 BUF_X1 _34513_ (.A(text_in[30]),
    .Z(_16935_));
 BUF_X1 _34514_ (.A(_00783_),
    .Z(_00184_));
 BUF_X1 _34515_ (.A(text_in[31]),
    .Z(_16936_));
 BUF_X1 _34516_ (.A(_00784_),
    .Z(_00185_));
 BUF_X1 _34517_ (.A(text_in[32]),
    .Z(_16937_));
 BUF_X1 _34518_ (.A(_00785_),
    .Z(_00186_));
 BUF_X1 _34519_ (.A(text_in[33]),
    .Z(_16938_));
 BUF_X1 _34520_ (.A(_00786_),
    .Z(_00187_));
 BUF_X1 _34521_ (.A(text_in[34]),
    .Z(_16939_));
 BUF_X1 _34522_ (.A(_00787_),
    .Z(_00188_));
 BUF_X1 _34523_ (.A(text_in[35]),
    .Z(_16940_));
 BUF_X1 _34524_ (.A(_00788_),
    .Z(_00189_));
 BUF_X1 _34525_ (.A(text_in[36]),
    .Z(_16941_));
 BUF_X1 _34526_ (.A(_00789_),
    .Z(_00190_));
 BUF_X1 _34527_ (.A(text_in[37]),
    .Z(_16942_));
 BUF_X1 _34528_ (.A(_00790_),
    .Z(_00191_));
 BUF_X1 _34529_ (.A(text_in[38]),
    .Z(_16943_));
 BUF_X1 _34530_ (.A(_00791_),
    .Z(_00192_));
 BUF_X1 _34531_ (.A(text_in[39]),
    .Z(_16944_));
 BUF_X1 _34532_ (.A(_00792_),
    .Z(_00193_));
 BUF_X1 _34533_ (.A(text_in[40]),
    .Z(_16946_));
 BUF_X1 _34534_ (.A(_00794_),
    .Z(_00195_));
 BUF_X1 _34535_ (.A(text_in[41]),
    .Z(_16947_));
 BUF_X1 _34536_ (.A(_00795_),
    .Z(_00196_));
 BUF_X1 _34537_ (.A(text_in[42]),
    .Z(_16948_));
 BUF_X1 _34538_ (.A(_00796_),
    .Z(_00197_));
 BUF_X1 _34539_ (.A(text_in[43]),
    .Z(_16949_));
 BUF_X1 _34540_ (.A(_00797_),
    .Z(_00198_));
 BUF_X1 _34541_ (.A(text_in[44]),
    .Z(_16950_));
 BUF_X1 _34542_ (.A(_00798_),
    .Z(_00199_));
 BUF_X1 _34543_ (.A(text_in[45]),
    .Z(_16951_));
 BUF_X1 _34544_ (.A(_00799_),
    .Z(_00200_));
 BUF_X1 _34545_ (.A(text_in[46]),
    .Z(_16952_));
 BUF_X1 _34546_ (.A(_00800_),
    .Z(_00201_));
 BUF_X1 _34547_ (.A(text_in[47]),
    .Z(_16953_));
 BUF_X1 _34548_ (.A(_00801_),
    .Z(_00202_));
 BUF_X1 _34549_ (.A(text_in[48]),
    .Z(_16954_));
 BUF_X1 _34550_ (.A(_00802_),
    .Z(_00203_));
 BUF_X1 _34551_ (.A(text_in[49]),
    .Z(_16955_));
 BUF_X1 _34552_ (.A(_00803_),
    .Z(_00204_));
 BUF_X1 _34553_ (.A(text_in[50]),
    .Z(_16957_));
 BUF_X1 _34554_ (.A(_00805_),
    .Z(_00206_));
 BUF_X1 _34555_ (.A(text_in[51]),
    .Z(_16958_));
 BUF_X1 _34556_ (.A(_00806_),
    .Z(_00207_));
 BUF_X1 _34557_ (.A(text_in[52]),
    .Z(_16959_));
 BUF_X1 _34558_ (.A(_00807_),
    .Z(_00208_));
 BUF_X1 _34559_ (.A(text_in[53]),
    .Z(_16960_));
 BUF_X1 _34560_ (.A(_00808_),
    .Z(_00209_));
 BUF_X1 _34561_ (.A(text_in[54]),
    .Z(_16961_));
 BUF_X1 _34562_ (.A(_00809_),
    .Z(_00210_));
 BUF_X1 _34563_ (.A(text_in[55]),
    .Z(_16962_));
 BUF_X1 _34564_ (.A(_00810_),
    .Z(_00211_));
 BUF_X1 _34565_ (.A(text_in[56]),
    .Z(_16963_));
 BUF_X1 _34566_ (.A(_00811_),
    .Z(_00212_));
 BUF_X1 _34567_ (.A(text_in[57]),
    .Z(_16964_));
 BUF_X1 _34568_ (.A(_00812_),
    .Z(_00213_));
 BUF_X1 _34569_ (.A(text_in[58]),
    .Z(_16965_));
 BUF_X1 _34570_ (.A(_00813_),
    .Z(_00214_));
 BUF_X1 _34571_ (.A(text_in[59]),
    .Z(_16966_));
 BUF_X1 _34572_ (.A(_00814_),
    .Z(_00215_));
 BUF_X1 _34573_ (.A(text_in[60]),
    .Z(_16968_));
 BUF_X1 _34574_ (.A(_00816_),
    .Z(_00217_));
 BUF_X1 _34575_ (.A(text_in[61]),
    .Z(_16969_));
 BUF_X1 _34576_ (.A(_00817_),
    .Z(_00218_));
 BUF_X1 _34577_ (.A(text_in[62]),
    .Z(_16970_));
 BUF_X1 _34578_ (.A(_00818_),
    .Z(_00219_));
 BUF_X1 _34579_ (.A(text_in[63]),
    .Z(_16971_));
 BUF_X1 _34580_ (.A(_00819_),
    .Z(_00220_));
 BUF_X1 _34581_ (.A(text_in[64]),
    .Z(_16972_));
 BUF_X1 _34582_ (.A(_00820_),
    .Z(_00221_));
 BUF_X1 _34583_ (.A(text_in[65]),
    .Z(_16973_));
 BUF_X1 _34584_ (.A(_00821_),
    .Z(_00222_));
 BUF_X1 _34585_ (.A(text_in[66]),
    .Z(_16974_));
 BUF_X1 _34586_ (.A(_00822_),
    .Z(_00223_));
 BUF_X1 _34587_ (.A(text_in[67]),
    .Z(_16975_));
 BUF_X1 _34588_ (.A(_00823_),
    .Z(_00224_));
 BUF_X1 _34589_ (.A(text_in[68]),
    .Z(_16976_));
 BUF_X1 _34590_ (.A(_00824_),
    .Z(_00225_));
 BUF_X1 _34591_ (.A(text_in[69]),
    .Z(_16977_));
 BUF_X1 _34592_ (.A(_00825_),
    .Z(_00226_));
 BUF_X1 _34593_ (.A(text_in[70]),
    .Z(_16979_));
 BUF_X1 _34594_ (.A(_00827_),
    .Z(_00228_));
 BUF_X1 _34595_ (.A(text_in[71]),
    .Z(_16980_));
 BUF_X1 _34596_ (.A(_00828_),
    .Z(_00229_));
 BUF_X1 _34597_ (.A(text_in[72]),
    .Z(_16981_));
 BUF_X1 _34598_ (.A(_00829_),
    .Z(_00230_));
 BUF_X1 _34599_ (.A(text_in[73]),
    .Z(_16982_));
 BUF_X1 _34600_ (.A(_00830_),
    .Z(_00231_));
 BUF_X1 _34601_ (.A(text_in[74]),
    .Z(_16983_));
 BUF_X1 _34602_ (.A(_00831_),
    .Z(_00232_));
 BUF_X1 _34603_ (.A(text_in[75]),
    .Z(_16984_));
 BUF_X1 _34604_ (.A(_00832_),
    .Z(_00233_));
 BUF_X1 _34605_ (.A(text_in[76]),
    .Z(_16985_));
 BUF_X1 _34606_ (.A(_00833_),
    .Z(_00234_));
 BUF_X1 _34607_ (.A(text_in[77]),
    .Z(_16986_));
 BUF_X1 _34608_ (.A(_00834_),
    .Z(_00235_));
 BUF_X1 _34609_ (.A(text_in[78]),
    .Z(_16987_));
 BUF_X1 _34610_ (.A(_00835_),
    .Z(_00236_));
 BUF_X1 _34611_ (.A(text_in[79]),
    .Z(_16988_));
 BUF_X1 _34612_ (.A(_00836_),
    .Z(_00237_));
 BUF_X1 _34613_ (.A(text_in[80]),
    .Z(_16990_));
 BUF_X1 _34614_ (.A(_00838_),
    .Z(_00239_));
 BUF_X1 _34615_ (.A(text_in[81]),
    .Z(_16991_));
 BUF_X1 _34616_ (.A(_00839_),
    .Z(_00240_));
 BUF_X1 _34617_ (.A(text_in[82]),
    .Z(_16992_));
 BUF_X1 _34618_ (.A(_00840_),
    .Z(_00241_));
 BUF_X1 _34619_ (.A(text_in[83]),
    .Z(_16993_));
 BUF_X1 _34620_ (.A(_00841_),
    .Z(_00242_));
 BUF_X1 _34621_ (.A(text_in[84]),
    .Z(_16994_));
 BUF_X1 _34622_ (.A(_00842_),
    .Z(_00243_));
 BUF_X1 _34623_ (.A(text_in[85]),
    .Z(_16995_));
 BUF_X1 _34624_ (.A(_00843_),
    .Z(_00244_));
 BUF_X1 _34625_ (.A(text_in[86]),
    .Z(_16996_));
 BUF_X1 _34626_ (.A(_00844_),
    .Z(_00245_));
 BUF_X1 _34627_ (.A(text_in[87]),
    .Z(_16997_));
 BUF_X1 _34628_ (.A(_00845_),
    .Z(_00246_));
 BUF_X1 _34629_ (.A(text_in[88]),
    .Z(_16998_));
 BUF_X1 _34630_ (.A(_00846_),
    .Z(_00247_));
 BUF_X1 _34631_ (.A(text_in[89]),
    .Z(_16999_));
 BUF_X1 _34632_ (.A(_00847_),
    .Z(_00248_));
 BUF_X1 _34633_ (.A(text_in[90]),
    .Z(_17001_));
 BUF_X1 _34634_ (.A(_00849_),
    .Z(_00250_));
 BUF_X1 _34635_ (.A(text_in[91]),
    .Z(_17002_));
 BUF_X1 _34636_ (.A(_00850_),
    .Z(_00251_));
 BUF_X1 _34637_ (.A(text_in[92]),
    .Z(_17003_));
 BUF_X1 _34638_ (.A(_00851_),
    .Z(_00252_));
 BUF_X1 _34639_ (.A(text_in[93]),
    .Z(_17004_));
 BUF_X1 _34640_ (.A(_00852_),
    .Z(_00253_));
 BUF_X1 _34641_ (.A(text_in[94]),
    .Z(_17005_));
 BUF_X1 _34642_ (.A(_00853_),
    .Z(_00254_));
 BUF_X1 _34643_ (.A(text_in[95]),
    .Z(_17006_));
 BUF_X1 _34644_ (.A(_00854_),
    .Z(_00255_));
 BUF_X1 _34645_ (.A(\sa00[5] ),
    .Z(_16761_));
 BUF_X1 _34646_ (.A(\sa00[4] ),
    .Z(_16760_));
 BUF_X1 _34647_ (.A(\sa00[7] ),
    .Z(_16763_));
 BUF_X1 _34648_ (.A(\sa00[6] ),
    .Z(_16762_));
 BUF_X1 _34649_ (.A(\sa00[1] ),
    .Z(_16757_));
 BUF_X1 _34650_ (.A(\sa00[0] ),
    .Z(_16756_));
 BUF_X1 _34651_ (.A(\sa00[2] ),
    .Z(_16758_));
 BUF_X1 _34652_ (.A(\sa00[3] ),
    .Z(_16759_));
 BUF_X1 _34653_ (.A(\sa11[5] ),
    .Z(_16801_));
 BUF_X1 _34654_ (.A(\sa11[4] ),
    .Z(_16800_));
 BUF_X1 _34655_ (.A(\sa11[7] ),
    .Z(_16803_));
 BUF_X1 _34656_ (.A(\sa11[6] ),
    .Z(_16802_));
 BUF_X1 _34657_ (.A(\sa11[1] ),
    .Z(_16797_));
 BUF_X1 _34658_ (.A(\sa11[0] ),
    .Z(_16796_));
 BUF_X1 _34659_ (.A(\sa11[2] ),
    .Z(_16798_));
 BUF_X1 _34660_ (.A(\sa11[3] ),
    .Z(_16799_));
 BUF_X1 _34661_ (.A(\sa22[5] ),
    .Z(_16841_));
 BUF_X1 _34662_ (.A(\sa22[4] ),
    .Z(_16840_));
 BUF_X1 _34663_ (.A(\sa22[7] ),
    .Z(_16843_));
 BUF_X1 _34664_ (.A(\sa22[6] ),
    .Z(_16842_));
 BUF_X1 _34665_ (.A(\sa22[1] ),
    .Z(_16837_));
 BUF_X1 _34666_ (.A(\sa22[0] ),
    .Z(_16836_));
 BUF_X1 _34667_ (.A(\sa22[2] ),
    .Z(_16838_));
 BUF_X1 _34668_ (.A(\sa22[3] ),
    .Z(_16839_));
 BUF_X1 _34669_ (.A(\sa33[0] ),
    .Z(_16876_));
 BUF_X1 _34670_ (.A(\sa33[1] ),
    .Z(_16877_));
 BUF_X1 _34671_ (.A(\sa33[3] ),
    .Z(_16879_));
 BUF_X1 _34672_ (.A(\sa33[2] ),
    .Z(_16878_));
 BUF_X1 _34673_ (.A(\sa33[5] ),
    .Z(_16881_));
 BUF_X1 _34674_ (.A(\sa33[4] ),
    .Z(_16880_));
 BUF_X1 _34675_ (.A(\sa33[6] ),
    .Z(_16882_));
 BUF_X1 _34676_ (.A(\sa33[7] ),
    .Z(_16883_));
 BUF_X1 _34677_ (.A(\text_in_r[96] ),
    .Z(_17135_));
 BUF_X1 _34678_ (.A(_00700_),
    .Z(_00101_));
 BUF_X1 _34679_ (.A(text_in[96]),
    .Z(_17007_));
 BUF_X1 _34680_ (.A(_00855_),
    .Z(_00256_));
 BUF_X1 _34681_ (.A(\text_in_r[97] ),
    .Z(_17136_));
 BUF_X1 _34682_ (.A(text_in[97]),
    .Z(_17008_));
 BUF_X1 _34683_ (.A(_00856_),
    .Z(_00257_));
 BUF_X1 _34684_ (.A(\text_in_r[98] ),
    .Z(_17137_));
 BUF_X1 _34685_ (.A(text_in[98]),
    .Z(_17009_));
 BUF_X1 _34686_ (.A(_00857_),
    .Z(_00258_));
 BUF_X1 _34687_ (.A(\text_in_r[99] ),
    .Z(_17138_));
 BUF_X1 _34688_ (.A(text_in[99]),
    .Z(_17010_));
 BUF_X1 _34689_ (.A(_00858_),
    .Z(_00259_));
 BUF_X1 _34690_ (.A(\text_in_r[100] ),
    .Z(_17013_));
 BUF_X1 _34691_ (.A(text_in[100]),
    .Z(_16885_));
 BUF_X1 _34692_ (.A(_00733_),
    .Z(_00134_));
 BUF_X1 _34693_ (.A(\text_in_r[101] ),
    .Z(_17014_));
 BUF_X1 _34694_ (.A(text_in[101]),
    .Z(_16886_));
 BUF_X1 _34695_ (.A(_00734_),
    .Z(_00135_));
 BUF_X1 _34696_ (.A(\text_in_r[102] ),
    .Z(_17015_));
 BUF_X1 _34697_ (.A(text_in[102]),
    .Z(_16887_));
 BUF_X1 _34698_ (.A(_00735_),
    .Z(_00136_));
 BUF_X1 _34699_ (.A(\text_in_r[103] ),
    .Z(_17016_));
 BUF_X1 _34700_ (.A(text_in[103]),
    .Z(_16888_));
 BUF_X1 _34701_ (.A(_00736_),
    .Z(_00137_));
 BUF_X1 _34702_ (.A(\text_in_r[104] ),
    .Z(_17017_));
 BUF_X1 _34703_ (.A(text_in[104]),
    .Z(_16889_));
 BUF_X1 _34704_ (.A(_00737_),
    .Z(_00138_));
 BUF_X1 _34705_ (.A(\text_in_r[105] ),
    .Z(_17018_));
 BUF_X1 _34706_ (.A(text_in[105]),
    .Z(_16890_));
 BUF_X1 _34707_ (.A(_00738_),
    .Z(_00139_));
 BUF_X1 _34708_ (.A(_00701_),
    .Z(_00102_));
 BUF_X1 _34709_ (.A(\text_in_r[106] ),
    .Z(_17019_));
 BUF_X1 _34710_ (.A(text_in[106]),
    .Z(_16891_));
 BUF_X1 _34711_ (.A(_00739_),
    .Z(_00140_));
 BUF_X1 _34712_ (.A(\text_in_r[107] ),
    .Z(_17020_));
 BUF_X1 _34713_ (.A(text_in[107]),
    .Z(_16892_));
 BUF_X1 _34714_ (.A(_00740_),
    .Z(_00141_));
 BUF_X1 _34715_ (.A(\text_in_r[108] ),
    .Z(_17021_));
 BUF_X1 _34716_ (.A(text_in[108]),
    .Z(_16893_));
 BUF_X1 _34717_ (.A(_00741_),
    .Z(_00142_));
 BUF_X1 _34718_ (.A(\text_in_r[109] ),
    .Z(_17022_));
 BUF_X1 _34719_ (.A(text_in[109]),
    .Z(_16894_));
 BUF_X1 _34720_ (.A(_00742_),
    .Z(_00143_));
 BUF_X1 _34721_ (.A(\text_in_r[110] ),
    .Z(_17024_));
 BUF_X1 _34722_ (.A(text_in[110]),
    .Z(_16896_));
 BUF_X1 _34723_ (.A(_00744_),
    .Z(_00145_));
 BUF_X1 _34724_ (.A(\text_in_r[111] ),
    .Z(_17025_));
 BUF_X1 _34725_ (.A(text_in[111]),
    .Z(_16897_));
 BUF_X1 _34726_ (.A(_00745_),
    .Z(_00146_));
 BUF_X1 _34727_ (.A(\text_in_r[112] ),
    .Z(_17026_));
 BUF_X1 _34728_ (.A(text_in[112]),
    .Z(_16898_));
 BUF_X1 _34729_ (.A(_00746_),
    .Z(_00147_));
 BUF_X1 _34730_ (.A(\text_in_r[113] ),
    .Z(_17027_));
 BUF_X1 _34731_ (.A(text_in[113]),
    .Z(_16899_));
 BUF_X1 _34732_ (.A(_00747_),
    .Z(_00148_));
 BUF_X1 _34733_ (.A(\text_in_r[114] ),
    .Z(_17028_));
 BUF_X1 _34734_ (.A(text_in[114]),
    .Z(_16900_));
 BUF_X1 _34735_ (.A(_00748_),
    .Z(_00149_));
 BUF_X1 _34736_ (.A(\text_in_r[115] ),
    .Z(_17029_));
 BUF_X1 _34737_ (.A(text_in[115]),
    .Z(_16901_));
 BUF_X1 _34738_ (.A(_00749_),
    .Z(_00150_));
 BUF_X1 _34739_ (.A(_00702_),
    .Z(_00103_));
 BUF_X1 _34740_ (.A(\text_in_r[116] ),
    .Z(_17030_));
 BUF_X1 _34741_ (.A(text_in[116]),
    .Z(_16902_));
 BUF_X1 _34742_ (.A(_00750_),
    .Z(_00151_));
 BUF_X1 _34743_ (.A(\text_in_r[117] ),
    .Z(_17031_));
 BUF_X1 _34744_ (.A(text_in[117]),
    .Z(_16903_));
 BUF_X1 _34745_ (.A(_00751_),
    .Z(_00152_));
 BUF_X1 _34746_ (.A(\text_in_r[118] ),
    .Z(_17032_));
 BUF_X1 _34747_ (.A(text_in[118]),
    .Z(_16904_));
 BUF_X1 _34748_ (.A(_00752_),
    .Z(_00153_));
 BUF_X1 _34749_ (.A(\text_in_r[119] ),
    .Z(_17033_));
 BUF_X1 _34750_ (.A(text_in[119]),
    .Z(_16905_));
 BUF_X1 _34751_ (.A(_00753_),
    .Z(_00154_));
 BUF_X1 _34752_ (.A(\text_in_r[120] ),
    .Z(_17035_));
 BUF_X1 _34753_ (.A(text_in[120]),
    .Z(_16907_));
 BUF_X1 _34754_ (.A(_00755_),
    .Z(_00156_));
 BUF_X1 _34755_ (.A(\text_in_r[121] ),
    .Z(_17036_));
 BUF_X1 _34756_ (.A(text_in[121]),
    .Z(_16908_));
 BUF_X1 _34757_ (.A(_00756_),
    .Z(_00157_));
 BUF_X1 _34758_ (.A(\text_in_r[122] ),
    .Z(_17037_));
 BUF_X1 _34759_ (.A(text_in[122]),
    .Z(_16909_));
 BUF_X1 _34760_ (.A(_00757_),
    .Z(_00158_));
 BUF_X1 _34761_ (.A(\text_in_r[123] ),
    .Z(_17038_));
 BUF_X1 _34762_ (.A(text_in[123]),
    .Z(_16910_));
 BUF_X1 _34763_ (.A(_00758_),
    .Z(_00159_));
 BUF_X1 _34764_ (.A(\text_in_r[124] ),
    .Z(_17039_));
 BUF_X1 _34765_ (.A(text_in[124]),
    .Z(_16911_));
 BUF_X1 _34766_ (.A(_00759_),
    .Z(_00160_));
 BUF_X1 _34767_ (.A(\text_in_r[125] ),
    .Z(_17040_));
 BUF_X1 _34768_ (.A(text_in[125]),
    .Z(_16912_));
 BUF_X1 _34769_ (.A(_00760_),
    .Z(_00161_));
 BUF_X1 _34770_ (.A(_00703_),
    .Z(_00104_));
 BUF_X1 _34771_ (.A(\text_in_r[126] ),
    .Z(_17041_));
 BUF_X1 _34772_ (.A(text_in[126]),
    .Z(_16913_));
 BUF_X1 _34773_ (.A(_00761_),
    .Z(_00162_));
 BUF_X1 _34774_ (.A(\text_in_r[127] ),
    .Z(_17042_));
 BUF_X1 _34775_ (.A(text_in[127]),
    .Z(_16914_));
 BUF_X1 _34776_ (.A(_00762_),
    .Z(_00163_));
 BUF_X1 _34777_ (.A(_00704_),
    .Z(_00105_));
 BUF_X1 _34778_ (.A(_00705_),
    .Z(_00106_));
 BUF_X1 _34779_ (.A(_00706_),
    .Z(_00107_));
 BUF_X1 _34780_ (.A(_00707_),
    .Z(_00108_));
 BUF_X1 _34781_ (.A(_00668_),
    .Z(_00069_));
 BUF_X1 _34782_ (.A(_00669_),
    .Z(_00070_));
 BUF_X1 _34783_ (.A(_00670_),
    .Z(_00071_));
 BUF_X1 _34784_ (.A(_00671_),
    .Z(_00072_));
 BUF_X1 _34785_ (.A(_00672_),
    .Z(_00073_));
 BUF_X1 _34786_ (.A(_00673_),
    .Z(_00074_));
 BUF_X1 _34787_ (.A(_00674_),
    .Z(_00075_));
 BUF_X1 _34788_ (.A(_00675_),
    .Z(_00076_));
 BUF_X1 _34789_ (.A(_00636_),
    .Z(_00037_));
 BUF_X1 _34790_ (.A(_00637_),
    .Z(_00038_));
 BUF_X1 _34791_ (.A(_00638_),
    .Z(_00039_));
 BUF_X1 _34792_ (.A(_00639_),
    .Z(_00040_));
 BUF_X1 _34793_ (.A(_00640_),
    .Z(_00041_));
 BUF_X1 _34794_ (.A(_00641_),
    .Z(_00042_));
 BUF_X1 _34795_ (.A(_00642_),
    .Z(_00043_));
 BUF_X1 _34796_ (.A(_00643_),
    .Z(_00044_));
 BUF_X1 _34797_ (.A(_00604_),
    .Z(_00005_));
 BUF_X1 _34798_ (.A(_00605_),
    .Z(_00006_));
 BUF_X1 _34799_ (.A(_00606_),
    .Z(_00007_));
 BUF_X1 _34800_ (.A(_00607_),
    .Z(_00008_));
 BUF_X1 _34801_ (.A(_00608_),
    .Z(_00009_));
 BUF_X1 _34802_ (.A(_00609_),
    .Z(_00010_));
 BUF_X1 _34803_ (.A(_00610_),
    .Z(_00011_));
 BUF_X1 _34804_ (.A(_00611_),
    .Z(_00012_));
 BUF_X1 _34805_ (.A(_00603_),
    .Z(_00004_));
 BUF_X1 _34806_ (.A(_00884_),
    .Z(_00285_));
 BUF_X1 _34807_ (.A(_00885_),
    .Z(_00286_));
 BUF_X1 _34808_ (.A(_00886_),
    .Z(_00287_));
 BUF_X1 _34809_ (.A(_00887_),
    .Z(_00288_));
 BUF_X1 _34810_ (.A(_00888_),
    .Z(_00289_));
 BUF_X1 _34811_ (.A(_00889_),
    .Z(_00290_));
 BUF_X1 _34812_ (.A(_00890_),
    .Z(_00291_));
 BUF_X1 _34813_ (.A(_00891_),
    .Z(_00292_));
 BUF_X1 _34814_ (.A(_00980_),
    .Z(_00381_));
 BUF_X1 _34815_ (.A(_00981_),
    .Z(_00382_));
 BUF_X1 _34816_ (.A(_00982_),
    .Z(_00383_));
 BUF_X1 _34817_ (.A(_00983_),
    .Z(_00384_));
 BUF_X1 _34818_ (.A(_00984_),
    .Z(_00385_));
 BUF_X1 _34819_ (.A(_00985_),
    .Z(_00386_));
 BUF_X1 _34820_ (.A(_00986_),
    .Z(_00387_));
 BUF_X1 _34821_ (.A(_00987_),
    .Z(_00388_));
 BUF_X1 _34822_ (.A(_00940_),
    .Z(_00341_));
 BUF_X1 _34823_ (.A(_00941_),
    .Z(_00342_));
 BUF_X1 _34824_ (.A(_00942_),
    .Z(_00343_));
 BUF_X1 _34825_ (.A(_00943_),
    .Z(_00344_));
 BUF_X1 _34826_ (.A(_00944_),
    .Z(_00345_));
 BUF_X1 _34827_ (.A(_00945_),
    .Z(_00346_));
 BUF_X1 _34828_ (.A(_00946_),
    .Z(_00347_));
 BUF_X1 _34829_ (.A(_00947_),
    .Z(_00348_));
 BUF_X1 _34830_ (.A(_00908_),
    .Z(_00309_));
 BUF_X1 _34831_ (.A(_00909_),
    .Z(_00310_));
 BUF_X1 _34832_ (.A(_00910_),
    .Z(_00311_));
 BUF_X1 _34833_ (.A(_00911_),
    .Z(_00312_));
 BUF_X1 _34834_ (.A(_00912_),
    .Z(_00313_));
 BUF_X1 _34835_ (.A(_00913_),
    .Z(_00314_));
 BUF_X1 _34836_ (.A(_00914_),
    .Z(_00315_));
 BUF_X1 _34837_ (.A(_00915_),
    .Z(_00316_));
 BUF_X1 _34838_ (.A(_00876_),
    .Z(_00277_));
 BUF_X1 _34839_ (.A(_00877_),
    .Z(_00278_));
 BUF_X1 _34840_ (.A(_00878_),
    .Z(_00279_));
 BUF_X1 _34841_ (.A(_00879_),
    .Z(_00280_));
 BUF_X1 _34842_ (.A(_00880_),
    .Z(_00281_));
 BUF_X1 _34843_ (.A(_00881_),
    .Z(_00282_));
 BUF_X1 _34844_ (.A(_00882_),
    .Z(_00283_));
 BUF_X1 _34845_ (.A(_00883_),
    .Z(_00284_));
 BUF_X1 _34846_ (.A(_00972_),
    .Z(_00373_));
 BUF_X1 _34847_ (.A(_00973_),
    .Z(_00374_));
 BUF_X1 _34848_ (.A(_00974_),
    .Z(_00375_));
 BUF_X1 _34849_ (.A(_00975_),
    .Z(_00376_));
 BUF_X1 _34850_ (.A(_00976_),
    .Z(_00377_));
 BUF_X1 _34851_ (.A(_00977_),
    .Z(_00378_));
 BUF_X1 _34852_ (.A(_00978_),
    .Z(_00379_));
 BUF_X1 _34853_ (.A(_00979_),
    .Z(_00380_));
 BUF_X1 _34854_ (.A(_00932_),
    .Z(_00333_));
 BUF_X1 _34855_ (.A(_00933_),
    .Z(_00334_));
 BUF_X1 _34856_ (.A(_00934_),
    .Z(_00335_));
 BUF_X1 _34857_ (.A(_00935_),
    .Z(_00336_));
 BUF_X1 _34858_ (.A(_00936_),
    .Z(_00337_));
 BUF_X1 _34859_ (.A(_00937_),
    .Z(_00338_));
 BUF_X1 _34860_ (.A(_00938_),
    .Z(_00339_));
 BUF_X1 _34861_ (.A(_00939_),
    .Z(_00340_));
 BUF_X1 _34862_ (.A(_00900_),
    .Z(_00301_));
 BUF_X1 _34863_ (.A(_00901_),
    .Z(_00302_));
 BUF_X1 _34864_ (.A(_00902_),
    .Z(_00303_));
 BUF_X1 _34865_ (.A(_00903_),
    .Z(_00304_));
 BUF_X1 _34866_ (.A(_00904_),
    .Z(_00305_));
 BUF_X1 _34867_ (.A(_00905_),
    .Z(_00306_));
 BUF_X1 _34868_ (.A(_00906_),
    .Z(_00307_));
 BUF_X1 _34869_ (.A(_00907_),
    .Z(_00308_));
 BUF_X1 _34870_ (.A(_00868_),
    .Z(_00269_));
 BUF_X1 _34871_ (.A(_00869_),
    .Z(_00270_));
 BUF_X1 _34872_ (.A(_00870_),
    .Z(_00271_));
 BUF_X1 _34873_ (.A(_00871_),
    .Z(_00272_));
 BUF_X1 _34874_ (.A(_00872_),
    .Z(_00273_));
 BUF_X1 _34875_ (.A(_00873_),
    .Z(_00274_));
 BUF_X1 _34876_ (.A(_00874_),
    .Z(_00275_));
 BUF_X1 _34877_ (.A(_00875_),
    .Z(_00276_));
 BUF_X1 _34878_ (.A(_00956_),
    .Z(_00357_));
 BUF_X1 _34879_ (.A(_00957_),
    .Z(_00358_));
 BUF_X1 _34880_ (.A(_00958_),
    .Z(_00359_));
 BUF_X1 _34881_ (.A(_00959_),
    .Z(_00360_));
 BUF_X1 _34882_ (.A(_00960_),
    .Z(_00361_));
 BUF_X1 _34883_ (.A(_00961_),
    .Z(_00362_));
 BUF_X1 _34884_ (.A(_00962_),
    .Z(_00363_));
 BUF_X1 _34885_ (.A(_00963_),
    .Z(_00364_));
 BUF_X1 _34886_ (.A(_00924_),
    .Z(_00325_));
 BUF_X1 _34887_ (.A(_00925_),
    .Z(_00326_));
 BUF_X1 _34888_ (.A(_00926_),
    .Z(_00327_));
 BUF_X1 _34889_ (.A(_00927_),
    .Z(_00328_));
 BUF_X1 _34890_ (.A(_00928_),
    .Z(_00329_));
 BUF_X1 _34891_ (.A(_00929_),
    .Z(_00330_));
 BUF_X1 _34892_ (.A(_00930_),
    .Z(_00331_));
 BUF_X1 _34893_ (.A(_00931_),
    .Z(_00332_));
 BUF_X1 _34894_ (.A(_00892_),
    .Z(_00293_));
 BUF_X1 _34895_ (.A(_00893_),
    .Z(_00294_));
 BUF_X1 _34896_ (.A(_00894_),
    .Z(_00295_));
 BUF_X1 _34897_ (.A(_00895_),
    .Z(_00296_));
 BUF_X1 _34898_ (.A(_00896_),
    .Z(_00297_));
 BUF_X1 _34899_ (.A(_00897_),
    .Z(_00298_));
 BUF_X1 _34900_ (.A(_00898_),
    .Z(_00299_));
 BUF_X1 _34901_ (.A(_00899_),
    .Z(_00300_));
 BUF_X1 _34902_ (.A(_00860_),
    .Z(_00261_));
 BUF_X1 _34903_ (.A(_00861_),
    .Z(_00262_));
 BUF_X1 _34904_ (.A(_00862_),
    .Z(_00263_));
 BUF_X1 _34905_ (.A(_00863_),
    .Z(_00264_));
 BUF_X1 _34906_ (.A(_00864_),
    .Z(_00265_));
 BUF_X1 _34907_ (.A(_00865_),
    .Z(_00266_));
 BUF_X1 _34908_ (.A(_00866_),
    .Z(_00267_));
 BUF_X1 _34909_ (.A(_00867_),
    .Z(_00268_));
 BUF_X1 _34910_ (.A(_00948_),
    .Z(_00349_));
 BUF_X1 _34911_ (.A(_00949_),
    .Z(_00350_));
 BUF_X1 _34912_ (.A(_00950_),
    .Z(_00351_));
 BUF_X1 _34913_ (.A(_00951_),
    .Z(_00352_));
 BUF_X1 _34914_ (.A(_00952_),
    .Z(_00353_));
 BUF_X1 _34915_ (.A(_00953_),
    .Z(_00354_));
 BUF_X1 _34916_ (.A(_00954_),
    .Z(_00355_));
 BUF_X1 _34917_ (.A(_00955_),
    .Z(_00356_));
 BUF_X1 _34918_ (.A(_00916_),
    .Z(_00317_));
 BUF_X1 _34919_ (.A(_00917_),
    .Z(_00318_));
 BUF_X1 _34920_ (.A(_00918_),
    .Z(_00319_));
 BUF_X1 _34921_ (.A(_00919_),
    .Z(_00320_));
 BUF_X1 _34922_ (.A(_00920_),
    .Z(_00321_));
 BUF_X1 _34923_ (.A(_00921_),
    .Z(_00322_));
 BUF_X1 _34924_ (.A(_00922_),
    .Z(_00323_));
 BUF_X1 _34925_ (.A(_00923_),
    .Z(_00324_));
 BUF_X1 _34926_ (.A(_00964_),
    .Z(_00365_));
 BUF_X1 _34927_ (.A(_00965_),
    .Z(_00366_));
 BUF_X1 _34928_ (.A(_00966_),
    .Z(_00367_));
 BUF_X1 _34929_ (.A(_00967_),
    .Z(_00368_));
 BUF_X1 _34930_ (.A(_00968_),
    .Z(_00369_));
 BUF_X1 _34931_ (.A(_00969_),
    .Z(_00370_));
 BUF_X1 _34932_ (.A(_00970_),
    .Z(_00371_));
 BUF_X1 _34933_ (.A(_00971_),
    .Z(_00372_));
 DFF_X1 _34934_ (.D(_00595_),
    .CK(clk),
    .Q(\u0.r0.rcnt[0] ),
    .QN(_17272_));
 DFF_X1 _34935_ (.D(_00596_),
    .CK(clk),
    .Q(\u0.r0.rcnt[1] ),
    .QN(_17273_));
 DFF_X1 _34936_ (.D(_00597_),
    .CK(clk),
    .Q(\u0.r0.rcnt[2] ),
    .QN(_17274_));
 DFF_X1 _34937_ (.D(_00598_),
    .CK(clk),
    .Q(\u0.r0.rcnt[3] ),
    .QN(_17275_));
 DFF_X1 _34938_ (.D(_00587_),
    .CK(clk),
    .Q(\u0.r0.out[24] ),
    .QN(_00414_));
 DFF_X1 _34939_ (.D(_00588_),
    .CK(clk),
    .Q(\u0.r0.out[25] ),
    .QN(_00416_));
 DFF_X1 _34940_ (.D(_00589_),
    .CK(clk),
    .Q(\u0.r0.out[26] ),
    .QN(_00418_));
 DFF_X1 _34941_ (.D(_00590_),
    .CK(clk),
    .Q(\u0.r0.out[27] ),
    .QN(_00420_));
 DFF_X1 _34942_ (.D(_00591_),
    .CK(clk),
    .Q(\u0.r0.out[28] ),
    .QN(_00422_));
 DFF_X1 _34943_ (.D(_00592_),
    .CK(clk),
    .Q(\u0.r0.out[29] ),
    .QN(_00424_));
 DFF_X1 _34944_ (.D(_00593_),
    .CK(clk),
    .Q(\u0.r0.out[30] ),
    .QN(_00426_));
 DFF_X1 _34945_ (.D(_00594_),
    .CK(clk),
    .Q(\u0.r0.out[31] ),
    .QN(_00428_));
 DFF_X1 _34946_ (.D(_00555_),
    .CK(clk),
    .Q(\u0.tmp_w[0] ),
    .QN(_17276_));
 DFF_X1 _34947_ (.D(_00566_),
    .CK(clk),
    .Q(\u0.tmp_w[1] ),
    .QN(_17277_));
 DFF_X1 _34948_ (.D(_00577_),
    .CK(clk),
    .Q(\u0.tmp_w[2] ),
    .QN(_17278_));
 DFF_X1 _34949_ (.D(_00580_),
    .CK(clk),
    .Q(\u0.tmp_w[3] ),
    .QN(_17279_));
 DFF_X1 _34950_ (.D(_00581_),
    .CK(clk),
    .Q(\u0.tmp_w[4] ),
    .QN(_17280_));
 DFF_X1 _34951_ (.D(_00582_),
    .CK(clk),
    .Q(\u0.tmp_w[5] ),
    .QN(_17281_));
 DFF_X1 _34952_ (.D(_00583_),
    .CK(clk),
    .Q(\u0.tmp_w[6] ),
    .QN(_17282_));
 DFF_X1 _34953_ (.D(_00584_),
    .CK(clk),
    .Q(\u0.tmp_w[7] ),
    .QN(_17283_));
 DFF_X1 _34954_ (.D(_00585_),
    .CK(clk),
    .Q(\u0.tmp_w[8] ),
    .QN(_00450_));
 DFF_X1 _34955_ (.D(_00586_),
    .CK(clk),
    .Q(\u0.tmp_w[9] ),
    .QN(_17284_));
 DFF_X1 _34956_ (.D(_00556_),
    .CK(clk),
    .Q(\u0.tmp_w[10] ),
    .QN(_17285_));
 DFF_X1 _34957_ (.D(_00557_),
    .CK(clk),
    .Q(\u0.tmp_w[11] ),
    .QN(_17286_));
 DFF_X1 _34958_ (.D(_00558_),
    .CK(clk),
    .Q(\u0.tmp_w[12] ),
    .QN(_17287_));
 DFF_X1 _34959_ (.D(_00559_),
    .CK(clk),
    .Q(\u0.tmp_w[13] ),
    .QN(_17288_));
 DFF_X1 _34960_ (.D(_00560_),
    .CK(clk),
    .Q(\u0.tmp_w[14] ),
    .QN(_17289_));
 DFF_X1 _34961_ (.D(_00561_),
    .CK(clk),
    .Q(\u0.tmp_w[15] ),
    .QN(_17290_));
 DFF_X1 _34962_ (.D(_00562_),
    .CK(clk),
    .Q(\u0.tmp_w[16] ),
    .QN(_00451_));
 DFF_X1 _34963_ (.D(_00563_),
    .CK(clk),
    .Q(\u0.tmp_w[17] ),
    .QN(_00452_));
 DFF_X1 _34964_ (.D(_00564_),
    .CK(clk),
    .Q(\u0.tmp_w[18] ),
    .QN(_17291_));
 DFF_X1 _34965_ (.D(_00565_),
    .CK(clk),
    .Q(\u0.tmp_w[19] ),
    .QN(_17292_));
 DFF_X1 _34966_ (.D(_00567_),
    .CK(clk),
    .Q(\u0.tmp_w[20] ),
    .QN(_17293_));
 DFF_X1 _34967_ (.D(_00568_),
    .CK(clk),
    .Q(\u0.tmp_w[21] ),
    .QN(_00453_));
 DFF_X1 _34968_ (.D(_00569_),
    .CK(clk),
    .Q(\u0.tmp_w[22] ),
    .QN(_00454_));
 DFF_X1 _34969_ (.D(_00570_),
    .CK(clk),
    .Q(\u0.tmp_w[23] ),
    .QN(_17294_));
 DFF_X1 _34970_ (.D(_00571_),
    .CK(clk),
    .Q(\u0.tmp_w[24] ),
    .QN(_00455_));
 DFF_X1 _34971_ (.D(_00572_),
    .CK(clk),
    .Q(\u0.tmp_w[25] ),
    .QN(_00456_));
 DFF_X1 _34972_ (.D(_00573_),
    .CK(clk),
    .Q(\u0.tmp_w[26] ),
    .QN(_17295_));
 DFF_X1 _34973_ (.D(_00574_),
    .CK(clk),
    .Q(\u0.tmp_w[27] ),
    .QN(_17296_));
 DFF_X1 _34974_ (.D(_00575_),
    .CK(clk),
    .Q(\u0.tmp_w[28] ),
    .QN(_17297_));
 DFF_X1 _34975_ (.D(_00576_),
    .CK(clk),
    .Q(\u0.tmp_w[29] ),
    .QN(_00457_));
 DFF_X1 _34976_ (.D(_00578_),
    .CK(clk),
    .Q(\u0.tmp_w[30] ),
    .QN(_00458_));
 DFF_X1 _34977_ (.D(_00579_),
    .CK(clk),
    .Q(\u0.tmp_w[31] ),
    .QN(_17298_));
 DFF_X1 _34978_ (.D(_00000_),
    .CK(clk),
    .Q(\dcnt[0] ),
    .QN(_17299_));
 DFF_X1 _34979_ (.D(_00001_),
    .CK(clk),
    .Q(\dcnt[1] ),
    .QN(_00446_));
 DFF_X1 _34980_ (.D(_00002_),
    .CK(clk),
    .Q(\dcnt[2] ),
    .QN(_00447_));
 DFF_X1 _34981_ (.D(_00003_),
    .CK(clk),
    .Q(\dcnt[3] ),
    .QN(_00448_));
 DFF_X1 _34982_ (.D(_00004_),
    .CK(clk),
    .Q(done),
    .QN(_17300_));
 DFF_X1 _34983_ (.D(_00133_),
    .CK(clk),
    .Q(\text_in_r[0] ),
    .QN(_17301_));
 DFF_X1 _34984_ (.D(_00172_),
    .CK(clk),
    .Q(\text_in_r[1] ),
    .QN(_17302_));
 DFF_X1 _34985_ (.D(_00183_),
    .CK(clk),
    .Q(\text_in_r[2] ),
    .QN(_17303_));
 DFF_X1 _34986_ (.D(_00194_),
    .CK(clk),
    .Q(\text_in_r[3] ),
    .QN(_17304_));
 DFF_X1 _34987_ (.D(_00205_),
    .CK(clk),
    .Q(\text_in_r[4] ),
    .QN(_17305_));
 DFF_X1 _34988_ (.D(_00216_),
    .CK(clk),
    .Q(\text_in_r[5] ),
    .QN(_17306_));
 DFF_X1 _34989_ (.D(_00227_),
    .CK(clk),
    .Q(\text_in_r[6] ),
    .QN(_17307_));
 DFF_X1 _34990_ (.D(_00238_),
    .CK(clk),
    .Q(\text_in_r[7] ),
    .QN(_17308_));
 DFF_X1 _34991_ (.D(_00249_),
    .CK(clk),
    .Q(\text_in_r[8] ),
    .QN(_17309_));
 DFF_X1 _34992_ (.D(_00260_),
    .CK(clk),
    .Q(\text_in_r[9] ),
    .QN(_17310_));
 DFF_X1 _34993_ (.D(_00144_),
    .CK(clk),
    .Q(\text_in_r[10] ),
    .QN(_17311_));
 DFF_X1 _34994_ (.D(_00155_),
    .CK(clk),
    .Q(\text_in_r[11] ),
    .QN(_17312_));
 DFF_X1 _34995_ (.D(_00164_),
    .CK(clk),
    .Q(\text_in_r[12] ),
    .QN(_17313_));
 DFF_X1 _34996_ (.D(_00165_),
    .CK(clk),
    .Q(\text_in_r[13] ),
    .QN(_17314_));
 DFF_X1 _34997_ (.D(_00166_),
    .CK(clk),
    .Q(\text_in_r[14] ),
    .QN(_17315_));
 DFF_X1 _34998_ (.D(_00167_),
    .CK(clk),
    .Q(\text_in_r[15] ),
    .QN(_17316_));
 DFF_X1 _34999_ (.D(_00168_),
    .CK(clk),
    .Q(\text_in_r[16] ),
    .QN(_17317_));
 DFF_X1 _35000_ (.D(_00169_),
    .CK(clk),
    .Q(\text_in_r[17] ),
    .QN(_17318_));
 DFF_X1 _35001_ (.D(_00170_),
    .CK(clk),
    .Q(\text_in_r[18] ),
    .QN(_17319_));
 DFF_X1 _35002_ (.D(_00171_),
    .CK(clk),
    .Q(\text_in_r[19] ),
    .QN(_17320_));
 DFF_X1 _35003_ (.D(_00173_),
    .CK(clk),
    .Q(\text_in_r[20] ),
    .QN(_17321_));
 DFF_X1 _35004_ (.D(_00174_),
    .CK(clk),
    .Q(\text_in_r[21] ),
    .QN(_17322_));
 DFF_X1 _35005_ (.D(_00175_),
    .CK(clk),
    .Q(\text_in_r[22] ),
    .QN(_17323_));
 DFF_X1 _35006_ (.D(_00176_),
    .CK(clk),
    .Q(\text_in_r[23] ),
    .QN(_17324_));
 DFF_X1 _35007_ (.D(_00177_),
    .CK(clk),
    .Q(\text_in_r[24] ),
    .QN(_17325_));
 DFF_X1 _35008_ (.D(_00178_),
    .CK(clk),
    .Q(\text_in_r[25] ),
    .QN(_17326_));
 DFF_X1 _35009_ (.D(_00179_),
    .CK(clk),
    .Q(\text_in_r[26] ),
    .QN(_17327_));
 DFF_X1 _35010_ (.D(_00180_),
    .CK(clk),
    .Q(\text_in_r[27] ),
    .QN(_17328_));
 DFF_X1 _35011_ (.D(_00181_),
    .CK(clk),
    .Q(\text_in_r[28] ),
    .QN(_17329_));
 DFF_X1 _35012_ (.D(_00182_),
    .CK(clk),
    .Q(\text_in_r[29] ),
    .QN(_17330_));
 DFF_X1 _35013_ (.D(_00184_),
    .CK(clk),
    .Q(\text_in_r[30] ),
    .QN(_17331_));
 DFF_X1 _35014_ (.D(_00185_),
    .CK(clk),
    .Q(\text_in_r[31] ),
    .QN(_17332_));
 DFF_X1 _35015_ (.D(_00186_),
    .CK(clk),
    .Q(\text_in_r[32] ),
    .QN(_17333_));
 DFF_X1 _35016_ (.D(_00187_),
    .CK(clk),
    .Q(\text_in_r[33] ),
    .QN(_17334_));
 DFF_X1 _35017_ (.D(_00188_),
    .CK(clk),
    .Q(\text_in_r[34] ),
    .QN(_17335_));
 DFF_X1 _35018_ (.D(_00189_),
    .CK(clk),
    .Q(\text_in_r[35] ),
    .QN(_17336_));
 DFF_X1 _35019_ (.D(_00190_),
    .CK(clk),
    .Q(\text_in_r[36] ),
    .QN(_17337_));
 DFF_X1 _35020_ (.D(_00191_),
    .CK(clk),
    .Q(\text_in_r[37] ),
    .QN(_17338_));
 DFF_X1 _35021_ (.D(_00192_),
    .CK(clk),
    .Q(\text_in_r[38] ),
    .QN(_17339_));
 DFF_X1 _35022_ (.D(_00193_),
    .CK(clk),
    .Q(\text_in_r[39] ),
    .QN(_17340_));
 DFF_X1 _35023_ (.D(_00195_),
    .CK(clk),
    .Q(\text_in_r[40] ),
    .QN(_17341_));
 DFF_X1 _35024_ (.D(_00196_),
    .CK(clk),
    .Q(\text_in_r[41] ),
    .QN(_17342_));
 DFF_X1 _35025_ (.D(_00197_),
    .CK(clk),
    .Q(\text_in_r[42] ),
    .QN(_17343_));
 DFF_X1 _35026_ (.D(_00198_),
    .CK(clk),
    .Q(\text_in_r[43] ),
    .QN(_17344_));
 DFF_X1 _35027_ (.D(_00199_),
    .CK(clk),
    .Q(\text_in_r[44] ),
    .QN(_17345_));
 DFF_X1 _35028_ (.D(_00200_),
    .CK(clk),
    .Q(\text_in_r[45] ),
    .QN(_17346_));
 DFF_X1 _35029_ (.D(_00201_),
    .CK(clk),
    .Q(\text_in_r[46] ),
    .QN(_17347_));
 DFF_X1 _35030_ (.D(_00202_),
    .CK(clk),
    .Q(\text_in_r[47] ),
    .QN(_17348_));
 DFF_X1 _35031_ (.D(_00203_),
    .CK(clk),
    .Q(\text_in_r[48] ),
    .QN(_17349_));
 DFF_X1 _35032_ (.D(_00204_),
    .CK(clk),
    .Q(\text_in_r[49] ),
    .QN(_17350_));
 DFF_X1 _35033_ (.D(_00206_),
    .CK(clk),
    .Q(\text_in_r[50] ),
    .QN(_17351_));
 DFF_X1 _35034_ (.D(_00207_),
    .CK(clk),
    .Q(\text_in_r[51] ),
    .QN(_17352_));
 DFF_X1 _35035_ (.D(_00208_),
    .CK(clk),
    .Q(\text_in_r[52] ),
    .QN(_17353_));
 DFF_X1 _35036_ (.D(_00209_),
    .CK(clk),
    .Q(\text_in_r[53] ),
    .QN(_17354_));
 DFF_X1 _35037_ (.D(_00210_),
    .CK(clk),
    .Q(\text_in_r[54] ),
    .QN(_17355_));
 DFF_X1 _35038_ (.D(_00211_),
    .CK(clk),
    .Q(\text_in_r[55] ),
    .QN(_17356_));
 DFF_X1 _35039_ (.D(_00212_),
    .CK(clk),
    .Q(\text_in_r[56] ),
    .QN(_17357_));
 DFF_X1 _35040_ (.D(_00213_),
    .CK(clk),
    .Q(\text_in_r[57] ),
    .QN(_17358_));
 DFF_X1 _35041_ (.D(_00214_),
    .CK(clk),
    .Q(\text_in_r[58] ),
    .QN(_17359_));
 DFF_X1 _35042_ (.D(_00215_),
    .CK(clk),
    .Q(\text_in_r[59] ),
    .QN(_17360_));
 DFF_X1 _35043_ (.D(_00217_),
    .CK(clk),
    .Q(\text_in_r[60] ),
    .QN(_17361_));
 DFF_X1 _35044_ (.D(_00218_),
    .CK(clk),
    .Q(\text_in_r[61] ),
    .QN(_17362_));
 DFF_X1 _35045_ (.D(_00219_),
    .CK(clk),
    .Q(\text_in_r[62] ),
    .QN(_17363_));
 DFF_X1 _35046_ (.D(_00220_),
    .CK(clk),
    .Q(\text_in_r[63] ),
    .QN(_17364_));
 DFF_X1 _35047_ (.D(_00221_),
    .CK(clk),
    .Q(\text_in_r[64] ),
    .QN(_17365_));
 DFF_X1 _35048_ (.D(_00222_),
    .CK(clk),
    .Q(\text_in_r[65] ),
    .QN(_17366_));
 DFF_X1 _35049_ (.D(_00223_),
    .CK(clk),
    .Q(\text_in_r[66] ),
    .QN(_17367_));
 DFF_X1 _35050_ (.D(_00224_),
    .CK(clk),
    .Q(\text_in_r[67] ),
    .QN(_17368_));
 DFF_X1 _35051_ (.D(_00225_),
    .CK(clk),
    .Q(\text_in_r[68] ),
    .QN(_17369_));
 DFF_X1 _35052_ (.D(_00226_),
    .CK(clk),
    .Q(\text_in_r[69] ),
    .QN(_17370_));
 DFF_X1 _35053_ (.D(_00228_),
    .CK(clk),
    .Q(\text_in_r[70] ),
    .QN(_17371_));
 DFF_X1 _35054_ (.D(_00229_),
    .CK(clk),
    .Q(\text_in_r[71] ),
    .QN(_17372_));
 DFF_X1 _35055_ (.D(_00230_),
    .CK(clk),
    .Q(\text_in_r[72] ),
    .QN(_17373_));
 DFF_X1 _35056_ (.D(_00231_),
    .CK(clk),
    .Q(\text_in_r[73] ),
    .QN(_17374_));
 DFF_X1 _35057_ (.D(_00232_),
    .CK(clk),
    .Q(\text_in_r[74] ),
    .QN(_17375_));
 DFF_X1 _35058_ (.D(_00233_),
    .CK(clk),
    .Q(\text_in_r[75] ),
    .QN(_17376_));
 DFF_X1 _35059_ (.D(_00234_),
    .CK(clk),
    .Q(\text_in_r[76] ),
    .QN(_17377_));
 DFF_X1 _35060_ (.D(_00235_),
    .CK(clk),
    .Q(\text_in_r[77] ),
    .QN(_17378_));
 DFF_X1 _35061_ (.D(_00236_),
    .CK(clk),
    .Q(\text_in_r[78] ),
    .QN(_17379_));
 DFF_X1 _35062_ (.D(_00237_),
    .CK(clk),
    .Q(\text_in_r[79] ),
    .QN(_17380_));
 DFF_X1 _35063_ (.D(_00239_),
    .CK(clk),
    .Q(\text_in_r[80] ),
    .QN(_17381_));
 DFF_X1 _35064_ (.D(_00240_),
    .CK(clk),
    .Q(\text_in_r[81] ),
    .QN(_17382_));
 DFF_X1 _35065_ (.D(_00241_),
    .CK(clk),
    .Q(\text_in_r[82] ),
    .QN(_17383_));
 DFF_X1 _35066_ (.D(_00242_),
    .CK(clk),
    .Q(\text_in_r[83] ),
    .QN(_17384_));
 DFF_X1 _35067_ (.D(_00243_),
    .CK(clk),
    .Q(\text_in_r[84] ),
    .QN(_17385_));
 DFF_X1 _35068_ (.D(_00244_),
    .CK(clk),
    .Q(\text_in_r[85] ),
    .QN(_17386_));
 DFF_X1 _35069_ (.D(_00245_),
    .CK(clk),
    .Q(\text_in_r[86] ),
    .QN(_17387_));
 DFF_X1 _35070_ (.D(_00246_),
    .CK(clk),
    .Q(\text_in_r[87] ),
    .QN(_17388_));
 DFF_X1 _35071_ (.D(_00247_),
    .CK(clk),
    .Q(\text_in_r[88] ),
    .QN(_17389_));
 DFF_X1 _35072_ (.D(_00248_),
    .CK(clk),
    .Q(\text_in_r[89] ),
    .QN(_17390_));
 DFF_X1 _35073_ (.D(_00250_),
    .CK(clk),
    .Q(\text_in_r[90] ),
    .QN(_17391_));
 DFF_X1 _35074_ (.D(_00251_),
    .CK(clk),
    .Q(\text_in_r[91] ),
    .QN(_17392_));
 DFF_X1 _35075_ (.D(_00252_),
    .CK(clk),
    .Q(\text_in_r[92] ),
    .QN(_17393_));
 DFF_X1 _35076_ (.D(_00253_),
    .CK(clk),
    .Q(\text_in_r[93] ),
    .QN(_17394_));
 DFF_X1 _35077_ (.D(_00254_),
    .CK(clk),
    .Q(\text_in_r[94] ),
    .QN(_17395_));
 DFF_X1 _35078_ (.D(_00255_),
    .CK(clk),
    .Q(\text_in_r[95] ),
    .QN(_17396_));
 DFF_X1 _35079_ (.D(_00256_),
    .CK(clk),
    .Q(\text_in_r[96] ),
    .QN(_17397_));
 DFF_X1 _35080_ (.D(_00257_),
    .CK(clk),
    .Q(\text_in_r[97] ),
    .QN(_17398_));
 DFF_X1 _35081_ (.D(_00258_),
    .CK(clk),
    .Q(\text_in_r[98] ),
    .QN(_17399_));
 DFF_X1 _35082_ (.D(_00259_),
    .CK(clk),
    .Q(\text_in_r[99] ),
    .QN(_17400_));
 DFF_X1 _35083_ (.D(_00134_),
    .CK(clk),
    .Q(\text_in_r[100] ),
    .QN(_17401_));
 DFF_X1 _35084_ (.D(_00135_),
    .CK(clk),
    .Q(\text_in_r[101] ),
    .QN(_17402_));
 DFF_X1 _35085_ (.D(_00136_),
    .CK(clk),
    .Q(\text_in_r[102] ),
    .QN(_17403_));
 DFF_X1 _35086_ (.D(_00137_),
    .CK(clk),
    .Q(\text_in_r[103] ),
    .QN(_17404_));
 DFF_X1 _35087_ (.D(_00138_),
    .CK(clk),
    .Q(\text_in_r[104] ),
    .QN(_17405_));
 DFF_X1 _35088_ (.D(_00139_),
    .CK(clk),
    .Q(\text_in_r[105] ),
    .QN(_17406_));
 DFF_X1 _35089_ (.D(_00140_),
    .CK(clk),
    .Q(\text_in_r[106] ),
    .QN(_17407_));
 DFF_X1 _35090_ (.D(_00141_),
    .CK(clk),
    .Q(\text_in_r[107] ),
    .QN(_17408_));
 DFF_X1 _35091_ (.D(_00142_),
    .CK(clk),
    .Q(\text_in_r[108] ),
    .QN(_17409_));
 DFF_X1 _35092_ (.D(_00143_),
    .CK(clk),
    .Q(\text_in_r[109] ),
    .QN(_17410_));
 DFF_X1 _35093_ (.D(_00145_),
    .CK(clk),
    .Q(\text_in_r[110] ),
    .QN(_17411_));
 DFF_X1 _35094_ (.D(_00146_),
    .CK(clk),
    .Q(\text_in_r[111] ),
    .QN(_17412_));
 DFF_X1 _35095_ (.D(_00147_),
    .CK(clk),
    .Q(\text_in_r[112] ),
    .QN(_17413_));
 DFF_X1 _35096_ (.D(_00148_),
    .CK(clk),
    .Q(\text_in_r[113] ),
    .QN(_17414_));
 DFF_X1 _35097_ (.D(_00149_),
    .CK(clk),
    .Q(\text_in_r[114] ),
    .QN(_17415_));
 DFF_X1 _35098_ (.D(_00150_),
    .CK(clk),
    .Q(\text_in_r[115] ),
    .QN(_17416_));
 DFF_X1 _35099_ (.D(_00151_),
    .CK(clk),
    .Q(\text_in_r[116] ),
    .QN(_17417_));
 DFF_X1 _35100_ (.D(_00152_),
    .CK(clk),
    .Q(\text_in_r[117] ),
    .QN(_17418_));
 DFF_X1 _35101_ (.D(_00153_),
    .CK(clk),
    .Q(\text_in_r[118] ),
    .QN(_17419_));
 DFF_X1 _35102_ (.D(_00154_),
    .CK(clk),
    .Q(\text_in_r[119] ),
    .QN(_17420_));
 DFF_X1 _35103_ (.D(_00156_),
    .CK(clk),
    .Q(\text_in_r[120] ),
    .QN(_17421_));
 DFF_X1 _35104_ (.D(_00157_),
    .CK(clk),
    .Q(\text_in_r[121] ),
    .QN(_17422_));
 DFF_X1 _35105_ (.D(_00158_),
    .CK(clk),
    .Q(\text_in_r[122] ),
    .QN(_17423_));
 DFF_X1 _35106_ (.D(_00159_),
    .CK(clk),
    .Q(\text_in_r[123] ),
    .QN(_17424_));
 DFF_X1 _35107_ (.D(_00160_),
    .CK(clk),
    .Q(\text_in_r[124] ),
    .QN(_17425_));
 DFF_X1 _35108_ (.D(_00161_),
    .CK(clk),
    .Q(\text_in_r[125] ),
    .QN(_17426_));
 DFF_X1 _35109_ (.D(_00162_),
    .CK(clk),
    .Q(\text_in_r[126] ),
    .QN(_17427_));
 DFF_X1 _35110_ (.D(_00163_),
    .CK(clk),
    .Q(\text_in_r[127] ),
    .QN(_17428_));
 DFF_X1 _35111_ (.D(ld),
    .CK(clk),
    .Q(ld_r),
    .QN(_17429_));
 DFF_X1 _35112_ (.D(_00125_),
    .CK(clk),
    .Q(\sa33[0] ),
    .QN(_17430_));
 DFF_X1 _35113_ (.D(_00126_),
    .CK(clk),
    .Q(\sa33[1] ),
    .QN(_17431_));
 DFF_X1 _35114_ (.D(_00127_),
    .CK(clk),
    .Q(\sa33[2] ),
    .QN(_17432_));
 DFF_X1 _35115_ (.D(_00128_),
    .CK(clk),
    .Q(\sa33[3] ),
    .QN(_17433_));
 DFF_X1 _35116_ (.D(_00129_),
    .CK(clk),
    .Q(\sa33[4] ),
    .QN(_17434_));
 DFF_X1 _35117_ (.D(_00130_),
    .CK(clk),
    .Q(\sa33[5] ),
    .QN(_17435_));
 DFF_X1 _35118_ (.D(_00131_),
    .CK(clk),
    .Q(\sa33[6] ),
    .QN(_17436_));
 DFF_X1 _35119_ (.D(_00132_),
    .CK(clk),
    .Q(\sa33[7] ),
    .QN(_17437_));
 DFF_X1 _35120_ (.D(_00093_),
    .CK(clk),
    .Q(\sa23[0] ),
    .QN(_17438_));
 DFF_X1 _35121_ (.D(_00094_),
    .CK(clk),
    .Q(\sa23[1] ),
    .QN(_17439_));
 DFF_X1 _35122_ (.D(_00095_),
    .CK(clk),
    .Q(\sa23[2] ),
    .QN(_17440_));
 DFF_X1 _35123_ (.D(_00096_),
    .CK(clk),
    .Q(\sa23[3] ),
    .QN(_17441_));
 DFF_X1 _35124_ (.D(_00097_),
    .CK(clk),
    .Q(\sa23[4] ),
    .QN(_17442_));
 DFF_X1 _35125_ (.D(_00098_),
    .CK(clk),
    .Q(\sa23[5] ),
    .QN(_17443_));
 DFF_X1 _35126_ (.D(_00099_),
    .CK(clk),
    .Q(\sa23[6] ),
    .QN(_17444_));
 DFF_X1 _35127_ (.D(_00100_),
    .CK(clk),
    .Q(\sa23[7] ),
    .QN(_17445_));
 DFF_X1 _35128_ (.D(_00061_),
    .CK(clk),
    .Q(\sa13[0] ),
    .QN(_17446_));
 DFF_X1 _35129_ (.D(_00062_),
    .CK(clk),
    .Q(\sa13[1] ),
    .QN(_17447_));
 DFF_X1 _35130_ (.D(_00063_),
    .CK(clk),
    .Q(\sa13[2] ),
    .QN(_17448_));
 DFF_X1 _35131_ (.D(_00064_),
    .CK(clk),
    .Q(\sa13[3] ),
    .QN(_17449_));
 DFF_X1 _35132_ (.D(_00065_),
    .CK(clk),
    .Q(\sa13[4] ),
    .QN(_17450_));
 DFF_X1 _35133_ (.D(_00066_),
    .CK(clk),
    .Q(\sa13[5] ),
    .QN(_17451_));
 DFF_X1 _35134_ (.D(_00067_),
    .CK(clk),
    .Q(\sa13[6] ),
    .QN(_17452_));
 DFF_X1 _35135_ (.D(_00068_),
    .CK(clk),
    .Q(\sa13[7] ),
    .QN(_17453_));
 DFF_X1 _35136_ (.D(_00029_),
    .CK(clk),
    .Q(\sa03[0] ),
    .QN(_17454_));
 DFF_X1 _35137_ (.D(_00030_),
    .CK(clk),
    .Q(\sa03[1] ),
    .QN(_17455_));
 DFF_X1 _35138_ (.D(_00031_),
    .CK(clk),
    .Q(\sa03[2] ),
    .QN(_17456_));
 DFF_X1 _35139_ (.D(_00032_),
    .CK(clk),
    .Q(\sa03[3] ),
    .QN(_17457_));
 DFF_X1 _35140_ (.D(_00033_),
    .CK(clk),
    .Q(\sa03[4] ),
    .QN(_17458_));
 DFF_X1 _35141_ (.D(_00034_),
    .CK(clk),
    .Q(\sa03[5] ),
    .QN(_17459_));
 DFF_X1 _35142_ (.D(_00035_),
    .CK(clk),
    .Q(\sa03[6] ),
    .QN(_17460_));
 DFF_X1 _35143_ (.D(_00036_),
    .CK(clk),
    .Q(\sa03[7] ),
    .QN(_17461_));
 DFF_X1 _35144_ (.D(_00117_),
    .CK(clk),
    .Q(\sa32[0] ),
    .QN(_17462_));
 DFF_X1 _35145_ (.D(_00118_),
    .CK(clk),
    .Q(\sa32[1] ),
    .QN(_17463_));
 DFF_X1 _35146_ (.D(_00119_),
    .CK(clk),
    .Q(\sa32[2] ),
    .QN(_17464_));
 DFF_X1 _35147_ (.D(_00120_),
    .CK(clk),
    .Q(\sa32[3] ),
    .QN(_17465_));
 DFF_X1 _35148_ (.D(_00121_),
    .CK(clk),
    .Q(\sa32[4] ),
    .QN(_17466_));
 DFF_X1 _35149_ (.D(_00122_),
    .CK(clk),
    .Q(\sa32[5] ),
    .QN(_17467_));
 DFF_X1 _35150_ (.D(_00123_),
    .CK(clk),
    .Q(\sa32[6] ),
    .QN(_17468_));
 DFF_X1 _35151_ (.D(_00124_),
    .CK(clk),
    .Q(\sa32[7] ),
    .QN(_17469_));
 DFF_X1 _35152_ (.D(_00085_),
    .CK(clk),
    .Q(\sa22[0] ),
    .QN(_17470_));
 DFF_X1 _35153_ (.D(_00086_),
    .CK(clk),
    .Q(\sa22[1] ),
    .QN(_17471_));
 DFF_X1 _35154_ (.D(_00087_),
    .CK(clk),
    .Q(\sa22[2] ),
    .QN(_17472_));
 DFF_X1 _35155_ (.D(_00088_),
    .CK(clk),
    .Q(\sa22[3] ),
    .QN(_17473_));
 DFF_X1 _35156_ (.D(_00089_),
    .CK(clk),
    .Q(\sa22[4] ),
    .QN(_17474_));
 DFF_X1 _35157_ (.D(_00090_),
    .CK(clk),
    .Q(\sa22[5] ),
    .QN(_17475_));
 DFF_X1 _35158_ (.D(_00091_),
    .CK(clk),
    .Q(\sa22[6] ),
    .QN(_17476_));
 DFF_X1 _35159_ (.D(_00092_),
    .CK(clk),
    .Q(\sa22[7] ),
    .QN(_17477_));
 DFF_X1 _35160_ (.D(_00053_),
    .CK(clk),
    .Q(\sa12[0] ),
    .QN(_17478_));
 DFF_X1 _35161_ (.D(_00054_),
    .CK(clk),
    .Q(\sa12[1] ),
    .QN(_17479_));
 DFF_X1 _35162_ (.D(_00055_),
    .CK(clk),
    .Q(\sa12[2] ),
    .QN(_17480_));
 DFF_X1 _35163_ (.D(_00056_),
    .CK(clk),
    .Q(\sa12[3] ),
    .QN(_17481_));
 DFF_X1 _35164_ (.D(_00057_),
    .CK(clk),
    .Q(\sa12[4] ),
    .QN(_17482_));
 DFF_X1 _35165_ (.D(_00058_),
    .CK(clk),
    .Q(\sa12[5] ),
    .QN(_17483_));
 DFF_X1 _35166_ (.D(_00059_),
    .CK(clk),
    .Q(\sa12[6] ),
    .QN(_17484_));
 DFF_X1 _35167_ (.D(_00060_),
    .CK(clk),
    .Q(\sa12[7] ),
    .QN(_17485_));
 DFF_X1 _35168_ (.D(_00021_),
    .CK(clk),
    .Q(\sa02[0] ),
    .QN(_17486_));
 DFF_X1 _35169_ (.D(_00022_),
    .CK(clk),
    .Q(\sa02[1] ),
    .QN(_17487_));
 DFF_X1 _35170_ (.D(_00023_),
    .CK(clk),
    .Q(\sa02[2] ),
    .QN(_17488_));
 DFF_X1 _35171_ (.D(_00024_),
    .CK(clk),
    .Q(\sa02[3] ),
    .QN(_17489_));
 DFF_X1 _35172_ (.D(_00025_),
    .CK(clk),
    .Q(\sa02[4] ),
    .QN(_17490_));
 DFF_X1 _35173_ (.D(_00026_),
    .CK(clk),
    .Q(\sa02[5] ),
    .QN(_17491_));
 DFF_X1 _35174_ (.D(_00027_),
    .CK(clk),
    .Q(\sa02[6] ),
    .QN(_17492_));
 DFF_X1 _35175_ (.D(_00028_),
    .CK(clk),
    .Q(\sa02[7] ),
    .QN(_17493_));
 DFF_X1 _35176_ (.D(_00109_),
    .CK(clk),
    .Q(\sa31[0] ),
    .QN(_17494_));
 DFF_X1 _35177_ (.D(_00110_),
    .CK(clk),
    .Q(\sa31[1] ),
    .QN(_17495_));
 DFF_X1 _35178_ (.D(_00111_),
    .CK(clk),
    .Q(\sa31[2] ),
    .QN(_17496_));
 DFF_X1 _35179_ (.D(_00112_),
    .CK(clk),
    .Q(\sa31[3] ),
    .QN(_17497_));
 DFF_X1 _35180_ (.D(_00113_),
    .CK(clk),
    .Q(\sa31[4] ),
    .QN(_17498_));
 DFF_X1 _35181_ (.D(_00114_),
    .CK(clk),
    .Q(\sa31[5] ),
    .QN(_17499_));
 DFF_X1 _35182_ (.D(_00115_),
    .CK(clk),
    .Q(\sa31[6] ),
    .QN(_17500_));
 DFF_X1 _35183_ (.D(_00116_),
    .CK(clk),
    .Q(\sa31[7] ),
    .QN(_17501_));
 DFF_X1 _35184_ (.D(_00077_),
    .CK(clk),
    .Q(\sa21[0] ),
    .QN(_17502_));
 DFF_X1 _35185_ (.D(_00078_),
    .CK(clk),
    .Q(\sa21[1] ),
    .QN(_17503_));
 DFF_X1 _35186_ (.D(_00079_),
    .CK(clk),
    .Q(\sa21[2] ),
    .QN(_17504_));
 DFF_X1 _35187_ (.D(_00080_),
    .CK(clk),
    .Q(\sa21[3] ),
    .QN(_17505_));
 DFF_X1 _35188_ (.D(_00081_),
    .CK(clk),
    .Q(\sa21[4] ),
    .QN(_17506_));
 DFF_X1 _35189_ (.D(_00082_),
    .CK(clk),
    .Q(\sa21[5] ),
    .QN(_17507_));
 DFF_X1 _35190_ (.D(_00083_),
    .CK(clk),
    .Q(\sa21[6] ),
    .QN(_17508_));
 DFF_X1 _35191_ (.D(_00084_),
    .CK(clk),
    .Q(\sa21[7] ),
    .QN(_17509_));
 DFF_X1 _35192_ (.D(_00045_),
    .CK(clk),
    .Q(\sa11[0] ),
    .QN(_17510_));
 DFF_X1 _35193_ (.D(_00046_),
    .CK(clk),
    .Q(\sa11[1] ),
    .QN(_17511_));
 DFF_X1 _35194_ (.D(_00047_),
    .CK(clk),
    .Q(\sa11[2] ),
    .QN(_17512_));
 DFF_X1 _35195_ (.D(_00048_),
    .CK(clk),
    .Q(\sa11[3] ),
    .QN(_17513_));
 DFF_X1 _35196_ (.D(_00049_),
    .CK(clk),
    .Q(\sa11[4] ),
    .QN(_17514_));
 DFF_X1 _35197_ (.D(_00050_),
    .CK(clk),
    .Q(\sa11[5] ),
    .QN(_17515_));
 DFF_X1 _35198_ (.D(_00051_),
    .CK(clk),
    .Q(\sa11[6] ),
    .QN(_17516_));
 DFF_X1 _35199_ (.D(_00052_),
    .CK(clk),
    .Q(\sa11[7] ),
    .QN(_17517_));
 DFF_X1 _35200_ (.D(_00013_),
    .CK(clk),
    .Q(\sa01[0] ),
    .QN(_17518_));
 DFF_X1 _35201_ (.D(_00014_),
    .CK(clk),
    .Q(\sa01[1] ),
    .QN(_17519_));
 DFF_X1 _35202_ (.D(_00015_),
    .CK(clk),
    .Q(\sa01[2] ),
    .QN(_17520_));
 DFF_X1 _35203_ (.D(_00016_),
    .CK(clk),
    .Q(\sa01[3] ),
    .QN(_17521_));
 DFF_X1 _35204_ (.D(_00017_),
    .CK(clk),
    .Q(\sa01[4] ),
    .QN(_17522_));
 DFF_X1 _35205_ (.D(_00018_),
    .CK(clk),
    .Q(\sa01[5] ),
    .QN(_17523_));
 DFF_X1 _35206_ (.D(_00019_),
    .CK(clk),
    .Q(\sa01[6] ),
    .QN(_17524_));
 DFF_X1 _35207_ (.D(_00020_),
    .CK(clk),
    .Q(\sa01[7] ),
    .QN(_17525_));
 DFF_X1 _35208_ (.D(_00101_),
    .CK(clk),
    .Q(\sa30[0] ),
    .QN(_17526_));
 DFF_X1 _35209_ (.D(_00102_),
    .CK(clk),
    .Q(\sa30[1] ),
    .QN(_17527_));
 DFF_X1 _35210_ (.D(_00103_),
    .CK(clk),
    .Q(\sa30[2] ),
    .QN(_17528_));
 DFF_X1 _35211_ (.D(_00104_),
    .CK(clk),
    .Q(\sa30[3] ),
    .QN(_17529_));
 DFF_X1 _35212_ (.D(_00105_),
    .CK(clk),
    .Q(\sa30[4] ),
    .QN(_17530_));
 DFF_X1 _35213_ (.D(_00106_),
    .CK(clk),
    .Q(\sa30[5] ),
    .QN(_17531_));
 DFF_X1 _35214_ (.D(_00107_),
    .CK(clk),
    .Q(\sa30[6] ),
    .QN(_17532_));
 DFF_X1 _35215_ (.D(_00108_),
    .CK(clk),
    .Q(\sa30[7] ),
    .QN(_17533_));
 DFF_X1 _35216_ (.D(_00069_),
    .CK(clk),
    .Q(\sa20[0] ),
    .QN(_17534_));
 DFF_X1 _35217_ (.D(_00070_),
    .CK(clk),
    .Q(\sa20[1] ),
    .QN(_17535_));
 DFF_X1 _35218_ (.D(_00071_),
    .CK(clk),
    .Q(\sa20[2] ),
    .QN(_17536_));
 DFF_X1 _35219_ (.D(_00072_),
    .CK(clk),
    .Q(\sa20[3] ),
    .QN(_17537_));
 DFF_X1 _35220_ (.D(_00073_),
    .CK(clk),
    .Q(\sa20[4] ),
    .QN(_17538_));
 DFF_X1 _35221_ (.D(_00074_),
    .CK(clk),
    .Q(\sa20[5] ),
    .QN(_17539_));
 DFF_X1 _35222_ (.D(_00075_),
    .CK(clk),
    .Q(\sa20[6] ),
    .QN(_17540_));
 DFF_X1 _35223_ (.D(_00076_),
    .CK(clk),
    .Q(\sa20[7] ),
    .QN(_17541_));
 DFF_X1 _35224_ (.D(_00037_),
    .CK(clk),
    .Q(\sa10[0] ),
    .QN(_17542_));
 DFF_X1 _35225_ (.D(_00038_),
    .CK(clk),
    .Q(\sa10[1] ),
    .QN(_17543_));
 DFF_X1 _35226_ (.D(_00039_),
    .CK(clk),
    .Q(\sa10[2] ),
    .QN(_17544_));
 DFF_X1 _35227_ (.D(_00040_),
    .CK(clk),
    .Q(\sa10[3] ),
    .QN(_17545_));
 DFF_X1 _35228_ (.D(_00041_),
    .CK(clk),
    .Q(\sa10[4] ),
    .QN(_17546_));
 DFF_X1 _35229_ (.D(_00042_),
    .CK(clk),
    .Q(\sa10[5] ),
    .QN(_17547_));
 DFF_X1 _35230_ (.D(_00043_),
    .CK(clk),
    .Q(\sa10[6] ),
    .QN(_17548_));
 DFF_X1 _35231_ (.D(_00044_),
    .CK(clk),
    .Q(\sa10[7] ),
    .QN(_17549_));
 DFF_X1 _35232_ (.D(_00005_),
    .CK(clk),
    .Q(\sa00[0] ),
    .QN(_17550_));
 DFF_X1 _35233_ (.D(_00006_),
    .CK(clk),
    .Q(\sa00[1] ),
    .QN(_17551_));
 DFF_X1 _35234_ (.D(_00007_),
    .CK(clk),
    .Q(\sa00[2] ),
    .QN(_17552_));
 DFF_X1 _35235_ (.D(_00008_),
    .CK(clk),
    .Q(\sa00[3] ),
    .QN(_17553_));
 DFF_X1 _35236_ (.D(_00009_),
    .CK(clk),
    .Q(\sa00[4] ),
    .QN(_17554_));
 DFF_X1 _35237_ (.D(_00010_),
    .CK(clk),
    .Q(\sa00[5] ),
    .QN(_17555_));
 DFF_X1 _35238_ (.D(_00011_),
    .CK(clk),
    .Q(\sa00[6] ),
    .QN(_17556_));
 DFF_X1 _35239_ (.D(_00012_),
    .CK(clk),
    .Q(\sa00[7] ),
    .QN(_17557_));
 DFF_X1 _35240_ (.D(_00285_),
    .CK(clk),
    .Q(text_out[120]),
    .QN(_17558_));
 DFF_X1 _35241_ (.D(_00286_),
    .CK(clk),
    .Q(text_out[121]),
    .QN(_17559_));
 DFF_X1 _35242_ (.D(_00287_),
    .CK(clk),
    .Q(text_out[122]),
    .QN(_17560_));
 DFF_X1 _35243_ (.D(_00288_),
    .CK(clk),
    .Q(text_out[123]),
    .QN(_17561_));
 DFF_X1 _35244_ (.D(_00289_),
    .CK(clk),
    .Q(text_out[124]),
    .QN(_17562_));
 DFF_X1 _35245_ (.D(_00290_),
    .CK(clk),
    .Q(text_out[125]),
    .QN(_17563_));
 DFF_X1 _35246_ (.D(_00291_),
    .CK(clk),
    .Q(text_out[126]),
    .QN(_17564_));
 DFF_X1 _35247_ (.D(_00292_),
    .CK(clk),
    .Q(text_out[127]),
    .QN(_17565_));
 DFF_X1 _35248_ (.D(_00381_),
    .CK(clk),
    .Q(text_out[88]),
    .QN(_17566_));
 DFF_X1 _35249_ (.D(_00382_),
    .CK(clk),
    .Q(text_out[89]),
    .QN(_17567_));
 DFF_X1 _35250_ (.D(_00383_),
    .CK(clk),
    .Q(text_out[90]),
    .QN(_17568_));
 DFF_X1 _35251_ (.D(_00384_),
    .CK(clk),
    .Q(text_out[91]),
    .QN(_17569_));
 DFF_X1 _35252_ (.D(_00385_),
    .CK(clk),
    .Q(text_out[92]),
    .QN(_17570_));
 DFF_X1 _35253_ (.D(_00386_),
    .CK(clk),
    .Q(text_out[93]),
    .QN(_17571_));
 DFF_X1 _35254_ (.D(_00387_),
    .CK(clk),
    .Q(text_out[94]),
    .QN(_17572_));
 DFF_X1 _35255_ (.D(_00388_),
    .CK(clk),
    .Q(text_out[95]),
    .QN(_17573_));
 DFF_X1 _35256_ (.D(_00341_),
    .CK(clk),
    .Q(text_out[56]),
    .QN(_17574_));
 DFF_X1 _35257_ (.D(_00342_),
    .CK(clk),
    .Q(text_out[57]),
    .QN(_17575_));
 DFF_X1 _35258_ (.D(_00343_),
    .CK(clk),
    .Q(text_out[58]),
    .QN(_17576_));
 DFF_X1 _35259_ (.D(_00344_),
    .CK(clk),
    .Q(text_out[59]),
    .QN(_17577_));
 DFF_X1 _35260_ (.D(_00345_),
    .CK(clk),
    .Q(text_out[60]),
    .QN(_17578_));
 DFF_X1 _35261_ (.D(_00346_),
    .CK(clk),
    .Q(text_out[61]),
    .QN(_17579_));
 DFF_X1 _35262_ (.D(_00347_),
    .CK(clk),
    .Q(text_out[62]),
    .QN(_17580_));
 DFF_X1 _35263_ (.D(_00348_),
    .CK(clk),
    .Q(text_out[63]),
    .QN(_17581_));
 DFF_X1 _35264_ (.D(_00309_),
    .CK(clk),
    .Q(text_out[24]),
    .QN(_17582_));
 DFF_X1 _35265_ (.D(_00310_),
    .CK(clk),
    .Q(text_out[25]),
    .QN(_17583_));
 DFF_X1 _35266_ (.D(_00311_),
    .CK(clk),
    .Q(text_out[26]),
    .QN(_17584_));
 DFF_X1 _35267_ (.D(_00312_),
    .CK(clk),
    .Q(text_out[27]),
    .QN(_17585_));
 DFF_X1 _35268_ (.D(_00313_),
    .CK(clk),
    .Q(text_out[28]),
    .QN(_17586_));
 DFF_X1 _35269_ (.D(_00314_),
    .CK(clk),
    .Q(text_out[29]),
    .QN(_17587_));
 DFF_X1 _35270_ (.D(_00315_),
    .CK(clk),
    .Q(text_out[30]),
    .QN(_17588_));
 DFF_X1 _35271_ (.D(_00316_),
    .CK(clk),
    .Q(text_out[31]),
    .QN(_17589_));
 DFF_X1 _35272_ (.D(_00277_),
    .CK(clk),
    .Q(text_out[112]),
    .QN(_17590_));
 DFF_X1 _35273_ (.D(_00278_),
    .CK(clk),
    .Q(text_out[113]),
    .QN(_17591_));
 DFF_X1 _35274_ (.D(_00279_),
    .CK(clk),
    .Q(text_out[114]),
    .QN(_17592_));
 DFF_X1 _35275_ (.D(_00280_),
    .CK(clk),
    .Q(text_out[115]),
    .QN(_17593_));
 DFF_X1 _35276_ (.D(_00281_),
    .CK(clk),
    .Q(text_out[116]),
    .QN(_17594_));
 DFF_X1 _35277_ (.D(_00282_),
    .CK(clk),
    .Q(text_out[117]),
    .QN(_17595_));
 DFF_X1 _35278_ (.D(_00283_),
    .CK(clk),
    .Q(text_out[118]),
    .QN(_17596_));
 DFF_X1 _35279_ (.D(_00284_),
    .CK(clk),
    .Q(text_out[119]),
    .QN(_17597_));
 DFF_X1 _35280_ (.D(_00373_),
    .CK(clk),
    .Q(text_out[80]),
    .QN(_17598_));
 DFF_X1 _35281_ (.D(_00374_),
    .CK(clk),
    .Q(text_out[81]),
    .QN(_17599_));
 DFF_X1 _35282_ (.D(_00375_),
    .CK(clk),
    .Q(text_out[82]),
    .QN(_17600_));
 DFF_X1 _35283_ (.D(_00376_),
    .CK(clk),
    .Q(text_out[83]),
    .QN(_17601_));
 DFF_X1 _35284_ (.D(_00377_),
    .CK(clk),
    .Q(text_out[84]),
    .QN(_17602_));
 DFF_X1 _35285_ (.D(_00378_),
    .CK(clk),
    .Q(text_out[85]),
    .QN(_17603_));
 DFF_X1 _35286_ (.D(_00379_),
    .CK(clk),
    .Q(text_out[86]),
    .QN(_17604_));
 DFF_X1 _35287_ (.D(_00380_),
    .CK(clk),
    .Q(text_out[87]),
    .QN(_17605_));
 DFF_X1 _35288_ (.D(_00333_),
    .CK(clk),
    .Q(text_out[48]),
    .QN(_17606_));
 DFF_X1 _35289_ (.D(_00334_),
    .CK(clk),
    .Q(text_out[49]),
    .QN(_17607_));
 DFF_X1 _35290_ (.D(_00335_),
    .CK(clk),
    .Q(text_out[50]),
    .QN(_17608_));
 DFF_X1 _35291_ (.D(_00336_),
    .CK(clk),
    .Q(text_out[51]),
    .QN(_17609_));
 DFF_X1 _35292_ (.D(_00337_),
    .CK(clk),
    .Q(text_out[52]),
    .QN(_17610_));
 DFF_X1 _35293_ (.D(_00338_),
    .CK(clk),
    .Q(text_out[53]),
    .QN(_17611_));
 DFF_X1 _35294_ (.D(_00339_),
    .CK(clk),
    .Q(text_out[54]),
    .QN(_17612_));
 DFF_X1 _35295_ (.D(_00340_),
    .CK(clk),
    .Q(text_out[55]),
    .QN(_17613_));
 DFF_X1 _35296_ (.D(_00301_),
    .CK(clk),
    .Q(text_out[16]),
    .QN(_17614_));
 DFF_X1 _35297_ (.D(_00302_),
    .CK(clk),
    .Q(text_out[17]),
    .QN(_17615_));
 DFF_X1 _35298_ (.D(_00303_),
    .CK(clk),
    .Q(text_out[18]),
    .QN(_17616_));
 DFF_X1 _35299_ (.D(_00304_),
    .CK(clk),
    .Q(text_out[19]),
    .QN(_17617_));
 DFF_X1 _35300_ (.D(_00305_),
    .CK(clk),
    .Q(text_out[20]),
    .QN(_17618_));
 DFF_X1 _35301_ (.D(_00306_),
    .CK(clk),
    .Q(text_out[21]),
    .QN(_17619_));
 DFF_X1 _35302_ (.D(_00307_),
    .CK(clk),
    .Q(text_out[22]),
    .QN(_17620_));
 DFF_X1 _35303_ (.D(_00308_),
    .CK(clk),
    .Q(text_out[23]),
    .QN(_17621_));
 DFF_X1 _35304_ (.D(_00269_),
    .CK(clk),
    .Q(text_out[104]),
    .QN(_17622_));
 DFF_X1 _35305_ (.D(_00270_),
    .CK(clk),
    .Q(text_out[105]),
    .QN(_17623_));
 DFF_X1 _35306_ (.D(_00271_),
    .CK(clk),
    .Q(text_out[106]),
    .QN(_17624_));
 DFF_X1 _35307_ (.D(_00272_),
    .CK(clk),
    .Q(text_out[107]),
    .QN(_17625_));
 DFF_X1 _35308_ (.D(_00273_),
    .CK(clk),
    .Q(text_out[108]),
    .QN(_17626_));
 DFF_X1 _35309_ (.D(_00274_),
    .CK(clk),
    .Q(text_out[109]),
    .QN(_17627_));
 DFF_X1 _35310_ (.D(_00275_),
    .CK(clk),
    .Q(text_out[110]),
    .QN(_17628_));
 DFF_X1 _35311_ (.D(_00276_),
    .CK(clk),
    .Q(text_out[111]),
    .QN(_17629_));
 DFF_X1 _35312_ (.D(_00357_),
    .CK(clk),
    .Q(text_out[72]),
    .QN(_17630_));
 DFF_X1 _35313_ (.D(_00358_),
    .CK(clk),
    .Q(text_out[73]),
    .QN(_17631_));
 DFF_X1 _35314_ (.D(_00359_),
    .CK(clk),
    .Q(text_out[74]),
    .QN(_17632_));
 DFF_X1 _35315_ (.D(_00360_),
    .CK(clk),
    .Q(text_out[75]),
    .QN(_17633_));
 DFF_X1 _35316_ (.D(_00361_),
    .CK(clk),
    .Q(text_out[76]),
    .QN(_17634_));
 DFF_X1 _35317_ (.D(_00362_),
    .CK(clk),
    .Q(text_out[77]),
    .QN(_17635_));
 DFF_X1 _35318_ (.D(_00363_),
    .CK(clk),
    .Q(text_out[78]),
    .QN(_17636_));
 DFF_X1 _35319_ (.D(_00364_),
    .CK(clk),
    .Q(text_out[79]),
    .QN(_17637_));
 DFF_X1 _35320_ (.D(_00325_),
    .CK(clk),
    .Q(text_out[40]),
    .QN(_17638_));
 DFF_X1 _35321_ (.D(_00326_),
    .CK(clk),
    .Q(text_out[41]),
    .QN(_17639_));
 DFF_X1 _35322_ (.D(_00327_),
    .CK(clk),
    .Q(text_out[42]),
    .QN(_17640_));
 DFF_X1 _35323_ (.D(_00328_),
    .CK(clk),
    .Q(text_out[43]),
    .QN(_17641_));
 DFF_X1 _35324_ (.D(_00329_),
    .CK(clk),
    .Q(text_out[44]),
    .QN(_17642_));
 DFF_X1 _35325_ (.D(_00330_),
    .CK(clk),
    .Q(text_out[45]),
    .QN(_17643_));
 DFF_X1 _35326_ (.D(_00331_),
    .CK(clk),
    .Q(text_out[46]),
    .QN(_17644_));
 DFF_X1 _35327_ (.D(_00332_),
    .CK(clk),
    .Q(text_out[47]),
    .QN(_17645_));
 DFF_X1 _35328_ (.D(_00293_),
    .CK(clk),
    .Q(text_out[8]),
    .QN(_17646_));
 DFF_X1 _35329_ (.D(_00294_),
    .CK(clk),
    .Q(text_out[9]),
    .QN(_17647_));
 DFF_X1 _35330_ (.D(_00295_),
    .CK(clk),
    .Q(text_out[10]),
    .QN(_17648_));
 DFF_X1 _35331_ (.D(_00296_),
    .CK(clk),
    .Q(text_out[11]),
    .QN(_17649_));
 DFF_X1 _35332_ (.D(_00297_),
    .CK(clk),
    .Q(text_out[12]),
    .QN(_17650_));
 DFF_X1 _35333_ (.D(_00298_),
    .CK(clk),
    .Q(text_out[13]),
    .QN(_17651_));
 DFF_X1 _35334_ (.D(_00299_),
    .CK(clk),
    .Q(text_out[14]),
    .QN(_17652_));
 DFF_X1 _35335_ (.D(_00300_),
    .CK(clk),
    .Q(text_out[15]),
    .QN(_17653_));
 DFF_X1 _35336_ (.D(_00261_),
    .CK(clk),
    .Q(text_out[96]),
    .QN(_17654_));
 DFF_X1 _35337_ (.D(_00262_),
    .CK(clk),
    .Q(text_out[97]),
    .QN(_17655_));
 DFF_X1 _35338_ (.D(_00263_),
    .CK(clk),
    .Q(text_out[98]),
    .QN(_17656_));
 DFF_X1 _35339_ (.D(_00264_),
    .CK(clk),
    .Q(text_out[99]),
    .QN(_17657_));
 DFF_X1 _35340_ (.D(_00265_),
    .CK(clk),
    .Q(text_out[100]),
    .QN(_17658_));
 DFF_X1 _35341_ (.D(_00266_),
    .CK(clk),
    .Q(text_out[101]),
    .QN(_17659_));
 DFF_X1 _35342_ (.D(_00267_),
    .CK(clk),
    .Q(text_out[102]),
    .QN(_17660_));
 DFF_X1 _35343_ (.D(_00268_),
    .CK(clk),
    .Q(text_out[103]),
    .QN(_17661_));
 DFF_X1 _35344_ (.D(_00349_),
    .CK(clk),
    .Q(text_out[64]),
    .QN(_17662_));
 DFF_X1 _35345_ (.D(_00350_),
    .CK(clk),
    .Q(text_out[65]),
    .QN(_17663_));
 DFF_X1 _35346_ (.D(_00351_),
    .CK(clk),
    .Q(text_out[66]),
    .QN(_17664_));
 DFF_X1 _35347_ (.D(_00352_),
    .CK(clk),
    .Q(text_out[67]),
    .QN(_17665_));
 DFF_X1 _35348_ (.D(_00353_),
    .CK(clk),
    .Q(text_out[68]),
    .QN(_17666_));
 DFF_X1 _35349_ (.D(_00354_),
    .CK(clk),
    .Q(text_out[69]),
    .QN(_17667_));
 DFF_X1 _35350_ (.D(_00355_),
    .CK(clk),
    .Q(text_out[70]),
    .QN(_17668_));
 DFF_X1 _35351_ (.D(_00356_),
    .CK(clk),
    .Q(text_out[71]),
    .QN(_17669_));
 DFF_X1 _35352_ (.D(_00317_),
    .CK(clk),
    .Q(text_out[32]),
    .QN(_17670_));
 DFF_X1 _35353_ (.D(_00318_),
    .CK(clk),
    .Q(text_out[33]),
    .QN(_17671_));
 DFF_X1 _35354_ (.D(_00319_),
    .CK(clk),
    .Q(text_out[34]),
    .QN(_17672_));
 DFF_X1 _35355_ (.D(_00320_),
    .CK(clk),
    .Q(text_out[35]),
    .QN(_17673_));
 DFF_X1 _35356_ (.D(_00321_),
    .CK(clk),
    .Q(text_out[36]),
    .QN(_17674_));
 DFF_X1 _35357_ (.D(_00322_),
    .CK(clk),
    .Q(text_out[37]),
    .QN(_17675_));
 DFF_X1 _35358_ (.D(_00323_),
    .CK(clk),
    .Q(text_out[38]),
    .QN(_17676_));
 DFF_X1 _35359_ (.D(_00324_),
    .CK(clk),
    .Q(text_out[39]),
    .QN(_17677_));
 DFF_X1 _35360_ (.D(_00365_),
    .CK(clk),
    .Q(text_out[0]),
    .QN(_17678_));
 DFF_X1 _35361_ (.D(_00366_),
    .CK(clk),
    .Q(text_out[1]),
    .QN(_17679_));
 DFF_X1 _35362_ (.D(_00367_),
    .CK(clk),
    .Q(text_out[2]),
    .QN(_17680_));
 DFF_X1 _35363_ (.D(_00368_),
    .CK(clk),
    .Q(text_out[3]),
    .QN(_17681_));
 DFF_X1 _35364_ (.D(_00369_),
    .CK(clk),
    .Q(text_out[4]),
    .QN(_17682_));
 DFF_X1 _35365_ (.D(_00370_),
    .CK(clk),
    .Q(text_out[5]),
    .QN(_17683_));
 DFF_X1 _35366_ (.D(_00371_),
    .CK(clk),
    .Q(text_out[6]),
    .QN(_17684_));
 DFF_X1 _35367_ (.D(_00372_),
    .CK(clk),
    .Q(text_out[7]),
    .QN(_17685_));
 DFF_X1 _35368_ (.D(_00459_),
    .CK(clk),
    .Q(\u0.w[0][0] ),
    .QN(_00389_));
 DFF_X1 _35369_ (.D(_00470_),
    .CK(clk),
    .Q(\u0.w[0][1] ),
    .QN(_00390_));
 DFF_X1 _35370_ (.D(_00481_),
    .CK(clk),
    .Q(\u0.w[0][2] ),
    .QN(_00392_));
 DFF_X1 _35371_ (.D(_00484_),
    .CK(clk),
    .Q(\u0.w[0][3] ),
    .QN(_00393_));
 DFF_X1 _35372_ (.D(_00485_),
    .CK(clk),
    .Q(\u0.w[0][4] ),
    .QN(_00394_));
 DFF_X1 _35373_ (.D(_00486_),
    .CK(clk),
    .Q(\u0.w[0][5] ),
    .QN(_00395_));
 DFF_X1 _35374_ (.D(_00487_),
    .CK(clk),
    .Q(\u0.w[0][6] ),
    .QN(_00396_));
 DFF_X1 _35375_ (.D(_00488_),
    .CK(clk),
    .Q(\u0.w[0][7] ),
    .QN(_00397_));
 DFF_X1 _35376_ (.D(_00489_),
    .CK(clk),
    .Q(\u0.w[0][8] ),
    .QN(_00398_));
 DFF_X1 _35377_ (.D(_00490_),
    .CK(clk),
    .Q(\u0.w[0][9] ),
    .QN(_00399_));
 DFF_X1 _35378_ (.D(_00460_),
    .CK(clk),
    .Q(\u0.w[0][10] ),
    .QN(_00400_));
 DFF_X1 _35379_ (.D(_00461_),
    .CK(clk),
    .Q(\u0.w[0][11] ),
    .QN(_00401_));
 DFF_X1 _35380_ (.D(_00462_),
    .CK(clk),
    .Q(\u0.w[0][12] ),
    .QN(_00402_));
 DFF_X1 _35381_ (.D(_00463_),
    .CK(clk),
    .Q(\u0.w[0][13] ),
    .QN(_00403_));
 DFF_X1 _35382_ (.D(_00464_),
    .CK(clk),
    .Q(\u0.w[0][14] ),
    .QN(_00404_));
 DFF_X1 _35383_ (.D(_00465_),
    .CK(clk),
    .Q(\u0.w[0][15] ),
    .QN(_00405_));
 DFF_X1 _35384_ (.D(_00466_),
    .CK(clk),
    .Q(\u0.w[0][16] ),
    .QN(_00406_));
 DFF_X1 _35385_ (.D(_00467_),
    .CK(clk),
    .Q(\u0.w[0][17] ),
    .QN(_00407_));
 DFF_X1 _35386_ (.D(_00468_),
    .CK(clk),
    .Q(\u0.w[0][18] ),
    .QN(_00408_));
 DFF_X1 _35387_ (.D(_00469_),
    .CK(clk),
    .Q(\u0.w[0][19] ),
    .QN(_00409_));
 DFF_X1 _35388_ (.D(_00471_),
    .CK(clk),
    .Q(\u0.w[0][20] ),
    .QN(_00410_));
 DFF_X1 _35389_ (.D(_00472_),
    .CK(clk),
    .Q(\u0.w[0][21] ),
    .QN(_00411_));
 DFF_X1 _35390_ (.D(_00473_),
    .CK(clk),
    .Q(\u0.w[0][22] ),
    .QN(_00412_));
 DFF_X1 _35391_ (.D(_00474_),
    .CK(clk),
    .Q(\u0.w[0][23] ),
    .QN(_00413_));
 DFF_X1 _35392_ (.D(_00475_),
    .CK(clk),
    .Q(\u0.w[0][24] ),
    .QN(_00415_));
 DFF_X1 _35393_ (.D(_00476_),
    .CK(clk),
    .Q(\u0.w[0][25] ),
    .QN(_00417_));
 DFF_X1 _35394_ (.D(_00477_),
    .CK(clk),
    .Q(\u0.w[0][26] ),
    .QN(_00419_));
 DFF_X1 _35395_ (.D(_00478_),
    .CK(clk),
    .Q(\u0.w[0][27] ),
    .QN(_00421_));
 DFF_X1 _35396_ (.D(_00479_),
    .CK(clk),
    .Q(\u0.w[0][28] ),
    .QN(_00423_));
 DFF_X1 _35397_ (.D(_00480_),
    .CK(clk),
    .Q(\u0.w[0][29] ),
    .QN(_00425_));
 DFF_X1 _35398_ (.D(_00482_),
    .CK(clk),
    .Q(\u0.w[0][30] ),
    .QN(_00427_));
 DFF_X1 _35399_ (.D(_00483_),
    .CK(clk),
    .Q(\u0.w[0][31] ),
    .QN(_00429_));
 DFF_X1 _35400_ (.D(_00491_),
    .CK(clk),
    .Q(\u0.w[1][0] ),
    .QN(_17686_));
 DFF_X1 _35401_ (.D(_00502_),
    .CK(clk),
    .Q(\u0.w[1][1] ),
    .QN(_17687_));
 DFF_X1 _35402_ (.D(_00513_),
    .CK(clk),
    .Q(\u0.w[1][2] ),
    .QN(_17688_));
 DFF_X1 _35403_ (.D(_00516_),
    .CK(clk),
    .Q(\u0.w[1][3] ),
    .QN(_17689_));
 DFF_X1 _35404_ (.D(_00517_),
    .CK(clk),
    .Q(\u0.w[1][4] ),
    .QN(_17690_));
 DFF_X1 _35405_ (.D(_00518_),
    .CK(clk),
    .Q(\u0.w[1][5] ),
    .QN(_17691_));
 DFF_X1 _35406_ (.D(_00519_),
    .CK(clk),
    .Q(\u0.w[1][6] ),
    .QN(_17692_));
 DFF_X1 _35407_ (.D(_00520_),
    .CK(clk),
    .Q(\u0.w[1][7] ),
    .QN(_17693_));
 DFF_X1 _35408_ (.D(_00521_),
    .CK(clk),
    .Q(\u0.w[1][8] ),
    .QN(_00438_));
 DFF_X1 _35409_ (.D(_00522_),
    .CK(clk),
    .Q(\u0.w[1][9] ),
    .QN(_17694_));
 DFF_X1 _35410_ (.D(_00492_),
    .CK(clk),
    .Q(\u0.w[1][10] ),
    .QN(_17695_));
 DFF_X1 _35411_ (.D(_00493_),
    .CK(clk),
    .Q(\u0.w[1][11] ),
    .QN(_17696_));
 DFF_X1 _35412_ (.D(_00494_),
    .CK(clk),
    .Q(\u0.w[1][12] ),
    .QN(_17697_));
 DFF_X1 _35413_ (.D(_00495_),
    .CK(clk),
    .Q(\u0.w[1][13] ),
    .QN(_17698_));
 DFF_X1 _35414_ (.D(_00496_),
    .CK(clk),
    .Q(\u0.w[1][14] ),
    .QN(_17699_));
 DFF_X1 _35415_ (.D(_00497_),
    .CK(clk),
    .Q(\u0.w[1][15] ),
    .QN(_17700_));
 DFF_X1 _35416_ (.D(_00498_),
    .CK(clk),
    .Q(\u0.w[1][16] ),
    .QN(_00439_));
 DFF_X1 _35417_ (.D(_00499_),
    .CK(clk),
    .Q(\u0.w[1][17] ),
    .QN(_00440_));
 DFF_X1 _35418_ (.D(_00500_),
    .CK(clk),
    .Q(\u0.w[1][18] ),
    .QN(_17701_));
 DFF_X1 _35419_ (.D(_00501_),
    .CK(clk),
    .Q(\u0.w[1][19] ),
    .QN(_17702_));
 DFF_X1 _35420_ (.D(_00503_),
    .CK(clk),
    .Q(\u0.w[1][20] ),
    .QN(_17703_));
 DFF_X1 _35421_ (.D(_00504_),
    .CK(clk),
    .Q(\u0.w[1][21] ),
    .QN(_00441_));
 DFF_X1 _35422_ (.D(_00505_),
    .CK(clk),
    .Q(\u0.w[1][22] ),
    .QN(_00442_));
 DFF_X1 _35423_ (.D(_00506_),
    .CK(clk),
    .Q(\u0.w[1][23] ),
    .QN(_17704_));
 DFF_X1 _35424_ (.D(_00507_),
    .CK(clk),
    .Q(\u0.w[1][24] ),
    .QN(_00443_));
 DFF_X1 _35425_ (.D(_00508_),
    .CK(clk),
    .Q(\u0.w[1][25] ),
    .QN(_00444_));
 DFF_X1 _35426_ (.D(_00509_),
    .CK(clk),
    .Q(\u0.w[1][26] ),
    .QN(_17705_));
 DFF_X1 _35427_ (.D(_00510_),
    .CK(clk),
    .Q(\u0.w[1][27] ),
    .QN(_17706_));
 DFF_X1 _35428_ (.D(_00511_),
    .CK(clk),
    .Q(\u0.w[1][28] ),
    .QN(_17707_));
 DFF_X1 _35429_ (.D(_00512_),
    .CK(clk),
    .Q(\u0.w[1][29] ),
    .QN(_00445_));
 DFF_X1 _35430_ (.D(_00514_),
    .CK(clk),
    .Q(\u0.w[1][30] ),
    .QN(_00449_));
 DFF_X1 _35431_ (.D(_00515_),
    .CK(clk),
    .Q(\u0.w[1][31] ),
    .QN(_17708_));
 DFF_X1 _35432_ (.D(_00523_),
    .CK(clk),
    .Q(\u0.w[2][0] ),
    .QN(_17709_));
 DFF_X1 _35433_ (.D(_00534_),
    .CK(clk),
    .Q(\u0.w[2][1] ),
    .QN(_17710_));
 DFF_X1 _35434_ (.D(_00545_),
    .CK(clk),
    .Q(\u0.w[2][2] ),
    .QN(_17711_));
 DFF_X1 _35435_ (.D(_00548_),
    .CK(clk),
    .Q(\u0.w[2][3] ),
    .QN(_17712_));
 DFF_X1 _35436_ (.D(_00549_),
    .CK(clk),
    .Q(\u0.w[2][4] ),
    .QN(_17713_));
 DFF_X1 _35437_ (.D(_00550_),
    .CK(clk),
    .Q(\u0.w[2][5] ),
    .QN(_17714_));
 DFF_X1 _35438_ (.D(_00551_),
    .CK(clk),
    .Q(\u0.w[2][6] ),
    .QN(_17715_));
 DFF_X1 _35439_ (.D(_00552_),
    .CK(clk),
    .Q(\u0.w[2][7] ),
    .QN(_17716_));
 DFF_X1 _35440_ (.D(_00553_),
    .CK(clk),
    .Q(\u0.w[2][8] ),
    .QN(_00391_));
 DFF_X1 _35441_ (.D(_00554_),
    .CK(clk),
    .Q(\u0.w[2][9] ),
    .QN(_17717_));
 DFF_X1 _35442_ (.D(_00524_),
    .CK(clk),
    .Q(\u0.w[2][10] ),
    .QN(_17718_));
 DFF_X1 _35443_ (.D(_00525_),
    .CK(clk),
    .Q(\u0.w[2][11] ),
    .QN(_17719_));
 DFF_X1 _35444_ (.D(_00526_),
    .CK(clk),
    .Q(\u0.w[2][12] ),
    .QN(_17720_));
 DFF_X1 _35445_ (.D(_00527_),
    .CK(clk),
    .Q(\u0.w[2][13] ),
    .QN(_17721_));
 DFF_X1 _35446_ (.D(_00528_),
    .CK(clk),
    .Q(\u0.w[2][14] ),
    .QN(_17722_));
 DFF_X1 _35447_ (.D(_00529_),
    .CK(clk),
    .Q(\u0.w[2][15] ),
    .QN(_17723_));
 DFF_X1 _35448_ (.D(_00530_),
    .CK(clk),
    .Q(\u0.w[2][16] ),
    .QN(_00430_));
 DFF_X1 _35449_ (.D(_00531_),
    .CK(clk),
    .Q(\u0.w[2][17] ),
    .QN(_00431_));
 DFF_X1 _35450_ (.D(_00532_),
    .CK(clk),
    .Q(\u0.w[2][18] ),
    .QN(_17724_));
 DFF_X1 _35451_ (.D(_00533_),
    .CK(clk),
    .Q(\u0.w[2][19] ),
    .QN(_17725_));
 DFF_X1 _35452_ (.D(_00535_),
    .CK(clk),
    .Q(\u0.w[2][20] ),
    .QN(_17726_));
 DFF_X1 _35453_ (.D(_00536_),
    .CK(clk),
    .Q(\u0.w[2][21] ),
    .QN(_00432_));
 DFF_X1 _35454_ (.D(_00537_),
    .CK(clk),
    .Q(\u0.w[2][22] ),
    .QN(_00433_));
 DFF_X1 _35455_ (.D(_00538_),
    .CK(clk),
    .Q(\u0.w[2][23] ),
    .QN(_17727_));
 DFF_X1 _35456_ (.D(_00539_),
    .CK(clk),
    .Q(\u0.w[2][24] ),
    .QN(_00434_));
 DFF_X1 _35457_ (.D(_00540_),
    .CK(clk),
    .Q(\u0.w[2][25] ),
    .QN(_00435_));
 DFF_X1 _35458_ (.D(_00541_),
    .CK(clk),
    .Q(\u0.w[2][26] ),
    .QN(_17728_));
 DFF_X1 _35459_ (.D(_00542_),
    .CK(clk),
    .Q(\u0.w[2][27] ),
    .QN(_17729_));
 DFF_X1 _35460_ (.D(_00543_),
    .CK(clk),
    .Q(\u0.w[2][28] ),
    .QN(_17730_));
 DFF_X1 _35461_ (.D(_00544_),
    .CK(clk),
    .Q(\u0.w[2][29] ),
    .QN(_00436_));
 DFF_X1 _35462_ (.D(_00546_),
    .CK(clk),
    .Q(\u0.w[2][30] ),
    .QN(_00437_));
 DFF_X1 _35463_ (.D(_00547_),
    .CK(clk),
    .Q(\u0.w[2][31] ),
    .QN(_17731_));
endmodule
