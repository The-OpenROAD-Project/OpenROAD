# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_io__top_ground_lvc_wpad
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 198 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    ANTENNAPARTIALMETALSIDEAREA  111.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 51.125000 1.270000 54.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.125000 75.000000 54.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    ANTENNAPARTIALMETALSIDEAREA  111.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 46.365000 1.270000 49.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 46.365000 75.000000 49.345000 ;
    END
  END AMUXBUS_B
  PIN G_PAD
    ANTENNAPARTIALMETALSIDEAREA  243.2170 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 31.695000 162.765000 52.340000 167.120000 ;
    END
  END G_PAD
  PIN BDY2_B2B
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 17.630000 5.115000 53.535000 9.540000 ;
        RECT 17.635000 5.110000 53.535000 5.115000 ;
        RECT 17.705000 5.040000 53.535000 5.110000 ;
        RECT 17.775000 4.970000 53.535000 5.040000 ;
        RECT 17.845000 4.900000 53.535000 4.970000 ;
        RECT 17.915000 4.830000 53.535000 4.900000 ;
        RECT 17.985000 4.760000 53.535000 4.830000 ;
        RECT 18.055000 4.690000 53.535000 4.760000 ;
        RECT 18.125000 4.620000 53.535000 4.690000 ;
        RECT 18.195000 4.550000 53.535000 4.620000 ;
        RECT 18.265000 4.480000 53.535000 4.550000 ;
        RECT 18.335000 4.410000 53.535000 4.480000 ;
        RECT 18.405000 4.340000 53.535000 4.410000 ;
        RECT 18.475000 4.270000 53.535000 4.340000 ;
        RECT 18.545000 4.200000 53.535000 4.270000 ;
        RECT 18.615000 4.130000 53.535000 4.200000 ;
        RECT 18.685000 4.060000 53.535000 4.130000 ;
        RECT 18.755000 3.990000 53.535000 4.060000 ;
        RECT 18.825000 3.920000 53.535000 3.990000 ;
        RECT 18.895000 3.850000 53.535000 3.920000 ;
        RECT 18.965000 3.780000 53.535000 3.850000 ;
        RECT 19.035000 3.710000 53.535000 3.780000 ;
        RECT 19.105000 3.640000 53.535000 3.710000 ;
        RECT 19.175000 3.570000 53.535000 3.640000 ;
        RECT 19.245000 3.500000 53.535000 3.570000 ;
        RECT 19.315000 3.430000 53.535000 3.500000 ;
        RECT 19.385000 3.360000 53.535000 3.430000 ;
        RECT 19.455000 3.290000 53.535000 3.360000 ;
        RECT 19.525000 3.220000 53.535000 3.290000 ;
        RECT 19.595000 3.150000 53.535000 3.220000 ;
        RECT 19.665000 3.080000 53.535000 3.150000 ;
        RECT 19.735000 3.010000 53.535000 3.080000 ;
        RECT 19.805000 2.940000 53.535000 3.010000 ;
        RECT 19.875000 2.870000 53.535000 2.940000 ;
        RECT 19.945000 2.800000 53.535000 2.870000 ;
        RECT 20.015000 2.730000 53.535000 2.800000 ;
        RECT 20.085000 2.660000 53.535000 2.730000 ;
        RECT 20.155000 2.590000 53.535000 2.660000 ;
        RECT 20.225000 2.520000 53.535000 2.590000 ;
        RECT 20.295000 2.450000 53.535000 2.520000 ;
        RECT 20.365000 2.380000 53.535000 2.450000 ;
        RECT 20.435000 2.310000 53.535000 2.380000 ;
        RECT 20.505000 2.240000 53.535000 2.310000 ;
        RECT 20.575000 2.170000 53.535000 2.240000 ;
        RECT 20.645000 2.100000 53.535000 2.170000 ;
        RECT 20.715000 2.030000 53.535000 2.100000 ;
        RECT 20.785000 1.960000 53.535000 2.030000 ;
        RECT 20.855000 1.890000 53.535000 1.960000 ;
        RECT 20.925000 0.000000 53.535000 1.820000 ;
        RECT 20.925000 1.820000 53.535000 1.890000 ;
    END
  END BDY2_B2B
  PIN DRN_LVC1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 15.605000  94.310000 23.935000  94.460000 ;
        RECT 15.605000  94.460000 23.785000  94.610000 ;
        RECT 15.605000  94.610000 23.635000  94.760000 ;
        RECT 15.605000  94.760000 23.485000  94.910000 ;
        RECT 15.605000  94.910000 23.335000  95.060000 ;
        RECT 15.605000  95.060000 23.185000  95.210000 ;
        RECT 15.605000  95.210000 23.035000  95.360000 ;
        RECT 15.605000  95.360000 22.885000  95.510000 ;
        RECT 15.605000  95.510000 22.735000  95.660000 ;
        RECT 15.605000  95.660000 22.585000  95.810000 ;
        RECT 15.605000  95.810000 22.435000  95.960000 ;
        RECT 15.605000  95.960000 22.285000  96.110000 ;
        RECT 15.605000  96.110000 22.135000  96.260000 ;
        RECT 15.605000  96.260000 21.985000  96.410000 ;
        RECT 15.605000  96.410000 21.835000  96.560000 ;
        RECT 15.605000  96.560000 21.685000  96.710000 ;
        RECT 15.605000  96.710000 21.605000  96.790000 ;
        RECT 15.605000  96.790000 21.605000 167.100000 ;
        RECT 15.605000 167.100000 21.605000 167.250000 ;
        RECT 15.605000 167.250000 21.755000 167.400000 ;
        RECT 15.605000 167.400000 21.905000 167.550000 ;
        RECT 15.605000 167.550000 22.055000 167.700000 ;
        RECT 15.605000 167.700000 22.205000 167.850000 ;
        RECT 15.605000 167.850000 22.355000 168.000000 ;
        RECT 15.605000 168.000000 22.505000 168.150000 ;
        RECT 15.605000 168.150000 22.655000 168.300000 ;
        RECT 15.605000 168.300000 22.805000 168.450000 ;
        RECT 15.605000 168.450000 22.955000 168.600000 ;
        RECT 15.605000 168.600000 23.105000 168.750000 ;
        RECT 15.605000 168.750000 23.255000 168.900000 ;
        RECT 15.605000 168.900000 23.405000 169.050000 ;
        RECT 15.605000 169.050000 23.555000 169.200000 ;
        RECT 15.605000 169.200000 23.705000 169.350000 ;
        RECT 15.605000 169.350000 23.855000 169.500000 ;
        RECT 15.605000 169.500000 24.005000 169.650000 ;
        RECT 15.605000 169.650000 24.155000 169.800000 ;
        RECT 15.605000 169.800000 24.305000 169.950000 ;
        RECT 15.605000 169.950000 24.455000 170.100000 ;
        RECT 15.605000 170.100000 24.605000 170.250000 ;
        RECT 15.605000 170.250000 24.755000 170.400000 ;
        RECT 15.605000 170.400000 24.905000 170.550000 ;
        RECT 15.605000 170.550000 25.055000 170.610000 ;
        RECT 15.605000 170.610000 25.115000 189.515000 ;
        RECT 15.715000  94.200000 24.085000  94.310000 ;
        RECT 15.865000  94.050000 24.195000  94.200000 ;
        RECT 16.015000  93.900000 24.345000  94.050000 ;
        RECT 16.165000  93.750000 24.495000  93.900000 ;
        RECT 16.315000  93.600000 24.645000  93.750000 ;
        RECT 16.465000  93.450000 24.795000  93.600000 ;
        RECT 16.615000  93.300000 24.945000  93.450000 ;
        RECT 16.765000  93.150000 25.095000  93.300000 ;
        RECT 16.915000  93.000000 25.245000  93.150000 ;
        RECT 17.065000  92.850000 25.395000  93.000000 ;
        RECT 17.215000  92.700000 25.545000  92.850000 ;
        RECT 17.365000  92.550000 25.695000  92.700000 ;
        RECT 17.515000  92.400000 25.845000  92.550000 ;
        RECT 17.665000  92.250000 25.995000  92.400000 ;
        RECT 17.815000  92.100000 26.145000  92.250000 ;
        RECT 17.965000  91.950000 26.295000  92.100000 ;
        RECT 18.115000  91.800000 26.445000  91.950000 ;
        RECT 18.265000  91.650000 26.595000  91.800000 ;
        RECT 18.415000  91.500000 26.745000  91.650000 ;
        RECT 18.565000  91.350000 26.895000  91.500000 ;
        RECT 18.715000  91.200000 27.045000  91.350000 ;
        RECT 18.865000  91.050000 27.195000  91.200000 ;
        RECT 19.015000  90.900000 27.345000  91.050000 ;
        RECT 19.165000  90.750000 27.495000  90.900000 ;
        RECT 19.315000  90.600000 27.645000  90.750000 ;
        RECT 19.465000  90.450000 27.795000  90.600000 ;
        RECT 19.615000  90.300000 27.945000  90.450000 ;
        RECT 19.765000  90.150000 28.095000  90.300000 ;
        RECT 19.915000  90.000000 28.245000  90.150000 ;
        RECT 20.065000  89.850000 28.395000  90.000000 ;
        RECT 20.215000  89.700000 28.545000  89.850000 ;
        RECT 20.365000  89.550000 28.695000  89.700000 ;
        RECT 20.515000  89.400000 28.845000  89.550000 ;
        RECT 20.665000  89.250000 28.995000  89.400000 ;
        RECT 20.815000  89.100000 29.145000  89.250000 ;
        RECT 20.965000  88.950000 29.295000  89.100000 ;
        RECT 21.115000  88.800000 29.445000  88.950000 ;
        RECT 21.265000  88.650000 29.595000  88.800000 ;
        RECT 21.415000  88.500000 29.745000  88.650000 ;
        RECT 21.565000  88.350000 29.895000  88.500000 ;
        RECT 21.715000  88.200000 30.045000  88.350000 ;
        RECT 21.865000  88.050000 30.195000  88.200000 ;
        RECT 22.015000  87.900000 30.345000  88.050000 ;
        RECT 22.165000  87.750000 30.495000  87.900000 ;
        RECT 22.315000  87.600000 30.645000  87.750000 ;
        RECT 22.465000  87.450000 30.795000  87.600000 ;
        RECT 22.615000  87.300000 30.945000  87.450000 ;
        RECT 22.765000  87.150000 31.095000  87.300000 ;
        RECT 22.915000  87.000000 31.245000  87.150000 ;
        RECT 23.065000  86.850000 31.395000  87.000000 ;
        RECT 23.215000  86.700000 31.545000  86.850000 ;
        RECT 23.365000  86.550000 31.695000  86.700000 ;
        RECT 23.515000  86.400000 31.845000  86.550000 ;
        RECT 23.665000  86.250000 31.995000  86.400000 ;
        RECT 23.670000  86.245000 32.145000  86.250000 ;
        RECT 23.760000  86.155000 32.145000  86.245000 ;
        RECT 23.850000  84.650000 32.165000  84.670000 ;
        RECT 23.850000  84.670000 32.145000  84.690000 ;
        RECT 23.850000  84.690000 32.145000  86.065000 ;
        RECT 23.850000  86.065000 32.145000  86.155000 ;
        RECT 23.920000  84.580000 32.185000  84.650000 ;
        RECT 24.070000  84.430000 32.255000  84.580000 ;
        RECT 24.220000  84.280000 32.405000  84.430000 ;
        RECT 24.370000  84.130000 32.555000  84.280000 ;
        RECT 24.520000  83.980000 32.705000  84.130000 ;
        RECT 24.650000  83.850000 48.870000  83.980000 ;
        RECT 24.800000  83.700000 48.870000  83.850000 ;
        RECT 24.950000  83.550000 48.870000  83.700000 ;
        RECT 25.100000  83.400000 48.870000  83.550000 ;
        RECT 25.250000  83.250000 48.870000  83.400000 ;
        RECT 25.400000  83.100000 48.870000  83.250000 ;
        RECT 25.550000  82.950000 48.870000  83.100000 ;
        RECT 25.700000  82.800000 48.870000  82.950000 ;
        RECT 25.850000  82.650000 48.870000  82.800000 ;
        RECT 26.000000   0.000000 36.880000  71.105000 ;
        RECT 26.000000  71.105000 36.880000  71.255000 ;
        RECT 26.000000  71.255000 37.030000  71.405000 ;
        RECT 26.000000  71.405000 37.180000  71.555000 ;
        RECT 26.000000  71.555000 37.330000  71.705000 ;
        RECT 26.000000  71.705000 37.480000  71.855000 ;
        RECT 26.000000  71.855000 37.630000  72.005000 ;
        RECT 26.000000  72.005000 37.780000  72.155000 ;
        RECT 26.000000  72.155000 37.930000  72.305000 ;
        RECT 26.000000  72.305000 38.080000  72.455000 ;
        RECT 26.000000  72.455000 38.230000  72.605000 ;
        RECT 26.000000  72.605000 38.380000  72.755000 ;
        RECT 26.000000  72.755000 38.530000  72.905000 ;
        RECT 26.000000  72.905000 38.680000  73.055000 ;
        RECT 26.000000  73.055000 38.830000  73.205000 ;
        RECT 26.000000  73.205000 38.980000  73.355000 ;
        RECT 26.000000  73.355000 39.130000  73.505000 ;
        RECT 26.000000  73.505000 39.280000  73.655000 ;
        RECT 26.000000  73.655000 39.430000  73.805000 ;
        RECT 26.000000  73.805000 39.580000  73.955000 ;
        RECT 26.000000  73.955000 39.730000  74.105000 ;
        RECT 26.000000  74.105000 39.880000  74.255000 ;
        RECT 26.000000  74.255000 40.030000  74.405000 ;
        RECT 26.000000  74.405000 40.180000  74.555000 ;
        RECT 26.000000  74.555000 40.330000  74.705000 ;
        RECT 26.000000  74.705000 40.480000  74.740000 ;
        RECT 26.000000  74.740000 46.795000  74.890000 ;
        RECT 26.000000  74.890000 46.945000  75.040000 ;
        RECT 26.000000  75.040000 47.095000  75.190000 ;
        RECT 26.000000  75.190000 47.245000  75.340000 ;
        RECT 26.000000  75.340000 47.395000  75.490000 ;
        RECT 26.000000  75.490000 47.545000  75.640000 ;
        RECT 26.000000  75.640000 47.695000  75.790000 ;
        RECT 26.000000  75.790000 47.845000  75.940000 ;
        RECT 26.000000  75.940000 47.995000  76.090000 ;
        RECT 26.000000  76.090000 48.145000  76.240000 ;
        RECT 26.000000  76.240000 48.295000  76.390000 ;
        RECT 26.000000  76.390000 48.445000  76.540000 ;
        RECT 26.000000  76.540000 48.595000  76.690000 ;
        RECT 26.000000  76.690000 48.745000  76.815000 ;
        RECT 26.000000  76.815000 48.870000  82.500000 ;
        RECT 26.000000  82.500000 48.870000  82.650000 ;
        RECT 26.035000  94.500000 32.035000 162.570000 ;
        RECT 26.035000 162.570000 32.035000 162.720000 ;
        RECT 26.035000 162.720000 32.185000 162.870000 ;
        RECT 26.035000 162.870000 32.335000 163.020000 ;
        RECT 26.035000 163.020000 32.485000 163.170000 ;
        RECT 26.035000 163.170000 32.635000 163.320000 ;
        RECT 26.035000 163.320000 32.785000 163.470000 ;
        RECT 26.035000 163.470000 32.935000 163.620000 ;
        RECT 26.035000 163.620000 33.085000 163.770000 ;
        RECT 26.035000 163.770000 33.235000 163.920000 ;
        RECT 26.035000 163.920000 33.385000 164.070000 ;
        RECT 26.035000 164.070000 33.535000 164.220000 ;
        RECT 26.035000 164.220000 33.685000 164.370000 ;
        RECT 26.035000 164.370000 33.835000 164.520000 ;
        RECT 26.035000 164.520000 33.985000 164.670000 ;
        RECT 26.035000 164.670000 34.135000 164.820000 ;
        RECT 26.035000 164.820000 34.285000 164.970000 ;
        RECT 26.035000 164.970000 34.435000 165.120000 ;
        RECT 26.035000 165.120000 34.585000 165.270000 ;
        RECT 26.035000 165.270000 34.735000 165.420000 ;
        RECT 26.035000 165.420000 34.885000 165.570000 ;
        RECT 26.035000 165.570000 35.035000 165.720000 ;
        RECT 26.035000 165.720000 35.185000 165.870000 ;
        RECT 26.035000 165.870000 35.335000 166.020000 ;
        RECT 26.035000 166.020000 35.485000 166.170000 ;
        RECT 26.035000 166.170000 35.635000 166.320000 ;
        RECT 26.035000 166.320000 35.785000 166.470000 ;
        RECT 26.035000 166.470000 35.935000 166.620000 ;
        RECT 26.035000 166.620000 36.085000 166.770000 ;
        RECT 26.035000 166.770000 36.235000 166.920000 ;
        RECT 26.035000 166.920000 36.385000 167.070000 ;
        RECT 26.035000 167.070000 36.535000 167.220000 ;
        RECT 26.035000 167.220000 36.685000 167.370000 ;
        RECT 26.035000 167.370000 36.835000 167.460000 ;
        RECT 26.035000 167.460000 36.925000 189.515000 ;
        RECT 26.095000  94.440000 32.035000  94.500000 ;
        RECT 26.245000  94.290000 32.035000  94.440000 ;
        RECT 26.395000  94.140000 32.035000  94.290000 ;
        RECT 26.545000  93.990000 32.035000  94.140000 ;
        RECT 26.695000  93.840000 32.035000  93.990000 ;
        RECT 26.845000  93.690000 32.035000  93.840000 ;
        RECT 26.995000  93.540000 32.035000  93.690000 ;
        RECT 27.145000  93.390000 32.035000  93.540000 ;
        RECT 27.160000  93.375000 32.035000  93.390000 ;
        RECT 27.310000  93.225000 32.050000  93.375000 ;
        RECT 27.460000  93.075000 32.200000  93.225000 ;
        RECT 27.610000  92.925000 32.350000  93.075000 ;
        RECT 27.760000  92.775000 32.500000  92.925000 ;
        RECT 27.910000  92.625000 32.650000  92.775000 ;
        RECT 28.060000  92.475000 32.800000  92.625000 ;
        RECT 28.210000  92.325000 32.950000  92.475000 ;
        RECT 28.360000  92.175000 33.100000  92.325000 ;
        RECT 28.510000  92.025000 33.250000  92.175000 ;
        RECT 28.660000  91.875000 33.400000  92.025000 ;
        RECT 28.810000  91.725000 33.550000  91.875000 ;
        RECT 28.960000  91.575000 33.700000  91.725000 ;
        RECT 29.110000  91.425000 33.850000  91.575000 ;
        RECT 29.260000  91.275000 34.000000  91.425000 ;
        RECT 29.410000  91.125000 34.150000  91.275000 ;
        RECT 29.560000  90.975000 34.300000  91.125000 ;
        RECT 29.710000  90.825000 34.450000  90.975000 ;
        RECT 29.860000  90.675000 34.600000  90.825000 ;
        RECT 30.010000  90.525000 34.750000  90.675000 ;
        RECT 30.160000  90.375000 34.900000  90.525000 ;
        RECT 30.175000  90.360000 42.385000  90.375000 ;
        RECT 30.325000  90.210000 42.235000  90.360000 ;
        RECT 30.475000  90.060000 42.085000  90.210000 ;
        RECT 30.625000  89.910000 41.935000  90.060000 ;
        RECT 30.775000  89.760000 41.785000  89.910000 ;
        RECT 30.925000  89.610000 41.635000  89.760000 ;
        RECT 31.075000  89.460000 41.485000  89.610000 ;
        RECT 31.225000  89.310000 41.335000  89.460000 ;
        RECT 31.375000  89.160000 41.185000  89.310000 ;
        RECT 31.525000  89.010000 41.035000  89.160000 ;
        RECT 31.675000  88.860000 40.885000  89.010000 ;
        RECT 31.825000  88.710000 40.735000  88.860000 ;
        RECT 31.975000  88.560000 40.585000  88.710000 ;
        RECT 32.125000  88.410000 40.435000  88.560000 ;
        RECT 32.275000  88.260000 40.285000  88.410000 ;
        RECT 32.425000  88.110000 40.135000  88.260000 ;
        RECT 32.575000  87.960000 39.985000  88.110000 ;
        RECT 32.725000  87.810000 39.835000  87.960000 ;
        RECT 32.875000  87.660000 39.685000  87.810000 ;
        RECT 33.025000  87.510000 39.535000  87.660000 ;
        RECT 33.175000  87.360000 39.385000  87.510000 ;
        RECT 33.305000  87.230000 39.385000  87.360000 ;
        RECT 33.455000  87.080000 39.385000  87.230000 ;
        RECT 33.605000  86.930000 39.385000  87.080000 ;
        RECT 33.755000  86.780000 39.385000  86.930000 ;
        RECT 33.905000  86.630000 39.385000  86.780000 ;
        RECT 33.945000  83.980000 39.945000  84.130000 ;
        RECT 34.055000  86.480000 39.385000  86.630000 ;
        RECT 34.095000  84.130000 39.795000  84.280000 ;
        RECT 34.205000  86.330000 39.385000  86.480000 ;
        RECT 34.245000  84.280000 39.645000  84.430000 ;
        RECT 34.355000  86.180000 39.385000  86.330000 ;
        RECT 34.395000  84.430000 39.495000  84.580000 ;
        RECT 34.505000  84.580000 39.385000  84.690000 ;
        RECT 34.505000  84.690000 39.385000  86.030000 ;
        RECT 34.505000  86.030000 39.385000  86.180000 ;
        RECT 37.945000  90.375000 42.400000  90.525000 ;
        RECT 37.945000 169.025000 48.835000 189.515000 ;
        RECT 38.035000 168.935000 48.835000 169.025000 ;
        RECT 38.095000  90.525000 42.550000  90.675000 ;
        RECT 38.185000 168.785000 48.835000 168.935000 ;
        RECT 38.245000  90.675000 42.700000  90.825000 ;
        RECT 38.335000 168.635000 48.835000 168.785000 ;
        RECT 38.395000  90.825000 42.850000  90.975000 ;
        RECT 38.485000 168.485000 48.835000 168.635000 ;
        RECT 38.545000  90.975000 43.000000  91.125000 ;
        RECT 38.635000 168.335000 48.835000 168.485000 ;
        RECT 38.695000  91.125000 43.150000  91.275000 ;
        RECT 38.785000 168.185000 48.835000 168.335000 ;
        RECT 38.845000  91.275000 43.300000  91.425000 ;
        RECT 38.935000 168.035000 48.835000 168.185000 ;
        RECT 38.995000  91.425000 43.450000  91.575000 ;
        RECT 39.085000 167.885000 48.835000 168.035000 ;
        RECT 39.145000  91.575000 43.600000  91.725000 ;
        RECT 39.235000 167.735000 48.835000 167.885000 ;
        RECT 39.295000  91.725000 43.750000  91.875000 ;
        RECT 39.385000 167.585000 48.835000 167.735000 ;
        RECT 39.445000  91.875000 43.900000  92.025000 ;
        RECT 39.535000 167.435000 48.835000 167.585000 ;
        RECT 39.595000  92.025000 44.050000  92.175000 ;
        RECT 39.685000 167.285000 48.835000 167.435000 ;
        RECT 39.745000  92.175000 44.200000  92.325000 ;
        RECT 39.835000 167.135000 48.835000 167.285000 ;
        RECT 39.895000  92.325000 44.350000  92.475000 ;
        RECT 39.985000 166.985000 48.835000 167.135000 ;
        RECT 40.045000  92.475000 44.500000  92.625000 ;
        RECT 40.135000 166.835000 48.835000 166.985000 ;
        RECT 40.195000  92.625000 44.650000  92.775000 ;
        RECT 40.285000 166.685000 48.835000 166.835000 ;
        RECT 40.345000  92.775000 44.800000  92.925000 ;
        RECT 40.435000 166.535000 48.835000 166.685000 ;
        RECT 40.495000  92.925000 44.950000  93.075000 ;
        RECT 40.585000 166.385000 48.835000 166.535000 ;
        RECT 40.645000  93.075000 45.100000  93.225000 ;
        RECT 40.735000 166.235000 48.835000 166.385000 ;
        RECT 40.795000  93.225000 45.250000  93.375000 ;
        RECT 40.885000 166.085000 48.835000 166.235000 ;
        RECT 40.945000  93.375000 45.400000  93.525000 ;
        RECT 41.035000 165.935000 48.835000 166.085000 ;
        RECT 41.050000  83.980000 48.870000  84.130000 ;
        RECT 41.095000  93.525000 45.550000  93.675000 ;
        RECT 41.185000 165.785000 48.835000 165.935000 ;
        RECT 41.200000  84.130000 48.870000  84.280000 ;
        RECT 41.245000  93.675000 45.700000  93.825000 ;
        RECT 41.335000 165.635000 48.835000 165.785000 ;
        RECT 41.350000  84.280000 48.870000  84.430000 ;
        RECT 41.395000  93.825000 45.850000  93.975000 ;
        RECT 41.485000 165.485000 48.835000 165.635000 ;
        RECT 41.500000  84.430000 48.870000  84.580000 ;
        RECT 41.545000  93.975000 46.000000  94.125000 ;
        RECT 41.610000  84.580000 48.870000  84.690000 ;
        RECT 41.610000  84.690000 48.870000  84.810000 ;
        RECT 41.610000  84.810000 48.870000  84.960000 ;
        RECT 41.610000  84.960000 49.020000  85.110000 ;
        RECT 41.610000  85.110000 49.170000  85.260000 ;
        RECT 41.610000  85.260000 49.320000  85.410000 ;
        RECT 41.610000  85.410000 49.470000  85.560000 ;
        RECT 41.610000  85.560000 49.620000  85.710000 ;
        RECT 41.610000  85.710000 49.770000  85.860000 ;
        RECT 41.610000  85.860000 49.920000  86.010000 ;
        RECT 41.610000  86.010000 50.070000  86.160000 ;
        RECT 41.610000  86.160000 50.220000  86.310000 ;
        RECT 41.610000  86.310000 50.370000  86.460000 ;
        RECT 41.610000  86.460000 50.520000  86.610000 ;
        RECT 41.610000  86.610000 50.670000  86.760000 ;
        RECT 41.610000  86.760000 50.820000  86.910000 ;
        RECT 41.610000  86.910000 50.970000  86.960000 ;
        RECT 41.610000  86.960000 51.020000  87.445000 ;
        RECT 41.635000 165.335000 48.835000 165.485000 ;
        RECT 41.695000  94.125000 46.150000  94.275000 ;
        RECT 41.760000  87.445000 51.020000  87.595000 ;
        RECT 41.785000 165.185000 48.835000 165.335000 ;
        RECT 41.845000  94.275000 46.300000  94.425000 ;
        RECT 41.910000  87.595000 51.020000  87.745000 ;
        RECT 41.935000 165.035000 48.835000 165.185000 ;
        RECT 41.995000  94.425000 46.450000  94.575000 ;
        RECT 42.060000  87.745000 51.020000  87.895000 ;
        RECT 42.085000 164.885000 48.835000 165.035000 ;
        RECT 42.145000  94.575000 46.600000  94.725000 ;
        RECT 42.210000  87.895000 51.020000  88.045000 ;
        RECT 42.235000 164.735000 48.835000 164.885000 ;
        RECT 42.295000  94.725000 46.750000  94.875000 ;
        RECT 42.360000  88.045000 51.020000  88.195000 ;
        RECT 42.385000 164.585000 48.835000 164.735000 ;
        RECT 42.445000  94.875000 46.900000  95.025000 ;
        RECT 42.510000  88.195000 51.020000  88.345000 ;
        RECT 42.535000 164.435000 48.835000 164.585000 ;
        RECT 42.540000  88.345000 51.020000  88.375000 ;
        RECT 42.595000  95.025000 47.050000  95.175000 ;
        RECT 42.685000 164.285000 48.835000 164.435000 ;
        RECT 42.690000  88.375000 51.020000  88.525000 ;
        RECT 42.745000  95.175000 47.200000  95.325000 ;
        RECT 42.835000  95.325000 47.350000  95.415000 ;
        RECT 42.835000  95.415000 47.440000  95.565000 ;
        RECT 42.835000  95.565000 47.590000  95.715000 ;
        RECT 42.835000  95.715000 47.740000  95.865000 ;
        RECT 42.835000  95.865000 47.890000  96.015000 ;
        RECT 42.835000  96.015000 48.040000  96.165000 ;
        RECT 42.835000  96.165000 48.190000  96.315000 ;
        RECT 42.835000  96.315000 48.340000  96.465000 ;
        RECT 42.835000  96.465000 48.490000  96.615000 ;
        RECT 42.835000  96.615000 48.640000  96.765000 ;
        RECT 42.835000  96.765000 48.790000  96.810000 ;
        RECT 42.835000  96.810000 48.835000 164.135000 ;
        RECT 42.835000 164.135000 48.835000 164.285000 ;
        RECT 42.840000  88.525000 51.170000  88.675000 ;
        RECT 42.990000  88.675000 51.320000  88.825000 ;
        RECT 43.140000  88.825000 51.470000  88.975000 ;
        RECT 43.290000  88.975000 51.620000  89.125000 ;
        RECT 43.440000  89.125000 51.770000  89.275000 ;
        RECT 43.590000  89.275000 51.920000  89.425000 ;
        RECT 43.740000  89.425000 52.070000  89.575000 ;
        RECT 43.890000  89.575000 52.220000  89.725000 ;
        RECT 44.040000  89.725000 52.370000  89.875000 ;
        RECT 44.190000  89.875000 52.520000  90.025000 ;
        RECT 44.340000  90.025000 52.670000  90.175000 ;
        RECT 44.490000  90.175000 52.820000  90.325000 ;
        RECT 44.640000  90.325000 52.970000  90.475000 ;
        RECT 44.790000  90.475000 53.120000  90.625000 ;
        RECT 44.940000  90.625000 53.270000  90.775000 ;
        RECT 45.090000  90.775000 53.420000  90.925000 ;
        RECT 45.240000  90.925000 53.570000  91.075000 ;
        RECT 45.390000  91.075000 53.720000  91.225000 ;
        RECT 45.540000  91.225000 53.870000  91.375000 ;
        RECT 45.690000  91.375000 54.020000  91.525000 ;
        RECT 45.840000  91.525000 54.170000  91.675000 ;
        RECT 45.990000  91.675000 54.320000  91.825000 ;
        RECT 46.140000  91.825000 54.470000  91.975000 ;
        RECT 46.290000  91.975000 54.620000  92.125000 ;
        RECT 46.440000  92.125000 54.770000  92.275000 ;
        RECT 46.590000  92.275000 54.920000  92.425000 ;
        RECT 46.740000  92.425000 55.070000  92.575000 ;
        RECT 46.890000  92.575000 55.220000  92.725000 ;
        RECT 47.040000  92.725000 55.370000  92.875000 ;
        RECT 47.190000  92.875000 55.520000  93.025000 ;
        RECT 47.340000  93.025000 55.670000  93.175000 ;
        RECT 47.490000  93.175000 55.820000  93.325000 ;
        RECT 47.640000  93.325000 55.970000  93.475000 ;
        RECT 47.790000  93.475000 56.120000  93.625000 ;
        RECT 47.940000  93.625000 56.270000  93.775000 ;
        RECT 48.090000  93.775000 56.420000  93.925000 ;
        RECT 48.240000  93.925000 56.570000  94.075000 ;
        RECT 48.390000  94.075000 56.720000  94.225000 ;
        RECT 48.540000  94.225000 56.870000  94.375000 ;
        RECT 48.690000  94.375000 57.020000  94.525000 ;
        RECT 48.840000  94.525000 57.170000  94.675000 ;
        RECT 48.990000  94.675000 57.320000  94.825000 ;
        RECT 49.140000  94.825000 57.470000  94.975000 ;
        RECT 49.290000  94.975000 57.620000  95.125000 ;
        RECT 49.440000  95.125000 57.770000  95.275000 ;
        RECT 49.590000  95.275000 57.920000  95.425000 ;
        RECT 49.740000  95.425000 58.070000  95.575000 ;
        RECT 49.870000 168.920000 60.330000 189.515000 ;
        RECT 49.890000  95.575000 58.220000  95.725000 ;
        RECT 49.980000 168.810000 60.330000 168.920000 ;
        RECT 50.040000  95.725000 58.370000  95.875000 ;
        RECT 50.130000 168.660000 60.330000 168.810000 ;
        RECT 50.190000  95.875000 58.520000  96.025000 ;
        RECT 50.280000 168.510000 60.330000 168.660000 ;
        RECT 50.340000  96.025000 58.670000  96.175000 ;
        RECT 50.430000 168.360000 60.330000 168.510000 ;
        RECT 50.490000  96.175000 58.820000  96.325000 ;
        RECT 50.580000 168.210000 60.330000 168.360000 ;
        RECT 50.640000  96.325000 58.970000  96.475000 ;
        RECT 50.730000 168.060000 60.330000 168.210000 ;
        RECT 50.790000  96.475000 59.120000  96.625000 ;
        RECT 50.880000 167.910000 60.330000 168.060000 ;
        RECT 50.940000  96.625000 59.270000  96.775000 ;
        RECT 51.030000 167.760000 60.330000 167.910000 ;
        RECT 51.090000  96.775000 59.420000  96.925000 ;
        RECT 51.180000 167.610000 60.330000 167.760000 ;
        RECT 51.240000  96.925000 59.570000  97.075000 ;
        RECT 51.330000 167.460000 60.330000 167.610000 ;
        RECT 51.390000  97.075000 59.720000  97.225000 ;
        RECT 51.480000 167.310000 60.330000 167.460000 ;
        RECT 51.540000  97.225000 59.870000  97.375000 ;
        RECT 51.630000 167.160000 60.330000 167.310000 ;
        RECT 51.690000  97.375000 60.020000  97.525000 ;
        RECT 51.780000 167.010000 60.330000 167.160000 ;
        RECT 51.840000  97.525000 60.170000  97.675000 ;
        RECT 51.850000  97.675000 60.320000  97.685000 ;
        RECT 51.930000 166.860000 60.330000 167.010000 ;
        RECT 52.000000  97.685000 60.330000  97.835000 ;
        RECT 52.080000 166.710000 60.330000 166.860000 ;
        RECT 52.150000  97.835000 60.330000  97.985000 ;
        RECT 52.230000 166.560000 60.330000 166.710000 ;
        RECT 52.300000  97.985000 60.330000  98.135000 ;
        RECT 52.380000 166.410000 60.330000 166.560000 ;
        RECT 52.450000  98.135000 60.330000  98.285000 ;
        RECT 52.530000 166.260000 60.330000 166.410000 ;
        RECT 52.600000  98.285000 60.330000  98.435000 ;
        RECT 52.680000 166.110000 60.330000 166.260000 ;
        RECT 52.750000  98.435000 60.330000  98.585000 ;
        RECT 52.830000 165.960000 60.330000 166.110000 ;
        RECT 52.900000  98.585000 60.330000  98.735000 ;
        RECT 52.980000 165.810000 60.330000 165.960000 ;
        RECT 53.050000  98.735000 60.330000  98.885000 ;
        RECT 53.130000 165.660000 60.330000 165.810000 ;
        RECT 53.200000  98.885000 60.330000  99.035000 ;
        RECT 53.280000 165.510000 60.330000 165.660000 ;
        RECT 53.350000  99.035000 60.330000  99.185000 ;
        RECT 53.430000 165.360000 60.330000 165.510000 ;
        RECT 53.500000  99.185000 60.330000  99.335000 ;
        RECT 53.580000 165.210000 60.330000 165.360000 ;
        RECT 53.650000  99.335000 60.330000  99.485000 ;
        RECT 53.730000 165.060000 60.330000 165.210000 ;
        RECT 53.800000  99.485000 60.330000  99.635000 ;
        RECT 53.880000 164.910000 60.330000 165.060000 ;
        RECT 53.950000  99.635000 60.330000  99.785000 ;
        RECT 54.030000 164.760000 60.330000 164.910000 ;
        RECT 54.100000  99.785000 60.330000  99.935000 ;
        RECT 54.180000 164.610000 60.330000 164.760000 ;
        RECT 54.250000  99.935000 60.330000 100.085000 ;
        RECT 54.330000 100.085000 60.330000 100.165000 ;
        RECT 54.330000 100.165000 60.330000 164.460000 ;
        RECT 54.330000 164.460000 60.330000 164.610000 ;
    END
  END DRN_LVC1
  PIN DRN_LVC2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 38.380000 0.000000 49.255000 69.490000 ;
    END
  END DRN_LVC2
  PIN G_CORE
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.500000  0.000000 24.500000  82.660000 ;
        RECT 0.500000 82.660000 24.350000  82.810000 ;
        RECT 0.500000 82.810000 24.200000  82.960000 ;
        RECT 0.500000 82.960000 24.050000  83.110000 ;
        RECT 0.500000 83.110000 23.900000  83.260000 ;
        RECT 0.500000 83.260000 23.750000  83.410000 ;
        RECT 0.500000 83.410000 23.600000  83.560000 ;
        RECT 0.500000 83.560000 23.450000  83.710000 ;
        RECT 0.500000 83.710000 23.300000  83.860000 ;
        RECT 0.500000 83.860000 23.150000  84.010000 ;
        RECT 0.500000 84.010000 23.000000  84.160000 ;
        RECT 0.500000 84.160000 22.850000  84.310000 ;
        RECT 0.500000 84.310000 22.700000  84.460000 ;
        RECT 0.500000 84.460000 22.550000  84.610000 ;
        RECT 0.500000 84.610000 22.400000  84.760000 ;
        RECT 0.500000 84.760000 22.250000  84.910000 ;
        RECT 0.500000 84.910000 22.100000  85.060000 ;
        RECT 0.500000 85.060000 21.950000  85.210000 ;
        RECT 0.500000 85.210000 21.800000  85.360000 ;
        RECT 0.500000 85.360000 21.650000  85.510000 ;
        RECT 0.500000 85.510000 21.500000  85.660000 ;
        RECT 0.500000 85.660000 21.350000  85.810000 ;
        RECT 0.500000 85.810000 21.200000  85.960000 ;
        RECT 0.500000 85.960000 21.050000  86.110000 ;
        RECT 0.500000 86.110000 20.900000  86.260000 ;
        RECT 0.500000 86.260000 20.750000  86.410000 ;
        RECT 0.500000 86.410000 20.600000  86.560000 ;
        RECT 0.500000 86.560000 20.450000  86.710000 ;
        RECT 0.500000 86.710000 20.300000  86.860000 ;
        RECT 0.500000 86.860000 20.150000  87.010000 ;
        RECT 0.500000 87.010000 20.000000  87.160000 ;
        RECT 0.500000 87.160000 19.850000  87.310000 ;
        RECT 0.500000 87.310000 19.700000  87.460000 ;
        RECT 0.500000 87.460000 19.550000  87.610000 ;
        RECT 0.500000 87.610000 19.400000  87.760000 ;
        RECT 0.500000 87.760000 19.250000  87.910000 ;
        RECT 0.500000 87.910000 19.100000  88.060000 ;
        RECT 0.500000 88.060000 18.950000  88.210000 ;
        RECT 0.500000 88.210000 18.800000  88.360000 ;
        RECT 0.500000 88.360000 18.650000  88.510000 ;
        RECT 0.500000 88.510000 18.500000  88.660000 ;
        RECT 0.500000 88.660000 18.350000  88.810000 ;
        RECT 0.500000 88.810000 18.200000  88.960000 ;
        RECT 0.500000 88.960000 18.050000  89.110000 ;
        RECT 0.500000 89.110000 17.900000  89.260000 ;
        RECT 0.500000 89.260000 17.750000  89.410000 ;
        RECT 0.500000 89.410000 17.600000  89.560000 ;
        RECT 0.500000 89.560000 17.450000  89.710000 ;
        RECT 0.500000 89.710000 17.300000  89.860000 ;
        RECT 0.500000 89.860000 17.150000  90.010000 ;
        RECT 0.500000 90.010000 17.000000  90.160000 ;
        RECT 0.500000 90.160000 16.850000  90.310000 ;
        RECT 0.500000 90.310000 16.700000  90.460000 ;
        RECT 0.500000 90.460000 16.550000  90.610000 ;
        RECT 0.500000 90.610000 16.400000  90.760000 ;
        RECT 0.500000 90.760000 16.250000  90.910000 ;
        RECT 0.500000 90.910000 16.100000  91.060000 ;
        RECT 0.500000 91.060000 15.950000  91.210000 ;
        RECT 0.500000 91.210000 15.800000  91.360000 ;
        RECT 0.500000 91.360000 15.650000  91.510000 ;
        RECT 0.500000 91.510000 15.500000  91.660000 ;
        RECT 0.500000 91.660000 15.350000  91.810000 ;
        RECT 0.500000 91.810000 15.200000  91.960000 ;
        RECT 0.500000 91.960000 15.050000  92.110000 ;
        RECT 0.500000 92.110000 14.900000  92.260000 ;
        RECT 0.500000 92.260000 14.750000  92.410000 ;
        RECT 0.500000 92.410000 14.600000  92.560000 ;
        RECT 0.500000 92.560000 14.450000  92.710000 ;
        RECT 0.500000 92.710000 14.300000  92.860000 ;
        RECT 0.500000 92.860000 14.150000  93.010000 ;
        RECT 0.500000 93.010000 14.000000  93.160000 ;
        RECT 0.500000 93.160000 13.850000  93.310000 ;
        RECT 0.500000 93.310000 13.700000  93.460000 ;
        RECT 0.500000 93.460000 13.550000  93.610000 ;
        RECT 0.500000 93.610000 13.400000  93.760000 ;
        RECT 0.500000 93.760000 13.250000  93.910000 ;
        RECT 0.500000 93.910000 13.100000  94.060000 ;
        RECT 0.500000 94.060000 12.950000  94.210000 ;
        RECT 0.500000 94.210000 12.900000  94.260000 ;
        RECT 0.500000 94.260000 12.900000 171.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755000  0.000000 74.700000  84.465000 ;
        RECT 50.905000 84.465000 74.700000  84.615000 ;
        RECT 51.055000 84.615000 74.700000  84.765000 ;
        RECT 51.205000 84.765000 74.700000  84.915000 ;
        RECT 51.355000 84.915000 74.700000  85.065000 ;
        RECT 51.505000 85.065000 74.700000  85.215000 ;
        RECT 51.655000 85.215000 74.700000  85.365000 ;
        RECT 51.805000 85.365000 74.700000  85.515000 ;
        RECT 51.955000 85.515000 74.700000  85.665000 ;
        RECT 52.105000 85.665000 74.700000  85.815000 ;
        RECT 52.255000 85.815000 74.700000  85.965000 ;
        RECT 52.405000 85.965000 74.700000  86.115000 ;
        RECT 52.555000 86.115000 74.700000  86.265000 ;
        RECT 52.705000 86.265000 74.700000  86.415000 ;
        RECT 52.855000 86.415000 74.700000  86.565000 ;
        RECT 53.005000 86.565000 74.700000  86.715000 ;
        RECT 53.155000 86.715000 74.700000  86.865000 ;
        RECT 53.305000 86.865000 74.700000  87.015000 ;
        RECT 53.455000 87.015000 74.700000  87.165000 ;
        RECT 53.605000 87.165000 74.700000  87.315000 ;
        RECT 53.755000 87.315000 74.700000  87.465000 ;
        RECT 53.905000 87.465000 74.700000  87.615000 ;
        RECT 54.055000 87.615000 74.700000  87.765000 ;
        RECT 54.205000 87.765000 74.700000  87.915000 ;
        RECT 54.355000 87.915000 74.700000  88.065000 ;
        RECT 54.505000 88.065000 74.700000  88.215000 ;
        RECT 54.655000 88.215000 74.700000  88.365000 ;
        RECT 54.805000 88.365000 74.700000  88.515000 ;
        RECT 54.955000 88.515000 74.700000  88.665000 ;
        RECT 55.105000 88.665000 74.700000  88.815000 ;
        RECT 55.255000 88.815000 74.700000  88.965000 ;
        RECT 55.405000 88.965000 74.700000  89.115000 ;
        RECT 55.555000 89.115000 74.700000  89.265000 ;
        RECT 55.705000 89.265000 74.700000  89.415000 ;
        RECT 55.855000 89.415000 74.700000  89.565000 ;
        RECT 56.005000 89.565000 74.700000  89.715000 ;
        RECT 56.155000 89.715000 74.700000  89.865000 ;
        RECT 56.305000 89.865000 74.700000  90.015000 ;
        RECT 56.455000 90.015000 74.700000  90.165000 ;
        RECT 56.605000 90.165000 74.700000  90.315000 ;
        RECT 56.755000 90.315000 74.700000  90.465000 ;
        RECT 56.905000 90.465000 74.700000  90.615000 ;
        RECT 57.055000 90.615000 74.700000  90.765000 ;
        RECT 57.205000 90.765000 74.700000  90.915000 ;
        RECT 57.355000 90.915000 74.700000  91.065000 ;
        RECT 57.505000 91.065000 74.700000  91.215000 ;
        RECT 57.655000 91.215000 74.700000  91.365000 ;
        RECT 57.805000 91.365000 74.700000  91.515000 ;
        RECT 57.955000 91.515000 74.700000  91.665000 ;
        RECT 58.105000 91.665000 74.700000  91.815000 ;
        RECT 58.255000 91.815000 74.700000  91.965000 ;
        RECT 58.405000 91.965000 74.700000  92.115000 ;
        RECT 58.555000 92.115000 74.700000  92.265000 ;
        RECT 58.705000 92.265000 74.700000  92.415000 ;
        RECT 58.855000 92.415000 74.700000  92.565000 ;
        RECT 59.005000 92.565000 74.700000  92.715000 ;
        RECT 59.155000 92.715000 74.700000  92.865000 ;
        RECT 59.305000 92.865000 74.700000  93.015000 ;
        RECT 59.455000 93.015000 74.700000  93.165000 ;
        RECT 59.605000 93.165000 74.700000  93.315000 ;
        RECT 59.755000 93.315000 74.700000  93.465000 ;
        RECT 59.905000 93.465000 74.700000  93.615000 ;
        RECT 60.055000 93.615000 74.700000  93.765000 ;
        RECT 60.205000 93.765000 74.700000  93.915000 ;
        RECT 60.355000 93.915000 74.700000  94.065000 ;
        RECT 60.505000 94.065000 74.700000  94.215000 ;
        RECT 60.655000 94.215000 74.700000  94.365000 ;
        RECT 60.805000 94.365000 74.700000  94.515000 ;
        RECT 60.955000 94.515000 74.700000  94.665000 ;
        RECT 61.105000 94.665000 74.700000  94.815000 ;
        RECT 61.255000 94.815000 74.700000  94.965000 ;
        RECT 61.405000 94.965000 74.700000  95.115000 ;
        RECT 61.555000 95.115000 74.700000  95.265000 ;
        RECT 61.705000 95.265000 74.700000  95.415000 ;
        RECT 61.855000 95.415000 74.700000  95.565000 ;
        RECT 62.005000 95.565000 74.700000  95.715000 ;
        RECT 62.045000 95.715000 74.700000  95.755000 ;
        RECT 62.045000 95.755000 74.700000 172.235000 ;
    END
  END G_CORE
  PIN OGC_LVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 26.210000 0.000000 27.700000 0.170000 ;
    END
  END OGC_LVC
  PIN SRC_BDY_LVC1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT  0.500000   0.000000 20.495000   1.485000 ;
        RECT  0.500000   1.485000 20.425000   1.555000 ;
        RECT  0.500000   1.555000 20.355000   1.625000 ;
        RECT  0.500000   1.625000 20.285000   1.695000 ;
        RECT  0.500000   1.695000 20.215000   1.765000 ;
        RECT  0.500000   1.765000 20.145000   1.835000 ;
        RECT  0.500000   1.835000 20.075000   1.905000 ;
        RECT  0.500000   1.905000 20.005000   1.975000 ;
        RECT  0.500000   1.975000 19.935000   2.045000 ;
        RECT  0.500000   2.045000 19.865000   2.115000 ;
        RECT  0.500000   2.115000 19.795000   2.185000 ;
        RECT  0.500000   2.185000 19.725000   2.255000 ;
        RECT  0.500000   2.255000 19.655000   2.325000 ;
        RECT  0.500000   2.325000 19.585000   2.395000 ;
        RECT  0.500000   2.395000 19.515000   2.465000 ;
        RECT  0.500000   2.465000 19.445000   2.535000 ;
        RECT  0.500000   2.535000 19.375000   2.605000 ;
        RECT  0.500000   2.605000 19.305000   2.675000 ;
        RECT  0.500000   2.675000 19.235000   2.745000 ;
        RECT  0.500000   2.745000 19.165000   2.815000 ;
        RECT  0.500000   2.815000 19.095000   2.885000 ;
        RECT  0.500000   2.885000 19.025000   2.955000 ;
        RECT  0.500000   2.955000 18.955000   3.025000 ;
        RECT  0.500000   3.025000 18.885000   3.095000 ;
        RECT  0.500000   3.095000 18.815000   3.165000 ;
        RECT  0.500000   3.165000 18.745000   3.235000 ;
        RECT  0.500000   3.235000 18.675000   3.305000 ;
        RECT  0.500000   3.305000 18.605000   3.375000 ;
        RECT  0.500000   3.375000 18.535000   3.445000 ;
        RECT  0.500000   3.445000 18.465000   3.515000 ;
        RECT  0.500000   3.515000 18.395000   3.585000 ;
        RECT  0.500000   3.585000 18.325000   3.655000 ;
        RECT  0.500000   3.655000 18.255000   3.725000 ;
        RECT  0.500000   3.725000 18.185000   3.795000 ;
        RECT  0.500000   3.795000 18.115000   3.865000 ;
        RECT  0.500000   3.865000 18.045000   3.935000 ;
        RECT  0.500000   3.935000 17.975000   4.005000 ;
        RECT  0.500000   4.005000 17.905000   4.075000 ;
        RECT  0.500000   4.075000 17.835000   4.145000 ;
        RECT  0.500000   4.145000 17.765000   4.215000 ;
        RECT  0.500000   4.215000 17.695000   4.285000 ;
        RECT  0.500000   4.285000 17.625000   4.355000 ;
        RECT  0.500000   4.355000 17.555000   4.425000 ;
        RECT  0.500000   4.425000 17.485000   4.495000 ;
        RECT  0.500000   4.495000 17.415000   4.565000 ;
        RECT  0.500000   4.565000 17.345000   4.635000 ;
        RECT  0.500000   4.635000 17.275000   4.705000 ;
        RECT  0.500000   4.705000 17.205000   4.775000 ;
        RECT  0.500000   4.775000 17.135000   4.845000 ;
        RECT  0.500000   4.845000 17.065000   4.915000 ;
        RECT  0.500000   4.915000 16.995000   4.985000 ;
        RECT  0.500000   4.985000 16.925000   5.055000 ;
        RECT  0.500000   5.055000 16.860000   5.120000 ;
        RECT  0.500000   5.120000 16.860000   7.655000 ;
        RECT  0.500000   7.655000 10.745000   7.725000 ;
        RECT  0.500000   7.725000 10.675000   7.795000 ;
        RECT  0.500000   7.795000 10.605000   7.865000 ;
        RECT  0.500000   7.865000 10.535000   7.935000 ;
        RECT  0.500000   7.935000 10.465000   8.005000 ;
        RECT  0.500000   8.005000 10.420000   8.050000 ;
        RECT  0.500000   8.050000 10.420000   9.820000 ;
        RECT  0.500000   9.820000 10.420000   9.890000 ;
        RECT  0.500000   9.890000 10.490000   9.960000 ;
        RECT  0.500000   9.960000 10.560000  10.030000 ;
        RECT  0.500000  10.030000 10.630000  10.100000 ;
        RECT  0.500000  10.100000 10.700000  10.170000 ;
        RECT  0.500000  10.170000 10.770000  10.215000 ;
        RECT  0.500000  10.215000 55.595000  17.080000 ;
        RECT  0.500000  17.080000 21.785000  17.150000 ;
        RECT  0.500000  17.150000 21.715000  17.220000 ;
        RECT  0.500000  17.220000 21.645000  17.290000 ;
        RECT  0.500000  17.290000 21.575000  17.360000 ;
        RECT  0.500000  17.360000 21.505000  17.430000 ;
        RECT  0.500000  17.430000 21.435000  17.500000 ;
        RECT  0.500000  17.500000 21.365000  17.570000 ;
        RECT  0.500000  17.570000 21.295000  17.640000 ;
        RECT  0.500000  17.640000 21.225000  17.710000 ;
        RECT  0.500000  17.710000 21.155000  17.780000 ;
        RECT  0.500000  17.780000 21.085000  17.850000 ;
        RECT  0.500000  17.850000 21.015000  17.920000 ;
        RECT  0.500000  17.920000 20.945000  17.990000 ;
        RECT  0.500000  17.990000 20.875000  18.060000 ;
        RECT  0.500000  18.060000 20.805000  18.130000 ;
        RECT  0.500000  18.130000 20.735000  18.200000 ;
        RECT  0.500000  18.200000 20.665000  18.270000 ;
        RECT  0.500000  18.270000 20.595000  18.340000 ;
        RECT  0.500000  18.340000 20.525000  18.410000 ;
        RECT  0.500000  18.410000 20.455000  18.480000 ;
        RECT  0.500000  18.480000 20.385000  18.550000 ;
        RECT  0.500000  18.550000 20.315000  18.620000 ;
        RECT  0.500000  18.620000 20.245000  18.690000 ;
        RECT  0.500000  18.690000 20.175000  18.760000 ;
        RECT  0.500000  18.760000 20.105000  18.830000 ;
        RECT  0.500000  18.830000 20.035000  18.900000 ;
        RECT  0.500000  18.900000 19.965000  18.970000 ;
        RECT  0.500000  18.970000 19.895000  19.040000 ;
        RECT  0.500000  19.040000 19.825000  19.110000 ;
        RECT  0.500000  19.110000 19.755000  19.180000 ;
        RECT  0.500000  19.180000 19.685000  19.250000 ;
        RECT  0.500000  19.250000 19.615000  19.320000 ;
        RECT  0.500000  19.320000 19.545000  19.390000 ;
        RECT  0.500000  19.390000 19.475000  19.460000 ;
        RECT  0.500000  19.460000 19.405000  19.530000 ;
        RECT  0.500000  19.530000 19.335000  19.600000 ;
        RECT  0.500000  19.600000 19.265000  19.670000 ;
        RECT  0.500000  19.670000 19.195000  19.740000 ;
        RECT  0.500000  19.740000 19.125000  19.810000 ;
        RECT  0.500000  19.810000 19.055000  19.880000 ;
        RECT  0.500000  19.880000 18.985000  19.950000 ;
        RECT  0.500000  19.950000 18.915000  20.020000 ;
        RECT  0.500000  20.020000 18.845000  20.090000 ;
        RECT  0.500000  20.090000 18.775000  20.160000 ;
        RECT  0.500000  20.160000 18.705000  20.230000 ;
        RECT  0.500000  20.230000 18.635000  20.300000 ;
        RECT  0.500000  20.300000 18.565000  20.370000 ;
        RECT  0.500000  20.370000 18.495000  20.440000 ;
        RECT  0.500000  20.440000 18.425000  20.510000 ;
        RECT  0.500000  20.510000 18.355000  20.580000 ;
        RECT  0.500000  20.580000 18.285000  20.650000 ;
        RECT  0.500000  20.650000 18.215000  20.720000 ;
        RECT  0.500000  20.720000 18.145000  20.790000 ;
        RECT  0.500000  20.790000 18.075000  20.860000 ;
        RECT  0.500000  20.860000 18.005000  20.930000 ;
        RECT  0.500000  20.930000 17.935000  21.000000 ;
        RECT  0.500000  21.000000 17.865000  21.070000 ;
        RECT  0.500000  21.070000 17.795000  21.140000 ;
        RECT  0.500000  21.140000 17.725000  21.210000 ;
        RECT  0.500000  21.210000 17.655000  21.280000 ;
        RECT  0.500000  21.280000 17.585000  21.350000 ;
        RECT  0.500000  21.350000 17.515000  21.420000 ;
        RECT  0.500000  21.420000 17.445000  21.490000 ;
        RECT  0.500000  21.490000 17.375000  21.560000 ;
        RECT  0.500000  21.560000 17.305000  21.630000 ;
        RECT  0.500000  21.630000 17.235000  21.700000 ;
        RECT  0.500000  21.700000 17.165000  21.770000 ;
        RECT  0.500000  21.770000 17.095000  21.840000 ;
        RECT  0.500000  21.840000 17.025000  21.910000 ;
        RECT  0.500000  21.910000 16.955000  21.980000 ;
        RECT  0.500000  21.980000 16.885000  22.050000 ;
        RECT  0.500000  22.050000 16.815000  22.120000 ;
        RECT  0.500000  22.120000 16.745000  22.190000 ;
        RECT  0.500000  22.190000 16.675000  22.260000 ;
        RECT  0.500000  22.260000 16.605000  22.330000 ;
        RECT  0.500000  22.330000 16.535000  22.400000 ;
        RECT  0.500000  22.400000 16.465000  22.470000 ;
        RECT  0.500000  22.470000 16.395000  22.540000 ;
        RECT  0.500000  22.540000 16.325000  22.610000 ;
        RECT  0.500000  22.610000 16.255000  22.680000 ;
        RECT  0.500000  22.680000 16.185000  22.750000 ;
        RECT  0.500000  22.750000 16.115000  22.820000 ;
        RECT  0.500000  22.820000 16.045000  22.890000 ;
        RECT  0.500000  22.890000 15.975000  22.960000 ;
        RECT  0.500000  22.960000 15.905000  23.030000 ;
        RECT  0.500000  23.030000 15.835000  23.100000 ;
        RECT  0.500000  23.100000 15.765000  23.170000 ;
        RECT  0.500000  23.170000 15.695000  23.240000 ;
        RECT  0.500000  23.240000 15.625000  23.310000 ;
        RECT  0.500000  23.310000 15.555000  23.380000 ;
        RECT  0.500000  23.380000 15.485000  23.450000 ;
        RECT  0.500000  23.450000 15.415000  23.520000 ;
        RECT  0.500000  23.520000 15.345000  23.590000 ;
        RECT  0.500000  23.590000 15.275000  23.660000 ;
        RECT  0.500000  23.660000 15.205000  23.730000 ;
        RECT  0.500000  23.730000 15.135000  23.800000 ;
        RECT  0.500000  23.800000 15.065000  23.870000 ;
        RECT  0.500000  23.870000 14.995000  23.940000 ;
        RECT  0.500000  23.940000 14.925000  24.010000 ;
        RECT  0.500000  24.010000 14.855000  24.080000 ;
        RECT  0.500000  24.080000 14.785000  24.150000 ;
        RECT  0.500000  24.150000 14.715000  24.220000 ;
        RECT  0.500000  24.220000 14.645000  24.290000 ;
        RECT  0.500000  24.290000 14.575000  24.360000 ;
        RECT  0.500000  24.360000 14.505000  24.430000 ;
        RECT  0.500000  24.430000 14.435000  24.500000 ;
        RECT  0.500000  24.500000 14.365000  24.570000 ;
        RECT  0.500000  24.570000 14.295000  24.640000 ;
        RECT  0.500000  24.640000 14.225000  24.710000 ;
        RECT  0.500000  24.710000 14.155000  24.780000 ;
        RECT  0.500000  24.780000 14.085000  24.850000 ;
        RECT  0.500000  24.850000 14.015000  24.920000 ;
        RECT  0.500000  24.920000 13.945000  24.990000 ;
        RECT  0.500000  24.990000 13.875000  25.060000 ;
        RECT  0.500000  25.060000 13.805000  25.130000 ;
        RECT  0.500000  25.130000 13.750000  25.185000 ;
        RECT  0.500000  25.185000 13.750000  74.295000 ;
        RECT  0.500000  74.295000 13.750000  74.365000 ;
        RECT  0.500000  74.365000 13.820000  74.435000 ;
        RECT  0.500000  74.435000 13.890000  74.505000 ;
        RECT  0.500000  74.505000 13.960000 129.935000 ;
        RECT  0.500000 129.935000 13.960000 130.005000 ;
        RECT  0.500000 130.005000 14.030000 130.075000 ;
        RECT  0.500000 130.075000 14.100000 130.145000 ;
        RECT  0.500000 130.145000 14.170000 130.215000 ;
        RECT  0.500000 130.215000 14.240000 130.285000 ;
        RECT  0.500000 130.285000 14.310000 130.355000 ;
        RECT  0.500000 130.355000 14.380000 130.425000 ;
        RECT  0.500000 130.425000 14.450000 130.495000 ;
        RECT  0.500000 130.495000 14.520000 130.565000 ;
        RECT  0.500000 130.565000 14.590000 130.635000 ;
        RECT  0.500000 130.635000 14.660000 130.705000 ;
        RECT  0.500000 130.705000 14.730000 130.775000 ;
        RECT  0.500000 130.775000 14.800000 130.845000 ;
        RECT  0.500000 130.845000 14.870000 130.915000 ;
        RECT  0.500000 130.915000 14.940000 130.985000 ;
        RECT  0.500000 130.985000 68.010000 133.630000 ;
        RECT  0.500000 133.630000 14.940000 133.700000 ;
        RECT  0.500000 133.700000 14.870000 133.770000 ;
        RECT  0.500000 133.770000 14.800000 133.840000 ;
        RECT  0.500000 133.840000 14.730000 133.910000 ;
        RECT  0.500000 133.910000 14.660000 133.980000 ;
        RECT  0.500000 133.980000 14.590000 134.050000 ;
        RECT  0.500000 134.050000 14.520000 134.120000 ;
        RECT  0.500000 134.120000 14.450000 134.190000 ;
        RECT  0.500000 134.190000 14.380000 134.260000 ;
        RECT  0.500000 134.260000 14.310000 134.330000 ;
        RECT  0.500000 134.330000 14.240000 134.400000 ;
        RECT  0.500000 134.400000 14.170000 134.470000 ;
        RECT  0.500000 134.470000 14.100000 134.540000 ;
        RECT  0.500000 134.540000 14.030000 134.610000 ;
        RECT  0.500000 134.610000 13.960000 134.680000 ;
        RECT  0.500000 134.680000 13.960000 139.940000 ;
        RECT  0.500000 139.940000 13.960000 140.010000 ;
        RECT  0.500000 140.010000 14.030000 140.080000 ;
        RECT  0.500000 140.080000 14.100000 140.150000 ;
        RECT  0.500000 140.150000 14.170000 140.220000 ;
        RECT  0.500000 140.220000 14.240000 140.290000 ;
        RECT  0.500000 140.290000 14.310000 140.360000 ;
        RECT  0.500000 140.360000 14.380000 140.430000 ;
        RECT  0.500000 140.430000 14.450000 140.500000 ;
        RECT  0.500000 140.500000 14.520000 140.570000 ;
        RECT  0.500000 140.570000 14.590000 140.640000 ;
        RECT  0.500000 140.640000 14.660000 140.710000 ;
        RECT  0.500000 140.710000 14.730000 140.780000 ;
        RECT  0.500000 140.780000 14.800000 140.850000 ;
        RECT  0.500000 140.850000 14.870000 140.920000 ;
        RECT  0.500000 140.920000 14.940000 140.990000 ;
        RECT  0.500000 140.990000 68.010000 143.630000 ;
        RECT  0.500000 143.630000 14.940000 143.700000 ;
        RECT  0.500000 143.700000 14.870000 143.770000 ;
        RECT  0.500000 143.770000 14.800000 143.840000 ;
        RECT  0.500000 143.840000 14.730000 143.910000 ;
        RECT  0.500000 143.910000 14.660000 143.980000 ;
        RECT  0.500000 143.980000 14.590000 144.050000 ;
        RECT  0.500000 144.050000 14.520000 144.120000 ;
        RECT  0.500000 144.120000 14.450000 144.190000 ;
        RECT  0.500000 144.190000 14.380000 144.260000 ;
        RECT  0.500000 144.260000 14.310000 144.330000 ;
        RECT  0.500000 144.330000 14.240000 144.400000 ;
        RECT  0.500000 144.400000 14.170000 144.470000 ;
        RECT  0.500000 144.470000 14.100000 144.540000 ;
        RECT  0.500000 144.540000 14.030000 144.610000 ;
        RECT  0.500000 144.610000 13.960000 144.680000 ;
        RECT  0.500000 144.680000 13.960000 149.940000 ;
        RECT  0.500000 149.940000 13.960000 150.010000 ;
        RECT  0.500000 150.010000 14.030000 150.080000 ;
        RECT  0.500000 150.080000 14.100000 150.150000 ;
        RECT  0.500000 150.150000 14.170000 150.220000 ;
        RECT  0.500000 150.220000 14.240000 150.290000 ;
        RECT  0.500000 150.290000 14.310000 150.360000 ;
        RECT  0.500000 150.360000 14.380000 150.430000 ;
        RECT  0.500000 150.430000 14.450000 150.500000 ;
        RECT  0.500000 150.500000 14.520000 150.570000 ;
        RECT  0.500000 150.570000 14.590000 150.640000 ;
        RECT  0.500000 150.640000 14.660000 150.710000 ;
        RECT  0.500000 150.710000 14.730000 150.780000 ;
        RECT  0.500000 150.780000 14.800000 150.850000 ;
        RECT  0.500000 150.850000 14.870000 150.920000 ;
        RECT  0.500000 150.920000 14.940000 150.990000 ;
        RECT  0.500000 150.990000 68.010000 153.630000 ;
        RECT  0.500000 153.630000 14.940000 153.700000 ;
        RECT  0.500000 153.700000 14.870000 153.770000 ;
        RECT  0.500000 153.770000 14.800000 153.840000 ;
        RECT  0.500000 153.840000 14.730000 153.910000 ;
        RECT  0.500000 153.910000 14.660000 153.980000 ;
        RECT  0.500000 153.980000 14.590000 154.050000 ;
        RECT  0.500000 154.050000 14.520000 154.120000 ;
        RECT  0.500000 154.120000 14.450000 154.190000 ;
        RECT  0.500000 154.190000 14.380000 154.260000 ;
        RECT  0.500000 154.260000 14.310000 154.330000 ;
        RECT  0.500000 154.330000 14.240000 154.400000 ;
        RECT  0.500000 154.400000 14.170000 154.470000 ;
        RECT  0.500000 154.470000 14.100000 154.540000 ;
        RECT  0.500000 154.540000 14.030000 154.610000 ;
        RECT  0.500000 154.610000 13.960000 154.680000 ;
        RECT  0.500000 154.680000 13.960000 159.940000 ;
        RECT  0.500000 159.940000 13.960000 160.010000 ;
        RECT  0.500000 160.010000 14.030000 160.080000 ;
        RECT  0.500000 160.080000 14.100000 160.150000 ;
        RECT  0.500000 160.150000 14.170000 160.220000 ;
        RECT  0.500000 160.220000 14.240000 160.290000 ;
        RECT  0.500000 160.290000 14.310000 160.360000 ;
        RECT  0.500000 160.360000 14.380000 160.430000 ;
        RECT  0.500000 160.430000 14.450000 160.500000 ;
        RECT  0.500000 160.500000 14.520000 160.570000 ;
        RECT  0.500000 160.570000 14.590000 160.640000 ;
        RECT  0.500000 160.640000 14.660000 160.710000 ;
        RECT  0.500000 160.710000 14.730000 160.780000 ;
        RECT  0.500000 160.780000 14.800000 160.850000 ;
        RECT  0.500000 160.850000 14.870000 160.920000 ;
        RECT  0.500000 160.920000 14.940000 160.990000 ;
        RECT  0.500000 160.990000 68.010000 163.630000 ;
        RECT  0.500000 163.630000 14.940000 163.700000 ;
        RECT  0.500000 163.700000 14.870000 163.770000 ;
        RECT  0.500000 163.770000 14.800000 163.840000 ;
        RECT  0.500000 163.840000 14.730000 163.910000 ;
        RECT  0.500000 163.910000 14.660000 163.980000 ;
        RECT  0.500000 163.980000 14.590000 164.050000 ;
        RECT  0.500000 164.050000 14.520000 164.120000 ;
        RECT  0.500000 164.120000 14.450000 164.190000 ;
        RECT  0.500000 164.190000 14.380000 164.260000 ;
        RECT  0.500000 164.260000 14.310000 164.330000 ;
        RECT  0.500000 164.330000 14.240000 164.400000 ;
        RECT  0.500000 164.400000 14.170000 164.470000 ;
        RECT  0.500000 164.470000 14.100000 164.540000 ;
        RECT  0.500000 164.540000 14.030000 164.610000 ;
        RECT  0.500000 164.610000 13.960000 164.680000 ;
        RECT  0.500000 164.680000 13.960000 169.940000 ;
        RECT  0.500000 169.940000 13.960000 170.010000 ;
        RECT  0.500000 170.010000 14.030000 170.080000 ;
        RECT  0.500000 170.080000 14.100000 170.150000 ;
        RECT  0.500000 170.150000 14.170000 170.220000 ;
        RECT  0.500000 170.220000 14.240000 170.290000 ;
        RECT  0.500000 170.290000 14.310000 170.360000 ;
        RECT  0.500000 170.360000 14.380000 170.430000 ;
        RECT  0.500000 170.430000 14.450000 170.500000 ;
        RECT  0.500000 170.500000 14.520000 170.570000 ;
        RECT  0.500000 170.570000 14.590000 170.640000 ;
        RECT  0.500000 170.640000 14.660000 170.710000 ;
        RECT  0.500000 170.710000 14.730000 170.780000 ;
        RECT  0.500000 170.780000 14.800000 170.850000 ;
        RECT  0.500000 170.850000 14.870000 170.920000 ;
        RECT  0.500000 170.920000 14.940000 170.990000 ;
        RECT  0.500000 170.990000 68.010000 173.630000 ;
        RECT  0.500000 173.630000 14.940000 173.700000 ;
        RECT  0.500000 173.700000 14.870000 173.770000 ;
        RECT  0.500000 173.770000 14.800000 173.840000 ;
        RECT  0.500000 173.840000 14.730000 173.910000 ;
        RECT  0.500000 173.910000 14.660000 173.980000 ;
        RECT  0.500000 173.980000 14.590000 174.050000 ;
        RECT  0.500000 174.050000 14.520000 174.120000 ;
        RECT  0.500000 174.120000 14.450000 174.190000 ;
        RECT  0.500000 174.190000 14.380000 174.260000 ;
        RECT  0.500000 174.260000 14.310000 174.330000 ;
        RECT  0.500000 174.330000 14.240000 174.400000 ;
        RECT  0.500000 174.400000 14.170000 174.470000 ;
        RECT  0.500000 174.470000 14.100000 174.540000 ;
        RECT  0.500000 174.540000 14.030000 174.610000 ;
        RECT  0.500000 174.610000 13.960000 174.680000 ;
        RECT  0.500000 174.680000 13.960000 179.940000 ;
        RECT  0.500000 179.940000 13.960000 180.010000 ;
        RECT  0.500000 180.010000 14.030000 180.080000 ;
        RECT  0.500000 180.080000 14.100000 180.150000 ;
        RECT  0.500000 180.150000 14.170000 180.220000 ;
        RECT  0.500000 180.220000 14.240000 180.290000 ;
        RECT  0.500000 180.290000 14.310000 180.360000 ;
        RECT  0.500000 180.360000 14.380000 180.430000 ;
        RECT  0.500000 180.430000 14.450000 180.500000 ;
        RECT  0.500000 180.500000 14.520000 180.570000 ;
        RECT  0.500000 180.570000 14.590000 180.640000 ;
        RECT  0.500000 180.640000 14.660000 180.710000 ;
        RECT  0.500000 180.710000 14.730000 180.780000 ;
        RECT  0.500000 180.780000 14.800000 180.850000 ;
        RECT  0.500000 180.850000 14.870000 180.920000 ;
        RECT  0.500000 180.920000 14.940000 180.990000 ;
        RECT  0.500000 180.990000 68.010000 183.630000 ;
        RECT  0.500000 183.630000 14.940000 183.700000 ;
        RECT  0.500000 183.700000 14.870000 183.770000 ;
        RECT  0.500000 183.770000 14.800000 183.840000 ;
        RECT  0.500000 183.840000 14.730000 183.910000 ;
        RECT  0.500000 183.910000 14.660000 183.980000 ;
        RECT  0.500000 183.980000 14.590000 184.050000 ;
        RECT  0.500000 184.050000 14.520000 184.120000 ;
        RECT  0.500000 184.120000 14.450000 184.190000 ;
        RECT  0.500000 184.190000 14.380000 184.260000 ;
        RECT  0.500000 184.260000 14.310000 184.330000 ;
        RECT  0.500000 184.330000 14.240000 184.400000 ;
        RECT  0.500000 184.400000 14.170000 184.470000 ;
        RECT  0.500000 184.470000 14.100000 184.540000 ;
        RECT  0.500000 184.540000 14.030000 184.610000 ;
        RECT  0.500000 184.610000 13.960000 184.680000 ;
        RECT  0.500000 184.680000 13.960000 189.940000 ;
        RECT  0.500000 189.940000 13.960000 190.010000 ;
        RECT  0.500000 190.010000 14.030000 190.080000 ;
        RECT  0.500000 190.080000 14.100000 190.150000 ;
        RECT  0.500000 190.150000 14.170000 190.220000 ;
        RECT  0.500000 190.220000 14.240000 190.290000 ;
        RECT  0.500000 190.290000 14.310000 190.360000 ;
        RECT  0.500000 190.360000 14.380000 190.430000 ;
        RECT  0.500000 190.430000 14.450000 190.500000 ;
        RECT  0.500000 190.500000 14.520000 190.570000 ;
        RECT  0.500000 190.570000 14.590000 190.640000 ;
        RECT  0.500000 190.640000 14.660000 190.710000 ;
        RECT  0.500000 190.710000 14.730000 190.780000 ;
        RECT  0.500000 190.780000 14.800000 190.850000 ;
        RECT  0.500000 190.850000 14.870000 190.920000 ;
        RECT  0.500000 190.920000 14.940000 190.990000 ;
        RECT  0.500000 190.990000 68.010000 193.630000 ;
        RECT 11.635000  10.210000 55.595000  10.215000 ;
        RECT 11.695000   7.655000 16.860000   7.725000 ;
        RECT 11.700000  10.145000 55.595000  10.210000 ;
        RECT 11.765000   7.725000 16.860000   7.795000 ;
        RECT 11.765000  10.080000 55.595000  10.145000 ;
        RECT 11.805000  10.040000 17.535000  10.080000 ;
        RECT 11.835000   7.795000 16.860000   7.865000 ;
        RECT 11.875000   9.970000 17.465000  10.040000 ;
        RECT 11.905000   7.865000 16.860000   7.935000 ;
        RECT 11.945000   9.900000 17.395000   9.970000 ;
        RECT 11.975000   7.935000 16.860000   8.005000 ;
        RECT 12.015000   8.005000 16.860000   8.045000 ;
        RECT 12.015000   8.045000 16.860000   9.365000 ;
        RECT 12.015000   9.365000 16.860000   9.435000 ;
        RECT 12.015000   9.435000 16.930000   9.505000 ;
        RECT 12.015000   9.505000 17.000000   9.575000 ;
        RECT 12.015000   9.575000 17.070000   9.645000 ;
        RECT 12.015000   9.645000 17.140000   9.715000 ;
        RECT 12.015000   9.715000 17.210000   9.785000 ;
        RECT 12.015000   9.785000 17.280000   9.830000 ;
        RECT 12.015000   9.830000 17.325000   9.900000 ;
    END
  END SRC_BDY_LVC1
  PIN SRC_BDY_LVC2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 16.135000 31.010000 74.700000 33.650000 ;
        RECT 16.135000 40.990000 74.700000 43.630000 ;
        RECT 16.135000 51.010000 74.700000 53.650000 ;
        RECT 16.135000 60.990000 74.700000 63.630000 ;
        RECT 16.135000 70.990000 74.700000 73.630000 ;
        RECT 54.095000  0.000000 74.700000  7.815000 ;
        RECT 54.095000 19.990000 74.700000 21.695000 ;
        RECT 54.150000 19.935000 74.700000 19.990000 ;
        RECT 54.165000  7.815000 74.700000  7.885000 ;
        RECT 54.220000 19.865000 74.700000 19.935000 ;
        RECT 54.235000  7.885000 74.700000  7.955000 ;
        RECT 54.290000 19.795000 74.700000 19.865000 ;
        RECT 54.305000  7.955000 74.700000  8.025000 ;
        RECT 54.360000 19.725000 74.700000 19.795000 ;
        RECT 54.375000  8.025000 74.700000  8.095000 ;
        RECT 54.430000 19.655000 74.700000 19.725000 ;
        RECT 54.445000  8.095000 74.700000  8.165000 ;
        RECT 54.500000 19.585000 74.700000 19.655000 ;
        RECT 54.515000  8.165000 74.700000  8.235000 ;
        RECT 54.570000 19.515000 74.700000 19.585000 ;
        RECT 54.585000  8.235000 74.700000  8.305000 ;
        RECT 54.640000 19.445000 74.700000 19.515000 ;
        RECT 54.655000  8.305000 74.700000  8.375000 ;
        RECT 54.710000 19.375000 74.700000 19.445000 ;
        RECT 54.725000  8.375000 74.700000  8.445000 ;
        RECT 54.780000 19.305000 74.700000 19.375000 ;
        RECT 54.795000  8.445000 74.700000  8.515000 ;
        RECT 54.850000 19.235000 74.700000 19.305000 ;
        RECT 54.865000  8.515000 74.700000  8.585000 ;
        RECT 54.920000 19.165000 74.700000 19.235000 ;
        RECT 54.935000  8.585000 74.700000  8.655000 ;
        RECT 54.990000 19.095000 74.700000 19.165000 ;
        RECT 55.005000  8.655000 74.700000  8.725000 ;
        RECT 55.060000 19.025000 74.700000 19.095000 ;
        RECT 55.075000  8.725000 74.700000  8.795000 ;
        RECT 55.130000 18.955000 74.700000 19.025000 ;
        RECT 55.145000  8.795000 74.700000  8.865000 ;
        RECT 55.200000 18.885000 74.700000 18.955000 ;
        RECT 55.215000  8.865000 74.700000  8.935000 ;
        RECT 55.270000 18.815000 74.700000 18.885000 ;
        RECT 55.285000  8.935000 74.700000  9.005000 ;
        RECT 55.340000 18.745000 74.700000 18.815000 ;
        RECT 55.355000  9.005000 74.700000  9.075000 ;
        RECT 55.410000 18.675000 74.700000 18.745000 ;
        RECT 55.425000  9.075000 74.700000  9.145000 ;
        RECT 55.480000 18.605000 74.700000 18.675000 ;
        RECT 55.495000  9.145000 74.700000  9.215000 ;
        RECT 55.550000 18.535000 74.700000 18.605000 ;
        RECT 55.565000  9.215000 74.700000  9.285000 ;
        RECT 55.620000 18.465000 74.700000 18.535000 ;
        RECT 55.635000  9.285000 74.700000  9.355000 ;
        RECT 55.690000 18.395000 74.700000 18.465000 ;
        RECT 55.705000  9.355000 74.700000  9.425000 ;
        RECT 55.760000 18.325000 74.700000 18.395000 ;
        RECT 55.775000  9.425000 74.700000  9.495000 ;
        RECT 55.830000 18.255000 74.700000 18.325000 ;
        RECT 55.845000  9.495000 74.700000  9.565000 ;
        RECT 55.900000 18.185000 74.700000 18.255000 ;
        RECT 55.915000  9.565000 74.700000  9.635000 ;
        RECT 55.970000 18.115000 74.700000 18.185000 ;
        RECT 55.985000  9.635000 74.700000  9.705000 ;
        RECT 56.040000 18.045000 74.700000 18.115000 ;
        RECT 56.055000  9.705000 74.700000  9.775000 ;
        RECT 56.110000 17.975000 74.700000 18.045000 ;
        RECT 56.125000  9.775000 74.700000  9.845000 ;
        RECT 56.180000 17.905000 74.700000 17.975000 ;
        RECT 56.195000  9.845000 74.700000  9.915000 ;
        RECT 56.250000  9.915000 74.700000  9.970000 ;
        RECT 56.250000  9.970000 74.700000 17.835000 ;
        RECT 56.250000 17.835000 74.700000 17.905000 ;
        RECT 62.325000 21.695000 74.700000 21.765000 ;
        RECT 62.395000 21.765000 74.700000 21.835000 ;
        RECT 62.465000 21.835000 74.700000 21.905000 ;
        RECT 62.535000 21.905000 74.700000 21.975000 ;
        RECT 62.605000 21.975000 74.700000 22.045000 ;
        RECT 62.675000 22.045000 74.700000 22.115000 ;
        RECT 62.745000 22.115000 74.700000 22.185000 ;
        RECT 62.815000 22.185000 74.700000 22.255000 ;
        RECT 62.885000 22.255000 74.700000 22.325000 ;
        RECT 62.955000 22.325000 74.700000 22.395000 ;
        RECT 63.025000 22.395000 74.700000 22.465000 ;
        RECT 63.095000 22.465000 74.700000 22.535000 ;
        RECT 63.165000 22.535000 74.700000 22.605000 ;
        RECT 63.235000 22.605000 74.700000 22.675000 ;
        RECT 63.305000 22.675000 74.700000 22.745000 ;
        RECT 63.375000 22.745000 74.700000 22.815000 ;
        RECT 63.445000 22.815000 74.700000 22.885000 ;
        RECT 63.515000 22.885000 74.700000 22.955000 ;
        RECT 63.585000 22.955000 74.700000 23.025000 ;
        RECT 63.655000 23.025000 74.700000 23.095000 ;
        RECT 63.725000 23.095000 74.700000 23.165000 ;
        RECT 63.795000 23.165000 74.700000 23.235000 ;
        RECT 63.865000 23.235000 74.700000 23.305000 ;
        RECT 63.935000 23.305000 74.700000 23.375000 ;
        RECT 64.005000 23.375000 74.700000 23.445000 ;
        RECT 64.075000 23.445000 74.700000 23.515000 ;
        RECT 64.145000 23.515000 74.700000 23.585000 ;
        RECT 64.215000 23.585000 74.700000 23.655000 ;
        RECT 64.285000 23.655000 74.700000 23.725000 ;
        RECT 64.355000 23.725000 74.700000 23.795000 ;
        RECT 64.425000 23.795000 74.700000 23.865000 ;
        RECT 64.495000 23.865000 74.700000 23.935000 ;
        RECT 64.565000 23.935000 74.700000 24.005000 ;
        RECT 64.635000 24.005000 74.700000 24.075000 ;
        RECT 64.705000 24.075000 74.700000 24.145000 ;
        RECT 64.775000 24.145000 74.700000 24.215000 ;
        RECT 64.845000 24.215000 74.700000 24.285000 ;
        RECT 64.880000 31.000000 74.700000 31.010000 ;
        RECT 64.915000 24.285000 74.700000 24.355000 ;
        RECT 64.950000 30.930000 74.700000 31.000000 ;
        RECT 64.950000 40.985000 74.700000 40.990000 ;
        RECT 64.950000 51.005000 74.700000 51.010000 ;
        RECT 64.985000 24.355000 74.700000 24.425000 ;
        RECT 65.015000 60.920000 74.700000 60.990000 ;
        RECT 65.015000 63.630000 74.700000 63.700000 ;
        RECT 65.015000 70.920000 74.700000 70.990000 ;
        RECT 65.020000 30.860000 74.700000 30.930000 ;
        RECT 65.020000 40.915000 74.700000 40.985000 ;
        RECT 65.020000 50.935000 74.700000 51.005000 ;
        RECT 65.030000 33.650000 74.700000 33.720000 ;
        RECT 65.030000 43.630000 74.700000 43.700000 ;
        RECT 65.030000 53.650000 74.700000 53.720000 ;
        RECT 65.055000 24.425000 74.700000 24.495000 ;
        RECT 65.085000 60.850000 74.700000 60.920000 ;
        RECT 65.085000 63.700000 74.700000 63.770000 ;
        RECT 65.085000 70.850000 74.700000 70.920000 ;
        RECT 65.090000 30.790000 74.700000 30.860000 ;
        RECT 65.090000 40.845000 74.700000 40.915000 ;
        RECT 65.090000 50.865000 74.700000 50.935000 ;
        RECT 65.100000 33.720000 74.700000 33.790000 ;
        RECT 65.100000 43.700000 74.700000 43.770000 ;
        RECT 65.100000 53.720000 74.700000 53.790000 ;
        RECT 65.125000 24.495000 74.700000 24.565000 ;
        RECT 65.155000 60.780000 74.700000 60.850000 ;
        RECT 65.155000 63.770000 74.700000 63.840000 ;
        RECT 65.155000 70.780000 74.700000 70.850000 ;
        RECT 65.160000 30.720000 74.700000 30.790000 ;
        RECT 65.160000 40.775000 74.700000 40.845000 ;
        RECT 65.160000 50.795000 74.700000 50.865000 ;
        RECT 65.170000 33.790000 74.700000 33.860000 ;
        RECT 65.170000 43.770000 74.700000 43.840000 ;
        RECT 65.170000 53.790000 74.700000 53.860000 ;
        RECT 65.195000 24.565000 74.700000 24.635000 ;
        RECT 65.225000 60.710000 74.700000 60.780000 ;
        RECT 65.225000 63.840000 74.700000 63.910000 ;
        RECT 65.225000 70.710000 74.700000 70.780000 ;
        RECT 65.230000 30.650000 74.700000 30.720000 ;
        RECT 65.230000 40.705000 74.700000 40.775000 ;
        RECT 65.230000 50.725000 74.700000 50.795000 ;
        RECT 65.240000 33.860000 74.700000 33.930000 ;
        RECT 65.240000 43.840000 74.700000 43.910000 ;
        RECT 65.240000 53.860000 74.700000 53.930000 ;
        RECT 65.265000 24.635000 74.700000 24.705000 ;
        RECT 65.270000 73.630000 68.740000 73.700000 ;
        RECT 65.295000 60.640000 74.700000 60.710000 ;
        RECT 65.295000 63.910000 74.700000 63.980000 ;
        RECT 65.295000 70.640000 74.700000 70.710000 ;
        RECT 65.300000 30.580000 74.700000 30.650000 ;
        RECT 65.300000 40.635000 74.700000 40.705000 ;
        RECT 65.300000 50.655000 74.700000 50.725000 ;
        RECT 65.310000 33.930000 74.700000 34.000000 ;
        RECT 65.310000 43.910000 74.700000 43.980000 ;
        RECT 65.310000 53.930000 74.700000 54.000000 ;
        RECT 65.335000 24.705000 74.700000 24.775000 ;
        RECT 65.340000 73.700000 68.670000 73.770000 ;
        RECT 65.365000 60.570000 74.700000 60.640000 ;
        RECT 65.365000 63.980000 74.700000 64.050000 ;
        RECT 65.365000 70.570000 74.700000 70.640000 ;
        RECT 65.370000 30.510000 74.700000 30.580000 ;
        RECT 65.370000 40.565000 74.700000 40.635000 ;
        RECT 65.370000 50.585000 74.700000 50.655000 ;
        RECT 65.380000 34.000000 74.700000 34.070000 ;
        RECT 65.380000 43.980000 74.700000 44.050000 ;
        RECT 65.380000 54.000000 74.700000 54.070000 ;
        RECT 65.405000 24.775000 74.700000 24.845000 ;
        RECT 65.410000 73.770000 68.600000 73.840000 ;
        RECT 65.435000 60.500000 74.700000 60.570000 ;
        RECT 65.435000 64.050000 74.700000 64.120000 ;
        RECT 65.435000 70.500000 74.700000 70.570000 ;
        RECT 65.440000 30.440000 74.700000 30.510000 ;
        RECT 65.440000 40.495000 74.700000 40.565000 ;
        RECT 65.440000 50.515000 74.700000 50.585000 ;
        RECT 65.450000 34.070000 74.700000 34.140000 ;
        RECT 65.450000 44.050000 74.700000 44.120000 ;
        RECT 65.450000 54.070000 74.700000 54.140000 ;
        RECT 65.475000 24.845000 74.700000 24.915000 ;
        RECT 65.480000 73.840000 68.530000 73.910000 ;
        RECT 65.505000 60.430000 74.700000 60.500000 ;
        RECT 65.505000 64.120000 74.700000 64.190000 ;
        RECT 65.505000 70.430000 74.700000 70.500000 ;
        RECT 65.510000 30.370000 74.700000 30.440000 ;
        RECT 65.510000 40.425000 74.700000 40.495000 ;
        RECT 65.510000 50.445000 74.700000 50.515000 ;
        RECT 65.520000 34.140000 74.700000 34.210000 ;
        RECT 65.520000 44.120000 74.700000 44.190000 ;
        RECT 65.520000 54.140000 74.700000 54.210000 ;
        RECT 65.545000 24.915000 74.700000 24.985000 ;
        RECT 65.550000 73.910000 68.460000 73.980000 ;
        RECT 65.575000 60.360000 74.700000 60.430000 ;
        RECT 65.575000 64.190000 74.700000 64.260000 ;
        RECT 65.575000 70.360000 74.700000 70.430000 ;
        RECT 65.580000 30.300000 74.700000 30.370000 ;
        RECT 65.580000 40.355000 74.700000 40.425000 ;
        RECT 65.580000 50.375000 74.700000 50.445000 ;
        RECT 65.590000 34.210000 74.700000 34.280000 ;
        RECT 65.590000 44.190000 74.700000 44.260000 ;
        RECT 65.590000 54.210000 74.700000 54.280000 ;
        RECT 65.615000 24.985000 74.700000 25.055000 ;
        RECT 65.620000 73.980000 68.390000 74.050000 ;
        RECT 65.645000 60.290000 74.700000 60.360000 ;
        RECT 65.645000 64.260000 74.700000 64.330000 ;
        RECT 65.645000 70.290000 74.700000 70.360000 ;
        RECT 65.650000 30.230000 74.700000 30.300000 ;
        RECT 65.650000 40.285000 74.700000 40.355000 ;
        RECT 65.650000 50.305000 74.700000 50.375000 ;
        RECT 65.660000 34.280000 74.700000 34.350000 ;
        RECT 65.660000 44.260000 74.700000 44.330000 ;
        RECT 65.660000 54.280000 74.700000 54.350000 ;
        RECT 65.685000 25.055000 74.700000 25.125000 ;
        RECT 65.690000 74.050000 68.320000 74.120000 ;
        RECT 65.715000 60.220000 74.700000 60.290000 ;
        RECT 65.715000 64.330000 74.700000 64.400000 ;
        RECT 65.715000 70.220000 74.700000 70.290000 ;
        RECT 65.720000 30.160000 74.700000 30.230000 ;
        RECT 65.720000 40.215000 74.700000 40.285000 ;
        RECT 65.720000 50.235000 74.700000 50.305000 ;
        RECT 65.730000 34.350000 74.700000 34.420000 ;
        RECT 65.730000 44.330000 74.700000 44.400000 ;
        RECT 65.730000 54.350000 74.700000 54.420000 ;
        RECT 65.755000 25.125000 74.700000 25.195000 ;
        RECT 65.760000 74.120000 68.250000 74.190000 ;
        RECT 65.785000 60.150000 74.700000 60.220000 ;
        RECT 65.785000 64.400000 74.700000 64.470000 ;
        RECT 65.785000 70.150000 74.700000 70.220000 ;
        RECT 65.790000 30.090000 74.700000 30.160000 ;
        RECT 65.790000 40.145000 74.700000 40.215000 ;
        RECT 65.790000 50.165000 74.700000 50.235000 ;
        RECT 65.800000 34.420000 74.700000 34.490000 ;
        RECT 65.800000 44.400000 74.700000 44.470000 ;
        RECT 65.800000 54.420000 74.700000 54.490000 ;
        RECT 65.825000 25.195000 74.700000 25.265000 ;
        RECT 65.830000 74.190000 68.180000 74.260000 ;
        RECT 65.855000 60.080000 74.700000 60.150000 ;
        RECT 65.855000 64.470000 74.700000 64.540000 ;
        RECT 65.855000 70.080000 74.700000 70.150000 ;
        RECT 65.860000 30.020000 74.700000 30.090000 ;
        RECT 65.860000 40.075000 74.700000 40.145000 ;
        RECT 65.860000 50.095000 74.700000 50.165000 ;
        RECT 65.870000 34.490000 74.700000 34.560000 ;
        RECT 65.870000 44.470000 74.700000 44.540000 ;
        RECT 65.870000 54.490000 74.700000 54.560000 ;
        RECT 65.895000 25.265000 74.700000 25.335000 ;
        RECT 65.900000 74.260000 68.110000 74.330000 ;
        RECT 65.925000 60.010000 74.700000 60.080000 ;
        RECT 65.925000 64.540000 74.700000 64.610000 ;
        RECT 65.925000 70.010000 74.700000 70.080000 ;
        RECT 65.930000 29.950000 74.700000 30.020000 ;
        RECT 65.930000 40.005000 74.700000 40.075000 ;
        RECT 65.930000 50.025000 74.700000 50.095000 ;
        RECT 65.940000 34.560000 74.700000 34.630000 ;
        RECT 65.940000 44.540000 74.700000 44.610000 ;
        RECT 65.940000 54.560000 74.700000 54.630000 ;
        RECT 65.965000 25.335000 74.700000 25.405000 ;
        RECT 65.970000 74.330000 68.040000 74.400000 ;
        RECT 65.995000 54.630000 74.700000 54.685000 ;
        RECT 65.995000 54.685000 74.700000 59.940000 ;
        RECT 65.995000 59.940000 74.700000 60.010000 ;
        RECT 65.995000 64.610000 74.700000 64.680000 ;
        RECT 65.995000 64.680000 74.700000 69.940000 ;
        RECT 65.995000 69.940000 74.700000 70.010000 ;
        RECT 66.000000 25.405000 74.700000 25.440000 ;
        RECT 66.000000 25.440000 74.700000 29.880000 ;
        RECT 66.000000 29.880000 74.700000 29.950000 ;
        RECT 66.000000 34.630000 74.700000 34.690000 ;
        RECT 66.000000 34.690000 74.700000 39.935000 ;
        RECT 66.000000 39.935000 74.700000 40.005000 ;
        RECT 66.000000 44.610000 74.700000 44.670000 ;
        RECT 66.000000 44.670000 74.700000 49.955000 ;
        RECT 66.000000 49.955000 74.700000 50.025000 ;
        RECT 66.000000 74.400000 68.010000 74.430000 ;
        RECT 66.000000 74.430000 68.010000 98.560000 ;
    END
  END SRC_BDY_LVC2
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 6.885000 1.270000 11.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 6.885000 75.000000 11.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 6.985000 1.270000 11.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 6.985000 75.000000 11.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 0.035000 1.270000 5.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 0.035000 75.000000 5.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 0.135000 1.270000 5.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 0.135000 75.000000 5.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 12.935000 0.965000 16.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035000 12.935000 75.000000 16.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 13.035000 0.965000 16.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 13.035000 75.000000 16.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 17.785000 1.270000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 68.035000 1.270000 93.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 17.785000 75.000000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 68.035000 75.000000 93.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 17.885000 1.270000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 68.035000 1.270000 92.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 17.885000 75.000000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 68.035000 75.000000 92.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 62.085000 1.270000 66.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 62.085000 75.000000 66.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 62.185000 1.270000 66.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 62.185000 75.000000 66.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 34.735000 1.270000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 45.735000 1.270000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 49.645000 1.270000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 54.405000 1.270000 54.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 34.735000 75.000000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 45.735000 75.000000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 49.645000 75.000000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 54.405000 75.000000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 34.840000 1.270000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 45.735000 1.270000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 34.840000 75.000000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 45.735000 75.000000 54.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 39.585000 1.270000 44.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 39.585000 75.000000 44.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 39.685000 1.270000 44.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 39.685000 75.000000 44.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 23.835000 1.270000 28.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 23.835000 75.000000 28.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 23.935000 1.270000 28.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 23.935000 75.000000 28.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 56.235000 1.270000 60.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 56.235000 75.000000 60.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 56.335000 1.270000 60.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 56.335000 75.000000 60.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 29.885000 1.270000 33.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 29.885000 75.000000 33.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 29.985000 1.270000 33.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 29.985000 75.000000 33.235000 ;
    END
  END VSWITCH
  OBS
    LAYER li1 ;
      RECT  0.240000  17.210000  2.995000  19.200000 ;
      RECT  1.350000   1.020000  7.110000   1.190000 ;
      RECT  1.350000   1.190000  1.520000  17.040000 ;
      RECT  1.350000  17.040000  7.110000  17.210000 ;
      RECT  1.760000  19.630000  9.385000  20.140000 ;
      RECT  1.760000  20.140000  2.685000  23.060000 ;
      RECT  1.845000   3.220000  2.015000   8.960000 ;
      RECT  1.845000   9.710000  2.015000  16.610000 ;
      RECT  2.070000   1.610000  6.390000   1.780000 ;
      RECT  2.070000   9.260000  6.390000   9.430000 ;
      RECT  2.305000   2.490000  2.475000   8.960000 ;
      RECT  2.305000  10.140000  2.475000  15.440000 ;
      RECT  2.765000   3.220000  2.935000   8.960000 ;
      RECT  2.765000   9.710000  2.935000  16.610000 ;
      RECT  3.225000   2.490000  3.395000   8.960000 ;
      RECT  3.225000  10.140000  3.395000  15.440000 ;
      RECT  3.685000   3.220000  3.855000   8.960000 ;
      RECT  3.685000   9.710000  3.855000  16.610000 ;
      RECT  4.145000   2.490000  4.315000   8.960000 ;
      RECT  4.145000  10.140000  4.315000  15.440000 ;
      RECT  4.605000   3.220000  4.775000   8.960000 ;
      RECT  4.605000   9.710000  4.775000  16.610000 ;
      RECT  4.975000  22.290000 10.650000  23.010000 ;
      RECT  5.065000   2.490000  5.235000   8.960000 ;
      RECT  5.065000  10.140000  5.235000  15.440000 ;
      RECT  5.525000   3.220000  5.695000   8.960000 ;
      RECT  5.525000   9.710000  5.695000  16.610000 ;
      RECT  5.890000  23.010000 10.650000  23.015000 ;
      RECT  5.985000   2.490000  6.155000   8.960000 ;
      RECT  5.985000  10.140000  6.155000  15.440000 ;
      RECT  6.445000   2.060000  6.615000   8.960000 ;
      RECT  6.445000   9.710000  6.615000  16.610000 ;
      RECT  6.940000   1.190000  7.110000  17.040000 ;
      RECT  8.340000 196.360000  8.670000 196.420000 ;
      RECT  8.345000   1.410000 16.655000  18.350000 ;
      RECT  8.420000 195.890000  8.590000 196.360000 ;
      RECT  9.155000 106.965000 10.280000 196.850000 ;
      RECT  9.155000 196.850000 69.720000 197.380000 ;
      RECT  9.185000  23.825000 69.720000  24.355000 ;
      RECT  9.185000  24.355000 10.280000  82.980000 ;
      RECT  9.185000  82.980000 21.740000  83.150000 ;
      RECT  9.185000  83.150000 10.280000  99.490000 ;
      RECT  9.730000  99.490000 10.280000 106.965000 ;
      RECT 10.920000  83.820000 11.830000  84.585000 ;
      RECT 11.065000 168.280000 12.220000 194.935000 ;
      RECT 11.065000 194.935000 68.495000 195.885000 ;
      RECT 11.095000 144.465000 21.490000 145.315000 ;
      RECT 11.095000 145.315000 12.220000 168.280000 ;
      RECT 11.275000  25.065000 68.140000  26.015000 ;
      RECT 11.275000  26.015000 12.220000  34.040000 ;
      RECT 11.275000  36.745000 12.220000  43.620000 ;
      RECT 11.275000  46.905000 12.220000  81.575000 ;
      RECT 11.275000  81.575000 23.280000  82.085000 ;
      RECT 11.370000  34.040000 12.220000  36.745000 ;
      RECT 11.370000  43.620000 12.220000  46.905000 ;
      RECT 12.405000 184.140000 66.575000 186.620000 ;
      RECT 12.430000 184.100000 66.575000 184.140000 ;
      RECT 12.750000  75.785000 12.920000  80.300000 ;
      RECT 12.975000  81.045000 66.655000  81.215000 ;
      RECT 13.060000  44.100000 65.590000  46.620000 ;
      RECT 13.060000  64.100000 65.590000  66.620000 ;
      RECT 13.190000  34.100000 65.590000  36.620000 ;
      RECT 13.190000  54.100000 65.590000  56.620000 ;
      RECT 13.335000 174.100000 65.590000 176.620000 ;
      RECT 13.365000 145.615000 14.305000 145.620000 ;
      RECT 13.365000 145.620000 65.590000 146.620000 ;
      RECT 13.365000 154.100000 65.590000 156.620000 ;
      RECT 13.365000 164.100000 65.590000 166.620000 ;
      RECT 13.395000  26.900000 13.925000  33.570000 ;
      RECT 13.395000  36.900000 13.925000  43.570000 ;
      RECT 13.395000  46.900000 13.925000  53.570000 ;
      RECT 13.395000  56.900000 13.925000  63.570000 ;
      RECT 13.395000  66.900000 13.925000  71.725000 ;
      RECT 13.395000 186.900000 13.925000 193.570000 ;
      RECT 14.360000 194.100000 65.590000 194.270000 ;
      RECT 14.780000  26.900000 15.310000  33.570000 ;
      RECT 14.780000  36.900000 15.310000  43.570000 ;
      RECT 14.780000  46.900000 15.310000  53.570000 ;
      RECT 14.780000  56.900000 15.310000  63.570000 ;
      RECT 14.780000  66.900000 15.310000  71.725000 ;
      RECT 14.780000 186.900000 15.310000 193.570000 ;
      RECT 14.790000  26.840000 15.300000  26.900000 ;
      RECT 14.790000  33.570000 15.300000  33.630000 ;
      RECT 14.790000  36.840000 15.300000  36.900000 ;
      RECT 14.790000  43.570000 15.300000  43.630000 ;
      RECT 14.790000  46.840000 15.300000  46.900000 ;
      RECT 14.790000  53.570000 15.300000  53.630000 ;
      RECT 14.790000  56.840000 15.300000  56.900000 ;
      RECT 14.790000  63.570000 15.300000  63.630000 ;
      RECT 14.790000  66.840000 15.300000  66.900000 ;
      RECT 14.790000 186.840000 15.300000 186.900000 ;
      RECT 14.790000 193.570000 15.300000 193.630000 ;
      RECT 15.865000 146.900000 16.395000 153.570000 ;
      RECT 15.865000 156.900000 16.395000 163.570000 ;
      RECT 15.865000 166.900000 16.395000 173.570000 ;
      RECT 16.165000  26.900000 16.695000  33.570000 ;
      RECT 16.165000  36.900000 16.695000  43.570000 ;
      RECT 16.165000  46.900000 16.695000  53.570000 ;
      RECT 16.165000  56.900000 16.695000  63.570000 ;
      RECT 16.165000  66.900000 16.695000  71.725000 ;
      RECT 16.165000 176.900000 16.695000 183.570000 ;
      RECT 16.165000 186.900000 16.695000 193.570000 ;
      RECT 17.000000  17.580000 56.200000  18.350000 ;
      RECT 17.030000  75.785000 17.200000  80.300000 ;
      RECT 17.550000  26.900000 18.080000  33.570000 ;
      RECT 17.550000  36.900000 18.080000  43.570000 ;
      RECT 17.550000  46.900000 18.080000  53.570000 ;
      RECT 17.550000  56.900000 18.080000  63.570000 ;
      RECT 17.550000  66.900000 18.080000  71.725000 ;
      RECT 17.550000 176.900000 18.080000 183.570000 ;
      RECT 17.550000 186.900000 18.080000 193.570000 ;
      RECT 17.560000  26.840000 18.070000  26.900000 ;
      RECT 17.560000  33.570000 18.070000  33.630000 ;
      RECT 17.560000  36.840000 18.070000  36.900000 ;
      RECT 17.560000  43.570000 18.070000  43.630000 ;
      RECT 17.560000  46.840000 18.070000  46.900000 ;
      RECT 17.560000  53.570000 18.070000  53.630000 ;
      RECT 17.560000  56.840000 18.070000  56.900000 ;
      RECT 17.560000  63.570000 18.070000  63.630000 ;
      RECT 17.560000  66.840000 18.070000  66.900000 ;
      RECT 17.560000 176.840000 18.070000 176.900000 ;
      RECT 17.560000 183.570000 18.070000 183.630000 ;
      RECT 17.560000 186.840000 18.070000 186.900000 ;
      RECT 17.560000 193.570000 18.070000 193.630000 ;
      RECT 17.955000 146.900000 18.485000 153.570000 ;
      RECT 17.955000 156.900000 18.485000 163.570000 ;
      RECT 17.955000 166.900000 18.485000 173.570000 ;
      RECT 17.965000 146.840000 18.475000 146.900000 ;
      RECT 17.965000 153.570000 18.475000 153.630000 ;
      RECT 17.965000 156.840000 18.475000 156.900000 ;
      RECT 17.965000 163.570000 18.475000 163.630000 ;
      RECT 17.965000 166.840000 18.475000 166.900000 ;
      RECT 17.965000 173.570000 18.475000 173.630000 ;
      RECT 18.935000  26.900000 19.465000  33.570000 ;
      RECT 18.935000  36.900000 19.465000  43.570000 ;
      RECT 18.935000  46.900000 19.465000  53.570000 ;
      RECT 18.935000  56.900000 19.465000  63.570000 ;
      RECT 18.935000  66.900000 19.465000  71.725000 ;
      RECT 18.935000 176.900000 19.465000 183.570000 ;
      RECT 18.935000 186.900000 19.465000 193.570000 ;
      RECT 19.495000  83.820000 20.405000  84.585000 ;
      RECT 20.045000 146.900000 20.575000 153.570000 ;
      RECT 20.045000 156.900000 20.575000 163.570000 ;
      RECT 20.045000 166.900000 20.575000 173.570000 ;
      RECT 20.320000  26.900000 20.850000  33.570000 ;
      RECT 20.320000  36.900000 20.850000  43.570000 ;
      RECT 20.320000  46.900000 20.850000  53.570000 ;
      RECT 20.320000  56.900000 20.850000  63.570000 ;
      RECT 20.320000  66.900000 20.850000  71.725000 ;
      RECT 20.320000 176.900000 20.850000 183.570000 ;
      RECT 20.320000 186.900000 20.850000 193.570000 ;
      RECT 20.330000  26.840000 20.840000  26.900000 ;
      RECT 20.330000  33.570000 20.840000  33.630000 ;
      RECT 20.330000  36.840000 20.840000  36.900000 ;
      RECT 20.330000  43.570000 20.840000  43.630000 ;
      RECT 20.330000  46.840000 20.840000  46.900000 ;
      RECT 20.330000  53.570000 20.840000  53.630000 ;
      RECT 20.330000  56.840000 20.840000  56.900000 ;
      RECT 20.330000  63.570000 20.840000  63.630000 ;
      RECT 20.330000  66.840000 20.840000  66.900000 ;
      RECT 20.330000 176.840000 20.840000 176.900000 ;
      RECT 20.330000 183.570000 20.840000 183.630000 ;
      RECT 20.330000 186.840000 20.840000 186.900000 ;
      RECT 20.330000 193.570000 20.840000 193.630000 ;
      RECT 20.640000 100.865000 68.495000 101.035000 ;
      RECT 20.640000 101.035000 21.490000 109.275000 ;
      RECT 20.640000 109.275000 68.495000 109.445000 ;
      RECT 20.640000 109.445000 21.490000 117.770000 ;
      RECT 20.640000 117.770000 68.495000 117.940000 ;
      RECT 20.640000 117.940000 21.490000 144.465000 ;
      RECT 21.570000  83.150000 21.740000  99.925000 ;
      RECT 21.570000  99.925000 69.720000 100.095000 ;
      RECT 21.660000 128.010000 65.590000 128.515000 ;
      RECT 21.690000 134.100000 65.590000 136.620000 ;
      RECT 21.705000  26.900000 22.235000  33.570000 ;
      RECT 21.705000  36.900000 22.235000  43.570000 ;
      RECT 21.705000  46.900000 22.235000  53.570000 ;
      RECT 21.705000  56.900000 22.235000  63.570000 ;
      RECT 21.705000  66.900000 22.235000  71.725000 ;
      RECT 21.705000 176.900000 22.235000 183.570000 ;
      RECT 21.705000 186.900000 22.235000 193.570000 ;
      RECT 22.135000 146.900000 22.665000 153.570000 ;
      RECT 22.135000 156.900000 22.665000 163.570000 ;
      RECT 22.135000 166.900000 22.665000 173.570000 ;
      RECT 22.145000 146.840000 22.655000 146.900000 ;
      RECT 22.145000 153.570000 22.655000 153.630000 ;
      RECT 22.145000 156.840000 22.655000 156.900000 ;
      RECT 22.145000 163.570000 22.655000 163.630000 ;
      RECT 22.145000 166.840000 22.655000 166.900000 ;
      RECT 22.145000 173.570000 22.655000 173.630000 ;
      RECT 22.430000  82.085000 23.280000  82.180000 ;
      RECT 22.430000  82.180000 68.140000  82.350000 ;
      RECT 22.430000  82.350000 23.280000  90.675000 ;
      RECT 22.430000  90.675000 68.140000  90.845000 ;
      RECT 22.430000  90.845000 23.280000  97.890000 ;
      RECT 22.770000  97.890000 23.280000  98.990000 ;
      RECT 22.770000  98.990000 68.140000  99.160000 ;
      RECT 23.090000  26.900000 23.620000  33.570000 ;
      RECT 23.090000  36.900000 23.620000  43.570000 ;
      RECT 23.090000  46.900000 23.620000  53.570000 ;
      RECT 23.090000  56.900000 23.620000  63.570000 ;
      RECT 23.090000  66.900000 23.620000  71.725000 ;
      RECT 23.090000 176.900000 23.620000 183.570000 ;
      RECT 23.090000 186.900000 23.620000 193.570000 ;
      RECT 23.100000  26.840000 23.610000  26.900000 ;
      RECT 23.100000  33.570000 23.610000  33.630000 ;
      RECT 23.100000  36.840000 23.610000  36.900000 ;
      RECT 23.100000  43.570000 23.610000  43.630000 ;
      RECT 23.100000  46.840000 23.610000  46.900000 ;
      RECT 23.100000  53.570000 23.610000  53.630000 ;
      RECT 23.100000  56.840000 23.610000  56.900000 ;
      RECT 23.100000  63.570000 23.610000  63.630000 ;
      RECT 23.100000  66.840000 23.610000  66.900000 ;
      RECT 23.100000 176.840000 23.610000 176.900000 ;
      RECT 23.100000 183.570000 23.610000 183.630000 ;
      RECT 23.100000 186.840000 23.610000 186.900000 ;
      RECT 23.100000 193.570000 23.610000 193.630000 ;
      RECT 23.405000 144.100000 65.590000 145.620000 ;
      RECT 23.635000 101.385000 24.045000 108.175000 ;
      RECT 23.635000 109.880000 24.045000 115.550000 ;
      RECT 23.635000 120.080000 24.045000 125.295000 ;
      RECT 23.685000  82.785000 24.215000  89.575000 ;
      RECT 23.685000  91.280000 24.215000  98.070000 ;
      RECT 23.805000 115.550000 24.045000 116.670000 ;
      RECT 23.805000 118.955000 24.045000 120.080000 ;
      RECT 23.805000 125.295000 24.045000 125.745000 ;
      RECT 24.225000 128.730000 24.755000 133.760000 ;
      RECT 24.225000 136.900000 24.755000 143.570000 ;
      RECT 24.225000 146.900000 24.755000 153.570000 ;
      RECT 24.225000 156.900000 24.755000 163.570000 ;
      RECT 24.225000 166.900000 24.755000 173.570000 ;
      RECT 24.475000  26.900000 25.005000  33.570000 ;
      RECT 24.475000  36.900000 25.005000  43.570000 ;
      RECT 24.475000  46.900000 25.005000  53.570000 ;
      RECT 24.475000  56.900000 25.005000  63.570000 ;
      RECT 24.475000  66.900000 25.005000  71.725000 ;
      RECT 24.475000 176.900000 25.005000 183.570000 ;
      RECT 24.475000 186.900000 25.005000 193.570000 ;
      RECT 24.615000  90.045000 66.655000  90.215000 ;
      RECT 24.615000  98.540000 66.655000  98.710000 ;
      RECT 24.670000 108.645000 66.655000 108.815000 ;
      RECT 24.670000 117.140000 66.655000 117.310000 ;
      RECT 24.670000 118.315000 66.655000 118.485000 ;
      RECT 25.310000  75.785000 25.480000  80.300000 ;
      RECT 25.310000  82.915000 25.480000  89.020000 ;
      RECT 25.310000  91.930000 25.480000  96.925000 ;
      RECT 25.365000 101.385000 25.535000 106.255000 ;
      RECT 25.365000 110.450000 25.535000 115.330000 ;
      RECT 25.365000 120.080000 25.535000 124.860000 ;
      RECT 25.860000  26.900000 26.390000  33.570000 ;
      RECT 25.860000  36.900000 26.390000  43.570000 ;
      RECT 25.860000  46.900000 26.390000  53.570000 ;
      RECT 25.860000  56.900000 26.390000  63.570000 ;
      RECT 25.860000  66.900000 26.390000  71.725000 ;
      RECT 25.860000 176.900000 26.390000 183.570000 ;
      RECT 25.860000 186.900000 26.390000 193.570000 ;
      RECT 25.870000  26.840000 26.380000  26.900000 ;
      RECT 25.870000  33.570000 26.380000  33.630000 ;
      RECT 25.870000  36.840000 26.380000  36.900000 ;
      RECT 25.870000  43.570000 26.380000  43.630000 ;
      RECT 25.870000  46.840000 26.380000  46.900000 ;
      RECT 25.870000  53.570000 26.380000  53.630000 ;
      RECT 25.870000  56.840000 26.380000  56.900000 ;
      RECT 25.870000  63.570000 26.380000  63.630000 ;
      RECT 25.870000  66.840000 26.380000  66.900000 ;
      RECT 25.870000 176.840000 26.380000 176.900000 ;
      RECT 25.870000 183.570000 26.380000 183.630000 ;
      RECT 25.870000 186.840000 26.380000 186.900000 ;
      RECT 25.870000 193.570000 26.380000 193.630000 ;
      RECT 26.315000 128.730000 26.845000 133.715000 ;
      RECT 26.315000 136.900000 26.845000 143.570000 ;
      RECT 26.315000 146.900000 26.845000 153.570000 ;
      RECT 26.315000 156.900000 26.845000 163.570000 ;
      RECT 26.315000 166.900000 26.845000 173.570000 ;
      RECT 26.325000 136.840000 26.835000 136.900000 ;
      RECT 26.325000 143.570000 26.835000 143.630000 ;
      RECT 26.325000 146.840000 26.835000 146.900000 ;
      RECT 26.325000 153.570000 26.835000 153.630000 ;
      RECT 26.325000 156.840000 26.835000 156.900000 ;
      RECT 26.325000 163.570000 26.835000 163.630000 ;
      RECT 26.325000 166.840000 26.835000 166.900000 ;
      RECT 26.325000 173.570000 26.835000 173.630000 ;
      RECT 27.245000  26.900000 27.775000  33.570000 ;
      RECT 27.245000  36.900000 27.775000  43.570000 ;
      RECT 27.245000  46.900000 27.775000  53.570000 ;
      RECT 27.245000  56.900000 27.775000  63.570000 ;
      RECT 27.245000  66.900000 27.775000  71.725000 ;
      RECT 27.245000 176.900000 27.775000 183.570000 ;
      RECT 27.245000 186.900000 27.775000 193.570000 ;
      RECT 28.405000 128.860000 28.935000 133.760000 ;
      RECT 28.405000 136.900000 28.935000 143.570000 ;
      RECT 28.405000 146.900000 28.935000 153.570000 ;
      RECT 28.405000 156.900000 28.935000 163.570000 ;
      RECT 28.405000 166.900000 28.935000 173.570000 ;
      RECT 28.630000  26.900000 29.160000  33.570000 ;
      RECT 28.630000  36.900000 29.160000  43.570000 ;
      RECT 28.630000  46.900000 29.160000  53.570000 ;
      RECT 28.630000  56.900000 29.160000  63.570000 ;
      RECT 28.630000  66.900000 29.160000  71.725000 ;
      RECT 28.630000 176.900000 29.160000 183.570000 ;
      RECT 28.630000 186.900000 29.160000 193.570000 ;
      RECT 28.640000  26.840000 29.150000  26.900000 ;
      RECT 28.640000  33.570000 29.150000  33.630000 ;
      RECT 28.640000  36.840000 29.150000  36.900000 ;
      RECT 28.640000  43.570000 29.150000  43.630000 ;
      RECT 28.640000  46.840000 29.150000  46.900000 ;
      RECT 28.640000  53.570000 29.150000  53.630000 ;
      RECT 28.640000  56.840000 29.150000  56.900000 ;
      RECT 28.640000  63.570000 29.150000  63.630000 ;
      RECT 28.640000  66.840000 29.150000  66.900000 ;
      RECT 28.640000 176.840000 29.150000 176.900000 ;
      RECT 28.640000 183.570000 29.150000 183.630000 ;
      RECT 28.640000 186.840000 29.150000 186.900000 ;
      RECT 28.640000 193.570000 29.150000 193.630000 ;
      RECT 30.015000  26.900000 30.545000  33.570000 ;
      RECT 30.015000  36.900000 30.545000  43.570000 ;
      RECT 30.015000  46.900000 30.545000  53.570000 ;
      RECT 30.015000  56.900000 30.545000  63.570000 ;
      RECT 30.015000  66.900000 30.545000  71.725000 ;
      RECT 30.015000 176.900000 30.545000 183.570000 ;
      RECT 30.015000 186.900000 30.545000 193.570000 ;
      RECT 30.495000 128.730000 31.025000 133.715000 ;
      RECT 30.495000 136.900000 31.025000 143.570000 ;
      RECT 30.495000 146.900000 31.025000 153.570000 ;
      RECT 30.495000 156.900000 31.025000 163.570000 ;
      RECT 30.495000 166.900000 31.025000 173.570000 ;
      RECT 30.505000 136.840000 31.015000 136.900000 ;
      RECT 30.505000 143.570000 31.015000 143.630000 ;
      RECT 30.505000 146.840000 31.015000 146.900000 ;
      RECT 30.505000 153.570000 31.015000 153.630000 ;
      RECT 30.505000 156.840000 31.015000 156.900000 ;
      RECT 30.505000 163.570000 31.015000 163.630000 ;
      RECT 30.505000 166.840000 31.015000 166.900000 ;
      RECT 30.505000 173.570000 31.015000 173.630000 ;
      RECT 31.400000  26.900000 31.930000  33.570000 ;
      RECT 31.400000  36.900000 31.930000  43.570000 ;
      RECT 31.400000  46.900000 31.930000  53.570000 ;
      RECT 31.400000  56.900000 31.930000  63.570000 ;
      RECT 31.400000  66.900000 31.930000  71.725000 ;
      RECT 31.400000 176.900000 31.930000 183.570000 ;
      RECT 31.400000 186.900000 31.930000 193.570000 ;
      RECT 31.410000  26.840000 31.920000  26.900000 ;
      RECT 31.410000  33.570000 31.920000  33.630000 ;
      RECT 31.410000  36.840000 31.920000  36.900000 ;
      RECT 31.410000  43.570000 31.920000  43.630000 ;
      RECT 31.410000  46.840000 31.920000  46.900000 ;
      RECT 31.410000  53.570000 31.920000  53.630000 ;
      RECT 31.410000  56.840000 31.920000  56.900000 ;
      RECT 31.410000  63.570000 31.920000  63.630000 ;
      RECT 31.410000  66.840000 31.920000  66.900000 ;
      RECT 31.410000 176.840000 31.920000 176.900000 ;
      RECT 31.410000 183.570000 31.920000 183.630000 ;
      RECT 31.410000 186.840000 31.920000 186.900000 ;
      RECT 31.410000 193.570000 31.920000 193.630000 ;
      RECT 32.585000 128.730000 33.115000 133.755000 ;
      RECT 32.585000 136.900000 33.115000 143.570000 ;
      RECT 32.585000 146.900000 33.115000 153.570000 ;
      RECT 32.585000 156.900000 33.115000 163.570000 ;
      RECT 32.585000 166.900000 33.115000 173.570000 ;
      RECT 32.785000  26.900000 33.315000  33.570000 ;
      RECT 32.785000  36.900000 33.315000  43.570000 ;
      RECT 32.785000  46.900000 33.315000  53.570000 ;
      RECT 32.785000  56.900000 33.315000  63.570000 ;
      RECT 32.785000  66.900000 33.315000  71.725000 ;
      RECT 32.785000 176.900000 33.315000 183.570000 ;
      RECT 32.785000 186.900000 33.315000 193.570000 ;
      RECT 33.590000  75.785000 33.760000  80.300000 ;
      RECT 33.590000  82.915000 33.760000  89.020000 ;
      RECT 33.590000  91.930000 33.760000  96.925000 ;
      RECT 33.590000 101.385000 33.760000 106.255000 ;
      RECT 33.590000 110.450000 33.760000 115.270000 ;
      RECT 33.595000 120.080000 33.765000 124.860000 ;
      RECT 34.170000  26.900000 34.700000  33.570000 ;
      RECT 34.170000  36.900000 34.700000  43.570000 ;
      RECT 34.170000  46.900000 34.700000  53.570000 ;
      RECT 34.170000  56.900000 34.700000  63.570000 ;
      RECT 34.170000  66.900000 34.700000  71.725000 ;
      RECT 34.170000 176.900000 34.700000 183.570000 ;
      RECT 34.170000 186.900000 34.700000 193.570000 ;
      RECT 34.180000  26.840000 34.690000  26.900000 ;
      RECT 34.180000  33.570000 34.690000  33.630000 ;
      RECT 34.180000  36.840000 34.690000  36.900000 ;
      RECT 34.180000  43.570000 34.690000  43.630000 ;
      RECT 34.180000  46.840000 34.690000  46.900000 ;
      RECT 34.180000  53.570000 34.690000  53.630000 ;
      RECT 34.180000  56.840000 34.690000  56.900000 ;
      RECT 34.180000  63.570000 34.690000  63.630000 ;
      RECT 34.180000  66.840000 34.690000  66.900000 ;
      RECT 34.180000 176.840000 34.690000 176.900000 ;
      RECT 34.180000 183.570000 34.690000 183.630000 ;
      RECT 34.180000 186.840000 34.690000 186.900000 ;
      RECT 34.180000 193.570000 34.690000 193.630000 ;
      RECT 34.675000 128.730000 35.205000 133.840000 ;
      RECT 34.675000 136.900000 35.205000 143.570000 ;
      RECT 34.675000 146.900000 35.205000 153.570000 ;
      RECT 34.675000 156.900000 35.205000 163.570000 ;
      RECT 34.675000 166.900000 35.205000 173.570000 ;
      RECT 34.685000 136.840000 35.195000 136.900000 ;
      RECT 34.685000 143.570000 35.195000 143.630000 ;
      RECT 34.685000 146.840000 35.195000 146.900000 ;
      RECT 34.685000 153.570000 35.195000 153.630000 ;
      RECT 34.685000 156.840000 35.195000 156.900000 ;
      RECT 34.685000 163.570000 35.195000 163.630000 ;
      RECT 34.685000 166.840000 35.195000 166.900000 ;
      RECT 34.685000 173.570000 35.195000 173.630000 ;
      RECT 35.555000  26.900000 36.085000  33.570000 ;
      RECT 35.555000  36.900000 36.085000  43.570000 ;
      RECT 35.555000  46.900000 36.085000  53.570000 ;
      RECT 35.555000  56.900000 36.085000  63.570000 ;
      RECT 35.555000  66.900000 36.085000  71.725000 ;
      RECT 35.555000 176.900000 36.085000 183.570000 ;
      RECT 35.555000 186.900000 36.085000 193.570000 ;
      RECT 36.765000 128.730000 37.295000 133.755000 ;
      RECT 36.765000 136.900000 37.295000 143.570000 ;
      RECT 36.765000 146.900000 37.295000 153.570000 ;
      RECT 36.765000 156.900000 37.295000 163.570000 ;
      RECT 36.765000 166.900000 37.295000 173.570000 ;
      RECT 36.940000  26.900000 37.470000  33.570000 ;
      RECT 36.940000  36.900000 37.470000  43.570000 ;
      RECT 36.940000  46.900000 37.470000  53.570000 ;
      RECT 36.940000  56.900000 37.470000  63.570000 ;
      RECT 36.940000  66.900000 37.470000  71.725000 ;
      RECT 36.940000 176.900000 37.470000 183.570000 ;
      RECT 36.940000 186.900000 37.470000 193.570000 ;
      RECT 36.950000  26.840000 37.460000  26.900000 ;
      RECT 36.950000  33.570000 37.460000  33.630000 ;
      RECT 36.950000  36.840000 37.460000  36.900000 ;
      RECT 36.950000  43.570000 37.460000  43.630000 ;
      RECT 36.950000  46.840000 37.460000  46.900000 ;
      RECT 36.950000  53.570000 37.460000  53.630000 ;
      RECT 36.950000  56.840000 37.460000  56.900000 ;
      RECT 36.950000  63.570000 37.460000  63.630000 ;
      RECT 36.950000  66.840000 37.460000  66.900000 ;
      RECT 36.950000 176.840000 37.460000 176.900000 ;
      RECT 36.950000 183.570000 37.460000 183.630000 ;
      RECT 36.950000 186.840000 37.460000 186.900000 ;
      RECT 36.950000 193.570000 37.460000 193.630000 ;
      RECT 38.325000  26.900000 38.855000  33.570000 ;
      RECT 38.325000  36.900000 38.855000  43.570000 ;
      RECT 38.325000  46.900000 38.855000  53.570000 ;
      RECT 38.325000  56.900000 38.855000  63.570000 ;
      RECT 38.325000  66.900000 38.855000  71.725000 ;
      RECT 38.325000 176.900000 38.855000 183.570000 ;
      RECT 38.325000 186.900000 38.855000 193.570000 ;
      RECT 38.855000 128.730000 39.385000 133.925000 ;
      RECT 38.855000 136.900000 39.385000 143.570000 ;
      RECT 38.855000 146.900000 39.385000 153.570000 ;
      RECT 38.855000 156.900000 39.385000 163.570000 ;
      RECT 38.855000 166.900000 39.385000 173.570000 ;
      RECT 38.865000 136.840000 39.375000 136.900000 ;
      RECT 38.865000 143.570000 39.375000 143.630000 ;
      RECT 38.865000 146.840000 39.375000 146.900000 ;
      RECT 38.865000 153.570000 39.375000 153.630000 ;
      RECT 38.865000 156.840000 39.375000 156.900000 ;
      RECT 38.865000 163.570000 39.375000 163.630000 ;
      RECT 38.865000 166.840000 39.375000 166.900000 ;
      RECT 38.865000 173.570000 39.375000 173.630000 ;
      RECT 39.710000  26.900000 40.240000  33.570000 ;
      RECT 39.710000  36.900000 40.240000  43.570000 ;
      RECT 39.710000  46.900000 40.240000  53.570000 ;
      RECT 39.710000  56.900000 40.240000  63.570000 ;
      RECT 39.710000  66.900000 40.240000  71.725000 ;
      RECT 39.710000 176.900000 40.240000 183.570000 ;
      RECT 39.710000 186.900000 40.240000 193.570000 ;
      RECT 39.720000  26.840000 40.230000  26.900000 ;
      RECT 39.720000  33.570000 40.230000  33.630000 ;
      RECT 39.720000  36.840000 40.230000  36.900000 ;
      RECT 39.720000  43.570000 40.230000  43.630000 ;
      RECT 39.720000  46.840000 40.230000  46.900000 ;
      RECT 39.720000  53.570000 40.230000  53.630000 ;
      RECT 39.720000  56.840000 40.230000  56.900000 ;
      RECT 39.720000  63.570000 40.230000  63.630000 ;
      RECT 39.720000  66.840000 40.230000  66.900000 ;
      RECT 39.720000 176.840000 40.230000 176.900000 ;
      RECT 39.720000 183.570000 40.230000 183.630000 ;
      RECT 39.720000 186.840000 40.230000 186.900000 ;
      RECT 39.720000 193.570000 40.230000 193.630000 ;
      RECT 40.945000 128.730000 41.475000 133.755000 ;
      RECT 40.945000 136.900000 41.475000 143.570000 ;
      RECT 40.945000 146.900000 41.475000 153.570000 ;
      RECT 40.945000 156.900000 41.475000 163.570000 ;
      RECT 40.945000 166.900000 41.475000 173.570000 ;
      RECT 41.095000  26.900000 41.625000  33.570000 ;
      RECT 41.095000  36.900000 41.625000  43.570000 ;
      RECT 41.095000  46.900000 41.625000  53.570000 ;
      RECT 41.095000  56.900000 41.625000  63.570000 ;
      RECT 41.095000  66.900000 41.625000  71.725000 ;
      RECT 41.095000 176.900000 41.625000 183.570000 ;
      RECT 41.095000 186.900000 41.625000 193.570000 ;
      RECT 41.870000  75.785000 42.040000  80.300000 ;
      RECT 41.870000  82.915000 42.040000  89.020000 ;
      RECT 41.870000  91.930000 42.040000  96.925000 ;
      RECT 41.870000 101.385000 42.040000 106.255000 ;
      RECT 41.870000 110.450000 42.040000 115.270000 ;
      RECT 41.870000 120.080000 42.040000 124.860000 ;
      RECT 42.480000  26.900000 43.010000  33.570000 ;
      RECT 42.480000  36.900000 43.010000  43.570000 ;
      RECT 42.480000  46.900000 43.010000  53.570000 ;
      RECT 42.480000  56.900000 43.010000  63.570000 ;
      RECT 42.480000  66.900000 43.010000  71.725000 ;
      RECT 42.480000 176.900000 43.010000 183.570000 ;
      RECT 42.480000 186.900000 43.010000 193.570000 ;
      RECT 42.490000  26.840000 43.000000  26.900000 ;
      RECT 42.490000  33.570000 43.000000  33.630000 ;
      RECT 42.490000  36.840000 43.000000  36.900000 ;
      RECT 42.490000  43.570000 43.000000  43.630000 ;
      RECT 42.490000  46.840000 43.000000  46.900000 ;
      RECT 42.490000  53.570000 43.000000  53.630000 ;
      RECT 42.490000  56.840000 43.000000  56.900000 ;
      RECT 42.490000  63.570000 43.000000  63.630000 ;
      RECT 42.490000  66.840000 43.000000  66.900000 ;
      RECT 42.490000 176.840000 43.000000 176.900000 ;
      RECT 42.490000 183.570000 43.000000 183.630000 ;
      RECT 42.490000 186.840000 43.000000 186.900000 ;
      RECT 42.490000 193.570000 43.000000 193.630000 ;
      RECT 43.035000 128.730000 43.565000 133.925000 ;
      RECT 43.035000 136.900000 43.565000 143.570000 ;
      RECT 43.035000 146.900000 43.565000 153.570000 ;
      RECT 43.035000 156.900000 43.565000 163.570000 ;
      RECT 43.035000 166.900000 43.565000 173.570000 ;
      RECT 43.045000 136.840000 43.555000 136.900000 ;
      RECT 43.045000 143.570000 43.555000 143.630000 ;
      RECT 43.045000 146.840000 43.555000 146.900000 ;
      RECT 43.045000 153.570000 43.555000 153.630000 ;
      RECT 43.045000 156.840000 43.555000 156.900000 ;
      RECT 43.045000 163.570000 43.555000 163.630000 ;
      RECT 43.045000 166.840000 43.555000 166.900000 ;
      RECT 43.045000 173.570000 43.555000 173.630000 ;
      RECT 43.865000  26.900000 44.395000  33.570000 ;
      RECT 43.865000  36.900000 44.395000  43.570000 ;
      RECT 43.865000  46.900000 44.395000  53.570000 ;
      RECT 43.865000  56.900000 44.395000  63.570000 ;
      RECT 43.865000  66.900000 44.395000  71.725000 ;
      RECT 43.865000 176.900000 44.395000 183.570000 ;
      RECT 43.865000 186.900000 44.395000 193.570000 ;
      RECT 45.125000 128.730000 45.655000 133.755000 ;
      RECT 45.125000 136.900000 45.655000 143.570000 ;
      RECT 45.125000 146.900000 45.655000 153.570000 ;
      RECT 45.125000 156.900000 45.655000 163.570000 ;
      RECT 45.125000 166.900000 45.655000 173.570000 ;
      RECT 45.250000  26.900000 45.780000  33.570000 ;
      RECT 45.250000  36.900000 45.780000  43.570000 ;
      RECT 45.250000  46.900000 45.780000  53.570000 ;
      RECT 45.250000  56.900000 45.780000  63.570000 ;
      RECT 45.250000  66.900000 45.780000  71.725000 ;
      RECT 45.250000 176.900000 45.780000 183.570000 ;
      RECT 45.250000 186.900000 45.780000 193.570000 ;
      RECT 45.260000  26.840000 45.770000  26.900000 ;
      RECT 45.260000  33.570000 45.770000  33.630000 ;
      RECT 45.260000  36.840000 45.770000  36.900000 ;
      RECT 45.260000  43.570000 45.770000  43.630000 ;
      RECT 45.260000  46.840000 45.770000  46.900000 ;
      RECT 45.260000  53.570000 45.770000  53.630000 ;
      RECT 45.260000  56.840000 45.770000  56.900000 ;
      RECT 45.260000  63.570000 45.770000  63.630000 ;
      RECT 45.260000  66.840000 45.770000  66.900000 ;
      RECT 45.260000 176.840000 45.770000 176.900000 ;
      RECT 45.260000 183.570000 45.770000 183.630000 ;
      RECT 45.260000 186.840000 45.770000 186.900000 ;
      RECT 45.260000 193.570000 45.770000 193.630000 ;
      RECT 46.635000  26.900000 47.165000  33.570000 ;
      RECT 46.635000  36.900000 47.165000  43.570000 ;
      RECT 46.635000  46.900000 47.165000  53.570000 ;
      RECT 46.635000  56.900000 47.165000  63.570000 ;
      RECT 46.635000  66.900000 47.165000  71.725000 ;
      RECT 46.635000 176.900000 47.165000 183.570000 ;
      RECT 46.635000 186.900000 47.165000 193.570000 ;
      RECT 47.215000 128.730000 47.745000 133.925000 ;
      RECT 47.215000 136.900000 47.745000 143.570000 ;
      RECT 47.215000 146.900000 47.745000 153.570000 ;
      RECT 47.215000 156.900000 47.745000 163.570000 ;
      RECT 47.215000 166.900000 47.745000 173.570000 ;
      RECT 47.225000 136.840000 47.735000 136.900000 ;
      RECT 47.225000 143.570000 47.735000 143.630000 ;
      RECT 47.225000 146.840000 47.735000 146.900000 ;
      RECT 47.225000 153.570000 47.735000 153.630000 ;
      RECT 47.225000 156.840000 47.735000 156.900000 ;
      RECT 47.225000 163.570000 47.735000 163.630000 ;
      RECT 47.225000 166.840000 47.735000 166.900000 ;
      RECT 47.225000 173.570000 47.735000 173.630000 ;
      RECT 48.020000  26.900000 48.550000  33.570000 ;
      RECT 48.020000  36.900000 48.550000  43.570000 ;
      RECT 48.020000  46.900000 48.550000  53.570000 ;
      RECT 48.020000  56.900000 48.550000  63.570000 ;
      RECT 48.020000  66.900000 48.550000  71.725000 ;
      RECT 48.020000 176.900000 48.550000 183.570000 ;
      RECT 48.020000 186.900000 48.550000 193.570000 ;
      RECT 48.030000  26.840000 48.540000  26.900000 ;
      RECT 48.030000  33.570000 48.540000  33.630000 ;
      RECT 48.030000  36.840000 48.540000  36.900000 ;
      RECT 48.030000  43.570000 48.540000  43.630000 ;
      RECT 48.030000  46.840000 48.540000  46.900000 ;
      RECT 48.030000  53.570000 48.540000  53.630000 ;
      RECT 48.030000  56.840000 48.540000  56.900000 ;
      RECT 48.030000  63.570000 48.540000  63.630000 ;
      RECT 48.030000  66.840000 48.540000  66.900000 ;
      RECT 48.030000 176.840000 48.540000 176.900000 ;
      RECT 48.030000 183.570000 48.540000 183.630000 ;
      RECT 48.030000 186.840000 48.540000 186.900000 ;
      RECT 48.030000 193.570000 48.540000 193.630000 ;
      RECT 49.305000 128.730000 49.835000 133.755000 ;
      RECT 49.305000 136.900000 49.835000 143.570000 ;
      RECT 49.305000 146.900000 49.835000 153.570000 ;
      RECT 49.305000 156.900000 49.835000 163.570000 ;
      RECT 49.305000 166.900000 49.835000 173.570000 ;
      RECT 49.405000  26.900000 49.935000  33.570000 ;
      RECT 49.405000  36.900000 49.935000  43.570000 ;
      RECT 49.405000  46.900000 49.935000  53.570000 ;
      RECT 49.405000  56.900000 49.935000  63.570000 ;
      RECT 49.405000  66.900000 49.935000  71.725000 ;
      RECT 49.405000 176.900000 49.935000 183.570000 ;
      RECT 49.405000 186.900000 49.935000 193.570000 ;
      RECT 50.150000  75.785000 50.320000  80.300000 ;
      RECT 50.150000  82.915000 50.320000  89.020000 ;
      RECT 50.150000  91.930000 50.320000  96.925000 ;
      RECT 50.150000 101.385000 50.320000 106.255000 ;
      RECT 50.150000 110.450000 50.320000 115.270000 ;
      RECT 50.150000 120.080000 50.320000 124.860000 ;
      RECT 50.790000  26.900000 51.320000  33.570000 ;
      RECT 50.790000  36.900000 51.320000  43.570000 ;
      RECT 50.790000  46.900000 51.320000  53.570000 ;
      RECT 50.790000  56.900000 51.320000  63.570000 ;
      RECT 50.790000  66.900000 51.320000  71.725000 ;
      RECT 50.790000 176.900000 51.320000 183.570000 ;
      RECT 50.790000 186.900000 51.320000 193.570000 ;
      RECT 50.800000  26.840000 51.310000  26.900000 ;
      RECT 50.800000  33.570000 51.310000  33.630000 ;
      RECT 50.800000  36.840000 51.310000  36.900000 ;
      RECT 50.800000  43.570000 51.310000  43.630000 ;
      RECT 50.800000  46.840000 51.310000  46.900000 ;
      RECT 50.800000  53.570000 51.310000  53.630000 ;
      RECT 50.800000  56.840000 51.310000  56.900000 ;
      RECT 50.800000  63.570000 51.310000  63.630000 ;
      RECT 50.800000  66.840000 51.310000  66.900000 ;
      RECT 50.800000 176.840000 51.310000 176.900000 ;
      RECT 50.800000 183.570000 51.310000 183.630000 ;
      RECT 50.800000 186.840000 51.310000 186.900000 ;
      RECT 50.800000 193.570000 51.310000 193.630000 ;
      RECT 51.395000 128.730000 51.925000 133.925000 ;
      RECT 51.395000 136.900000 51.925000 143.570000 ;
      RECT 51.395000 146.900000 51.925000 153.570000 ;
      RECT 51.395000 156.900000 51.925000 163.570000 ;
      RECT 51.395000 166.900000 51.925000 173.570000 ;
      RECT 51.405000 136.840000 51.915000 136.900000 ;
      RECT 51.405000 143.570000 51.915000 143.630000 ;
      RECT 51.405000 146.840000 51.915000 146.900000 ;
      RECT 51.405000 153.570000 51.915000 153.630000 ;
      RECT 51.405000 156.840000 51.915000 156.900000 ;
      RECT 51.405000 163.570000 51.915000 163.630000 ;
      RECT 51.405000 166.840000 51.915000 166.900000 ;
      RECT 51.405000 173.570000 51.915000 173.630000 ;
      RECT 52.175000  26.900000 52.705000  33.570000 ;
      RECT 52.175000  36.900000 52.705000  43.570000 ;
      RECT 52.175000  46.900000 52.705000  53.570000 ;
      RECT 52.175000  56.900000 52.705000  63.570000 ;
      RECT 52.175000  66.900000 52.705000  71.725000 ;
      RECT 52.175000 176.900000 52.705000 183.570000 ;
      RECT 52.175000 186.900000 52.705000 193.570000 ;
      RECT 53.485000 128.730000 54.015000 133.755000 ;
      RECT 53.485000 136.900000 54.015000 143.570000 ;
      RECT 53.485000 146.900000 54.015000 153.570000 ;
      RECT 53.485000 156.900000 54.015000 163.570000 ;
      RECT 53.485000 166.900000 54.015000 173.570000 ;
      RECT 53.560000  26.900000 54.090000  33.570000 ;
      RECT 53.560000  36.900000 54.090000  43.570000 ;
      RECT 53.560000  46.900000 54.090000  53.570000 ;
      RECT 53.560000  56.900000 54.090000  63.570000 ;
      RECT 53.560000  66.900000 54.090000  71.725000 ;
      RECT 53.560000 176.900000 54.090000 183.570000 ;
      RECT 53.560000 186.900000 54.090000 193.570000 ;
      RECT 53.570000  26.840000 54.080000  26.900000 ;
      RECT 53.570000  33.570000 54.080000  33.630000 ;
      RECT 53.570000  36.840000 54.080000  36.900000 ;
      RECT 53.570000  43.570000 54.080000  43.630000 ;
      RECT 53.570000  46.840000 54.080000  46.900000 ;
      RECT 53.570000  53.570000 54.080000  53.630000 ;
      RECT 53.570000  56.840000 54.080000  56.900000 ;
      RECT 53.570000  63.570000 54.080000  63.630000 ;
      RECT 53.570000  66.840000 54.080000  66.900000 ;
      RECT 53.570000 176.840000 54.080000 176.900000 ;
      RECT 53.570000 183.570000 54.080000 183.630000 ;
      RECT 53.570000 186.840000 54.080000 186.900000 ;
      RECT 53.570000 193.570000 54.080000 193.630000 ;
      RECT 54.945000  26.900000 55.475000  33.570000 ;
      RECT 54.945000  36.900000 55.475000  43.570000 ;
      RECT 54.945000  46.900000 55.475000  53.570000 ;
      RECT 54.945000  56.900000 55.475000  63.570000 ;
      RECT 54.945000  66.900000 55.475000  71.725000 ;
      RECT 54.945000 176.900000 55.475000 183.570000 ;
      RECT 54.945000 186.900000 55.475000 193.570000 ;
      RECT 55.575000 128.730000 56.105000 133.925000 ;
      RECT 55.575000 136.900000 56.105000 143.570000 ;
      RECT 55.575000 146.900000 56.105000 153.570000 ;
      RECT 55.575000 156.900000 56.105000 163.570000 ;
      RECT 55.575000 166.900000 56.105000 173.570000 ;
      RECT 55.585000 136.840000 56.095000 136.900000 ;
      RECT 55.585000 143.570000 56.095000 143.630000 ;
      RECT 55.585000 146.840000 56.095000 146.900000 ;
      RECT 55.585000 153.570000 56.095000 153.630000 ;
      RECT 55.585000 156.840000 56.095000 156.900000 ;
      RECT 55.585000 163.570000 56.095000 163.630000 ;
      RECT 55.585000 166.840000 56.095000 166.900000 ;
      RECT 55.585000 173.570000 56.095000 173.630000 ;
      RECT 56.330000  26.900000 56.860000  33.570000 ;
      RECT 56.330000  36.900000 56.860000  43.570000 ;
      RECT 56.330000  46.900000 56.860000  53.570000 ;
      RECT 56.330000  56.900000 56.860000  63.570000 ;
      RECT 56.330000  66.900000 56.860000  71.725000 ;
      RECT 56.330000 176.900000 56.860000 183.570000 ;
      RECT 56.330000 186.900000 56.860000 193.570000 ;
      RECT 56.340000  26.840000 56.850000  26.900000 ;
      RECT 56.340000  33.570000 56.850000  33.630000 ;
      RECT 56.340000  36.840000 56.850000  36.900000 ;
      RECT 56.340000  43.570000 56.850000  43.630000 ;
      RECT 56.340000  46.840000 56.850000  46.900000 ;
      RECT 56.340000  53.570000 56.850000  53.630000 ;
      RECT 56.340000  56.840000 56.850000  56.900000 ;
      RECT 56.340000  63.570000 56.850000  63.630000 ;
      RECT 56.340000  66.840000 56.850000  66.900000 ;
      RECT 56.340000 176.840000 56.850000 176.900000 ;
      RECT 56.340000 183.570000 56.850000 183.630000 ;
      RECT 56.340000 186.840000 56.850000 186.900000 ;
      RECT 56.340000 193.570000 56.850000 193.630000 ;
      RECT 56.980000  16.365000 57.510000  16.895000 ;
      RECT 57.665000 128.730000 58.195000 133.755000 ;
      RECT 57.665000 136.900000 58.195000 143.570000 ;
      RECT 57.665000 146.900000 58.195000 153.570000 ;
      RECT 57.665000 156.900000 58.195000 163.570000 ;
      RECT 57.665000 166.900000 58.195000 173.570000 ;
      RECT 57.715000  26.900000 58.245000  33.570000 ;
      RECT 57.715000  36.900000 58.245000  43.570000 ;
      RECT 57.715000  46.900000 58.245000  53.570000 ;
      RECT 57.715000  56.900000 58.245000  63.570000 ;
      RECT 57.715000  66.900000 58.245000  71.725000 ;
      RECT 57.715000 176.900000 58.245000 183.570000 ;
      RECT 57.715000 186.900000 58.245000 193.570000 ;
      RECT 58.430000  75.785000 58.600000  80.300000 ;
      RECT 58.430000  82.915000 58.600000  89.020000 ;
      RECT 58.430000  91.930000 58.600000  96.925000 ;
      RECT 58.430000 101.385000 58.600000 106.255000 ;
      RECT 58.430000 110.450000 58.600000 115.270000 ;
      RECT 58.430000 120.080000 58.600000 124.860000 ;
      RECT 59.100000  26.900000 59.630000  33.570000 ;
      RECT 59.100000  36.900000 59.630000  43.570000 ;
      RECT 59.100000  46.900000 59.630000  53.570000 ;
      RECT 59.100000  56.900000 59.630000  63.570000 ;
      RECT 59.100000  66.900000 59.630000  71.725000 ;
      RECT 59.100000 176.900000 59.630000 183.570000 ;
      RECT 59.100000 186.900000 59.630000 193.570000 ;
      RECT 59.110000  26.840000 59.620000  26.900000 ;
      RECT 59.110000  33.570000 59.620000  33.630000 ;
      RECT 59.110000  36.840000 59.620000  36.900000 ;
      RECT 59.110000  43.570000 59.620000  43.630000 ;
      RECT 59.110000  46.840000 59.620000  46.900000 ;
      RECT 59.110000  53.570000 59.620000  53.630000 ;
      RECT 59.110000  56.840000 59.620000  56.900000 ;
      RECT 59.110000  63.570000 59.620000  63.630000 ;
      RECT 59.110000  66.840000 59.620000  66.900000 ;
      RECT 59.110000 176.840000 59.620000 176.900000 ;
      RECT 59.110000 183.570000 59.620000 183.630000 ;
      RECT 59.110000 186.840000 59.620000 186.900000 ;
      RECT 59.110000 193.570000 59.620000 193.630000 ;
      RECT 59.755000 128.730000 60.285000 133.925000 ;
      RECT 59.755000 136.900000 60.285000 143.570000 ;
      RECT 59.755000 146.900000 60.285000 153.570000 ;
      RECT 59.755000 156.900000 60.285000 163.570000 ;
      RECT 59.755000 166.900000 60.285000 173.570000 ;
      RECT 59.765000 136.840000 60.275000 136.900000 ;
      RECT 59.765000 143.570000 60.275000 143.630000 ;
      RECT 59.765000 146.840000 60.275000 146.900000 ;
      RECT 59.765000 153.570000 60.275000 153.630000 ;
      RECT 59.765000 156.840000 60.275000 156.900000 ;
      RECT 59.765000 163.570000 60.275000 163.630000 ;
      RECT 59.765000 166.840000 60.275000 166.900000 ;
      RECT 59.765000 173.570000 60.275000 173.630000 ;
      RECT 60.485000  26.900000 61.015000  33.570000 ;
      RECT 60.485000  36.900000 61.015000  43.570000 ;
      RECT 60.485000  46.900000 61.015000  53.570000 ;
      RECT 60.485000  56.900000 61.015000  63.570000 ;
      RECT 60.485000  66.900000 61.015000  71.725000 ;
      RECT 60.485000 176.900000 61.015000 183.570000 ;
      RECT 60.485000 186.900000 61.015000 193.570000 ;
      RECT 61.845000 128.730000 62.375000 133.755000 ;
      RECT 61.845000 136.900000 62.375000 143.570000 ;
      RECT 61.845000 146.900000 62.375000 153.570000 ;
      RECT 61.845000 156.900000 62.375000 163.570000 ;
      RECT 61.845000 166.900000 62.375000 173.570000 ;
      RECT 61.870000  26.900000 62.400000  33.570000 ;
      RECT 61.870000  36.900000 62.400000  43.570000 ;
      RECT 61.870000  46.900000 62.400000  53.570000 ;
      RECT 61.870000  56.900000 62.400000  63.570000 ;
      RECT 61.870000  66.900000 62.400000  71.725000 ;
      RECT 61.870000 176.900000 62.400000 183.570000 ;
      RECT 61.870000 186.900000 62.400000 193.570000 ;
      RECT 61.880000  26.840000 62.390000  26.900000 ;
      RECT 61.880000  33.570000 62.390000  33.630000 ;
      RECT 61.880000  36.840000 62.390000  36.900000 ;
      RECT 61.880000  43.570000 62.390000  43.630000 ;
      RECT 61.880000  46.840000 62.390000  46.900000 ;
      RECT 61.880000  53.570000 62.390000  53.630000 ;
      RECT 61.880000  56.840000 62.390000  56.900000 ;
      RECT 61.880000  63.570000 62.390000  63.630000 ;
      RECT 61.880000  66.840000 62.390000  66.900000 ;
      RECT 61.880000 176.840000 62.390000 176.900000 ;
      RECT 61.880000 183.570000 62.390000 183.630000 ;
      RECT 61.880000 186.840000 62.390000 186.900000 ;
      RECT 61.880000 193.570000 62.390000 193.630000 ;
      RECT 63.255000  26.900000 63.785000  33.570000 ;
      RECT 63.255000  36.900000 63.785000  43.570000 ;
      RECT 63.255000  46.900000 63.785000  53.570000 ;
      RECT 63.255000  56.900000 63.785000  63.570000 ;
      RECT 63.255000  66.900000 63.785000  71.725000 ;
      RECT 63.255000 176.900000 63.785000 183.570000 ;
      RECT 63.255000 186.900000 63.785000 193.570000 ;
      RECT 63.935000 128.730000 64.465000 133.925000 ;
      RECT 63.935000 136.900000 64.465000 143.570000 ;
      RECT 63.935000 146.900000 64.465000 153.570000 ;
      RECT 63.935000 156.900000 64.465000 163.570000 ;
      RECT 63.935000 166.900000 64.465000 173.570000 ;
      RECT 63.945000 136.840000 64.455000 136.900000 ;
      RECT 63.945000 143.570000 64.455000 143.630000 ;
      RECT 63.945000 146.840000 64.455000 146.900000 ;
      RECT 63.945000 153.570000 64.455000 153.630000 ;
      RECT 63.945000 156.840000 64.455000 156.900000 ;
      RECT 63.945000 163.570000 64.455000 163.630000 ;
      RECT 63.945000 166.840000 64.455000 166.900000 ;
      RECT 63.945000 173.570000 64.455000 173.630000 ;
      RECT 64.640000  26.900000 65.170000  33.570000 ;
      RECT 64.640000  36.900000 65.170000  43.570000 ;
      RECT 64.640000  46.900000 65.170000  53.570000 ;
      RECT 64.640000  56.900000 65.170000  63.570000 ;
      RECT 64.640000  66.900000 65.170000  71.725000 ;
      RECT 64.640000 176.900000 65.170000 183.570000 ;
      RECT 64.640000 186.900000 65.170000 193.570000 ;
      RECT 64.650000  26.840000 65.160000  26.900000 ;
      RECT 64.650000  33.570000 65.160000  33.630000 ;
      RECT 64.650000  36.840000 65.160000  36.900000 ;
      RECT 64.650000  43.570000 65.160000  43.630000 ;
      RECT 64.650000  46.840000 65.160000  46.900000 ;
      RECT 64.650000  53.570000 65.160000  53.630000 ;
      RECT 64.650000  56.840000 65.160000  56.900000 ;
      RECT 64.650000  63.570000 65.160000  63.630000 ;
      RECT 64.650000  66.840000 65.160000  66.900000 ;
      RECT 64.650000 176.840000 65.160000 176.900000 ;
      RECT 64.650000 183.570000 65.160000 183.630000 ;
      RECT 64.650000 186.840000 65.160000 186.900000 ;
      RECT 64.650000 193.570000 65.160000 193.630000 ;
      RECT 66.025000  26.900000 66.555000  33.570000 ;
      RECT 66.025000  36.900000 66.555000  43.570000 ;
      RECT 66.025000  46.900000 66.555000  53.570000 ;
      RECT 66.025000  56.900000 66.555000  63.570000 ;
      RECT 66.025000  66.900000 66.555000  71.725000 ;
      RECT 66.025000 128.730000 66.555000 133.755000 ;
      RECT 66.025000 136.900000 66.555000 143.570000 ;
      RECT 66.025000 146.900000 66.555000 153.570000 ;
      RECT 66.025000 156.900000 66.555000 163.570000 ;
      RECT 66.025000 166.900000 66.555000 173.570000 ;
      RECT 66.025000 176.900000 66.555000 183.570000 ;
      RECT 66.025000 186.900000 66.555000 193.570000 ;
      RECT 66.700000   1.205000 67.230000   1.735000 ;
      RECT 66.710000  75.785000 66.880000  80.535000 ;
      RECT 66.710000  82.785000 66.880000  89.375000 ;
      RECT 66.710000  91.280000 66.880000  97.870000 ;
      RECT 66.710000 101.385000 66.880000 106.255000 ;
      RECT 66.710000 110.450000 66.880000 115.270000 ;
      RECT 66.710000 120.080000 66.880000 124.860000 ;
      RECT 67.290000  26.015000 68.140000  82.180000 ;
      RECT 67.290000  82.350000 68.140000  90.675000 ;
      RECT 67.290000  90.845000 68.140000  98.990000 ;
      RECT 67.575000 101.035000 68.495000 109.275000 ;
      RECT 67.575000 109.445000 68.495000 117.770000 ;
      RECT 67.575000 117.940000 68.495000 194.935000 ;
      RECT 67.610000   1.080000 73.375000   1.250000 ;
      RECT 67.615000   1.250000 67.785000  17.100000 ;
      RECT 67.615000  17.100000 73.375000  17.270000 ;
      RECT 68.110000   3.280000 68.280000   9.020000 ;
      RECT 68.110000   9.770000 68.280000  16.670000 ;
      RECT 68.335000   1.670000 72.655000   1.840000 ;
      RECT 68.335000   9.320000 72.655000   9.490000 ;
      RECT 68.570000   2.550000 68.740000   9.020000 ;
      RECT 68.570000  10.200000 68.740000  15.660000 ;
      RECT 69.030000   3.280000 69.200000   9.020000 ;
      RECT 69.030000   9.770000 69.200000  16.670000 ;
      RECT 69.190000  24.355000 69.720000  99.925000 ;
      RECT 69.190000 100.095000 69.720000 196.850000 ;
      RECT 69.490000   2.550000 69.660000   9.020000 ;
      RECT 69.490000  10.200000 69.660000  15.660000 ;
      RECT 69.530000  19.010000 70.265000  19.610000 ;
      RECT 69.950000   3.280000 70.120000   9.020000 ;
      RECT 69.950000   9.770000 70.120000  16.670000 ;
      RECT 70.410000   2.550000 70.580000   9.020000 ;
      RECT 70.410000  10.200000 70.580000  15.660000 ;
      RECT 70.495000  17.960000 71.095000  18.695000 ;
      RECT 70.870000   3.280000 71.040000   9.020000 ;
      RECT 70.870000   9.770000 71.040000  16.670000 ;
      RECT 71.330000   2.550000 71.500000   9.020000 ;
      RECT 71.330000  10.200000 71.500000  15.660000 ;
      RECT 71.790000   3.280000 71.960000   9.020000 ;
      RECT 71.790000   9.770000 71.960000  16.670000 ;
      RECT 72.250000   2.550000 72.420000   9.020000 ;
      RECT 72.250000  10.200000 72.420000  15.660000 ;
      RECT 72.710000   2.120000 72.880000   9.020000 ;
      RECT 72.710000   9.770000 72.880000  16.670000 ;
      RECT 73.205000   1.250000 73.375000  17.100000 ;
      RECT 73.875000 196.920000 74.755000 197.780000 ;
    LAYER met1 ;
      RECT  0.000000   0.000000 25.930000   0.295000 ;
      RECT  0.000000   0.000000 26.070000   0.310000 ;
      RECT  0.000000   0.295000 25.930000   0.310000 ;
      RECT  0.000000   0.310000 25.945000   0.325000 ;
      RECT  0.000000   0.310000 75.000000 198.000000 ;
      RECT  0.000000   0.325000 75.000000   3.330000 ;
      RECT  0.000000   3.330000  3.005000 194.995000 ;
      RECT  0.000000 194.995000 75.000000 198.000000 ;
      RECT  3.000000   3.002000 24.390000   3.070000 ;
      RECT  3.000000   3.002000 24.390000   3.070000 ;
      RECT  3.000000   3.070000 24.460000   3.140000 ;
      RECT  3.000000   3.070000 24.460000   3.140000 ;
      RECT  3.000000   3.140000 24.530000   3.210000 ;
      RECT  3.000000   3.140000 24.530000   3.210000 ;
      RECT  3.000000   3.210000 24.600000   3.280000 ;
      RECT  3.000000   3.210000 24.600000   3.280000 ;
      RECT  3.000000   3.280000 24.670000   3.325000 ;
      RECT  3.000000   3.280000 24.670000   3.325000 ;
      RECT  3.000000   3.325000 72.000000 195.000000 ;
      RECT 27.840000   0.000000 75.000000   0.310000 ;
      RECT 27.950000   0.320000 75.000000   0.325000 ;
      RECT 27.965000   0.305000 75.000000   0.320000 ;
      RECT 27.980000   0.000000 75.000000   0.290000 ;
      RECT 27.980000   0.290000 75.000000   0.305000 ;
      RECT 30.950000   3.000000 72.000000   6.330000 ;
      RECT 71.995000   3.330000 75.000000 194.995000 ;
    LAYER met2 ;
      RECT  0.000000   0.000000  0.220000 193.910000 ;
      RECT  0.000000   0.000000  0.220000 193.910000 ;
      RECT  0.000000 193.910000 75.000000 198.000000 ;
      RECT  0.000000 193.910000 75.000000 198.000000 ;
      RECT 10.700000   8.165000 11.735000   9.705000 ;
      RECT 10.700000   8.165000 11.735000   9.705000 ;
      RECT 10.700000   9.705000 11.735000   9.715000 ;
      RECT 10.705000   8.160000 11.735000   8.165000 ;
      RECT 10.705000   8.160000 11.735000   8.165000 ;
      RECT 10.705000   9.705000 11.735000   9.710000 ;
      RECT 10.710000   9.710000 11.735000   9.715000 ;
      RECT 10.710000   9.715000 11.515000   9.935000 ;
      RECT 10.720000   8.145000 11.720000   8.160000 ;
      RECT 10.780000   9.715000 11.665000   9.785000 ;
      RECT 10.790000   8.075000 11.650000   8.145000 ;
      RECT 10.850000   9.785000 11.595000   9.855000 ;
      RECT 10.860000   8.005000 11.580000   8.075000 ;
      RECT 10.920000   9.855000 11.525000   9.925000 ;
      RECT 10.930000   7.935000 11.510000   8.005000 ;
      RECT 10.930000   7.935000 11.735000   8.160000 ;
      RECT 10.930000   9.925000 11.515000   9.935000 ;
      RECT 14.030000  25.300000 65.465000  25.370000 ;
      RECT 14.030000  25.300000 65.465000  25.370000 ;
      RECT 14.030000  25.300000 65.860000  25.500000 ;
      RECT 14.030000  25.370000 65.535000  25.440000 ;
      RECT 14.030000  25.370000 65.535000  25.440000 ;
      RECT 14.030000  25.440000 65.605000  25.510000 ;
      RECT 14.030000  25.440000 65.605000  25.510000 ;
      RECT 14.030000  25.500000 65.860000  29.820000 ;
      RECT 14.030000  25.510000 65.675000  25.555000 ;
      RECT 14.030000  25.510000 65.675000  25.555000 ;
      RECT 14.030000  25.555000 65.720000  29.765000 ;
      RECT 14.030000  29.765000 65.650000  29.835000 ;
      RECT 14.030000  29.765000 65.650000  29.835000 ;
      RECT 14.030000  29.820000 64.810000  30.870000 ;
      RECT 14.030000  29.835000 65.580000  29.905000 ;
      RECT 14.030000  29.835000 65.580000  29.905000 ;
      RECT 14.030000  29.905000 65.510000  29.975000 ;
      RECT 14.030000  29.905000 65.510000  29.975000 ;
      RECT 14.030000  29.975000 65.440000  30.045000 ;
      RECT 14.030000  29.975000 65.440000  30.045000 ;
      RECT 14.030000  30.045000 65.370000  30.115000 ;
      RECT 14.030000  30.045000 65.370000  30.115000 ;
      RECT 14.030000  30.115000 65.300000  30.185000 ;
      RECT 14.030000  30.115000 65.300000  30.185000 ;
      RECT 14.030000  30.185000 65.230000  30.255000 ;
      RECT 14.030000  30.185000 65.230000  30.255000 ;
      RECT 14.030000  30.255000 65.160000  30.325000 ;
      RECT 14.030000  30.255000 65.160000  30.325000 ;
      RECT 14.030000  30.325000 65.090000  30.395000 ;
      RECT 14.030000  30.325000 65.090000  30.395000 ;
      RECT 14.030000  30.395000 65.020000  30.465000 ;
      RECT 14.030000  30.395000 65.020000  30.465000 ;
      RECT 14.030000  30.465000 64.950000  30.535000 ;
      RECT 14.030000  30.465000 64.950000  30.535000 ;
      RECT 14.030000  30.535000 64.880000  30.605000 ;
      RECT 14.030000  30.535000 64.880000  30.605000 ;
      RECT 14.030000  30.605000 64.810000  30.675000 ;
      RECT 14.030000  30.605000 64.810000  30.675000 ;
      RECT 14.030000  30.675000 64.755000  30.730000 ;
      RECT 14.030000  30.675000 64.755000  30.730000 ;
      RECT 14.030000  30.730000 15.855000  33.930000 ;
      RECT 14.030000  30.870000 15.995000  33.790000 ;
      RECT 14.030000  33.790000 65.860000  34.750000 ;
      RECT 14.030000  33.930000 64.845000  34.000000 ;
      RECT 14.030000  33.930000 64.845000  34.000000 ;
      RECT 14.030000  34.000000 64.915000  34.070000 ;
      RECT 14.030000  34.000000 64.915000  34.070000 ;
      RECT 14.030000  34.070000 64.985000  34.140000 ;
      RECT 14.030000  34.070000 64.985000  34.140000 ;
      RECT 14.030000  34.140000 65.055000  34.210000 ;
      RECT 14.030000  34.140000 65.055000  34.210000 ;
      RECT 14.030000  34.210000 65.125000  34.280000 ;
      RECT 14.030000  34.210000 65.125000  34.280000 ;
      RECT 14.030000  34.280000 65.195000  34.350000 ;
      RECT 14.030000  34.280000 65.195000  34.350000 ;
      RECT 14.030000  34.350000 65.265000  34.420000 ;
      RECT 14.030000  34.350000 65.265000  34.420000 ;
      RECT 14.030000  34.420000 65.335000  34.490000 ;
      RECT 14.030000  34.420000 65.335000  34.490000 ;
      RECT 14.030000  34.490000 65.405000  34.560000 ;
      RECT 14.030000  34.490000 65.405000  34.560000 ;
      RECT 14.030000  34.560000 65.475000  34.630000 ;
      RECT 14.030000  34.560000 65.475000  34.630000 ;
      RECT 14.030000  34.630000 65.545000  34.700000 ;
      RECT 14.030000  34.630000 65.545000  34.700000 ;
      RECT 14.030000  34.700000 65.615000  34.770000 ;
      RECT 14.030000  34.700000 65.615000  34.770000 ;
      RECT 14.030000  34.750000 65.860000  39.875000 ;
      RECT 14.030000  34.770000 65.685000  34.805000 ;
      RECT 14.030000  34.770000 65.685000  34.805000 ;
      RECT 14.030000  34.805000 65.720000  39.820000 ;
      RECT 14.030000  39.820000 65.650000  39.890000 ;
      RECT 14.030000  39.820000 65.650000  39.890000 ;
      RECT 14.030000  39.875000 64.885000  40.850000 ;
      RECT 14.030000  39.890000 65.580000  39.960000 ;
      RECT 14.030000  39.890000 65.580000  39.960000 ;
      RECT 14.030000  39.960000 65.510000  40.030000 ;
      RECT 14.030000  39.960000 65.510000  40.030000 ;
      RECT 14.030000  40.030000 65.440000  40.100000 ;
      RECT 14.030000  40.030000 65.440000  40.100000 ;
      RECT 14.030000  40.100000 65.370000  40.170000 ;
      RECT 14.030000  40.100000 65.370000  40.170000 ;
      RECT 14.030000  40.170000 65.300000  40.240000 ;
      RECT 14.030000  40.170000 65.300000  40.240000 ;
      RECT 14.030000  40.240000 65.230000  40.310000 ;
      RECT 14.030000  40.240000 65.230000  40.310000 ;
      RECT 14.030000  40.310000 65.160000  40.380000 ;
      RECT 14.030000  40.310000 65.160000  40.380000 ;
      RECT 14.030000  40.380000 65.090000  40.450000 ;
      RECT 14.030000  40.380000 65.090000  40.450000 ;
      RECT 14.030000  40.450000 65.020000  40.520000 ;
      RECT 14.030000  40.450000 65.020000  40.520000 ;
      RECT 14.030000  40.520000 64.950000  40.590000 ;
      RECT 14.030000  40.520000 64.950000  40.590000 ;
      RECT 14.030000  40.590000 64.880000  40.660000 ;
      RECT 14.030000  40.590000 64.880000  40.660000 ;
      RECT 14.030000  40.660000 64.830000  40.710000 ;
      RECT 14.030000  40.660000 64.830000  40.710000 ;
      RECT 14.030000  40.710000 15.855000  43.910000 ;
      RECT 14.030000  40.850000 15.995000  43.770000 ;
      RECT 14.030000  43.770000 65.860000  44.730000 ;
      RECT 14.030000  43.910000 64.845000  43.980000 ;
      RECT 14.030000  43.910000 64.845000  43.980000 ;
      RECT 14.030000  43.980000 64.915000  44.050000 ;
      RECT 14.030000  43.980000 64.915000  44.050000 ;
      RECT 14.030000  44.050000 64.985000  44.120000 ;
      RECT 14.030000  44.050000 64.985000  44.120000 ;
      RECT 14.030000  44.120000 65.055000  44.190000 ;
      RECT 14.030000  44.120000 65.055000  44.190000 ;
      RECT 14.030000  44.190000 65.125000  44.260000 ;
      RECT 14.030000  44.190000 65.125000  44.260000 ;
      RECT 14.030000  44.260000 65.195000  44.330000 ;
      RECT 14.030000  44.260000 65.195000  44.330000 ;
      RECT 14.030000  44.330000 65.265000  44.400000 ;
      RECT 14.030000  44.330000 65.265000  44.400000 ;
      RECT 14.030000  44.400000 65.335000  44.470000 ;
      RECT 14.030000  44.400000 65.335000  44.470000 ;
      RECT 14.030000  44.470000 65.405000  44.540000 ;
      RECT 14.030000  44.470000 65.405000  44.540000 ;
      RECT 14.030000  44.540000 65.475000  44.610000 ;
      RECT 14.030000  44.540000 65.475000  44.610000 ;
      RECT 14.030000  44.610000 65.545000  44.680000 ;
      RECT 14.030000  44.610000 65.545000  44.680000 ;
      RECT 14.030000  44.680000 65.615000  44.750000 ;
      RECT 14.030000  44.680000 65.615000  44.750000 ;
      RECT 14.030000  44.730000 65.860000  49.895000 ;
      RECT 14.030000  44.750000 65.685000  44.785000 ;
      RECT 14.030000  44.750000 65.685000  44.785000 ;
      RECT 14.030000  44.785000 65.720000  49.840000 ;
      RECT 14.030000  49.840000 65.650000  49.910000 ;
      RECT 14.030000  49.840000 65.650000  49.910000 ;
      RECT 14.030000  49.895000 64.885000  50.870000 ;
      RECT 14.030000  49.910000 65.580000  49.980000 ;
      RECT 14.030000  49.910000 65.580000  49.980000 ;
      RECT 14.030000  49.980000 65.510000  50.050000 ;
      RECT 14.030000  49.980000 65.510000  50.050000 ;
      RECT 14.030000  50.050000 65.440000  50.120000 ;
      RECT 14.030000  50.050000 65.440000  50.120000 ;
      RECT 14.030000  50.120000 65.370000  50.190000 ;
      RECT 14.030000  50.120000 65.370000  50.190000 ;
      RECT 14.030000  50.190000 65.300000  50.260000 ;
      RECT 14.030000  50.190000 65.300000  50.260000 ;
      RECT 14.030000  50.260000 65.230000  50.330000 ;
      RECT 14.030000  50.260000 65.230000  50.330000 ;
      RECT 14.030000  50.330000 65.160000  50.400000 ;
      RECT 14.030000  50.330000 65.160000  50.400000 ;
      RECT 14.030000  50.400000 65.090000  50.470000 ;
      RECT 14.030000  50.400000 65.090000  50.470000 ;
      RECT 14.030000  50.470000 65.020000  50.540000 ;
      RECT 14.030000  50.470000 65.020000  50.540000 ;
      RECT 14.030000  50.540000 64.950000  50.610000 ;
      RECT 14.030000  50.540000 64.950000  50.610000 ;
      RECT 14.030000  50.610000 64.880000  50.680000 ;
      RECT 14.030000  50.610000 64.880000  50.680000 ;
      RECT 14.030000  50.680000 64.830000  50.730000 ;
      RECT 14.030000  50.680000 64.830000  50.730000 ;
      RECT 14.030000  50.730000 15.855000  53.930000 ;
      RECT 14.030000  50.870000 15.995000  53.790000 ;
      RECT 14.030000  53.790000 65.855000  54.745000 ;
      RECT 14.030000  53.930000 64.845000  54.000000 ;
      RECT 14.030000  53.930000 64.845000  54.000000 ;
      RECT 14.030000  54.000000 64.915000  54.070000 ;
      RECT 14.030000  54.000000 64.915000  54.070000 ;
      RECT 14.030000  54.070000 64.985000  54.140000 ;
      RECT 14.030000  54.070000 64.985000  54.140000 ;
      RECT 14.030000  54.140000 65.055000  54.210000 ;
      RECT 14.030000  54.140000 65.055000  54.210000 ;
      RECT 14.030000  54.210000 65.125000  54.280000 ;
      RECT 14.030000  54.210000 65.125000  54.280000 ;
      RECT 14.030000  54.280000 65.195000  54.350000 ;
      RECT 14.030000  54.280000 65.195000  54.350000 ;
      RECT 14.030000  54.350000 65.265000  54.420000 ;
      RECT 14.030000  54.350000 65.265000  54.420000 ;
      RECT 14.030000  54.420000 65.335000  54.490000 ;
      RECT 14.030000  54.420000 65.335000  54.490000 ;
      RECT 14.030000  54.490000 65.405000  54.560000 ;
      RECT 14.030000  54.490000 65.405000  54.560000 ;
      RECT 14.030000  54.560000 65.475000  54.630000 ;
      RECT 14.030000  54.560000 65.475000  54.630000 ;
      RECT 14.030000  54.630000 65.545000  54.700000 ;
      RECT 14.030000  54.630000 65.545000  54.700000 ;
      RECT 14.030000  54.700000 65.615000  54.770000 ;
      RECT 14.030000  54.700000 65.615000  54.770000 ;
      RECT 14.030000  54.745000 65.855000  59.880000 ;
      RECT 14.030000  54.770000 65.685000  54.800000 ;
      RECT 14.030000  54.770000 65.685000  54.800000 ;
      RECT 14.030000  54.800000 65.715000  59.825000 ;
      RECT 14.030000  59.825000 65.645000  59.895000 ;
      RECT 14.030000  59.825000 65.645000  59.895000 ;
      RECT 14.030000  59.880000 64.885000  60.850000 ;
      RECT 14.030000  59.895000 65.575000  59.965000 ;
      RECT 14.030000  59.895000 65.575000  59.965000 ;
      RECT 14.030000  59.965000 65.505000  60.035000 ;
      RECT 14.030000  59.965000 65.505000  60.035000 ;
      RECT 14.030000  60.035000 65.435000  60.105000 ;
      RECT 14.030000  60.035000 65.435000  60.105000 ;
      RECT 14.030000  60.105000 65.365000  60.175000 ;
      RECT 14.030000  60.105000 65.365000  60.175000 ;
      RECT 14.030000  60.175000 65.295000  60.245000 ;
      RECT 14.030000  60.175000 65.295000  60.245000 ;
      RECT 14.030000  60.245000 65.225000  60.315000 ;
      RECT 14.030000  60.245000 65.225000  60.315000 ;
      RECT 14.030000  60.315000 65.155000  60.385000 ;
      RECT 14.030000  60.315000 65.155000  60.385000 ;
      RECT 14.030000  60.385000 65.085000  60.455000 ;
      RECT 14.030000  60.385000 65.085000  60.455000 ;
      RECT 14.030000  60.455000 65.015000  60.525000 ;
      RECT 14.030000  60.455000 65.015000  60.525000 ;
      RECT 14.030000  60.525000 64.945000  60.595000 ;
      RECT 14.030000  60.525000 64.945000  60.595000 ;
      RECT 14.030000  60.595000 64.875000  60.665000 ;
      RECT 14.030000  60.595000 64.875000  60.665000 ;
      RECT 14.030000  60.665000 64.830000  60.710000 ;
      RECT 14.030000  60.665000 64.830000  60.710000 ;
      RECT 14.030000  60.710000 15.855000  63.910000 ;
      RECT 14.030000  60.850000 15.995000  63.770000 ;
      RECT 14.030000  63.770000 65.855000  64.735000 ;
      RECT 14.030000  63.910000 64.830000  63.980000 ;
      RECT 14.030000  63.910000 64.830000  63.980000 ;
      RECT 14.030000  63.980000 64.900000  64.050000 ;
      RECT 14.030000  63.980000 64.900000  64.050000 ;
      RECT 14.030000  64.050000 64.970000  64.120000 ;
      RECT 14.030000  64.050000 64.970000  64.120000 ;
      RECT 14.030000  64.120000 65.040000  64.190000 ;
      RECT 14.030000  64.120000 65.040000  64.190000 ;
      RECT 14.030000  64.190000 65.110000  64.260000 ;
      RECT 14.030000  64.190000 65.110000  64.260000 ;
      RECT 14.030000  64.260000 65.180000  64.330000 ;
      RECT 14.030000  64.260000 65.180000  64.330000 ;
      RECT 14.030000  64.330000 65.250000  64.400000 ;
      RECT 14.030000  64.330000 65.250000  64.400000 ;
      RECT 14.030000  64.400000 65.320000  64.470000 ;
      RECT 14.030000  64.400000 65.320000  64.470000 ;
      RECT 14.030000  64.470000 65.390000  64.540000 ;
      RECT 14.030000  64.470000 65.390000  64.540000 ;
      RECT 14.030000  64.540000 65.460000  64.610000 ;
      RECT 14.030000  64.540000 65.460000  64.610000 ;
      RECT 14.030000  64.610000 65.530000  64.680000 ;
      RECT 14.030000  64.610000 65.530000  64.680000 ;
      RECT 14.030000  64.680000 65.600000  64.750000 ;
      RECT 14.030000  64.680000 65.600000  64.750000 ;
      RECT 14.030000  64.735000 65.855000  69.880000 ;
      RECT 14.030000  64.750000 65.670000  64.795000 ;
      RECT 14.030000  64.750000 65.670000  64.795000 ;
      RECT 14.030000  64.795000 65.715000  69.825000 ;
      RECT 14.030000  69.825000 65.645000  69.895000 ;
      RECT 14.030000  69.825000 65.645000  69.895000 ;
      RECT 14.030000  69.880000 64.885000  70.850000 ;
      RECT 14.030000  69.895000 65.575000  69.965000 ;
      RECT 14.030000  69.895000 65.575000  69.965000 ;
      RECT 14.030000  69.965000 65.505000  70.035000 ;
      RECT 14.030000  69.965000 65.505000  70.035000 ;
      RECT 14.030000  70.035000 65.435000  70.105000 ;
      RECT 14.030000  70.035000 65.435000  70.105000 ;
      RECT 14.030000  70.105000 65.365000  70.175000 ;
      RECT 14.030000  70.105000 65.365000  70.175000 ;
      RECT 14.030000  70.175000 65.295000  70.245000 ;
      RECT 14.030000  70.175000 65.295000  70.245000 ;
      RECT 14.030000  70.245000 65.225000  70.315000 ;
      RECT 14.030000  70.245000 65.225000  70.315000 ;
      RECT 14.030000  70.315000 65.155000  70.385000 ;
      RECT 14.030000  70.315000 65.155000  70.385000 ;
      RECT 14.030000  70.385000 65.085000  70.455000 ;
      RECT 14.030000  70.385000 65.085000  70.455000 ;
      RECT 14.030000  70.455000 65.015000  70.525000 ;
      RECT 14.030000  70.455000 65.015000  70.525000 ;
      RECT 14.030000  70.525000 64.945000  70.595000 ;
      RECT 14.030000  70.525000 64.945000  70.595000 ;
      RECT 14.030000  70.595000 64.875000  70.665000 ;
      RECT 14.030000  70.595000 64.875000  70.665000 ;
      RECT 14.030000  70.665000 64.830000  70.710000 ;
      RECT 14.030000  70.665000 64.830000  70.710000 ;
      RECT 14.030000  70.710000 15.855000  73.910000 ;
      RECT 14.030000  70.850000 15.995000  73.770000 ;
      RECT 14.030000  73.770000 65.550000  74.180000 ;
      RECT 14.030000  73.910000 65.085000  73.980000 ;
      RECT 14.030000  73.980000 65.155000  74.050000 ;
      RECT 14.030000  74.050000 65.225000  74.120000 ;
      RECT 14.030000  74.120000 65.295000  74.180000 ;
      RECT 14.030000  74.180000 65.760000  74.390000 ;
      RECT 14.065000  25.265000 65.430000  25.300000 ;
      RECT 14.065000  25.265000 65.430000  25.300000 ;
      RECT 14.100000  74.180000 65.350000  74.250000 ;
      RECT 14.135000  25.195000 65.360000  25.265000 ;
      RECT 14.135000  25.195000 65.360000  25.265000 ;
      RECT 14.170000  74.250000 65.425000  74.320000 ;
      RECT 14.205000  25.125000 65.290000  25.195000 ;
      RECT 14.205000  25.125000 65.290000  25.195000 ;
      RECT 14.240000  73.910000 65.085000  73.980000 ;
      RECT 14.240000  73.910000 65.085000  73.980000 ;
      RECT 14.240000  73.980000 65.155000  74.050000 ;
      RECT 14.240000  73.980000 65.155000  74.050000 ;
      RECT 14.240000  74.050000 65.225000  74.120000 ;
      RECT 14.240000  74.050000 65.225000  74.120000 ;
      RECT 14.240000  74.120000 65.295000  74.180000 ;
      RECT 14.240000  74.120000 65.295000  74.180000 ;
      RECT 14.240000  74.180000 65.350000  74.250000 ;
      RECT 14.240000  74.180000 65.350000  74.250000 ;
      RECT 14.240000  74.250000 65.425000  74.320000 ;
      RECT 14.240000  74.250000 65.425000  74.320000 ;
      RECT 14.240000  74.320000 65.495000  74.390000 ;
      RECT 14.240000  74.320000 65.495000  74.390000 ;
      RECT 14.240000  74.320000 65.495000  74.390000 ;
      RECT 14.240000  74.390000 65.565000  74.460000 ;
      RECT 14.240000  74.390000 65.565000  74.460000 ;
      RECT 14.240000  74.390000 65.860000  74.490000 ;
      RECT 14.240000  74.460000 65.635000  74.530000 ;
      RECT 14.240000  74.460000 65.635000  74.530000 ;
      RECT 14.240000  74.490000 65.860000  98.700000 ;
      RECT 14.240000  74.530000 65.705000  74.545000 ;
      RECT 14.240000  74.530000 65.705000  74.545000 ;
      RECT 14.240000  74.545000 65.720000  98.840000 ;
      RECT 14.240000  98.700000 75.000000 129.820000 ;
      RECT 14.240000  98.840000 75.000000 129.820000 ;
      RECT 14.240000 129.820000 75.000000 130.705000 ;
      RECT 14.240000 134.795000 75.000000 139.825000 ;
      RECT 14.240000 134.795000 75.000000 139.825000 ;
      RECT 14.240000 139.825000 75.000000 140.710000 ;
      RECT 14.240000 144.795000 75.000000 149.825000 ;
      RECT 14.240000 144.795000 75.000000 149.825000 ;
      RECT 14.240000 149.825000 75.000000 150.710000 ;
      RECT 14.240000 154.795000 75.000000 159.825000 ;
      RECT 14.240000 154.795000 75.000000 159.825000 ;
      RECT 14.240000 159.825000 75.000000 160.710000 ;
      RECT 14.240000 164.795000 75.000000 169.825000 ;
      RECT 14.240000 164.795000 75.000000 169.825000 ;
      RECT 14.240000 169.825000 75.000000 170.710000 ;
      RECT 14.240000 174.795000 75.000000 179.825000 ;
      RECT 14.240000 174.795000 75.000000 179.825000 ;
      RECT 14.240000 179.825000 75.000000 180.710000 ;
      RECT 14.240000 184.795000 75.000000 189.825000 ;
      RECT 14.240000 184.795000 75.000000 189.825000 ;
      RECT 14.240000 189.825000 75.000000 190.710000 ;
      RECT 14.275000  25.055000 65.220000  25.125000 ;
      RECT 14.275000  25.055000 65.220000  25.125000 ;
      RECT 14.285000 134.750000 75.000000 134.795000 ;
      RECT 14.285000 134.750000 75.000000 134.795000 ;
      RECT 14.285000 144.750000 75.000000 144.795000 ;
      RECT 14.285000 144.750000 75.000000 144.795000 ;
      RECT 14.285000 154.750000 75.000000 154.795000 ;
      RECT 14.285000 154.750000 75.000000 154.795000 ;
      RECT 14.285000 164.750000 75.000000 164.795000 ;
      RECT 14.285000 164.750000 75.000000 164.795000 ;
      RECT 14.285000 174.750000 75.000000 174.795000 ;
      RECT 14.285000 174.750000 75.000000 174.795000 ;
      RECT 14.285000 184.750000 75.000000 184.795000 ;
      RECT 14.285000 184.750000 75.000000 184.795000 ;
      RECT 14.310000 129.820000 75.000000 129.890000 ;
      RECT 14.310000 129.820000 75.000000 129.890000 ;
      RECT 14.310000 139.825000 75.000000 139.895000 ;
      RECT 14.310000 139.825000 75.000000 139.895000 ;
      RECT 14.310000 149.825000 75.000000 149.895000 ;
      RECT 14.310000 149.825000 75.000000 149.895000 ;
      RECT 14.310000 159.825000 75.000000 159.895000 ;
      RECT 14.310000 159.825000 75.000000 159.895000 ;
      RECT 14.310000 169.825000 75.000000 169.895000 ;
      RECT 14.310000 169.825000 75.000000 169.895000 ;
      RECT 14.310000 179.825000 75.000000 179.895000 ;
      RECT 14.310000 179.825000 75.000000 179.895000 ;
      RECT 14.310000 189.825000 75.000000 189.895000 ;
      RECT 14.310000 189.825000 75.000000 189.895000 ;
      RECT 14.345000  24.985000 65.150000  25.055000 ;
      RECT 14.345000  24.985000 65.150000  25.055000 ;
      RECT 14.355000 134.680000 75.000000 134.750000 ;
      RECT 14.355000 134.680000 75.000000 134.750000 ;
      RECT 14.355000 144.680000 75.000000 144.750000 ;
      RECT 14.355000 144.680000 75.000000 144.750000 ;
      RECT 14.355000 154.680000 75.000000 154.750000 ;
      RECT 14.355000 154.680000 75.000000 154.750000 ;
      RECT 14.355000 164.680000 75.000000 164.750000 ;
      RECT 14.355000 164.680000 75.000000 164.750000 ;
      RECT 14.355000 174.680000 75.000000 174.750000 ;
      RECT 14.355000 174.680000 75.000000 174.750000 ;
      RECT 14.355000 184.680000 75.000000 184.750000 ;
      RECT 14.355000 184.680000 75.000000 184.750000 ;
      RECT 14.380000 129.890000 75.000000 129.960000 ;
      RECT 14.380000 129.890000 75.000000 129.960000 ;
      RECT 14.380000 139.895000 75.000000 139.965000 ;
      RECT 14.380000 139.895000 75.000000 139.965000 ;
      RECT 14.380000 149.895000 75.000000 149.965000 ;
      RECT 14.380000 149.895000 75.000000 149.965000 ;
      RECT 14.380000 159.895000 75.000000 159.965000 ;
      RECT 14.380000 159.895000 75.000000 159.965000 ;
      RECT 14.380000 169.895000 75.000000 169.965000 ;
      RECT 14.380000 169.895000 75.000000 169.965000 ;
      RECT 14.380000 179.895000 75.000000 179.965000 ;
      RECT 14.380000 179.895000 75.000000 179.965000 ;
      RECT 14.380000 189.895000 75.000000 189.965000 ;
      RECT 14.380000 189.895000 75.000000 189.965000 ;
      RECT 14.415000  24.915000 65.080000  24.985000 ;
      RECT 14.415000  24.915000 65.080000  24.985000 ;
      RECT 14.425000 134.610000 75.000000 134.680000 ;
      RECT 14.425000 134.610000 75.000000 134.680000 ;
      RECT 14.425000 144.610000 75.000000 144.680000 ;
      RECT 14.425000 144.610000 75.000000 144.680000 ;
      RECT 14.425000 154.610000 75.000000 154.680000 ;
      RECT 14.425000 154.610000 75.000000 154.680000 ;
      RECT 14.425000 164.610000 75.000000 164.680000 ;
      RECT 14.425000 164.610000 75.000000 164.680000 ;
      RECT 14.425000 174.610000 75.000000 174.680000 ;
      RECT 14.425000 174.610000 75.000000 174.680000 ;
      RECT 14.425000 184.610000 75.000000 184.680000 ;
      RECT 14.425000 184.610000 75.000000 184.680000 ;
      RECT 14.450000 129.960000 75.000000 130.030000 ;
      RECT 14.450000 129.960000 75.000000 130.030000 ;
      RECT 14.450000 139.965000 75.000000 140.035000 ;
      RECT 14.450000 139.965000 75.000000 140.035000 ;
      RECT 14.450000 149.965000 75.000000 150.035000 ;
      RECT 14.450000 149.965000 75.000000 150.035000 ;
      RECT 14.450000 159.965000 75.000000 160.035000 ;
      RECT 14.450000 159.965000 75.000000 160.035000 ;
      RECT 14.450000 169.965000 75.000000 170.035000 ;
      RECT 14.450000 169.965000 75.000000 170.035000 ;
      RECT 14.450000 179.965000 75.000000 180.035000 ;
      RECT 14.450000 179.965000 75.000000 180.035000 ;
      RECT 14.450000 189.965000 75.000000 190.035000 ;
      RECT 14.450000 189.965000 75.000000 190.035000 ;
      RECT 14.485000  24.845000 65.010000  24.915000 ;
      RECT 14.485000  24.845000 65.010000  24.915000 ;
      RECT 14.495000 134.540000 75.000000 134.610000 ;
      RECT 14.495000 134.540000 75.000000 134.610000 ;
      RECT 14.495000 144.540000 75.000000 144.610000 ;
      RECT 14.495000 144.540000 75.000000 144.610000 ;
      RECT 14.495000 154.540000 75.000000 154.610000 ;
      RECT 14.495000 154.540000 75.000000 154.610000 ;
      RECT 14.495000 164.540000 75.000000 164.610000 ;
      RECT 14.495000 164.540000 75.000000 164.610000 ;
      RECT 14.495000 174.540000 75.000000 174.610000 ;
      RECT 14.495000 174.540000 75.000000 174.610000 ;
      RECT 14.495000 184.540000 75.000000 184.610000 ;
      RECT 14.495000 184.540000 75.000000 184.610000 ;
      RECT 14.520000 130.030000 75.000000 130.100000 ;
      RECT 14.520000 130.030000 75.000000 130.100000 ;
      RECT 14.520000 140.035000 75.000000 140.105000 ;
      RECT 14.520000 140.035000 75.000000 140.105000 ;
      RECT 14.520000 150.035000 75.000000 150.105000 ;
      RECT 14.520000 150.035000 75.000000 150.105000 ;
      RECT 14.520000 160.035000 75.000000 160.105000 ;
      RECT 14.520000 160.035000 75.000000 160.105000 ;
      RECT 14.520000 170.035000 75.000000 170.105000 ;
      RECT 14.520000 170.035000 75.000000 170.105000 ;
      RECT 14.520000 180.035000 75.000000 180.105000 ;
      RECT 14.520000 180.035000 75.000000 180.105000 ;
      RECT 14.520000 190.035000 75.000000 190.105000 ;
      RECT 14.520000 190.035000 75.000000 190.105000 ;
      RECT 14.555000  24.775000 64.940000  24.845000 ;
      RECT 14.555000  24.775000 64.940000  24.845000 ;
      RECT 14.565000 134.470000 75.000000 134.540000 ;
      RECT 14.565000 134.470000 75.000000 134.540000 ;
      RECT 14.565000 144.470000 75.000000 144.540000 ;
      RECT 14.565000 144.470000 75.000000 144.540000 ;
      RECT 14.565000 154.470000 75.000000 154.540000 ;
      RECT 14.565000 154.470000 75.000000 154.540000 ;
      RECT 14.565000 164.470000 75.000000 164.540000 ;
      RECT 14.565000 164.470000 75.000000 164.540000 ;
      RECT 14.565000 174.470000 75.000000 174.540000 ;
      RECT 14.565000 174.470000 75.000000 174.540000 ;
      RECT 14.565000 184.470000 75.000000 184.540000 ;
      RECT 14.565000 184.470000 75.000000 184.540000 ;
      RECT 14.590000 130.100000 75.000000 130.170000 ;
      RECT 14.590000 130.100000 75.000000 130.170000 ;
      RECT 14.590000 140.105000 75.000000 140.175000 ;
      RECT 14.590000 140.105000 75.000000 140.175000 ;
      RECT 14.590000 150.105000 75.000000 150.175000 ;
      RECT 14.590000 150.105000 75.000000 150.175000 ;
      RECT 14.590000 160.105000 75.000000 160.175000 ;
      RECT 14.590000 160.105000 75.000000 160.175000 ;
      RECT 14.590000 170.105000 75.000000 170.175000 ;
      RECT 14.590000 170.105000 75.000000 170.175000 ;
      RECT 14.590000 180.105000 75.000000 180.175000 ;
      RECT 14.590000 180.105000 75.000000 180.175000 ;
      RECT 14.590000 190.105000 75.000000 190.175000 ;
      RECT 14.590000 190.105000 75.000000 190.175000 ;
      RECT 14.625000  24.705000 64.870000  24.775000 ;
      RECT 14.625000  24.705000 64.870000  24.775000 ;
      RECT 14.635000 134.400000 75.000000 134.470000 ;
      RECT 14.635000 134.400000 75.000000 134.470000 ;
      RECT 14.635000 144.400000 75.000000 144.470000 ;
      RECT 14.635000 144.400000 75.000000 144.470000 ;
      RECT 14.635000 154.400000 75.000000 154.470000 ;
      RECT 14.635000 154.400000 75.000000 154.470000 ;
      RECT 14.635000 164.400000 75.000000 164.470000 ;
      RECT 14.635000 164.400000 75.000000 164.470000 ;
      RECT 14.635000 174.400000 75.000000 174.470000 ;
      RECT 14.635000 174.400000 75.000000 174.470000 ;
      RECT 14.635000 184.400000 75.000000 184.470000 ;
      RECT 14.635000 184.400000 75.000000 184.470000 ;
      RECT 14.660000 130.170000 75.000000 130.240000 ;
      RECT 14.660000 130.170000 75.000000 130.240000 ;
      RECT 14.660000 140.175000 75.000000 140.245000 ;
      RECT 14.660000 140.175000 75.000000 140.245000 ;
      RECT 14.660000 150.175000 75.000000 150.245000 ;
      RECT 14.660000 150.175000 75.000000 150.245000 ;
      RECT 14.660000 160.175000 75.000000 160.245000 ;
      RECT 14.660000 160.175000 75.000000 160.245000 ;
      RECT 14.660000 170.175000 75.000000 170.245000 ;
      RECT 14.660000 170.175000 75.000000 170.245000 ;
      RECT 14.660000 180.175000 75.000000 180.245000 ;
      RECT 14.660000 180.175000 75.000000 180.245000 ;
      RECT 14.660000 190.175000 75.000000 190.245000 ;
      RECT 14.660000 190.175000 75.000000 190.245000 ;
      RECT 14.695000  24.635000 64.800000  24.705000 ;
      RECT 14.695000  24.635000 64.800000  24.705000 ;
      RECT 14.705000 134.330000 75.000000 134.400000 ;
      RECT 14.705000 134.330000 75.000000 134.400000 ;
      RECT 14.705000 144.330000 75.000000 144.400000 ;
      RECT 14.705000 144.330000 75.000000 144.400000 ;
      RECT 14.705000 154.330000 75.000000 154.400000 ;
      RECT 14.705000 154.330000 75.000000 154.400000 ;
      RECT 14.705000 164.330000 75.000000 164.400000 ;
      RECT 14.705000 164.330000 75.000000 164.400000 ;
      RECT 14.705000 174.330000 75.000000 174.400000 ;
      RECT 14.705000 174.330000 75.000000 174.400000 ;
      RECT 14.705000 184.330000 75.000000 184.400000 ;
      RECT 14.705000 184.330000 75.000000 184.400000 ;
      RECT 14.730000 130.240000 75.000000 130.310000 ;
      RECT 14.730000 130.240000 75.000000 130.310000 ;
      RECT 14.730000 140.245000 75.000000 140.315000 ;
      RECT 14.730000 140.245000 75.000000 140.315000 ;
      RECT 14.730000 150.245000 75.000000 150.315000 ;
      RECT 14.730000 150.245000 75.000000 150.315000 ;
      RECT 14.730000 160.245000 75.000000 160.315000 ;
      RECT 14.730000 160.245000 75.000000 160.315000 ;
      RECT 14.730000 170.245000 75.000000 170.315000 ;
      RECT 14.730000 170.245000 75.000000 170.315000 ;
      RECT 14.730000 180.245000 75.000000 180.315000 ;
      RECT 14.730000 180.245000 75.000000 180.315000 ;
      RECT 14.730000 190.245000 75.000000 190.315000 ;
      RECT 14.730000 190.245000 75.000000 190.315000 ;
      RECT 14.765000  24.565000 64.730000  24.635000 ;
      RECT 14.765000  24.565000 64.730000  24.635000 ;
      RECT 14.775000 134.260000 75.000000 134.330000 ;
      RECT 14.775000 134.260000 75.000000 134.330000 ;
      RECT 14.775000 144.260000 75.000000 144.330000 ;
      RECT 14.775000 144.260000 75.000000 144.330000 ;
      RECT 14.775000 154.260000 75.000000 154.330000 ;
      RECT 14.775000 154.260000 75.000000 154.330000 ;
      RECT 14.775000 164.260000 75.000000 164.330000 ;
      RECT 14.775000 164.260000 75.000000 164.330000 ;
      RECT 14.775000 174.260000 75.000000 174.330000 ;
      RECT 14.775000 174.260000 75.000000 174.330000 ;
      RECT 14.775000 184.260000 75.000000 184.330000 ;
      RECT 14.775000 184.260000 75.000000 184.330000 ;
      RECT 14.800000 130.310000 75.000000 130.380000 ;
      RECT 14.800000 130.310000 75.000000 130.380000 ;
      RECT 14.800000 140.315000 75.000000 140.385000 ;
      RECT 14.800000 140.315000 75.000000 140.385000 ;
      RECT 14.800000 150.315000 75.000000 150.385000 ;
      RECT 14.800000 150.315000 75.000000 150.385000 ;
      RECT 14.800000 160.315000 75.000000 160.385000 ;
      RECT 14.800000 160.315000 75.000000 160.385000 ;
      RECT 14.800000 170.315000 75.000000 170.385000 ;
      RECT 14.800000 170.315000 75.000000 170.385000 ;
      RECT 14.800000 180.315000 75.000000 180.385000 ;
      RECT 14.800000 180.315000 75.000000 180.385000 ;
      RECT 14.800000 190.315000 75.000000 190.385000 ;
      RECT 14.800000 190.315000 75.000000 190.385000 ;
      RECT 14.835000  24.495000 64.660000  24.565000 ;
      RECT 14.835000  24.495000 64.660000  24.565000 ;
      RECT 14.845000 134.190000 75.000000 134.260000 ;
      RECT 14.845000 134.190000 75.000000 134.260000 ;
      RECT 14.845000 144.190000 75.000000 144.260000 ;
      RECT 14.845000 144.190000 75.000000 144.260000 ;
      RECT 14.845000 154.190000 75.000000 154.260000 ;
      RECT 14.845000 154.190000 75.000000 154.260000 ;
      RECT 14.845000 164.190000 75.000000 164.260000 ;
      RECT 14.845000 164.190000 75.000000 164.260000 ;
      RECT 14.845000 174.190000 75.000000 174.260000 ;
      RECT 14.845000 174.190000 75.000000 174.260000 ;
      RECT 14.845000 184.190000 75.000000 184.260000 ;
      RECT 14.845000 184.190000 75.000000 184.260000 ;
      RECT 14.870000 130.380000 75.000000 130.450000 ;
      RECT 14.870000 130.380000 75.000000 130.450000 ;
      RECT 14.870000 140.385000 75.000000 140.455000 ;
      RECT 14.870000 140.385000 75.000000 140.455000 ;
      RECT 14.870000 150.385000 75.000000 150.455000 ;
      RECT 14.870000 150.385000 75.000000 150.455000 ;
      RECT 14.870000 160.385000 75.000000 160.455000 ;
      RECT 14.870000 160.385000 75.000000 160.455000 ;
      RECT 14.870000 170.385000 75.000000 170.455000 ;
      RECT 14.870000 170.385000 75.000000 170.455000 ;
      RECT 14.870000 180.385000 75.000000 180.455000 ;
      RECT 14.870000 180.385000 75.000000 180.455000 ;
      RECT 14.870000 190.385000 75.000000 190.455000 ;
      RECT 14.870000 190.385000 75.000000 190.455000 ;
      RECT 14.905000  24.425000 64.590000  24.495000 ;
      RECT 14.905000  24.425000 64.590000  24.495000 ;
      RECT 14.915000 134.120000 75.000000 134.190000 ;
      RECT 14.915000 134.120000 75.000000 134.190000 ;
      RECT 14.915000 144.120000 75.000000 144.190000 ;
      RECT 14.915000 144.120000 75.000000 144.190000 ;
      RECT 14.915000 154.120000 75.000000 154.190000 ;
      RECT 14.915000 154.120000 75.000000 154.190000 ;
      RECT 14.915000 164.120000 75.000000 164.190000 ;
      RECT 14.915000 164.120000 75.000000 164.190000 ;
      RECT 14.915000 174.120000 75.000000 174.190000 ;
      RECT 14.915000 174.120000 75.000000 174.190000 ;
      RECT 14.915000 184.120000 75.000000 184.190000 ;
      RECT 14.915000 184.120000 75.000000 184.190000 ;
      RECT 14.940000 130.450000 75.000000 130.520000 ;
      RECT 14.940000 130.450000 75.000000 130.520000 ;
      RECT 14.940000 140.455000 75.000000 140.525000 ;
      RECT 14.940000 140.455000 75.000000 140.525000 ;
      RECT 14.940000 150.455000 75.000000 150.525000 ;
      RECT 14.940000 150.455000 75.000000 150.525000 ;
      RECT 14.940000 160.455000 75.000000 160.525000 ;
      RECT 14.940000 160.455000 75.000000 160.525000 ;
      RECT 14.940000 170.455000 75.000000 170.525000 ;
      RECT 14.940000 170.455000 75.000000 170.525000 ;
      RECT 14.940000 180.455000 75.000000 180.525000 ;
      RECT 14.940000 180.455000 75.000000 180.525000 ;
      RECT 14.940000 190.455000 75.000000 190.525000 ;
      RECT 14.940000 190.455000 75.000000 190.525000 ;
      RECT 14.975000  24.355000 64.520000  24.425000 ;
      RECT 14.975000  24.355000 64.520000  24.425000 ;
      RECT 14.985000 134.050000 75.000000 134.120000 ;
      RECT 14.985000 134.050000 75.000000 134.120000 ;
      RECT 14.985000 144.050000 75.000000 144.120000 ;
      RECT 14.985000 144.050000 75.000000 144.120000 ;
      RECT 14.985000 154.050000 75.000000 154.120000 ;
      RECT 14.985000 154.050000 75.000000 154.120000 ;
      RECT 14.985000 164.050000 75.000000 164.120000 ;
      RECT 14.985000 164.050000 75.000000 164.120000 ;
      RECT 14.985000 174.050000 75.000000 174.120000 ;
      RECT 14.985000 174.050000 75.000000 174.120000 ;
      RECT 14.985000 184.050000 75.000000 184.120000 ;
      RECT 14.985000 184.050000 75.000000 184.120000 ;
      RECT 15.010000 130.520000 75.000000 130.590000 ;
      RECT 15.010000 130.520000 75.000000 130.590000 ;
      RECT 15.010000 140.525000 75.000000 140.595000 ;
      RECT 15.010000 140.525000 75.000000 140.595000 ;
      RECT 15.010000 150.525000 75.000000 150.595000 ;
      RECT 15.010000 150.525000 75.000000 150.595000 ;
      RECT 15.010000 160.525000 75.000000 160.595000 ;
      RECT 15.010000 160.525000 75.000000 160.595000 ;
      RECT 15.010000 170.525000 75.000000 170.595000 ;
      RECT 15.010000 170.525000 75.000000 170.595000 ;
      RECT 15.010000 180.525000 75.000000 180.595000 ;
      RECT 15.010000 180.525000 75.000000 180.595000 ;
      RECT 15.010000 190.525000 75.000000 190.595000 ;
      RECT 15.010000 190.525000 75.000000 190.595000 ;
      RECT 15.045000  24.285000 64.450000  24.355000 ;
      RECT 15.045000  24.285000 64.450000  24.355000 ;
      RECT 15.055000 133.980000 75.000000 134.050000 ;
      RECT 15.055000 133.980000 75.000000 134.050000 ;
      RECT 15.055000 143.980000 75.000000 144.050000 ;
      RECT 15.055000 143.980000 75.000000 144.050000 ;
      RECT 15.055000 153.980000 75.000000 154.050000 ;
      RECT 15.055000 153.980000 75.000000 154.050000 ;
      RECT 15.055000 163.980000 75.000000 164.050000 ;
      RECT 15.055000 163.980000 75.000000 164.050000 ;
      RECT 15.055000 173.980000 75.000000 174.050000 ;
      RECT 15.055000 173.980000 75.000000 174.050000 ;
      RECT 15.055000 183.980000 75.000000 184.050000 ;
      RECT 15.055000 183.980000 75.000000 184.050000 ;
      RECT 15.080000 130.590000 75.000000 130.660000 ;
      RECT 15.080000 130.590000 75.000000 130.660000 ;
      RECT 15.080000 140.595000 75.000000 140.665000 ;
      RECT 15.080000 140.595000 75.000000 140.665000 ;
      RECT 15.080000 150.595000 75.000000 150.665000 ;
      RECT 15.080000 150.595000 75.000000 150.665000 ;
      RECT 15.080000 160.595000 75.000000 160.665000 ;
      RECT 15.080000 160.595000 75.000000 160.665000 ;
      RECT 15.080000 170.595000 75.000000 170.665000 ;
      RECT 15.080000 170.595000 75.000000 170.665000 ;
      RECT 15.080000 180.595000 75.000000 180.665000 ;
      RECT 15.080000 180.595000 75.000000 180.665000 ;
      RECT 15.080000 190.595000 75.000000 190.665000 ;
      RECT 15.080000 190.595000 75.000000 190.665000 ;
      RECT 15.115000  24.215000 64.380000  24.285000 ;
      RECT 15.115000  24.215000 64.380000  24.285000 ;
      RECT 15.125000 130.660000 75.000000 130.705000 ;
      RECT 15.125000 130.660000 75.000000 130.705000 ;
      RECT 15.125000 133.910000 75.000000 133.980000 ;
      RECT 15.125000 133.910000 75.000000 133.980000 ;
      RECT 15.125000 133.910000 75.000000 134.795000 ;
      RECT 15.125000 140.665000 75.000000 140.710000 ;
      RECT 15.125000 140.665000 75.000000 140.710000 ;
      RECT 15.125000 143.910000 75.000000 143.980000 ;
      RECT 15.125000 143.910000 75.000000 143.980000 ;
      RECT 15.125000 143.910000 75.000000 144.795000 ;
      RECT 15.125000 150.665000 75.000000 150.710000 ;
      RECT 15.125000 150.665000 75.000000 150.710000 ;
      RECT 15.125000 153.910000 75.000000 153.980000 ;
      RECT 15.125000 153.910000 75.000000 153.980000 ;
      RECT 15.125000 153.910000 75.000000 154.795000 ;
      RECT 15.125000 160.665000 75.000000 160.710000 ;
      RECT 15.125000 160.665000 75.000000 160.710000 ;
      RECT 15.125000 163.910000 75.000000 163.980000 ;
      RECT 15.125000 163.910000 75.000000 163.980000 ;
      RECT 15.125000 163.910000 75.000000 164.795000 ;
      RECT 15.125000 170.665000 75.000000 170.710000 ;
      RECT 15.125000 170.665000 75.000000 170.710000 ;
      RECT 15.125000 173.910000 75.000000 173.980000 ;
      RECT 15.125000 173.910000 75.000000 173.980000 ;
      RECT 15.125000 173.910000 75.000000 174.795000 ;
      RECT 15.125000 180.665000 75.000000 180.710000 ;
      RECT 15.125000 180.665000 75.000000 180.710000 ;
      RECT 15.125000 183.910000 75.000000 183.980000 ;
      RECT 15.125000 183.910000 75.000000 183.980000 ;
      RECT 15.125000 183.910000 75.000000 184.795000 ;
      RECT 15.125000 190.665000 75.000000 190.710000 ;
      RECT 15.125000 190.665000 75.000000 190.710000 ;
      RECT 15.185000  24.145000 64.310000  24.215000 ;
      RECT 15.185000  24.145000 64.310000  24.215000 ;
      RECT 15.255000  24.075000 64.240000  24.145000 ;
      RECT 15.255000  24.075000 64.240000  24.145000 ;
      RECT 15.325000  24.005000 64.170000  24.075000 ;
      RECT 15.325000  24.005000 64.170000  24.075000 ;
      RECT 15.395000  23.935000 64.100000  24.005000 ;
      RECT 15.395000  23.935000 64.100000  24.005000 ;
      RECT 15.465000  23.865000 64.030000  23.935000 ;
      RECT 15.465000  23.865000 64.030000  23.935000 ;
      RECT 15.520000 130.705000 75.000000 130.845000 ;
      RECT 15.520000 140.710000 75.000000 140.850000 ;
      RECT 15.520000 150.710000 75.000000 150.850000 ;
      RECT 15.520000 160.710000 75.000000 160.850000 ;
      RECT 15.520000 170.710000 75.000000 170.850000 ;
      RECT 15.520000 180.710000 75.000000 180.850000 ;
      RECT 15.520000 190.710000 75.000000 190.850000 ;
      RECT 15.535000  23.795000 63.960000  23.865000 ;
      RECT 15.535000  23.795000 63.960000  23.865000 ;
      RECT 15.605000  23.725000 63.890000  23.795000 ;
      RECT 15.605000  23.725000 63.890000  23.795000 ;
      RECT 15.660000 133.770000 75.000000 133.910000 ;
      RECT 15.660000 143.770000 75.000000 143.910000 ;
      RECT 15.660000 153.770000 75.000000 153.910000 ;
      RECT 15.660000 163.770000 75.000000 163.910000 ;
      RECT 15.660000 173.770000 75.000000 173.910000 ;
      RECT 15.660000 183.770000 75.000000 183.910000 ;
      RECT 15.675000  23.655000 63.820000  23.725000 ;
      RECT 15.675000  23.655000 63.820000  23.725000 ;
      RECT 15.745000  23.585000 63.750000  23.655000 ;
      RECT 15.745000  23.585000 63.750000  23.655000 ;
      RECT 15.815000  23.515000 63.680000  23.585000 ;
      RECT 15.815000  23.515000 63.680000  23.585000 ;
      RECT 15.885000  23.445000 63.610000  23.515000 ;
      RECT 15.885000  23.445000 63.610000  23.515000 ;
      RECT 15.955000  23.375000 63.540000  23.445000 ;
      RECT 15.955000  23.375000 63.540000  23.445000 ;
      RECT 16.025000  23.305000 63.470000  23.375000 ;
      RECT 16.025000  23.305000 63.470000  23.375000 ;
      RECT 16.095000  23.235000 63.400000  23.305000 ;
      RECT 16.095000  23.235000 63.400000  23.305000 ;
      RECT 16.165000  23.165000 63.330000  23.235000 ;
      RECT 16.165000  23.165000 63.330000  23.235000 ;
      RECT 16.235000  23.095000 63.260000  23.165000 ;
      RECT 16.235000  23.095000 63.260000  23.165000 ;
      RECT 16.305000  23.025000 63.190000  23.095000 ;
      RECT 16.305000  23.025000 63.190000  23.095000 ;
      RECT 16.375000  22.955000 63.120000  23.025000 ;
      RECT 16.375000  22.955000 63.120000  23.025000 ;
      RECT 16.445000  22.885000 63.050000  22.955000 ;
      RECT 16.445000  22.885000 63.050000  22.955000 ;
      RECT 16.515000  22.815000 62.980000  22.885000 ;
      RECT 16.515000  22.815000 62.980000  22.885000 ;
      RECT 16.585000  22.745000 62.910000  22.815000 ;
      RECT 16.585000  22.745000 62.910000  22.815000 ;
      RECT 16.655000  22.675000 62.840000  22.745000 ;
      RECT 16.655000  22.675000 62.840000  22.745000 ;
      RECT 16.725000  22.605000 62.770000  22.675000 ;
      RECT 16.725000  22.605000 62.770000  22.675000 ;
      RECT 16.795000  22.535000 62.700000  22.605000 ;
      RECT 16.795000  22.535000 62.700000  22.605000 ;
      RECT 16.865000  22.465000 62.630000  22.535000 ;
      RECT 16.865000  22.465000 62.630000  22.535000 ;
      RECT 16.935000  22.395000 62.560000  22.465000 ;
      RECT 16.935000  22.395000 62.560000  22.465000 ;
      RECT 17.005000  22.325000 62.490000  22.395000 ;
      RECT 17.005000  22.325000 62.490000  22.395000 ;
      RECT 17.075000  22.255000 62.420000  22.325000 ;
      RECT 17.075000  22.255000 62.420000  22.325000 ;
      RECT 17.140000   5.235000 17.350000   9.250000 ;
      RECT 17.140000   5.235000 17.490000   9.250000 ;
      RECT 17.140000   9.250000 17.490000   9.600000 ;
      RECT 17.145000  22.185000 62.350000  22.255000 ;
      RECT 17.145000  22.185000 62.350000  22.255000 ;
      RECT 17.210000   5.165000 17.350000   5.235000 ;
      RECT 17.210000   9.250000 17.350000   9.320000 ;
      RECT 17.215000  22.115000 62.280000  22.185000 ;
      RECT 17.215000  22.115000 62.280000  22.185000 ;
      RECT 17.280000   5.095000 17.350000   5.165000 ;
      RECT 17.280000   9.320000 17.350000   9.390000 ;
      RECT 17.285000  22.045000 62.210000  22.115000 ;
      RECT 17.285000  22.045000 62.210000  22.115000 ;
      RECT 17.320000   5.055000 17.490000   5.235000 ;
      RECT 17.355000  21.975000 62.140000  22.045000 ;
      RECT 17.355000  21.975000 62.140000  22.045000 ;
      RECT 17.425000  21.905000 53.815000  21.975000 ;
      RECT 17.425000  21.905000 53.815000  21.975000 ;
      RECT 17.495000  21.835000 53.815000  21.905000 ;
      RECT 17.495000  21.835000 53.815000  21.905000 ;
      RECT 17.495000  21.835000 65.660000  25.300000 ;
      RECT 17.565000  21.765000 53.815000  21.835000 ;
      RECT 17.565000  21.765000 53.815000  21.835000 ;
      RECT 17.570000   9.680000 55.880000   9.800000 ;
      RECT 17.635000  21.695000 53.815000  21.765000 ;
      RECT 17.635000  21.695000 53.815000  21.765000 ;
      RECT 17.705000  21.625000 53.815000  21.695000 ;
      RECT 17.705000  21.625000 53.815000  21.695000 ;
      RECT 17.775000  21.555000 53.815000  21.625000 ;
      RECT 17.775000  21.555000 53.815000  21.625000 ;
      RECT 17.845000  21.485000 53.815000  21.555000 ;
      RECT 17.845000  21.485000 53.815000  21.555000 ;
      RECT 17.915000  21.415000 53.815000  21.485000 ;
      RECT 17.915000  21.415000 53.815000  21.485000 ;
      RECT 17.985000  21.345000 53.815000  21.415000 ;
      RECT 17.985000  21.345000 53.815000  21.415000 ;
      RECT 18.055000  21.275000 53.815000  21.345000 ;
      RECT 18.055000  21.275000 53.815000  21.345000 ;
      RECT 18.125000  21.205000 53.815000  21.275000 ;
      RECT 18.125000  21.205000 53.815000  21.275000 ;
      RECT 18.195000  21.135000 53.815000  21.205000 ;
      RECT 18.195000  21.135000 53.815000  21.205000 ;
      RECT 18.265000  21.065000 53.815000  21.135000 ;
      RECT 18.265000  21.065000 53.815000  21.135000 ;
      RECT 18.335000  20.995000 53.815000  21.065000 ;
      RECT 18.335000  20.995000 53.815000  21.065000 ;
      RECT 18.405000  20.925000 53.815000  20.995000 ;
      RECT 18.405000  20.925000 53.815000  20.995000 ;
      RECT 18.475000  20.855000 53.815000  20.925000 ;
      RECT 18.475000  20.855000 53.815000  20.925000 ;
      RECT 18.545000  20.785000 53.815000  20.855000 ;
      RECT 18.545000  20.785000 53.815000  20.855000 ;
      RECT 18.580000 193.770000 75.000000 193.910000 ;
      RECT 18.615000  20.715000 53.815000  20.785000 ;
      RECT 18.615000  20.715000 53.815000  20.785000 ;
      RECT 18.685000  20.645000 53.815000  20.715000 ;
      RECT 18.685000  20.645000 53.815000  20.715000 ;
      RECT 18.755000  20.575000 53.815000  20.645000 ;
      RECT 18.755000  20.575000 53.815000  20.645000 ;
      RECT 18.825000  20.505000 53.815000  20.575000 ;
      RECT 18.825000  20.505000 53.815000  20.575000 ;
      RECT 18.895000  20.435000 53.815000  20.505000 ;
      RECT 18.895000  20.435000 53.815000  20.505000 ;
      RECT 18.965000  20.365000 53.815000  20.435000 ;
      RECT 18.965000  20.365000 53.815000  20.435000 ;
      RECT 19.035000  20.295000 53.815000  20.365000 ;
      RECT 19.035000  20.295000 53.815000  20.365000 ;
      RECT 19.105000  20.225000 53.815000  20.295000 ;
      RECT 19.105000  20.225000 53.815000  20.295000 ;
      RECT 19.175000  20.155000 53.815000  20.225000 ;
      RECT 19.175000  20.155000 53.815000  20.225000 ;
      RECT 19.245000  20.085000 53.815000  20.155000 ;
      RECT 19.245000  20.085000 53.815000  20.155000 ;
      RECT 19.315000  20.015000 53.815000  20.085000 ;
      RECT 19.315000  20.015000 53.815000  20.085000 ;
      RECT 19.385000  19.945000 53.815000  20.015000 ;
      RECT 19.385000  19.945000 53.815000  20.015000 ;
      RECT 19.400000  19.930000 53.955000  21.835000 ;
      RECT 19.455000  19.875000 53.815000  19.945000 ;
      RECT 19.455000  19.875000 53.815000  19.945000 ;
      RECT 19.510000  19.820000 53.815000  19.875000 ;
      RECT 19.510000  19.820000 53.815000  19.875000 ;
      RECT 19.580000  19.750000 53.870000  19.820000 ;
      RECT 19.580000  19.750000 53.870000  19.820000 ;
      RECT 19.650000  19.680000 53.940000  19.750000 ;
      RECT 19.650000  19.680000 53.940000  19.750000 ;
      RECT 19.720000  19.610000 54.010000  19.680000 ;
      RECT 19.720000  19.610000 54.010000  19.680000 ;
      RECT 19.790000  19.540000 54.080000  19.610000 ;
      RECT 19.790000  19.540000 54.080000  19.610000 ;
      RECT 19.860000  19.470000 54.150000  19.540000 ;
      RECT 19.860000  19.470000 54.150000  19.540000 ;
      RECT 19.930000  19.400000 54.220000  19.470000 ;
      RECT 19.930000  19.400000 54.220000  19.470000 ;
      RECT 20.000000  19.330000 54.290000  19.400000 ;
      RECT 20.000000  19.330000 54.290000  19.400000 ;
      RECT 20.070000  19.260000 54.360000  19.330000 ;
      RECT 20.070000  19.260000 54.360000  19.330000 ;
      RECT 20.140000  19.190000 54.430000  19.260000 ;
      RECT 20.140000  19.190000 54.430000  19.260000 ;
      RECT 20.210000  19.120000 54.500000  19.190000 ;
      RECT 20.210000  19.120000 54.500000  19.190000 ;
      RECT 20.280000  19.050000 54.570000  19.120000 ;
      RECT 20.280000  19.050000 54.570000  19.120000 ;
      RECT 20.350000  18.980000 54.640000  19.050000 ;
      RECT 20.350000  18.980000 54.640000  19.050000 ;
      RECT 20.420000  18.910000 54.710000  18.980000 ;
      RECT 20.420000  18.910000 54.710000  18.980000 ;
      RECT 20.490000  18.840000 54.780000  18.910000 ;
      RECT 20.490000  18.840000 54.780000  18.910000 ;
      RECT 20.560000  18.770000 54.850000  18.840000 ;
      RECT 20.560000  18.770000 54.850000  18.840000 ;
      RECT 20.630000  18.700000 54.920000  18.770000 ;
      RECT 20.630000  18.700000 54.920000  18.770000 ;
      RECT 20.700000  18.630000 54.990000  18.700000 ;
      RECT 20.700000  18.630000 54.990000  18.700000 ;
      RECT 20.770000  18.560000 55.060000  18.630000 ;
      RECT 20.770000  18.560000 55.060000  18.630000 ;
      RECT 20.775000   0.000000 20.785000   1.600000 ;
      RECT 20.775000   1.600000 20.785000   1.760000 ;
      RECT 20.840000  18.490000 55.130000  18.560000 ;
      RECT 20.840000  18.490000 55.130000  18.560000 ;
      RECT 20.910000  18.420000 55.200000  18.490000 ;
      RECT 20.910000  18.420000 55.200000  18.490000 ;
      RECT 20.980000  18.350000 55.270000  18.420000 ;
      RECT 20.980000  18.350000 55.270000  18.420000 ;
      RECT 21.050000  18.280000 55.340000  18.350000 ;
      RECT 21.050000  18.280000 55.340000  18.350000 ;
      RECT 21.120000  18.210000 55.410000  18.280000 ;
      RECT 21.120000  18.210000 55.410000  18.280000 ;
      RECT 21.190000  18.140000 55.480000  18.210000 ;
      RECT 21.190000  18.140000 55.480000  18.210000 ;
      RECT 21.260000  18.070000 55.550000  18.140000 ;
      RECT 21.260000  18.070000 55.550000  18.140000 ;
      RECT 21.330000  18.000000 55.620000  18.070000 ;
      RECT 21.330000  18.000000 55.620000  18.070000 ;
      RECT 21.400000  17.930000 55.690000  18.000000 ;
      RECT 21.400000  17.930000 55.690000  18.000000 ;
      RECT 21.470000  17.860000 55.760000  17.930000 ;
      RECT 21.470000  17.860000 55.760000  17.930000 ;
      RECT 21.540000  17.790000 55.830000  17.860000 ;
      RECT 21.540000  17.790000 55.830000  17.860000 ;
      RECT 21.555000  17.775000 53.955000  19.930000 ;
      RECT 21.610000  17.720000 55.900000  17.790000 ;
      RECT 21.610000  17.720000 55.900000  17.790000 ;
      RECT 21.620000  17.710000 55.970000  17.720000 ;
      RECT 21.620000  17.710000 55.970000  17.720000 ;
      RECT 21.690000  17.640000 55.970000  17.710000 ;
      RECT 21.690000  17.640000 55.970000  17.710000 ;
      RECT 21.760000  17.570000 55.970000  17.640000 ;
      RECT 21.760000  17.570000 55.970000  17.640000 ;
      RECT 21.830000  17.500000 55.970000  17.570000 ;
      RECT 21.830000  17.500000 55.970000  17.570000 ;
      RECT 21.900000  17.430000 55.970000  17.500000 ;
      RECT 21.900000  17.430000 55.970000  17.500000 ;
      RECT 21.970000  17.360000 55.970000  17.430000 ;
      RECT 21.970000  17.360000 55.970000  17.430000 ;
      RECT 21.970000  17.360000 56.110000  17.775000 ;
      RECT 53.675000   0.000000 53.955000   7.875000 ;
      RECT 53.675000   7.875000 55.760000   9.680000 ;
      RECT 53.815000   8.000000 53.885000   8.070000 ;
      RECT 53.815000   8.070000 53.955000   8.140000 ;
      RECT 53.815000   8.140000 54.025000   8.210000 ;
      RECT 53.815000   8.210000 54.095000   8.280000 ;
      RECT 53.815000   8.280000 54.165000   8.350000 ;
      RECT 53.815000   8.350000 54.235000   8.420000 ;
      RECT 53.815000   8.420000 54.305000   8.490000 ;
      RECT 53.815000   8.490000 54.375000   8.560000 ;
      RECT 53.815000   8.560000 54.445000   8.630000 ;
      RECT 53.815000   8.630000 54.515000   8.700000 ;
      RECT 53.815000   8.700000 54.585000   8.770000 ;
      RECT 53.815000   8.770000 54.655000   8.840000 ;
      RECT 53.815000   8.840000 54.725000   8.910000 ;
      RECT 53.815000   8.910000 54.795000   8.980000 ;
      RECT 53.815000   8.980000 54.865000   9.050000 ;
      RECT 53.815000   9.050000 54.935000   9.120000 ;
      RECT 53.815000   9.120000 55.005000   9.190000 ;
      RECT 53.815000   9.190000 55.075000   9.260000 ;
      RECT 53.815000   9.260000 55.145000   9.330000 ;
      RECT 53.815000   9.330000 55.215000   9.400000 ;
      RECT 53.815000   9.400000 55.285000   9.470000 ;
      RECT 53.815000   9.470000 55.355000   9.540000 ;
      RECT 53.815000   9.540000 55.425000   9.610000 ;
      RECT 53.815000   9.610000 55.495000   9.680000 ;
      RECT 53.815000   9.680000 55.565000   9.750000 ;
      RECT 53.815000   9.750000 55.635000   9.800000 ;
      RECT 55.875000   9.800000 56.110000  10.030000 ;
      RECT 55.875000  10.030000 56.110000  17.360000 ;
      RECT 68.150000  74.490000 75.000000  98.700000 ;
      RECT 68.150000 130.845000 75.000000 133.770000 ;
      RECT 68.150000 140.850000 75.000000 143.770000 ;
      RECT 68.150000 150.850000 75.000000 153.770000 ;
      RECT 68.150000 160.850000 75.000000 163.770000 ;
      RECT 68.150000 170.850000 75.000000 173.770000 ;
      RECT 68.150000 180.850000 75.000000 183.770000 ;
      RECT 68.150000 190.850000 75.000000 193.770000 ;
      RECT 68.290000  74.545000 75.000000  98.840000 ;
      RECT 68.290000 130.705000 75.000000 133.910000 ;
      RECT 68.290000 140.710000 75.000000 143.910000 ;
      RECT 68.290000 150.710000 75.000000 153.910000 ;
      RECT 68.290000 160.710000 75.000000 163.910000 ;
      RECT 68.290000 170.710000 75.000000 173.910000 ;
      RECT 68.290000 180.710000 75.000000 183.910000 ;
      RECT 68.290000 190.710000 75.000000 193.910000 ;
      RECT 68.295000  74.540000 75.000000  74.545000 ;
      RECT 68.295000  74.540000 75.000000  74.545000 ;
      RECT 68.365000  74.470000 75.000000  74.540000 ;
      RECT 68.365000  74.470000 75.000000  74.540000 ;
      RECT 68.435000  74.400000 75.000000  74.470000 ;
      RECT 68.435000  74.400000 75.000000  74.470000 ;
      RECT 68.505000  74.330000 75.000000  74.400000 ;
      RECT 68.505000  74.330000 75.000000  74.400000 ;
      RECT 68.575000  74.260000 75.000000  74.330000 ;
      RECT 68.575000  74.260000 75.000000  74.330000 ;
      RECT 68.645000  74.190000 75.000000  74.260000 ;
      RECT 68.645000  74.190000 75.000000  74.260000 ;
      RECT 68.715000  74.120000 75.000000  74.190000 ;
      RECT 68.715000  74.120000 75.000000  74.190000 ;
      RECT 68.785000  74.050000 75.000000  74.120000 ;
      RECT 68.785000  74.050000 75.000000  74.120000 ;
      RECT 68.855000  73.980000 75.000000  74.050000 ;
      RECT 68.855000  73.980000 75.000000  74.050000 ;
      RECT 68.865000  73.770000 75.000000  74.490000 ;
      RECT 68.925000  73.910000 75.000000  73.980000 ;
      RECT 68.925000  73.910000 75.000000  73.980000 ;
      RECT 74.840000   0.000000 75.000000  73.770000 ;
    LAYER met3 ;
      RECT  0.000000   0.000000  0.200000 171.495000 ;
      RECT  0.000000 171.495000 15.205000 189.915000 ;
      RECT  0.000000 171.595000 15.205000 189.915000 ;
      RECT  0.000000 171.595000 15.205000 198.000000 ;
      RECT  0.000000 189.915000 75.000000 198.000000 ;
      RECT  0.000000 189.915000 75.000000 198.000000 ;
      RECT 13.200000  94.385000 15.205000 171.495000 ;
      RECT 13.300000  94.425000 15.205000 171.595000 ;
      RECT 13.440000  94.145000 15.205000  94.385000 ;
      RECT 13.440000  94.285000 15.205000  94.425000 ;
      RECT 13.580000  94.145000 15.205000  94.285000 ;
      RECT 13.725000  94.000000 15.205000  94.145000 ;
      RECT 13.875000  93.850000 15.350000  94.000000 ;
      RECT 14.025000  93.700000 15.500000  93.850000 ;
      RECT 14.175000  93.550000 15.650000  93.700000 ;
      RECT 14.325000  93.400000 15.800000  93.550000 ;
      RECT 14.475000  93.250000 15.950000  93.400000 ;
      RECT 14.625000  93.100000 16.100000  93.250000 ;
      RECT 14.775000  92.950000 16.250000  93.100000 ;
      RECT 14.925000  92.800000 16.400000  92.950000 ;
      RECT 15.075000  92.650000 16.550000  92.800000 ;
      RECT 15.225000  92.500000 16.700000  92.650000 ;
      RECT 15.375000  92.350000 16.850000  92.500000 ;
      RECT 15.525000  92.200000 17.000000  92.350000 ;
      RECT 15.675000  92.050000 17.150000  92.200000 ;
      RECT 15.825000  91.900000 17.300000  92.050000 ;
      RECT 15.975000  91.750000 17.450000  91.900000 ;
      RECT 16.125000  91.600000 17.600000  91.750000 ;
      RECT 16.275000  91.450000 17.750000  91.600000 ;
      RECT 16.425000  91.300000 17.900000  91.450000 ;
      RECT 16.575000  91.150000 18.050000  91.300000 ;
      RECT 16.725000  91.000000 18.200000  91.150000 ;
      RECT 16.875000  90.850000 18.350000  91.000000 ;
      RECT 17.025000  90.700000 18.500000  90.850000 ;
      RECT 17.175000  90.550000 18.650000  90.700000 ;
      RECT 17.325000  90.400000 18.800000  90.550000 ;
      RECT 17.475000  90.250000 18.950000  90.400000 ;
      RECT 17.625000  90.100000 19.100000  90.250000 ;
      RECT 17.775000  89.950000 19.250000  90.100000 ;
      RECT 17.925000  89.800000 19.400000  89.950000 ;
      RECT 18.075000  89.650000 19.550000  89.800000 ;
      RECT 18.225000  89.500000 19.700000  89.650000 ;
      RECT 18.375000  89.350000 19.850000  89.500000 ;
      RECT 18.525000  89.200000 20.000000  89.350000 ;
      RECT 18.675000  89.050000 20.150000  89.200000 ;
      RECT 18.825000  88.900000 20.300000  89.050000 ;
      RECT 18.975000  88.750000 20.450000  88.900000 ;
      RECT 19.125000  88.600000 20.600000  88.750000 ;
      RECT 19.275000  88.450000 20.750000  88.600000 ;
      RECT 19.425000  88.300000 20.900000  88.450000 ;
      RECT 19.575000  88.150000 21.050000  88.300000 ;
      RECT 19.725000  88.000000 21.200000  88.150000 ;
      RECT 19.875000  87.850000 21.350000  88.000000 ;
      RECT 20.025000  87.700000 21.500000  87.850000 ;
      RECT 20.175000  87.550000 21.650000  87.700000 ;
      RECT 20.325000  87.400000 21.800000  87.550000 ;
      RECT 20.475000  87.250000 21.950000  87.400000 ;
      RECT 20.625000  87.100000 22.100000  87.250000 ;
      RECT 20.775000  86.950000 22.250000  87.100000 ;
      RECT 20.925000  86.800000 22.400000  86.950000 ;
      RECT 21.075000  86.650000 22.550000  86.800000 ;
      RECT 21.225000  86.500000 22.700000  86.650000 ;
      RECT 21.375000  86.350000 22.850000  86.500000 ;
      RECT 21.525000  86.200000 23.000000  86.350000 ;
      RECT 21.675000  86.050000 23.150000  86.200000 ;
      RECT 21.825000  85.900000 23.300000  86.050000 ;
      RECT 21.950000  85.775000 23.450000  85.900000 ;
      RECT 22.005000  96.955000 25.635000 166.935000 ;
      RECT 22.005000  96.955000 25.635000 166.935000 ;
      RECT 22.005000 166.935000 25.635000 170.445000 ;
      RECT 22.075000  96.885000 25.635000  96.955000 ;
      RECT 22.100000  85.625000 23.450000  85.775000 ;
      RECT 22.155000 166.935000 25.635000 167.085000 ;
      RECT 22.225000  96.735000 25.635000  96.885000 ;
      RECT 22.250000  85.475000 23.450000  85.625000 ;
      RECT 22.305000 167.085000 25.635000 167.235000 ;
      RECT 22.375000  96.585000 25.635000  96.735000 ;
      RECT 22.400000  85.325000 23.450000  85.475000 ;
      RECT 22.455000 167.235000 25.635000 167.385000 ;
      RECT 22.525000  96.435000 25.635000  96.585000 ;
      RECT 22.550000  85.175000 23.450000  85.325000 ;
      RECT 22.605000 167.385000 25.635000 167.535000 ;
      RECT 22.675000  96.285000 25.635000  96.435000 ;
      RECT 22.700000  85.025000 23.450000  85.175000 ;
      RECT 22.755000 167.535000 25.635000 167.685000 ;
      RECT 22.825000  96.135000 25.635000  96.285000 ;
      RECT 22.850000  84.875000 23.450000  85.025000 ;
      RECT 22.905000 167.685000 25.635000 167.835000 ;
      RECT 22.975000  95.985000 25.635000  96.135000 ;
      RECT 23.000000  84.725000 23.450000  84.875000 ;
      RECT 23.055000 167.835000 25.635000 167.985000 ;
      RECT 23.100000  84.485000 23.450000  85.900000 ;
      RECT 23.125000  95.835000 25.635000  95.985000 ;
      RECT 23.150000  84.575000 23.450000  84.725000 ;
      RECT 23.205000 167.985000 25.635000 168.135000 ;
      RECT 23.275000  95.685000 25.635000  95.835000 ;
      RECT 23.300000  84.425000 23.450000  84.575000 ;
      RECT 23.355000 168.135000 25.635000 168.285000 ;
      RECT 23.425000  95.535000 25.635000  95.685000 ;
      RECT 23.505000 168.285000 25.635000 168.435000 ;
      RECT 23.575000  95.385000 25.635000  95.535000 ;
      RECT 23.655000 168.435000 25.635000 168.585000 ;
      RECT 23.725000  95.235000 25.635000  95.385000 ;
      RECT 23.805000 168.585000 25.635000 168.735000 ;
      RECT 23.875000  95.085000 25.635000  95.235000 ;
      RECT 23.955000 168.735000 25.635000 168.885000 ;
      RECT 24.025000  94.935000 25.635000  95.085000 ;
      RECT 24.105000 168.885000 25.635000 169.035000 ;
      RECT 24.175000  94.785000 25.635000  94.935000 ;
      RECT 24.255000 169.035000 25.635000 169.185000 ;
      RECT 24.325000  94.635000 25.635000  94.785000 ;
      RECT 24.405000 169.185000 25.635000 169.335000 ;
      RECT 24.475000  94.485000 25.635000  94.635000 ;
      RECT 24.555000 169.335000 25.635000 169.485000 ;
      RECT 24.625000  94.335000 25.635000  94.485000 ;
      RECT 24.625000  94.335000 25.635000  96.955000 ;
      RECT 24.705000 169.485000 25.635000 169.635000 ;
      RECT 24.745000  94.215000 25.635000  94.335000 ;
      RECT 24.800000   0.000000 25.600000  82.335000 ;
      RECT 24.800000  82.335000 25.150000  82.785000 ;
      RECT 24.855000 169.635000 25.635000 169.785000 ;
      RECT 24.895000  94.065000 25.755000  94.215000 ;
      RECT 24.900000   0.000000 25.600000  82.335000 ;
      RECT 24.900000  82.335000 25.450000  82.485000 ;
      RECT 24.900000  82.485000 25.300000  82.635000 ;
      RECT 24.900000  82.635000 25.150000  82.785000 ;
      RECT 24.900000  82.785000 25.000000  82.935000 ;
      RECT 25.005000 169.785000 25.635000 169.935000 ;
      RECT 25.045000  93.915000 25.905000  94.065000 ;
      RECT 25.155000 169.935000 25.635000 170.085000 ;
      RECT 25.195000  93.765000 26.055000  93.915000 ;
      RECT 25.305000 170.085000 25.635000 170.235000 ;
      RECT 25.345000  93.615000 26.205000  93.765000 ;
      RECT 25.455000 170.235000 25.635000 170.385000 ;
      RECT 25.495000  93.465000 26.355000  93.615000 ;
      RECT 25.515000 170.445000 25.635000 189.915000 ;
      RECT 25.605000 170.385000 25.635000 170.535000 ;
      RECT 25.645000  93.315000 26.505000  93.465000 ;
      RECT 25.795000  93.165000 26.655000  93.315000 ;
      RECT 25.945000  93.015000 26.805000  93.165000 ;
      RECT 26.095000  92.865000 26.955000  93.015000 ;
      RECT 26.245000  92.715000 27.105000  92.865000 ;
      RECT 26.395000  92.565000 27.255000  92.715000 ;
      RECT 26.545000  92.415000 27.405000  92.565000 ;
      RECT 26.695000  92.265000 27.555000  92.415000 ;
      RECT 26.845000  92.115000 27.705000  92.265000 ;
      RECT 26.995000  91.965000 27.855000  92.115000 ;
      RECT 27.145000  91.815000 28.005000  91.965000 ;
      RECT 27.295000  91.665000 28.155000  91.815000 ;
      RECT 27.445000  91.515000 28.305000  91.665000 ;
      RECT 27.595000  91.365000 28.455000  91.515000 ;
      RECT 27.745000  91.215000 28.605000  91.365000 ;
      RECT 27.895000  91.065000 28.755000  91.215000 ;
      RECT 28.045000  90.915000 28.905000  91.065000 ;
      RECT 28.195000  90.765000 29.055000  90.915000 ;
      RECT 28.345000  90.615000 29.205000  90.765000 ;
      RECT 28.495000  90.465000 29.355000  90.615000 ;
      RECT 28.645000  90.315000 29.505000  90.465000 ;
      RECT 28.795000  90.165000 29.655000  90.315000 ;
      RECT 28.945000  90.015000 29.805000  90.165000 ;
      RECT 29.095000  89.865000 29.955000  90.015000 ;
      RECT 29.245000  89.715000 30.105000  89.865000 ;
      RECT 29.395000  89.565000 30.255000  89.715000 ;
      RECT 29.545000  89.415000 30.405000  89.565000 ;
      RECT 29.695000  89.265000 30.555000  89.415000 ;
      RECT 29.845000  89.115000 30.705000  89.265000 ;
      RECT 29.995000  88.965000 30.855000  89.115000 ;
      RECT 30.145000  88.815000 31.005000  88.965000 ;
      RECT 30.295000  88.665000 31.155000  88.815000 ;
      RECT 30.445000  88.515000 31.305000  88.665000 ;
      RECT 30.595000  88.365000 31.455000  88.515000 ;
      RECT 30.745000  88.215000 31.605000  88.365000 ;
      RECT 30.895000  88.065000 31.755000  88.215000 ;
      RECT 31.045000  87.915000 31.905000  88.065000 ;
      RECT 31.195000  87.765000 32.055000  87.915000 ;
      RECT 31.345000  87.615000 32.205000  87.765000 ;
      RECT 31.495000  87.465000 32.355000  87.615000 ;
      RECT 31.645000  87.315000 32.505000  87.465000 ;
      RECT 31.795000  87.165000 32.655000  87.315000 ;
      RECT 31.945000  87.015000 32.805000  87.165000 ;
      RECT 32.095000  86.865000 32.955000  87.015000 ;
      RECT 32.245000  86.715000 33.105000  86.865000 ;
      RECT 32.395000  86.565000 33.255000  86.715000 ;
      RECT 32.435000  93.555000 40.410000  93.705000 ;
      RECT 32.435000  93.555000 42.435000  95.580000 ;
      RECT 32.435000  93.705000 40.560000  93.855000 ;
      RECT 32.435000  93.855000 40.710000  94.005000 ;
      RECT 32.435000  94.005000 40.860000  94.155000 ;
      RECT 32.435000  94.155000 41.010000  94.305000 ;
      RECT 32.435000  94.305000 41.160000  94.455000 ;
      RECT 32.435000  94.455000 41.310000  94.605000 ;
      RECT 32.435000  94.605000 41.460000  94.755000 ;
      RECT 32.435000  94.755000 41.610000  94.905000 ;
      RECT 32.435000  94.905000 41.760000  95.055000 ;
      RECT 32.435000  95.055000 41.910000  95.205000 ;
      RECT 32.435000  95.205000 42.060000  95.355000 ;
      RECT 32.435000  95.355000 42.210000  95.505000 ;
      RECT 32.435000  95.505000 42.360000  95.580000 ;
      RECT 32.435000  95.580000 35.440000 159.400000 ;
      RECT 32.435000  95.580000 42.435000 162.405000 ;
      RECT 32.435000 159.400000 36.680000 162.405000 ;
      RECT 32.435000 162.405000 42.435000 163.970000 ;
      RECT 32.515000  93.475000 40.330000  93.555000 ;
      RECT 32.545000  84.855000 34.105000  85.865000 ;
      RECT 32.545000  84.855000 34.105000  85.865000 ;
      RECT 32.545000  85.865000 33.555000  86.415000 ;
      RECT 32.545000  85.865000 33.955000  86.015000 ;
      RECT 32.545000  86.015000 33.805000  86.165000 ;
      RECT 32.545000  86.165000 33.655000  86.315000 ;
      RECT 32.545000  86.315000 33.555000  86.415000 ;
      RECT 32.545000  86.415000 33.405000  86.565000 ;
      RECT 32.570000  84.830000 34.080000  84.855000 ;
      RECT 32.585000 162.405000 42.435000 162.555000 ;
      RECT 32.665000  93.325000 40.180000  93.475000 ;
      RECT 32.720000  84.680000 33.930000  84.830000 ;
      RECT 32.735000 162.555000 42.435000 162.705000 ;
      RECT 32.815000  93.175000 40.030000  93.325000 ;
      RECT 32.870000  84.530000 33.780000  84.680000 ;
      RECT 32.885000 162.705000 42.435000 162.855000 ;
      RECT 32.965000  93.025000 39.880000  93.175000 ;
      RECT 33.020000  84.380000 33.630000  84.530000 ;
      RECT 33.020000  84.380000 34.105000  84.855000 ;
      RECT 33.035000 162.855000 42.435000 163.005000 ;
      RECT 33.115000  92.875000 39.730000  93.025000 ;
      RECT 33.185000 163.005000 42.435000 163.155000 ;
      RECT 33.265000  92.725000 39.580000  92.875000 ;
      RECT 33.335000 163.155000 42.435000 163.305000 ;
      RECT 33.415000  92.575000 39.430000  92.725000 ;
      RECT 33.485000 163.305000 42.435000 163.455000 ;
      RECT 33.565000  92.425000 39.280000  92.575000 ;
      RECT 33.635000 163.455000 42.435000 163.605000 ;
      RECT 33.715000  92.275000 39.130000  92.425000 ;
      RECT 33.785000 163.605000 42.435000 163.755000 ;
      RECT 33.865000  92.125000 38.980000  92.275000 ;
      RECT 33.935000 163.755000 42.435000 163.905000 ;
      RECT 34.000000 163.905000 42.435000 163.970000 ;
      RECT 34.000000 163.970000 39.110000 167.295000 ;
      RECT 34.015000  91.975000 38.830000  92.125000 ;
      RECT 34.150000 163.970000 42.285000 164.120000 ;
      RECT 34.165000  91.825000 38.680000  91.975000 ;
      RECT 34.300000 164.120000 42.135000 164.270000 ;
      RECT 34.315000  91.675000 38.530000  91.825000 ;
      RECT 34.450000 164.270000 41.985000 164.420000 ;
      RECT 34.465000  91.525000 38.380000  91.675000 ;
      RECT 34.600000 164.420000 41.835000 164.570000 ;
      RECT 34.615000  91.375000 38.230000  91.525000 ;
      RECT 34.750000 164.570000 41.685000 164.720000 ;
      RECT 34.765000  91.225000 38.080000  91.375000 ;
      RECT 34.900000 164.720000 41.535000 164.870000 ;
      RECT 34.915000  91.075000 37.930000  91.225000 ;
      RECT 35.050000 164.870000 41.385000 165.020000 ;
      RECT 35.065000  90.925000 37.780000  91.075000 ;
      RECT 35.200000 165.020000 41.235000 165.170000 ;
      RECT 35.215000  90.775000 37.630000  90.925000 ;
      RECT 35.215000  90.775000 40.410000  93.555000 ;
      RECT 35.350000 165.170000 41.085000 165.320000 ;
      RECT 35.435000  94.800000 37.410000  94.950000 ;
      RECT 35.435000  94.800000 37.410000  94.950000 ;
      RECT 35.435000  94.950000 37.560000  95.100000 ;
      RECT 35.435000  94.950000 37.560000  95.100000 ;
      RECT 35.435000  95.100000 37.710000  95.250000 ;
      RECT 35.435000  95.100000 37.710000  95.250000 ;
      RECT 35.435000  95.250000 37.860000  95.400000 ;
      RECT 35.435000  95.250000 37.860000  95.400000 ;
      RECT 35.435000  95.400000 38.010000  95.550000 ;
      RECT 35.435000  95.400000 38.010000  95.550000 ;
      RECT 35.435000  95.550000 38.160000  95.700000 ;
      RECT 35.435000  95.550000 38.160000  95.700000 ;
      RECT 35.435000  95.700000 38.310000  95.850000 ;
      RECT 35.435000  95.700000 38.310000  95.850000 ;
      RECT 35.435000  95.850000 38.460000  96.000000 ;
      RECT 35.435000  95.850000 38.460000  96.000000 ;
      RECT 35.435000  96.000000 38.610000  96.150000 ;
      RECT 35.435000  96.000000 38.610000  96.150000 ;
      RECT 35.435000  96.150000 38.760000  96.300000 ;
      RECT 35.435000  96.150000 38.760000  96.300000 ;
      RECT 35.435000  96.300000 38.910000  96.450000 ;
      RECT 35.435000  96.300000 38.910000  96.450000 ;
      RECT 35.435000  96.450000 39.060000  96.600000 ;
      RECT 35.435000  96.450000 39.060000  96.600000 ;
      RECT 35.435000  96.600000 39.210000  96.750000 ;
      RECT 35.435000  96.600000 39.210000  96.750000 ;
      RECT 35.435000  96.750000 39.360000  96.825000 ;
      RECT 35.435000  96.750000 39.360000  96.825000 ;
      RECT 35.435000  96.825000 39.435000 161.160000 ;
      RECT 35.500000 165.320000 40.935000 165.470000 ;
      RECT 35.520000  94.715000 37.325000  94.800000 ;
      RECT 35.520000  94.715000 37.325000  94.800000 ;
      RECT 35.585000 161.160000 39.435000 161.310000 ;
      RECT 35.585000 161.160000 39.435000 161.310000 ;
      RECT 35.650000 165.470000 40.785000 165.620000 ;
      RECT 35.670000  94.565000 37.175000  94.715000 ;
      RECT 35.670000  94.565000 37.175000  94.715000 ;
      RECT 35.735000 161.310000 39.435000 161.460000 ;
      RECT 35.735000 161.310000 39.435000 161.460000 ;
      RECT 35.800000 165.620000 40.635000 165.770000 ;
      RECT 35.820000  94.415000 37.025000  94.565000 ;
      RECT 35.820000  94.415000 37.025000  94.565000 ;
      RECT 35.885000 161.460000 39.435000 161.610000 ;
      RECT 35.885000 161.460000 39.435000 161.610000 ;
      RECT 35.950000 165.770000 40.485000 165.920000 ;
      RECT 35.975000  94.265000 36.875000  94.415000 ;
      RECT 35.975000  94.265000 36.875000  94.415000 ;
      RECT 36.035000 161.610000 39.435000 161.760000 ;
      RECT 36.035000 161.610000 39.435000 161.760000 ;
      RECT 36.100000 165.920000 40.335000 166.070000 ;
      RECT 36.125000  94.115000 36.725000  94.265000 ;
      RECT 36.125000  94.115000 36.725000  94.265000 ;
      RECT 36.185000 161.760000 39.435000 161.910000 ;
      RECT 36.185000 161.760000 39.435000 161.910000 ;
      RECT 36.250000 166.070000 40.185000 166.220000 ;
      RECT 36.275000  93.965000 36.575000  94.115000 ;
      RECT 36.275000  93.965000 36.575000  94.115000 ;
      RECT 36.335000 161.910000 39.435000 162.060000 ;
      RECT 36.335000 161.910000 39.435000 162.060000 ;
      RECT 36.400000 166.220000 40.035000 166.370000 ;
      RECT 36.485000 162.060000 39.435000 162.210000 ;
      RECT 36.485000 162.060000 39.435000 162.210000 ;
      RECT 36.550000 166.370000 39.885000 166.520000 ;
      RECT 36.635000 162.210000 39.435000 162.360000 ;
      RECT 36.635000 162.210000 39.435000 162.360000 ;
      RECT 36.700000 166.520000 39.735000 166.670000 ;
      RECT 36.785000 162.360000 39.435000 162.510000 ;
      RECT 36.785000 162.360000 39.435000 162.510000 ;
      RECT 36.850000 166.670000 39.585000 166.820000 ;
      RECT 36.935000 162.510000 39.435000 162.660000 ;
      RECT 36.935000 162.510000 39.435000 162.660000 ;
      RECT 37.000000 162.660000 39.435000 162.725000 ;
      RECT 37.000000 162.660000 39.435000 162.725000 ;
      RECT 37.000000 166.820000 39.435000 166.970000 ;
      RECT 37.150000 162.725000 39.285000 162.875000 ;
      RECT 37.150000 162.725000 39.285000 162.875000 ;
      RECT 37.150000 166.970000 39.285000 167.120000 ;
      RECT 37.280000   0.000000 37.980000  69.890000 ;
      RECT 37.280000   0.000000 37.980000  69.890000 ;
      RECT 37.280000  69.890000 50.355000  70.940000 ;
      RECT 37.280000  69.890000 50.355000  74.340000 ;
      RECT 37.280000  69.890000 50.455000  70.940000 ;
      RECT 37.280000  70.940000 50.455000  74.340000 ;
      RECT 37.300000 162.875000 39.135000 163.025000 ;
      RECT 37.300000 162.875000 39.135000 163.025000 ;
      RECT 37.300000 167.120000 39.135000 167.270000 ;
      RECT 37.325000 167.270000 39.110000 167.295000 ;
      RECT 37.325000 167.295000 37.545000 168.860000 ;
      RECT 37.325000 167.295000 38.960000 167.445000 ;
      RECT 37.325000 167.445000 38.810000 167.595000 ;
      RECT 37.325000 167.595000 38.660000 167.745000 ;
      RECT 37.325000 167.745000 38.510000 167.895000 ;
      RECT 37.325000 167.895000 38.360000 168.045000 ;
      RECT 37.325000 168.045000 38.210000 168.195000 ;
      RECT 37.325000 168.195000 38.060000 168.345000 ;
      RECT 37.325000 168.345000 37.910000 168.495000 ;
      RECT 37.325000 168.495000 37.760000 168.645000 ;
      RECT 37.325000 168.645000 37.610000 168.795000 ;
      RECT 37.325000 168.795000 37.460000 168.945000 ;
      RECT 37.325000 168.860000 37.545000 189.915000 ;
      RECT 37.430000  70.940000 50.355000  71.090000 ;
      RECT 37.430000  70.940000 50.355000  71.090000 ;
      RECT 37.450000 163.025000 38.985000 163.175000 ;
      RECT 37.450000 163.025000 38.985000 163.175000 ;
      RECT 37.580000  71.090000 50.355000  71.240000 ;
      RECT 37.580000  71.090000 50.355000  71.240000 ;
      RECT 37.600000 163.175000 38.835000 163.325000 ;
      RECT 37.600000 163.175000 38.835000 163.325000 ;
      RECT 37.730000  71.240000 50.355000  71.390000 ;
      RECT 37.730000  71.240000 50.355000  71.390000 ;
      RECT 37.750000 163.325000 38.685000 163.475000 ;
      RECT 37.750000 163.325000 38.685000 163.475000 ;
      RECT 37.880000  71.390000 50.355000  71.540000 ;
      RECT 37.880000  71.390000 50.355000  71.540000 ;
      RECT 37.900000 163.475000 38.535000 163.625000 ;
      RECT 37.900000 163.475000 38.535000 163.625000 ;
      RECT 38.030000  71.540000 50.355000  71.690000 ;
      RECT 38.030000  71.540000 50.355000  71.690000 ;
      RECT 38.050000 163.625000 38.385000 163.775000 ;
      RECT 38.050000 163.625000 38.385000 163.775000 ;
      RECT 38.180000  71.690000 50.355000  71.840000 ;
      RECT 38.180000  71.690000 50.355000  71.840000 ;
      RECT 38.190000  95.580000 42.435000  98.585000 ;
      RECT 38.200000 163.775000 38.235000 163.925000 ;
      RECT 38.200000 163.775000 38.235000 163.925000 ;
      RECT 38.215000 163.925000 38.220000 163.940000 ;
      RECT 38.215000 163.925000 38.220000 163.940000 ;
      RECT 38.330000  71.840000 50.355000  71.990000 ;
      RECT 38.330000  71.840000 50.355000  71.990000 ;
      RECT 38.480000  71.990000 50.355000  72.140000 ;
      RECT 38.480000  71.990000 50.355000  72.140000 ;
      RECT 38.630000  72.140000 50.355000  72.290000 ;
      RECT 38.630000  72.140000 50.355000  72.290000 ;
      RECT 38.780000  72.290000 50.355000  72.440000 ;
      RECT 38.780000  72.290000 50.355000  72.440000 ;
      RECT 38.930000  72.440000 50.355000  72.590000 ;
      RECT 38.930000  72.440000 50.355000  72.590000 ;
      RECT 39.080000  72.590000 50.355000  72.740000 ;
      RECT 39.080000  72.590000 50.355000  72.740000 ;
      RECT 39.230000  72.740000 50.355000  72.890000 ;
      RECT 39.230000  72.740000 50.355000  72.890000 ;
      RECT 39.380000  72.890000 50.355000  73.040000 ;
      RECT 39.380000  72.890000 50.355000  73.040000 ;
      RECT 39.430000  98.585000 42.435000 162.405000 ;
      RECT 39.530000  73.040000 50.355000  73.190000 ;
      RECT 39.530000  73.040000 50.355000  73.190000 ;
      RECT 39.680000  73.190000 50.355000  73.340000 ;
      RECT 39.680000  73.190000 50.355000  73.340000 ;
      RECT 39.785000  84.855000 41.210000  87.195000 ;
      RECT 39.785000  84.855000 41.210000  87.195000 ;
      RECT 39.785000  87.195000 41.210000  87.610000 ;
      RECT 39.810000  84.830000 41.185000  84.855000 ;
      RECT 39.830000  73.340000 50.355000  73.490000 ;
      RECT 39.830000  73.340000 50.355000  73.490000 ;
      RECT 39.935000  87.195000 41.210000  87.345000 ;
      RECT 39.960000  84.680000 41.035000  84.830000 ;
      RECT 39.980000  73.490000 50.355000  73.640000 ;
      RECT 39.980000  73.490000 50.355000  73.640000 ;
      RECT 40.085000  87.345000 41.210000  87.495000 ;
      RECT 40.110000  84.530000 40.885000  84.680000 ;
      RECT 40.130000  73.640000 50.355000  73.790000 ;
      RECT 40.130000  73.640000 50.355000  73.790000 ;
      RECT 40.200000  87.495000 41.210000  87.610000 ;
      RECT 40.200000  87.610000 50.245000  96.645000 ;
      RECT 40.260000  84.380000 40.735000  84.530000 ;
      RECT 40.260000  84.380000 41.210000  84.855000 ;
      RECT 40.280000  73.790000 50.355000  73.940000 ;
      RECT 40.280000  73.790000 50.355000  73.940000 ;
      RECT 40.350000  87.610000 41.210000  87.760000 ;
      RECT 40.430000  73.940000 50.355000  74.090000 ;
      RECT 40.430000  73.940000 50.355000  74.090000 ;
      RECT 40.500000  87.760000 41.360000  87.910000 ;
      RECT 40.580000  74.090000 50.355000  74.240000 ;
      RECT 40.580000  74.090000 50.355000  74.240000 ;
      RECT 40.650000  87.910000 41.510000  88.060000 ;
      RECT 40.680000  74.240000 50.355000  74.340000 ;
      RECT 40.680000  74.240000 50.355000  74.340000 ;
      RECT 40.800000  88.060000 41.660000  88.210000 ;
      RECT 40.950000  88.210000 41.810000  88.360000 ;
      RECT 41.100000  88.360000 41.960000  88.510000 ;
      RECT 41.250000  88.510000 42.110000  88.660000 ;
      RECT 41.400000  88.660000 42.260000  88.810000 ;
      RECT 41.550000  88.810000 42.410000  88.960000 ;
      RECT 41.700000  88.960000 42.560000  89.110000 ;
      RECT 41.850000  89.110000 42.710000  89.260000 ;
      RECT 42.000000  89.260000 42.860000  89.410000 ;
      RECT 42.150000  89.410000 43.010000  89.560000 ;
      RECT 42.300000  89.560000 43.160000  89.710000 ;
      RECT 42.450000  89.710000 43.310000  89.860000 ;
      RECT 42.600000  89.860000 43.460000  90.010000 ;
      RECT 42.750000  90.010000 43.610000  90.160000 ;
      RECT 42.900000  90.160000 43.760000  90.310000 ;
      RECT 43.050000  90.310000 43.910000  90.460000 ;
      RECT 43.200000  90.460000 44.060000  90.610000 ;
      RECT 43.350000  90.610000 44.210000  90.760000 ;
      RECT 43.500000  90.760000 44.360000  90.910000 ;
      RECT 43.650000  90.910000 44.510000  91.060000 ;
      RECT 43.800000  91.060000 44.660000  91.210000 ;
      RECT 43.950000  91.210000 44.810000  91.360000 ;
      RECT 44.100000  91.360000 44.960000  91.510000 ;
      RECT 44.250000  91.510000 45.110000  91.660000 ;
      RECT 44.400000  91.660000 45.260000  91.810000 ;
      RECT 44.550000  91.810000 45.410000  91.960000 ;
      RECT 44.700000  91.960000 45.560000  92.110000 ;
      RECT 44.850000  92.110000 45.710000  92.260000 ;
      RECT 45.000000  92.260000 45.860000  92.410000 ;
      RECT 45.150000  92.410000 46.010000  92.560000 ;
      RECT 45.300000  92.560000 46.160000  92.710000 ;
      RECT 45.450000  92.710000 46.310000  92.860000 ;
      RECT 45.600000  92.860000 46.460000  93.010000 ;
      RECT 45.750000  93.010000 46.610000  93.160000 ;
      RECT 45.900000  93.160000 46.760000  93.310000 ;
      RECT 46.050000  93.310000 46.910000  93.460000 ;
      RECT 46.200000  93.460000 47.060000  93.610000 ;
      RECT 46.350000  93.610000 47.210000  93.760000 ;
      RECT 46.500000  93.760000 47.360000  93.910000 ;
      RECT 46.650000  93.910000 47.510000  94.060000 ;
      RECT 46.800000  94.060000 47.660000  94.210000 ;
      RECT 46.950000  94.210000 47.810000  94.360000 ;
      RECT 46.960000  74.340000 50.455000  76.650000 ;
      RECT 47.100000  94.360000 47.960000  94.510000 ;
      RECT 47.110000  74.340000 50.355000  74.490000 ;
      RECT 47.110000  74.340000 50.355000  74.490000 ;
      RECT 47.250000  94.510000 48.110000  94.660000 ;
      RECT 47.260000  74.490000 50.355000  74.640000 ;
      RECT 47.260000  74.490000 50.355000  74.640000 ;
      RECT 47.400000  94.660000 48.260000  94.810000 ;
      RECT 47.410000  74.640000 50.355000  74.790000 ;
      RECT 47.410000  74.640000 50.355000  74.790000 ;
      RECT 47.550000  94.810000 48.410000  94.960000 ;
      RECT 47.560000  74.790000 50.355000  74.940000 ;
      RECT 47.560000  74.790000 50.355000  74.940000 ;
      RECT 47.700000  94.960000 48.560000  95.110000 ;
      RECT 47.710000  74.940000 50.355000  75.090000 ;
      RECT 47.710000  74.940000 50.355000  75.090000 ;
      RECT 47.850000  95.110000 48.710000  95.260000 ;
      RECT 47.860000  75.090000 50.355000  75.240000 ;
      RECT 47.860000  75.090000 50.355000  75.240000 ;
      RECT 48.000000  95.260000 48.860000  95.410000 ;
      RECT 48.010000  75.240000 50.355000  75.390000 ;
      RECT 48.010000  75.240000 50.355000  75.390000 ;
      RECT 48.150000  95.410000 49.010000  95.560000 ;
      RECT 48.160000  75.390000 50.355000  75.540000 ;
      RECT 48.160000  75.390000 50.355000  75.540000 ;
      RECT 48.300000  95.560000 49.160000  95.710000 ;
      RECT 48.310000  75.540000 50.355000  75.690000 ;
      RECT 48.310000  75.540000 50.355000  75.690000 ;
      RECT 48.450000  95.710000 49.310000  95.860000 ;
      RECT 48.460000  75.690000 50.355000  75.840000 ;
      RECT 48.460000  75.690000 50.355000  75.840000 ;
      RECT 48.600000  95.860000 49.460000  96.010000 ;
      RECT 48.610000  75.840000 50.355000  75.990000 ;
      RECT 48.610000  75.840000 50.355000  75.990000 ;
      RECT 48.750000  96.010000 49.610000  96.160000 ;
      RECT 48.760000  75.990000 50.355000  76.140000 ;
      RECT 48.760000  75.990000 50.355000  76.140000 ;
      RECT 48.900000  96.160000 49.760000  96.310000 ;
      RECT 48.910000  76.140000 50.355000  76.290000 ;
      RECT 48.910000  76.140000 50.355000  76.290000 ;
      RECT 49.050000  96.310000 49.910000  96.460000 ;
      RECT 49.060000  76.290000 50.355000  76.440000 ;
      RECT 49.060000  76.290000 50.355000  76.440000 ;
      RECT 49.200000  96.460000 50.060000  96.610000 ;
      RECT 49.210000  76.440000 50.355000  76.590000 ;
      RECT 49.210000  76.440000 50.355000  76.590000 ;
      RECT 49.235000  96.610000 50.210000  96.645000 ;
      RECT 49.235000  96.645000 50.245000  96.795000 ;
      RECT 49.235000  96.645000 53.930000 100.330000 ;
      RECT 49.235000  96.795000 50.395000  96.945000 ;
      RECT 49.235000  96.945000 50.545000  97.095000 ;
      RECT 49.235000  97.095000 50.695000  97.245000 ;
      RECT 49.235000  97.245000 50.845000  97.395000 ;
      RECT 49.235000  97.395000 50.995000  97.545000 ;
      RECT 49.235000  97.545000 51.145000  97.695000 ;
      RECT 49.235000  97.695000 51.295000  97.845000 ;
      RECT 49.235000  97.845000 51.445000  97.995000 ;
      RECT 49.235000  97.995000 51.595000  98.145000 ;
      RECT 49.235000  98.145000 51.745000  98.295000 ;
      RECT 49.235000  98.295000 51.895000  98.445000 ;
      RECT 49.235000  98.445000 52.045000  98.595000 ;
      RECT 49.235000  98.595000 52.195000  98.745000 ;
      RECT 49.235000  98.745000 52.345000  98.895000 ;
      RECT 49.235000  98.895000 52.495000  99.045000 ;
      RECT 49.235000  99.045000 52.645000  99.195000 ;
      RECT 49.235000  99.195000 52.795000  99.345000 ;
      RECT 49.235000  99.345000 52.945000  99.495000 ;
      RECT 49.235000  99.495000 53.095000  99.645000 ;
      RECT 49.235000  99.645000 53.245000  99.795000 ;
      RECT 49.235000  99.795000 53.395000  99.945000 ;
      RECT 49.235000  99.945000 53.545000 100.095000 ;
      RECT 49.235000 100.095000 53.695000 100.245000 ;
      RECT 49.235000 100.245000 53.845000 100.330000 ;
      RECT 49.235000 100.330000 53.930000 164.295000 ;
      RECT 49.235000 100.330000 53.930000 164.295000 ;
      RECT 49.235000 164.295000 49.470000 168.755000 ;
      RECT 49.235000 164.295000 53.780000 164.445000 ;
      RECT 49.235000 164.445000 53.630000 164.595000 ;
      RECT 49.235000 164.595000 53.480000 164.745000 ;
      RECT 49.235000 164.745000 53.330000 164.895000 ;
      RECT 49.235000 164.895000 53.180000 165.045000 ;
      RECT 49.235000 165.045000 53.030000 165.195000 ;
      RECT 49.235000 165.195000 52.880000 165.345000 ;
      RECT 49.235000 165.345000 52.730000 165.495000 ;
      RECT 49.235000 165.495000 52.580000 165.645000 ;
      RECT 49.235000 165.645000 52.430000 165.795000 ;
      RECT 49.235000 165.795000 52.280000 165.945000 ;
      RECT 49.235000 165.945000 52.130000 166.095000 ;
      RECT 49.235000 166.095000 51.980000 166.245000 ;
      RECT 49.235000 166.245000 51.830000 166.395000 ;
      RECT 49.235000 166.395000 51.680000 166.545000 ;
      RECT 49.235000 166.545000 51.530000 166.695000 ;
      RECT 49.235000 166.695000 51.380000 166.845000 ;
      RECT 49.235000 166.845000 51.230000 166.995000 ;
      RECT 49.235000 166.995000 51.080000 167.145000 ;
      RECT 49.235000 167.145000 50.930000 167.295000 ;
      RECT 49.235000 167.295000 50.780000 167.445000 ;
      RECT 49.235000 167.445000 50.630000 167.595000 ;
      RECT 49.235000 167.595000 50.480000 167.745000 ;
      RECT 49.235000 167.745000 50.330000 167.895000 ;
      RECT 49.235000 167.895000 50.180000 168.045000 ;
      RECT 49.235000 168.045000 50.030000 168.195000 ;
      RECT 49.235000 168.195000 49.880000 168.345000 ;
      RECT 49.235000 168.345000 49.730000 168.495000 ;
      RECT 49.235000 168.495000 49.580000 168.645000 ;
      RECT 49.235000 168.645000 49.430000 168.795000 ;
      RECT 49.235000 168.755000 49.470000 189.915000 ;
      RECT 49.235000 168.795000 49.280000 168.945000 ;
      RECT 49.270000  76.590000 50.355000  76.650000 ;
      RECT 49.270000  76.590000 50.355000  76.650000 ;
      RECT 49.270000  76.650000 50.455000  84.590000 ;
      RECT 49.270000  77.735000 50.355000  84.630000 ;
      RECT 49.270000  84.590000 50.510000  84.645000 ;
      RECT 49.270000  84.630000 50.355000  84.635000 ;
      RECT 49.270000  84.635000 50.360000  84.640000 ;
      RECT 49.270000  84.640000 50.365000  84.645000 ;
      RECT 49.270000  84.645000 52.660000  86.795000 ;
      RECT 49.420000  76.650000 50.355000  76.800000 ;
      RECT 49.420000  76.650000 50.355000  76.800000 ;
      RECT 49.420000  84.645000 50.370000  84.795000 ;
      RECT 49.570000  76.800000 50.355000  76.950000 ;
      RECT 49.570000  76.800000 50.355000  76.950000 ;
      RECT 49.570000  84.795000 50.520000  84.945000 ;
      RECT 49.655000   0.000000 50.355000  69.890000 ;
      RECT 49.655000   0.000000 50.455000  69.890000 ;
      RECT 49.720000  76.950000 50.355000  77.100000 ;
      RECT 49.720000  76.950000 50.355000  77.100000 ;
      RECT 49.720000  84.945000 50.670000  85.095000 ;
      RECT 49.870000  77.100000 50.355000  77.250000 ;
      RECT 49.870000  77.100000 50.355000  77.250000 ;
      RECT 49.870000  85.095000 50.820000  85.245000 ;
      RECT 50.020000  77.250000 50.355000  77.400000 ;
      RECT 50.020000  77.250000 50.355000  77.400000 ;
      RECT 50.020000  85.245000 50.970000  85.395000 ;
      RECT 50.170000  77.400000 50.355000  77.550000 ;
      RECT 50.170000  77.400000 50.355000  77.550000 ;
      RECT 50.170000  85.395000 51.120000  85.545000 ;
      RECT 50.320000  77.550000 50.355000  77.700000 ;
      RECT 50.320000  77.550000 50.355000  77.700000 ;
      RECT 50.320000  85.545000 51.270000  85.695000 ;
      RECT 50.470000  85.695000 51.420000  85.845000 ;
      RECT 50.620000  85.845000 51.570000  85.995000 ;
      RECT 50.770000  85.995000 51.720000  86.145000 ;
      RECT 50.920000  86.145000 51.870000  86.295000 ;
      RECT 51.070000  86.295000 52.020000  86.445000 ;
      RECT 51.220000  86.445000 52.170000  86.595000 ;
      RECT 51.370000  86.595000 52.320000  86.745000 ;
      RECT 51.420000  86.745000 52.470000  86.795000 ;
      RECT 51.420000  86.795000 52.520000  86.945000 ;
      RECT 51.420000  86.795000 54.075000  88.210000 ;
      RECT 51.420000  86.945000 52.670000  87.095000 ;
      RECT 51.420000  87.095000 52.820000  87.245000 ;
      RECT 51.420000  87.245000 52.970000  87.395000 ;
      RECT 51.420000  87.395000 53.120000  87.545000 ;
      RECT 51.420000  87.545000 53.270000  87.695000 ;
      RECT 51.420000  87.695000 53.420000  87.845000 ;
      RECT 51.420000  87.845000 53.570000  87.995000 ;
      RECT 51.420000  87.995000 53.720000  88.145000 ;
      RECT 51.420000  88.145000 53.870000  88.210000 ;
      RECT 51.420000  88.210000 61.745000  95.880000 ;
      RECT 51.570000  88.210000 53.935000  88.360000 ;
      RECT 51.720000  88.360000 54.085000  88.510000 ;
      RECT 51.870000  88.510000 54.235000  88.660000 ;
      RECT 52.020000  88.660000 54.385000  88.810000 ;
      RECT 52.170000  88.810000 54.535000  88.960000 ;
      RECT 52.320000  88.960000 54.685000  89.110000 ;
      RECT 52.470000  89.110000 54.835000  89.260000 ;
      RECT 52.620000  89.260000 54.985000  89.410000 ;
      RECT 52.770000  89.410000 55.135000  89.560000 ;
      RECT 52.920000  89.560000 55.285000  89.710000 ;
      RECT 53.070000  89.710000 55.435000  89.860000 ;
      RECT 53.220000  89.860000 55.585000  90.010000 ;
      RECT 53.370000  90.010000 55.735000  90.160000 ;
      RECT 53.520000  90.160000 55.885000  90.310000 ;
      RECT 53.670000  90.310000 56.035000  90.460000 ;
      RECT 53.820000  90.460000 56.185000  90.610000 ;
      RECT 53.970000  90.610000 56.335000  90.760000 ;
      RECT 54.120000  90.760000 56.485000  90.910000 ;
      RECT 54.270000  90.910000 56.635000  91.060000 ;
      RECT 54.420000  91.060000 56.785000  91.210000 ;
      RECT 54.570000  91.210000 56.935000  91.360000 ;
      RECT 54.720000  91.360000 57.085000  91.510000 ;
      RECT 54.870000  91.510000 57.235000  91.660000 ;
      RECT 55.020000  91.660000 57.385000  91.810000 ;
      RECT 55.170000  91.810000 57.535000  91.960000 ;
      RECT 55.320000  91.960000 57.685000  92.110000 ;
      RECT 55.470000  92.110000 57.835000  92.260000 ;
      RECT 55.620000  92.260000 57.985000  92.410000 ;
      RECT 55.770000  92.410000 58.135000  92.560000 ;
      RECT 55.920000  92.560000 58.285000  92.710000 ;
      RECT 56.070000  92.710000 58.435000  92.860000 ;
      RECT 56.220000  92.860000 58.585000  93.010000 ;
      RECT 56.370000  93.010000 58.735000  93.160000 ;
      RECT 56.520000  93.160000 58.885000  93.310000 ;
      RECT 56.670000  93.310000 59.035000  93.460000 ;
      RECT 56.820000  93.460000 59.185000  93.610000 ;
      RECT 56.970000  93.610000 59.335000  93.760000 ;
      RECT 57.120000  93.760000 59.485000  93.910000 ;
      RECT 57.270000  93.910000 59.635000  94.060000 ;
      RECT 57.420000  94.060000 59.785000  94.210000 ;
      RECT 57.570000  94.210000 59.935000  94.360000 ;
      RECT 57.720000  94.360000 60.085000  94.510000 ;
      RECT 57.870000  94.510000 60.235000  94.660000 ;
      RECT 58.020000  94.660000 60.385000  94.810000 ;
      RECT 58.170000  94.810000 60.535000  94.960000 ;
      RECT 58.320000  94.960000 60.685000  95.110000 ;
      RECT 58.470000  95.110000 60.835000  95.260000 ;
      RECT 58.620000  95.260000 60.985000  95.410000 ;
      RECT 58.770000  95.410000 61.135000  95.560000 ;
      RECT 58.920000  95.560000 61.285000  95.710000 ;
      RECT 59.070000  95.710000 61.435000  95.860000 ;
      RECT 59.090000  95.880000 61.745000  97.520000 ;
      RECT 59.130000  95.860000 61.585000  95.920000 ;
      RECT 59.280000  95.920000 61.645000  96.070000 ;
      RECT 59.430000  96.070000 61.645000  96.220000 ;
      RECT 59.580000  96.220000 61.645000  96.370000 ;
      RECT 59.730000  96.370000 61.645000  96.520000 ;
      RECT 59.880000  96.520000 61.645000  96.670000 ;
      RECT 60.030000  96.670000 61.645000  96.820000 ;
      RECT 60.180000  96.820000 61.645000  96.970000 ;
      RECT 60.330000  96.970000 61.645000  97.120000 ;
      RECT 60.480000  97.120000 61.645000  97.270000 ;
      RECT 60.630000  97.270000 61.645000  97.420000 ;
      RECT 60.730000  97.420000 61.645000  97.520000 ;
      RECT 60.730000  97.520000 61.645000 172.635000 ;
      RECT 60.730000  97.520000 61.745000 172.535000 ;
      RECT 60.730000 172.535000 75.000000 189.915000 ;
      RECT 60.730000 172.635000 75.000000 189.915000 ;
      RECT 60.730000 172.635000 75.000000 198.000000 ;
    LAYER met4 ;
      RECT  4.820000 102.300000  7.470000 164.545000 ;
      RECT  5.440000 101.650000  5.945000 102.180000 ;
      RECT  5.440000 164.605000  5.945000 165.135000 ;
      RECT  6.070000 101.090000  8.445000 102.160000 ;
      RECT  6.070000 164.625000  8.445000 165.695000 ;
      RECT  6.555000 100.535000  7.060000 101.065000 ;
      RECT  6.555000 165.720000  7.060000 166.250000 ;
      RECT  7.350000  99.950000  9.725000 101.020000 ;
      RECT  7.350000 165.765000  9.725000 166.835000 ;
      RECT  7.535000 102.245000  8.040000 102.775000 ;
      RECT  7.535000 164.010000  8.040000 164.540000 ;
      RECT  7.750000  99.340000  8.255000  99.870000 ;
      RECT  7.750000 166.915000  8.255000 167.445000 ;
      RECT  8.340000  98.810000 10.715000  99.880000 ;
      RECT  8.415000 166.915000 10.700000 167.865000 ;
      RECT  8.650000 101.130000  9.155000 101.660000 ;
      RECT  8.650000 165.125000  9.155000 165.655000 ;
      RECT  8.825000  98.265000  9.330000  98.795000 ;
      RECT  8.825000 167.990000  9.330000 168.520000 ;
      RECT  9.460000  97.645000 11.835000  98.715000 ;
      RECT  9.460000 168.025000 11.835000 169.095000 ;
      RECT  9.845000  99.935000 10.350000 100.465000 ;
      RECT  9.845000 166.320000 10.350000 166.850000 ;
      RECT  9.985000  97.070000 10.490000  97.600000 ;
      RECT  9.985000 169.150000 10.490000 169.680000 ;
      RECT 10.595000  96.475000 11.850000  96.480000 ;
      RECT 10.595000  96.480000 11.835000  97.545000 ;
      RECT 10.610000 169.340000 11.745000 170.260000 ;
      RECT 10.920000  98.860000 11.425000  99.390000 ;
      RECT 10.920000 167.395000 11.425000 167.925000 ;
      RECT 11.095000  95.950000 11.850000  96.475000 ;
      RECT 11.095000 170.260000 11.850000 170.790000 ;
      RECT 11.965000  95.795000 12.835000  98.295000 ;
      RECT 11.965000 168.490000 12.835000 170.990000 ;
      RECT 25.035000  17.815000 25.465000  22.250000 ;
      RECT 25.035000  39.785000 25.365000  41.435000 ;
      RECT 62.225000  95.795000 63.095000  98.295000 ;
      RECT 62.225000 168.490000 63.095000 170.990000 ;
      RECT 63.225000  96.475000 64.465000  97.545000 ;
      RECT 63.225000  97.645000 65.600000  98.715000 ;
      RECT 63.225000 169.160000 64.465000 170.230000 ;
      RECT 63.235000 168.165000 65.495000 169.005000 ;
      RECT 63.635000  98.860000 64.140000  99.390000 ;
      RECT 63.635000 167.395000 64.140000 167.925000 ;
      RECT 64.345000  98.810000 66.720000  99.880000 ;
      RECT 64.345000 166.905000 66.720000 167.975000 ;
      RECT 64.570000  97.070000 65.075000  97.600000 ;
      RECT 64.570000 169.150000 65.075000 169.680000 ;
      RECT 64.710000  99.935000 65.215000 100.465000 ;
      RECT 64.710000 166.320000 65.215000 166.850000 ;
      RECT 65.335000  99.950000 67.710000 101.020000 ;
      RECT 65.335000 165.765000 67.710000 166.835000 ;
      RECT 65.730000  98.265000 66.235000  98.795000 ;
      RECT 65.730000 167.990000 66.235000 168.520000 ;
      RECT 65.905000 101.130000 66.410000 101.660000 ;
      RECT 65.905000 165.125000 66.410000 165.655000 ;
      RECT 66.615000 101.090000 68.990000 102.160000 ;
      RECT 66.615000 164.625000 68.990000 165.695000 ;
      RECT 66.805000  99.340000 67.310000  99.870000 ;
      RECT 66.805000 166.915000 67.310000 167.445000 ;
      RECT 67.020000 102.245000 70.110000 102.775000 ;
      RECT 67.020000 164.010000 70.165000 164.350000 ;
      RECT 67.020000 164.350000 67.525000 164.540000 ;
      RECT 67.515000 103.000000 70.165000 164.010000 ;
      RECT 68.000000 100.535000 68.505000 101.065000 ;
      RECT 68.000000 165.720000 68.505000 166.250000 ;
      RECT 69.115000 101.650000 69.620000 102.180000 ;
      RECT 69.115000 164.605000 69.620000 165.135000 ;
  END
END sky130_fd_io__top_ground_lvc_wpad
END LIBRARY
