VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

SITE asap7sc7p5t_pg
 CLASS CORE ;
 SIZE 0.054 BY 0.540 ;
 SYMMETRY X Y ;
END asap7sc7p5t_pg

MACRO DFFHQNH2V2Xx1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNH2V2Xx1_ASAP7_75t_L 0 0 ;
  SIZE 2.16 BY 0.54 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t_pg ;
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.314 0.126 1.37 0.144 ;
        RECT 1.314 0.225 1.351 0.243 ;
        RECT 1.314 0.027 1.351 0.045 ;
        RECT 1.314 0.027 1.332 0.243 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.314 0.396 1.37 0.414 ;
        RECT 1.314 0.495 1.351 0.513 ;
        RECT 1.314 0.297 1.351 0.315 ;
        RECT 1.314 0.297 1.332 0.513 ;
    END
  END D1
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.809 0.225 0.846 0.243 ;
        RECT 0.828 0.027 0.846 0.243 ;
        RECT 0.79 0.126 0.846 0.144 ;
        RECT 0.809 0.027 0.846 0.045 ;
    END
  END D2
  PIN D3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.809 0.495 0.846 0.513 ;
        RECT 0.828 0.297 0.846 0.513 ;
        RECT 0.79 0.396 0.846 0.414 ;
        RECT 0.809 0.297 0.846 0.315 ;
    END
  END D3
  PIN QN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.092 0.225 2.142 0.243 ;
        RECT 2.124 0.027 2.142 0.243 ;
        RECT 2.092 0.027 2.142 0.045 ;
    END
  END QN0
  PIN QN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.092 0.495 2.142 0.513 ;
        RECT 2.124 0.297 2.142 0.513 ;
        RECT 2.092 0.297 2.142 0.315 ;
    END
  END QN1
  PIN QN2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.225 0.068 0.243 ;
        RECT 0.018 0.027 0.068 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END QN2
  PIN QN3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.495 0.068 0.513 ;
        RECT 0.018 0.297 0.068 0.315 ;
        RECT 0.018 0.297 0.036 0.513 ;
    END
  END QN3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 2.16 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 2.16 0.009 ;
        RECT 0 0.531 2.16 0.549 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 0.958 0.07 1.202 0.088 ;
        RECT 0.958 0.452 1.202 0.47 ;
      LAYER M3 ;
        RECT 1.017 0.05 1.035 0.492 ;
      LAYER M1 ;
        RECT 1.179 0.164 1.197 0.236 ;
        RECT 1.152 0.07 1.197 0.106 ;
        RECT 1.179 0.034 1.197 0.106 ;
        RECT 1.152 0.164 1.197 0.2 ;
        RECT 1.152 0.07 1.17 0.2 ;
        RECT 1.179 0.434 1.197 0.506 ;
        RECT 1.152 0.34 1.197 0.376 ;
        RECT 1.179 0.304 1.197 0.376 ;
        RECT 1.152 0.434 1.197 0.47 ;
        RECT 1.152 0.34 1.17 0.47 ;
        RECT 0.963 0.164 1.008 0.2 ;
        RECT 0.99 0.07 1.008 0.2 ;
        RECT 0.963 0.07 1.008 0.106 ;
        RECT 0.963 0.164 0.981 0.236 ;
        RECT 0.963 0.034 0.981 0.106 ;
        RECT 0.963 0.434 1.008 0.47 ;
        RECT 0.99 0.34 1.008 0.47 ;
        RECT 0.963 0.34 1.008 0.376 ;
        RECT 0.963 0.434 0.981 0.506 ;
        RECT 0.963 0.304 0.981 0.376 ;
      LAYER V2 ;
        RECT 1.017 0.452 1.035 0.47 ;
        RECT 1.017 0.07 1.035 0.088 ;
      LAYER V1 ;
        RECT 0.963 0.452 0.981 0.47 ;
        RECT 0.963 0.07 0.981 0.088 ;
        RECT 1.179 0.452 1.197 0.47 ;
        RECT 1.179 0.07 1.197 0.088 ;
    END
  END CLK
  OBS
    LAYER M1 ;
      RECT 1.93 0.225 2.034 0.243 ;
      RECT 2.016 0.027 2.034 0.243 ;
      RECT 1.854 0.027 1.872 0.119 ;
      RECT 1.854 0.027 2.034 0.045 ;
      RECT 1.854 0.495 2.034 0.513 ;
      RECT 2.016 0.297 2.034 0.513 ;
      RECT 1.854 0.421 1.872 0.513 ;
      RECT 1.93 0.297 2.034 0.315 ;
      RECT 1.768 0.224 1.818 0.242 ;
      RECT 1.8 0.027 1.818 0.242 ;
      RECT 1.8 0.153 1.98 0.171 ;
      RECT 1.962 0.117 1.98 0.171 ;
      RECT 1.908 0.117 1.926 0.171 ;
      RECT 1.714 0.027 1.818 0.045 ;
      RECT 1.714 0.495 1.818 0.513 ;
      RECT 1.8 0.298 1.818 0.513 ;
      RECT 1.962 0.369 1.98 0.423 ;
      RECT 1.908 0.369 1.926 0.423 ;
      RECT 1.8 0.369 1.98 0.387 ;
      RECT 1.768 0.298 1.818 0.316 ;
      RECT 1.656 0.225 1.71 0.243 ;
      RECT 1.692 0.081 1.71 0.243 ;
      RECT 1.576 0.081 1.71 0.099 ;
      RECT 1.665 0.045 1.683 0.099 ;
      RECT 1.665 0.441 1.683 0.495 ;
      RECT 1.576 0.441 1.71 0.459 ;
      RECT 1.692 0.297 1.71 0.459 ;
      RECT 1.656 0.297 1.71 0.315 ;
      RECT 1.444 0.225 1.548 0.243 ;
      RECT 1.53 0.027 1.548 0.243 ;
      RECT 1.53 0.122 1.656 0.14 ;
      RECT 1.498 0.027 1.548 0.045 ;
      RECT 1.498 0.495 1.548 0.513 ;
      RECT 1.53 0.297 1.548 0.513 ;
      RECT 1.53 0.4 1.656 0.418 ;
      RECT 1.444 0.297 1.548 0.315 ;
      RECT 1.395 0.126 1.413 0.203 ;
      RECT 1.395 0.126 1.447 0.144 ;
      RECT 1.395 0.396 1.447 0.414 ;
      RECT 1.395 0.337 1.413 0.414 ;
      RECT 1.228 0.225 1.278 0.243 ;
      RECT 1.26 0.027 1.278 0.243 ;
      RECT 1.228 0.027 1.278 0.045 ;
      RECT 1.228 0.495 1.278 0.513 ;
      RECT 1.26 0.297 1.278 0.513 ;
      RECT 1.228 0.297 1.278 0.315 ;
      RECT 1.089 0.225 1.148 0.243 ;
      RECT 1.089 0.027 1.107 0.243 ;
      RECT 1.089 0.144 1.127 0.162 ;
      RECT 1.089 0.027 1.148 0.045 ;
      RECT 1.089 0.495 1.148 0.513 ;
      RECT 1.089 0.297 1.107 0.513 ;
      RECT 1.089 0.378 1.127 0.396 ;
      RECT 1.089 0.297 1.148 0.315 ;
      RECT 1.012 0.225 1.071 0.243 ;
      RECT 1.053 0.027 1.071 0.243 ;
      RECT 1.033 0.144 1.071 0.162 ;
      RECT 1.012 0.027 1.071 0.045 ;
      RECT 1.012 0.495 1.071 0.513 ;
      RECT 1.053 0.297 1.071 0.513 ;
      RECT 1.033 0.378 1.071 0.396 ;
      RECT 1.012 0.297 1.071 0.315 ;
      RECT 0.882 0.225 0.932 0.243 ;
      RECT 0.882 0.027 0.9 0.243 ;
      RECT 0.882 0.027 0.932 0.045 ;
      RECT 0.882 0.495 0.932 0.513 ;
      RECT 0.882 0.297 0.9 0.513 ;
      RECT 0.882 0.297 0.932 0.315 ;
      RECT 0.747 0.126 0.765 0.203 ;
      RECT 0.713 0.126 0.765 0.144 ;
      RECT 0.713 0.396 0.765 0.414 ;
      RECT 0.747 0.337 0.765 0.414 ;
      RECT 0.612 0.225 0.716 0.243 ;
      RECT 0.612 0.027 0.63 0.243 ;
      RECT 0.504 0.122 0.63 0.14 ;
      RECT 0.612 0.027 0.662 0.045 ;
      RECT 0.612 0.495 0.662 0.513 ;
      RECT 0.612 0.297 0.63 0.513 ;
      RECT 0.504 0.4 0.63 0.418 ;
      RECT 0.612 0.297 0.716 0.315 ;
      RECT 0.45 0.225 0.504 0.243 ;
      RECT 0.45 0.081 0.468 0.243 ;
      RECT 0.45 0.081 0.584 0.099 ;
      RECT 0.477 0.045 0.495 0.099 ;
      RECT 0.477 0.441 0.495 0.495 ;
      RECT 0.45 0.441 0.584 0.459 ;
      RECT 0.45 0.297 0.468 0.459 ;
      RECT 0.45 0.297 0.504 0.315 ;
      RECT 0.342 0.224 0.392 0.242 ;
      RECT 0.342 0.027 0.36 0.242 ;
      RECT 0.18 0.153 0.36 0.171 ;
      RECT 0.234 0.117 0.252 0.171 ;
      RECT 0.18 0.117 0.198 0.171 ;
      RECT 0.342 0.027 0.446 0.045 ;
      RECT 0.342 0.495 0.446 0.513 ;
      RECT 0.342 0.298 0.36 0.513 ;
      RECT 0.234 0.369 0.252 0.423 ;
      RECT 0.18 0.369 0.198 0.423 ;
      RECT 0.18 0.369 0.36 0.387 ;
      RECT 0.342 0.298 0.392 0.316 ;
      RECT 0.126 0.225 0.23 0.243 ;
      RECT 0.126 0.027 0.144 0.243 ;
      RECT 0.288 0.027 0.306 0.119 ;
      RECT 0.126 0.027 0.306 0.045 ;
      RECT 0.126 0.495 0.306 0.513 ;
      RECT 0.288 0.421 0.306 0.513 ;
      RECT 0.126 0.297 0.144 0.513 ;
      RECT 0.126 0.297 0.23 0.315 ;
      RECT 2.07 0.09 2.088 0.167 ;
      RECT 2.07 0.373 2.088 0.45 ;
      RECT 1.746 0.101 1.764 0.167 ;
      RECT 1.746 0.373 1.764 0.439 ;
      RECT 1.584 0.165 1.602 0.203 ;
      RECT 1.584 0.337 1.602 0.375 ;
      RECT 1.476 0.106 1.494 0.167 ;
      RECT 1.476 0.373 1.494 0.434 ;
      RECT 1.222 0.106 1.24 0.167 ;
      RECT 1.222 0.373 1.24 0.434 ;
      RECT 0.92 0.106 0.938 0.167 ;
      RECT 0.92 0.373 0.938 0.434 ;
      RECT 0.666 0.106 0.684 0.167 ;
      RECT 0.666 0.373 0.684 0.434 ;
      RECT 0.558 0.165 0.576 0.203 ;
      RECT 0.558 0.337 0.576 0.375 ;
      RECT 0.396 0.101 0.414 0.167 ;
      RECT 0.396 0.373 0.414 0.439 ;
      RECT 0.072 0.09 0.09 0.167 ;
      RECT 0.072 0.373 0.09 0.45 ;
    LAYER M2 ;
      RECT 1.957 0.144 2.093 0.162 ;
      RECT 1.957 0.378 2.093 0.396 ;
      RECT 1.099 0.144 1.769 0.162 ;
      RECT 1.099 0.378 1.769 0.396 ;
      RECT 1.255 0.18 1.607 0.198 ;
      RECT 1.255 0.342 1.607 0.36 ;
      RECT 0.391 0.144 1.061 0.162 ;
      RECT 0.391 0.378 1.061 0.396 ;
      RECT 0.553 0.18 0.905 0.198 ;
      RECT 0.553 0.342 0.905 0.36 ;
      RECT 0.067 0.144 0.203 0.162 ;
      RECT 0.067 0.378 0.203 0.396 ;
    LAYER V1 ;
      RECT 2.07 0.144 2.088 0.162 ;
      RECT 2.07 0.378 2.088 0.396 ;
      RECT 1.962 0.144 1.98 0.162 ;
      RECT 1.962 0.378 1.98 0.396 ;
      RECT 1.746 0.144 1.764 0.162 ;
      RECT 1.746 0.378 1.764 0.396 ;
      RECT 1.584 0.18 1.602 0.198 ;
      RECT 1.584 0.342 1.602 0.36 ;
      RECT 1.476 0.144 1.494 0.162 ;
      RECT 1.476 0.378 1.494 0.396 ;
      RECT 1.395 0.18 1.413 0.198 ;
      RECT 1.395 0.342 1.413 0.36 ;
      RECT 1.26 0.18 1.278 0.198 ;
      RECT 1.26 0.342 1.278 0.36 ;
      RECT 1.222 0.144 1.24 0.162 ;
      RECT 1.222 0.378 1.24 0.396 ;
      RECT 1.104 0.144 1.122 0.162 ;
      RECT 1.104 0.378 1.122 0.396 ;
      RECT 1.038 0.144 1.056 0.162 ;
      RECT 1.038 0.378 1.056 0.396 ;
      RECT 0.92 0.144 0.938 0.162 ;
      RECT 0.92 0.378 0.938 0.396 ;
      RECT 0.882 0.18 0.9 0.198 ;
      RECT 0.882 0.342 0.9 0.36 ;
      RECT 0.747 0.18 0.765 0.198 ;
      RECT 0.747 0.342 0.765 0.36 ;
      RECT 0.666 0.144 0.684 0.162 ;
      RECT 0.666 0.378 0.684 0.396 ;
      RECT 0.558 0.18 0.576 0.198 ;
      RECT 0.558 0.342 0.576 0.36 ;
      RECT 0.396 0.144 0.414 0.162 ;
      RECT 0.396 0.378 0.414 0.396 ;
      RECT 0.18 0.144 0.198 0.162 ;
      RECT 0.18 0.378 0.198 0.396 ;
      RECT 0.072 0.144 0.09 0.162 ;
      RECT 0.072 0.378 0.09 0.396 ;
  END
END DFFHQNH2V2Xx1_ASAP7_75t_L

MACRO DFFHQNH2V2Xx1_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNH2V2Xx1_ASAP7_75t_R 0 0 ;
  SIZE 2.16 BY 0.54 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t_pg ;
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.314 0.126 1.37 0.144 ;
        RECT 1.314 0.225 1.351 0.243 ;
        RECT 1.314 0.027 1.351 0.045 ;
        RECT 1.314 0.027 1.332 0.243 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.314 0.396 1.37 0.414 ;
        RECT 1.314 0.495 1.351 0.513 ;
        RECT 1.314 0.297 1.351 0.315 ;
        RECT 1.314 0.297 1.332 0.513 ;
    END
  END D1
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.809 0.225 0.846 0.243 ;
        RECT 0.828 0.027 0.846 0.243 ;
        RECT 0.79 0.126 0.846 0.144 ;
        RECT 0.809 0.027 0.846 0.045 ;
    END
  END D2
  PIN D3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.809 0.495 0.846 0.513 ;
        RECT 0.828 0.297 0.846 0.513 ;
        RECT 0.79 0.396 0.846 0.414 ;
        RECT 0.809 0.297 0.846 0.315 ;
    END
  END D3
  PIN QN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.092 0.225 2.142 0.243 ;
        RECT 2.124 0.027 2.142 0.243 ;
        RECT 2.092 0.027 2.142 0.045 ;
    END
  END QN0
  PIN QN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.092 0.495 2.142 0.513 ;
        RECT 2.124 0.297 2.142 0.513 ;
        RECT 2.092 0.297 2.142 0.315 ;
    END
  END QN1
  PIN QN2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.225 0.068 0.243 ;
        RECT 0.018 0.027 0.068 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END QN2
  PIN QN3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.495 0.068 0.513 ;
        RECT 0.018 0.297 0.068 0.315 ;
        RECT 0.018 0.297 0.036 0.513 ;
    END
  END QN3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 2.16 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 2.16 0.009 ;
        RECT 0 0.531 2.16 0.549 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 0.958 0.07 1.202 0.088 ;
        RECT 0.958 0.452 1.202 0.47 ;
      LAYER M3 ;
        RECT 1.017 0.05 1.035 0.492 ;
      LAYER M1 ;
        RECT 1.179 0.164 1.197 0.236 ;
        RECT 1.152 0.07 1.197 0.106 ;
        RECT 1.179 0.034 1.197 0.106 ;
        RECT 1.152 0.164 1.197 0.2 ;
        RECT 1.152 0.07 1.17 0.2 ;
        RECT 1.179 0.434 1.197 0.506 ;
        RECT 1.152 0.34 1.197 0.376 ;
        RECT 1.179 0.304 1.197 0.376 ;
        RECT 1.152 0.434 1.197 0.47 ;
        RECT 1.152 0.34 1.17 0.47 ;
        RECT 0.963 0.164 1.008 0.2 ;
        RECT 0.99 0.07 1.008 0.2 ;
        RECT 0.963 0.07 1.008 0.106 ;
        RECT 0.963 0.164 0.981 0.236 ;
        RECT 0.963 0.034 0.981 0.106 ;
        RECT 0.963 0.434 1.008 0.47 ;
        RECT 0.99 0.34 1.008 0.47 ;
        RECT 0.963 0.34 1.008 0.376 ;
        RECT 0.963 0.434 0.981 0.506 ;
        RECT 0.963 0.304 0.981 0.376 ;
      LAYER V2 ;
        RECT 1.017 0.452 1.035 0.47 ;
        RECT 1.017 0.07 1.035 0.088 ;
      LAYER V1 ;
        RECT 0.963 0.452 0.981 0.47 ;
        RECT 0.963 0.07 0.981 0.088 ;
        RECT 1.179 0.452 1.197 0.47 ;
        RECT 1.179 0.07 1.197 0.088 ;
    END
  END CLK
  OBS
    LAYER M1 ;
      RECT 1.93 0.225 2.034 0.243 ;
      RECT 2.016 0.027 2.034 0.243 ;
      RECT 1.854 0.027 1.872 0.119 ;
      RECT 1.854 0.027 2.034 0.045 ;
      RECT 1.854 0.495 2.034 0.513 ;
      RECT 2.016 0.297 2.034 0.513 ;
      RECT 1.854 0.421 1.872 0.513 ;
      RECT 1.93 0.297 2.034 0.315 ;
      RECT 1.768 0.224 1.818 0.242 ;
      RECT 1.8 0.027 1.818 0.242 ;
      RECT 1.8 0.153 1.98 0.171 ;
      RECT 1.962 0.117 1.98 0.171 ;
      RECT 1.908 0.117 1.926 0.171 ;
      RECT 1.714 0.027 1.818 0.045 ;
      RECT 1.714 0.495 1.818 0.513 ;
      RECT 1.8 0.298 1.818 0.513 ;
      RECT 1.962 0.369 1.98 0.423 ;
      RECT 1.908 0.369 1.926 0.423 ;
      RECT 1.8 0.369 1.98 0.387 ;
      RECT 1.768 0.298 1.818 0.316 ;
      RECT 1.656 0.225 1.71 0.243 ;
      RECT 1.692 0.081 1.71 0.243 ;
      RECT 1.576 0.081 1.71 0.099 ;
      RECT 1.665 0.045 1.683 0.099 ;
      RECT 1.665 0.441 1.683 0.495 ;
      RECT 1.576 0.441 1.71 0.459 ;
      RECT 1.692 0.297 1.71 0.459 ;
      RECT 1.656 0.297 1.71 0.315 ;
      RECT 1.444 0.225 1.548 0.243 ;
      RECT 1.53 0.027 1.548 0.243 ;
      RECT 1.53 0.122 1.656 0.14 ;
      RECT 1.498 0.027 1.548 0.045 ;
      RECT 1.498 0.495 1.548 0.513 ;
      RECT 1.53 0.297 1.548 0.513 ;
      RECT 1.53 0.4 1.656 0.418 ;
      RECT 1.444 0.297 1.548 0.315 ;
      RECT 1.395 0.126 1.413 0.203 ;
      RECT 1.395 0.126 1.447 0.144 ;
      RECT 1.395 0.396 1.447 0.414 ;
      RECT 1.395 0.337 1.413 0.414 ;
      RECT 1.228 0.225 1.278 0.243 ;
      RECT 1.26 0.027 1.278 0.243 ;
      RECT 1.228 0.027 1.278 0.045 ;
      RECT 1.228 0.495 1.278 0.513 ;
      RECT 1.26 0.297 1.278 0.513 ;
      RECT 1.228 0.297 1.278 0.315 ;
      RECT 1.089 0.225 1.148 0.243 ;
      RECT 1.089 0.027 1.107 0.243 ;
      RECT 1.089 0.144 1.127 0.162 ;
      RECT 1.089 0.027 1.148 0.045 ;
      RECT 1.089 0.495 1.148 0.513 ;
      RECT 1.089 0.297 1.107 0.513 ;
      RECT 1.089 0.378 1.127 0.396 ;
      RECT 1.089 0.297 1.148 0.315 ;
      RECT 1.012 0.225 1.071 0.243 ;
      RECT 1.053 0.027 1.071 0.243 ;
      RECT 1.033 0.144 1.071 0.162 ;
      RECT 1.012 0.027 1.071 0.045 ;
      RECT 1.012 0.495 1.071 0.513 ;
      RECT 1.053 0.297 1.071 0.513 ;
      RECT 1.033 0.378 1.071 0.396 ;
      RECT 1.012 0.297 1.071 0.315 ;
      RECT 0.882 0.225 0.932 0.243 ;
      RECT 0.882 0.027 0.9 0.243 ;
      RECT 0.882 0.027 0.932 0.045 ;
      RECT 0.882 0.495 0.932 0.513 ;
      RECT 0.882 0.297 0.9 0.513 ;
      RECT 0.882 0.297 0.932 0.315 ;
      RECT 0.747 0.126 0.765 0.203 ;
      RECT 0.713 0.126 0.765 0.144 ;
      RECT 0.713 0.396 0.765 0.414 ;
      RECT 0.747 0.337 0.765 0.414 ;
      RECT 0.612 0.225 0.716 0.243 ;
      RECT 0.612 0.027 0.63 0.243 ;
      RECT 0.504 0.122 0.63 0.14 ;
      RECT 0.612 0.027 0.662 0.045 ;
      RECT 0.612 0.495 0.662 0.513 ;
      RECT 0.612 0.297 0.63 0.513 ;
      RECT 0.504 0.4 0.63 0.418 ;
      RECT 0.612 0.297 0.716 0.315 ;
      RECT 0.45 0.225 0.504 0.243 ;
      RECT 0.45 0.081 0.468 0.243 ;
      RECT 0.45 0.081 0.584 0.099 ;
      RECT 0.477 0.045 0.495 0.099 ;
      RECT 0.477 0.441 0.495 0.495 ;
      RECT 0.45 0.441 0.584 0.459 ;
      RECT 0.45 0.297 0.468 0.459 ;
      RECT 0.45 0.297 0.504 0.315 ;
      RECT 0.342 0.224 0.392 0.242 ;
      RECT 0.342 0.027 0.36 0.242 ;
      RECT 0.18 0.153 0.36 0.171 ;
      RECT 0.234 0.117 0.252 0.171 ;
      RECT 0.18 0.117 0.198 0.171 ;
      RECT 0.342 0.027 0.446 0.045 ;
      RECT 0.342 0.495 0.446 0.513 ;
      RECT 0.342 0.298 0.36 0.513 ;
      RECT 0.234 0.369 0.252 0.423 ;
      RECT 0.18 0.369 0.198 0.423 ;
      RECT 0.18 0.369 0.36 0.387 ;
      RECT 0.342 0.298 0.392 0.316 ;
      RECT 0.126 0.225 0.23 0.243 ;
      RECT 0.126 0.027 0.144 0.243 ;
      RECT 0.288 0.027 0.306 0.119 ;
      RECT 0.126 0.027 0.306 0.045 ;
      RECT 0.126 0.495 0.306 0.513 ;
      RECT 0.288 0.421 0.306 0.513 ;
      RECT 0.126 0.297 0.144 0.513 ;
      RECT 0.126 0.297 0.23 0.315 ;
      RECT 2.07 0.09 2.088 0.167 ;
      RECT 2.07 0.373 2.088 0.45 ;
      RECT 1.746 0.101 1.764 0.167 ;
      RECT 1.746 0.373 1.764 0.439 ;
      RECT 1.584 0.165 1.602 0.203 ;
      RECT 1.584 0.337 1.602 0.375 ;
      RECT 1.476 0.106 1.494 0.167 ;
      RECT 1.476 0.373 1.494 0.434 ;
      RECT 1.222 0.106 1.24 0.167 ;
      RECT 1.222 0.373 1.24 0.434 ;
      RECT 0.92 0.106 0.938 0.167 ;
      RECT 0.92 0.373 0.938 0.434 ;
      RECT 0.666 0.106 0.684 0.167 ;
      RECT 0.666 0.373 0.684 0.434 ;
      RECT 0.558 0.165 0.576 0.203 ;
      RECT 0.558 0.337 0.576 0.375 ;
      RECT 0.396 0.101 0.414 0.167 ;
      RECT 0.396 0.373 0.414 0.439 ;
      RECT 0.072 0.09 0.09 0.167 ;
      RECT 0.072 0.373 0.09 0.45 ;
    LAYER M2 ;
      RECT 1.957 0.144 2.093 0.162 ;
      RECT 1.957 0.378 2.093 0.396 ;
      RECT 1.099 0.144 1.769 0.162 ;
      RECT 1.099 0.378 1.769 0.396 ;
      RECT 1.255 0.18 1.607 0.198 ;
      RECT 1.255 0.342 1.607 0.36 ;
      RECT 0.391 0.144 1.061 0.162 ;
      RECT 0.391 0.378 1.061 0.396 ;
      RECT 0.553 0.18 0.905 0.198 ;
      RECT 0.553 0.342 0.905 0.36 ;
      RECT 0.067 0.144 0.203 0.162 ;
      RECT 0.067 0.378 0.203 0.396 ;
    LAYER V1 ;
      RECT 2.07 0.144 2.088 0.162 ;
      RECT 2.07 0.378 2.088 0.396 ;
      RECT 1.962 0.144 1.98 0.162 ;
      RECT 1.962 0.378 1.98 0.396 ;
      RECT 1.746 0.144 1.764 0.162 ;
      RECT 1.746 0.378 1.764 0.396 ;
      RECT 1.584 0.18 1.602 0.198 ;
      RECT 1.584 0.342 1.602 0.36 ;
      RECT 1.476 0.144 1.494 0.162 ;
      RECT 1.476 0.378 1.494 0.396 ;
      RECT 1.395 0.18 1.413 0.198 ;
      RECT 1.395 0.342 1.413 0.36 ;
      RECT 1.26 0.18 1.278 0.198 ;
      RECT 1.26 0.342 1.278 0.36 ;
      RECT 1.222 0.144 1.24 0.162 ;
      RECT 1.222 0.378 1.24 0.396 ;
      RECT 1.104 0.144 1.122 0.162 ;
      RECT 1.104 0.378 1.122 0.396 ;
      RECT 1.038 0.144 1.056 0.162 ;
      RECT 1.038 0.378 1.056 0.396 ;
      RECT 0.92 0.144 0.938 0.162 ;
      RECT 0.92 0.378 0.938 0.396 ;
      RECT 0.882 0.18 0.9 0.198 ;
      RECT 0.882 0.342 0.9 0.36 ;
      RECT 0.747 0.18 0.765 0.198 ;
      RECT 0.747 0.342 0.765 0.36 ;
      RECT 0.666 0.144 0.684 0.162 ;
      RECT 0.666 0.378 0.684 0.396 ;
      RECT 0.558 0.18 0.576 0.198 ;
      RECT 0.558 0.342 0.576 0.36 ;
      RECT 0.396 0.144 0.414 0.162 ;
      RECT 0.396 0.378 0.414 0.396 ;
      RECT 0.18 0.144 0.198 0.162 ;
      RECT 0.18 0.378 0.198 0.396 ;
      RECT 0.072 0.144 0.09 0.162 ;
      RECT 0.072 0.378 0.09 0.396 ;
  END
END DFFHQNH2V2Xx1_ASAP7_75t_R

MACRO DFFHQNH2V2Xx1_ASAP7_75t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNH2V2Xx1_ASAP7_75t_SL 0 0 ;
  SIZE 2.16 BY 0.54 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t_pg ;
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.314 0.126 1.37 0.144 ;
        RECT 1.314 0.225 1.351 0.243 ;
        RECT 1.314 0.027 1.351 0.045 ;
        RECT 1.314 0.027 1.332 0.243 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.314 0.396 1.37 0.414 ;
        RECT 1.314 0.495 1.351 0.513 ;
        RECT 1.314 0.297 1.351 0.315 ;
        RECT 1.314 0.297 1.332 0.513 ;
    END
  END D1
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.809 0.225 0.846 0.243 ;
        RECT 0.828 0.027 0.846 0.243 ;
        RECT 0.79 0.126 0.846 0.144 ;
        RECT 0.809 0.027 0.846 0.045 ;
    END
  END D2
  PIN D3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.809 0.495 0.846 0.513 ;
        RECT 0.828 0.297 0.846 0.513 ;
        RECT 0.79 0.396 0.846 0.414 ;
        RECT 0.809 0.297 0.846 0.315 ;
    END
  END D3
  PIN QN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.092 0.225 2.142 0.243 ;
        RECT 2.124 0.027 2.142 0.243 ;
        RECT 2.092 0.027 2.142 0.045 ;
    END
  END QN0
  PIN QN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.092 0.495 2.142 0.513 ;
        RECT 2.124 0.297 2.142 0.513 ;
        RECT 2.092 0.297 2.142 0.315 ;
    END
  END QN1
  PIN QN2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.225 0.068 0.243 ;
        RECT 0.018 0.027 0.068 0.045 ;
        RECT 0.018 0.027 0.036 0.243 ;
    END
  END QN2
  PIN QN3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.495 0.068 0.513 ;
        RECT 0.018 0.297 0.068 0.315 ;
        RECT 0.018 0.297 0.036 0.513 ;
    END
  END QN3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 2.16 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 2.16 0.009 ;
        RECT 0 0.531 2.16 0.549 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 0.958 0.07 1.202 0.088 ;
        RECT 0.958 0.452 1.202 0.47 ;
      LAYER M3 ;
        RECT 1.017 0.05 1.035 0.492 ;
      LAYER M1 ;
        RECT 1.179 0.164 1.197 0.236 ;
        RECT 1.152 0.07 1.197 0.106 ;
        RECT 1.179 0.034 1.197 0.106 ;
        RECT 1.152 0.164 1.197 0.2 ;
        RECT 1.152 0.07 1.17 0.2 ;
        RECT 1.179 0.434 1.197 0.506 ;
        RECT 1.152 0.34 1.197 0.376 ;
        RECT 1.179 0.304 1.197 0.376 ;
        RECT 1.152 0.434 1.197 0.47 ;
        RECT 1.152 0.34 1.17 0.47 ;
        RECT 0.963 0.164 1.008 0.2 ;
        RECT 0.99 0.07 1.008 0.2 ;
        RECT 0.963 0.07 1.008 0.106 ;
        RECT 0.963 0.164 0.981 0.236 ;
        RECT 0.963 0.034 0.981 0.106 ;
        RECT 0.963 0.434 1.008 0.47 ;
        RECT 0.99 0.34 1.008 0.47 ;
        RECT 0.963 0.34 1.008 0.376 ;
        RECT 0.963 0.434 0.981 0.506 ;
        RECT 0.963 0.304 0.981 0.376 ;
      LAYER V2 ;
        RECT 1.017 0.452 1.035 0.47 ;
        RECT 1.017 0.07 1.035 0.088 ;
      LAYER V1 ;
        RECT 0.963 0.452 0.981 0.47 ;
        RECT 0.963 0.07 0.981 0.088 ;
        RECT 1.179 0.452 1.197 0.47 ;
        RECT 1.179 0.07 1.197 0.088 ;
    END
  END CLK
  OBS
    LAYER M1 ;
      RECT 1.93 0.225 2.034 0.243 ;
      RECT 2.016 0.027 2.034 0.243 ;
      RECT 1.854 0.027 1.872 0.119 ;
      RECT 1.854 0.027 2.034 0.045 ;
      RECT 1.854 0.495 2.034 0.513 ;
      RECT 2.016 0.297 2.034 0.513 ;
      RECT 1.854 0.421 1.872 0.513 ;
      RECT 1.93 0.297 2.034 0.315 ;
      RECT 1.768 0.224 1.818 0.242 ;
      RECT 1.8 0.027 1.818 0.242 ;
      RECT 1.8 0.153 1.98 0.171 ;
      RECT 1.962 0.117 1.98 0.171 ;
      RECT 1.908 0.117 1.926 0.171 ;
      RECT 1.714 0.027 1.818 0.045 ;
      RECT 1.714 0.495 1.818 0.513 ;
      RECT 1.8 0.298 1.818 0.513 ;
      RECT 1.962 0.369 1.98 0.423 ;
      RECT 1.908 0.369 1.926 0.423 ;
      RECT 1.8 0.369 1.98 0.387 ;
      RECT 1.768 0.298 1.818 0.316 ;
      RECT 1.656 0.225 1.71 0.243 ;
      RECT 1.692 0.081 1.71 0.243 ;
      RECT 1.576 0.081 1.71 0.099 ;
      RECT 1.665 0.045 1.683 0.099 ;
      RECT 1.665 0.441 1.683 0.495 ;
      RECT 1.576 0.441 1.71 0.459 ;
      RECT 1.692 0.297 1.71 0.459 ;
      RECT 1.656 0.297 1.71 0.315 ;
      RECT 1.444 0.225 1.548 0.243 ;
      RECT 1.53 0.027 1.548 0.243 ;
      RECT 1.53 0.122 1.656 0.14 ;
      RECT 1.498 0.027 1.548 0.045 ;
      RECT 1.498 0.495 1.548 0.513 ;
      RECT 1.53 0.297 1.548 0.513 ;
      RECT 1.53 0.4 1.656 0.418 ;
      RECT 1.444 0.297 1.548 0.315 ;
      RECT 1.395 0.126 1.413 0.203 ;
      RECT 1.395 0.126 1.447 0.144 ;
      RECT 1.395 0.396 1.447 0.414 ;
      RECT 1.395 0.337 1.413 0.414 ;
      RECT 1.228 0.225 1.278 0.243 ;
      RECT 1.26 0.027 1.278 0.243 ;
      RECT 1.228 0.027 1.278 0.045 ;
      RECT 1.228 0.495 1.278 0.513 ;
      RECT 1.26 0.297 1.278 0.513 ;
      RECT 1.228 0.297 1.278 0.315 ;
      RECT 1.089 0.225 1.148 0.243 ;
      RECT 1.089 0.027 1.107 0.243 ;
      RECT 1.089 0.144 1.127 0.162 ;
      RECT 1.089 0.027 1.148 0.045 ;
      RECT 1.089 0.495 1.148 0.513 ;
      RECT 1.089 0.297 1.107 0.513 ;
      RECT 1.089 0.378 1.127 0.396 ;
      RECT 1.089 0.297 1.148 0.315 ;
      RECT 1.012 0.225 1.071 0.243 ;
      RECT 1.053 0.027 1.071 0.243 ;
      RECT 1.033 0.144 1.071 0.162 ;
      RECT 1.012 0.027 1.071 0.045 ;
      RECT 1.012 0.495 1.071 0.513 ;
      RECT 1.053 0.297 1.071 0.513 ;
      RECT 1.033 0.378 1.071 0.396 ;
      RECT 1.012 0.297 1.071 0.315 ;
      RECT 0.882 0.225 0.932 0.243 ;
      RECT 0.882 0.027 0.9 0.243 ;
      RECT 0.882 0.027 0.932 0.045 ;
      RECT 0.882 0.495 0.932 0.513 ;
      RECT 0.882 0.297 0.9 0.513 ;
      RECT 0.882 0.297 0.932 0.315 ;
      RECT 0.747 0.126 0.765 0.203 ;
      RECT 0.713 0.126 0.765 0.144 ;
      RECT 0.713 0.396 0.765 0.414 ;
      RECT 0.747 0.337 0.765 0.414 ;
      RECT 0.612 0.225 0.716 0.243 ;
      RECT 0.612 0.027 0.63 0.243 ;
      RECT 0.504 0.122 0.63 0.14 ;
      RECT 0.612 0.027 0.662 0.045 ;
      RECT 0.612 0.495 0.662 0.513 ;
      RECT 0.612 0.297 0.63 0.513 ;
      RECT 0.504 0.4 0.63 0.418 ;
      RECT 0.612 0.297 0.716 0.315 ;
      RECT 0.45 0.225 0.504 0.243 ;
      RECT 0.45 0.081 0.468 0.243 ;
      RECT 0.45 0.081 0.584 0.099 ;
      RECT 0.477 0.045 0.495 0.099 ;
      RECT 0.477 0.441 0.495 0.495 ;
      RECT 0.45 0.441 0.584 0.459 ;
      RECT 0.45 0.297 0.468 0.459 ;
      RECT 0.45 0.297 0.504 0.315 ;
      RECT 0.342 0.224 0.392 0.242 ;
      RECT 0.342 0.027 0.36 0.242 ;
      RECT 0.18 0.153 0.36 0.171 ;
      RECT 0.234 0.117 0.252 0.171 ;
      RECT 0.18 0.117 0.198 0.171 ;
      RECT 0.342 0.027 0.446 0.045 ;
      RECT 0.342 0.495 0.446 0.513 ;
      RECT 0.342 0.298 0.36 0.513 ;
      RECT 0.234 0.369 0.252 0.423 ;
      RECT 0.18 0.369 0.198 0.423 ;
      RECT 0.18 0.369 0.36 0.387 ;
      RECT 0.342 0.298 0.392 0.316 ;
      RECT 0.126 0.225 0.23 0.243 ;
      RECT 0.126 0.027 0.144 0.243 ;
      RECT 0.288 0.027 0.306 0.119 ;
      RECT 0.126 0.027 0.306 0.045 ;
      RECT 0.126 0.495 0.306 0.513 ;
      RECT 0.288 0.421 0.306 0.513 ;
      RECT 0.126 0.297 0.144 0.513 ;
      RECT 0.126 0.297 0.23 0.315 ;
      RECT 2.07 0.09 2.088 0.167 ;
      RECT 2.07 0.373 2.088 0.45 ;
      RECT 1.746 0.101 1.764 0.167 ;
      RECT 1.746 0.373 1.764 0.439 ;
      RECT 1.584 0.165 1.602 0.203 ;
      RECT 1.584 0.337 1.602 0.375 ;
      RECT 1.476 0.106 1.494 0.167 ;
      RECT 1.476 0.373 1.494 0.434 ;
      RECT 1.222 0.106 1.24 0.167 ;
      RECT 1.222 0.373 1.24 0.434 ;
      RECT 0.92 0.106 0.938 0.167 ;
      RECT 0.92 0.373 0.938 0.434 ;
      RECT 0.666 0.106 0.684 0.167 ;
      RECT 0.666 0.373 0.684 0.434 ;
      RECT 0.558 0.165 0.576 0.203 ;
      RECT 0.558 0.337 0.576 0.375 ;
      RECT 0.396 0.101 0.414 0.167 ;
      RECT 0.396 0.373 0.414 0.439 ;
      RECT 0.072 0.09 0.09 0.167 ;
      RECT 0.072 0.373 0.09 0.45 ;
    LAYER M2 ;
      RECT 1.957 0.144 2.093 0.162 ;
      RECT 1.957 0.378 2.093 0.396 ;
      RECT 1.099 0.144 1.769 0.162 ;
      RECT 1.099 0.378 1.769 0.396 ;
      RECT 1.255 0.18 1.607 0.198 ;
      RECT 1.255 0.342 1.607 0.36 ;
      RECT 0.391 0.144 1.061 0.162 ;
      RECT 0.391 0.378 1.061 0.396 ;
      RECT 0.553 0.18 0.905 0.198 ;
      RECT 0.553 0.342 0.905 0.36 ;
      RECT 0.067 0.144 0.203 0.162 ;
      RECT 0.067 0.378 0.203 0.396 ;
    LAYER V1 ;
      RECT 2.07 0.144 2.088 0.162 ;
      RECT 2.07 0.378 2.088 0.396 ;
      RECT 1.962 0.144 1.98 0.162 ;
      RECT 1.962 0.378 1.98 0.396 ;
      RECT 1.746 0.144 1.764 0.162 ;
      RECT 1.746 0.378 1.764 0.396 ;
      RECT 1.584 0.18 1.602 0.198 ;
      RECT 1.584 0.342 1.602 0.36 ;
      RECT 1.476 0.144 1.494 0.162 ;
      RECT 1.476 0.378 1.494 0.396 ;
      RECT 1.395 0.18 1.413 0.198 ;
      RECT 1.395 0.342 1.413 0.36 ;
      RECT 1.26 0.18 1.278 0.198 ;
      RECT 1.26 0.342 1.278 0.36 ;
      RECT 1.222 0.144 1.24 0.162 ;
      RECT 1.222 0.378 1.24 0.396 ;
      RECT 1.104 0.144 1.122 0.162 ;
      RECT 1.104 0.378 1.122 0.396 ;
      RECT 1.038 0.144 1.056 0.162 ;
      RECT 1.038 0.378 1.056 0.396 ;
      RECT 0.92 0.144 0.938 0.162 ;
      RECT 0.92 0.378 0.938 0.396 ;
      RECT 0.882 0.18 0.9 0.198 ;
      RECT 0.882 0.342 0.9 0.36 ;
      RECT 0.747 0.18 0.765 0.198 ;
      RECT 0.747 0.342 0.765 0.36 ;
      RECT 0.666 0.144 0.684 0.162 ;
      RECT 0.666 0.378 0.684 0.396 ;
      RECT 0.558 0.18 0.576 0.198 ;
      RECT 0.558 0.342 0.576 0.36 ;
      RECT 0.396 0.144 0.414 0.162 ;
      RECT 0.396 0.378 0.414 0.396 ;
      RECT 0.18 0.144 0.198 0.162 ;
      RECT 0.18 0.378 0.198 0.396 ;
      RECT 0.072 0.144 0.09 0.162 ;
      RECT 0.072 0.378 0.09 0.396 ;
  END
END DFFHQNH2V2Xx1_ASAP7_75t_SL

MACRO DFFHQNH2V2Xx2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNH2V2Xx2_ASAP7_75t_L 0 0 ;
  SIZE 2.268 BY 0.54 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t_pg ;
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.126 1.424 0.144 ;
        RECT 1.368 0.225 1.405 0.243 ;
        RECT 1.368 0.027 1.405 0.045 ;
        RECT 1.368 0.027 1.386 0.243 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.396 1.424 0.414 ;
        RECT 1.368 0.495 1.405 0.513 ;
        RECT 1.368 0.297 1.405 0.315 ;
        RECT 1.368 0.297 1.386 0.513 ;
    END
  END D1
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.863 0.225 0.9 0.243 ;
        RECT 0.882 0.027 0.9 0.243 ;
        RECT 0.844 0.126 0.9 0.144 ;
        RECT 0.863 0.027 0.9 0.045 ;
    END
  END D2
  PIN D3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.863 0.495 0.9 0.513 ;
        RECT 0.882 0.297 0.9 0.513 ;
        RECT 0.844 0.396 0.9 0.414 ;
        RECT 0.863 0.297 0.9 0.315 ;
    END
  END D3
  PIN QN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.146 0.216 2.251 0.234 ;
        RECT 2.233 0.036 2.251 0.234 ;
        RECT 2.146 0.036 2.251 0.054 ;
    END
  END QN0
  PIN QN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.146 0.486 2.251 0.504 ;
        RECT 2.233 0.306 2.251 0.504 ;
        RECT 2.146 0.306 2.251 0.324 ;
    END
  END QN1
  PIN QN2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.017 0.216 0.122 0.234 ;
        RECT 0.017 0.036 0.122 0.054 ;
        RECT 0.017 0.036 0.035 0.234 ;
    END
  END QN2
  PIN QN3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.017 0.486 0.122 0.504 ;
        RECT 0.017 0.306 0.122 0.324 ;
        RECT 0.017 0.306 0.035 0.504 ;
    END
  END QN3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 2.268 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 2.268 0.009 ;
        RECT 0 0.531 2.268 0.549 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 1.012 0.07 1.256 0.088 ;
        RECT 1.012 0.452 1.256 0.47 ;
      LAYER M3 ;
        RECT 1.071 0.05 1.089 0.492 ;
      LAYER M1 ;
        RECT 1.233 0.164 1.251 0.236 ;
        RECT 1.206 0.07 1.251 0.106 ;
        RECT 1.233 0.034 1.251 0.106 ;
        RECT 1.206 0.164 1.251 0.2 ;
        RECT 1.206 0.07 1.224 0.2 ;
        RECT 1.233 0.434 1.251 0.506 ;
        RECT 1.206 0.34 1.251 0.376 ;
        RECT 1.233 0.304 1.251 0.376 ;
        RECT 1.206 0.434 1.251 0.47 ;
        RECT 1.206 0.34 1.224 0.47 ;
        RECT 1.017 0.164 1.062 0.2 ;
        RECT 1.044 0.07 1.062 0.2 ;
        RECT 1.017 0.07 1.062 0.106 ;
        RECT 1.017 0.164 1.035 0.236 ;
        RECT 1.017 0.034 1.035 0.106 ;
        RECT 1.017 0.434 1.062 0.47 ;
        RECT 1.044 0.34 1.062 0.47 ;
        RECT 1.017 0.34 1.062 0.376 ;
        RECT 1.017 0.434 1.035 0.506 ;
        RECT 1.017 0.304 1.035 0.376 ;
      LAYER V2 ;
        RECT 1.071 0.452 1.089 0.47 ;
        RECT 1.071 0.07 1.089 0.088 ;
      LAYER V1 ;
        RECT 1.017 0.452 1.035 0.47 ;
        RECT 1.017 0.07 1.035 0.088 ;
        RECT 1.233 0.452 1.251 0.47 ;
        RECT 1.233 0.07 1.251 0.088 ;
    END
  END CLK
  OBS
    LAYER M1 ;
      RECT 1.984 0.225 2.088 0.243 ;
      RECT 2.07 0.027 2.088 0.243 ;
      RECT 1.908 0.027 1.926 0.119 ;
      RECT 1.908 0.027 2.088 0.045 ;
      RECT 1.908 0.495 2.088 0.513 ;
      RECT 2.07 0.297 2.088 0.513 ;
      RECT 1.908 0.421 1.926 0.513 ;
      RECT 1.984 0.297 2.088 0.315 ;
      RECT 1.822 0.224 1.872 0.242 ;
      RECT 1.854 0.027 1.872 0.242 ;
      RECT 1.854 0.153 2.034 0.171 ;
      RECT 2.016 0.117 2.034 0.171 ;
      RECT 1.962 0.117 1.98 0.171 ;
      RECT 1.768 0.027 1.872 0.045 ;
      RECT 1.768 0.495 1.872 0.513 ;
      RECT 1.854 0.298 1.872 0.513 ;
      RECT 2.016 0.369 2.034 0.423 ;
      RECT 1.962 0.369 1.98 0.423 ;
      RECT 1.854 0.369 2.034 0.387 ;
      RECT 1.822 0.298 1.872 0.316 ;
      RECT 1.71 0.225 1.764 0.243 ;
      RECT 1.746 0.081 1.764 0.243 ;
      RECT 1.63 0.081 1.764 0.099 ;
      RECT 1.719 0.045 1.737 0.099 ;
      RECT 1.719 0.441 1.737 0.495 ;
      RECT 1.63 0.441 1.764 0.459 ;
      RECT 1.746 0.297 1.764 0.459 ;
      RECT 1.71 0.297 1.764 0.315 ;
      RECT 1.498 0.225 1.602 0.243 ;
      RECT 1.584 0.027 1.602 0.243 ;
      RECT 1.584 0.122 1.71 0.14 ;
      RECT 1.552 0.027 1.602 0.045 ;
      RECT 1.552 0.495 1.602 0.513 ;
      RECT 1.584 0.297 1.602 0.513 ;
      RECT 1.584 0.4 1.71 0.418 ;
      RECT 1.498 0.297 1.602 0.315 ;
      RECT 1.449 0.126 1.467 0.203 ;
      RECT 1.449 0.126 1.501 0.144 ;
      RECT 1.449 0.396 1.501 0.414 ;
      RECT 1.449 0.337 1.467 0.414 ;
      RECT 1.282 0.225 1.332 0.243 ;
      RECT 1.314 0.027 1.332 0.243 ;
      RECT 1.282 0.027 1.332 0.045 ;
      RECT 1.282 0.495 1.332 0.513 ;
      RECT 1.314 0.297 1.332 0.513 ;
      RECT 1.282 0.297 1.332 0.315 ;
      RECT 1.143 0.225 1.202 0.243 ;
      RECT 1.143 0.027 1.161 0.243 ;
      RECT 1.143 0.144 1.181 0.162 ;
      RECT 1.143 0.027 1.202 0.045 ;
      RECT 1.143 0.495 1.202 0.513 ;
      RECT 1.143 0.297 1.161 0.513 ;
      RECT 1.143 0.378 1.181 0.396 ;
      RECT 1.143 0.297 1.202 0.315 ;
      RECT 1.066 0.225 1.125 0.243 ;
      RECT 1.107 0.027 1.125 0.243 ;
      RECT 1.087 0.144 1.125 0.162 ;
      RECT 1.066 0.027 1.125 0.045 ;
      RECT 1.066 0.495 1.125 0.513 ;
      RECT 1.107 0.297 1.125 0.513 ;
      RECT 1.087 0.378 1.125 0.396 ;
      RECT 1.066 0.297 1.125 0.315 ;
      RECT 0.936 0.225 0.986 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.936 0.027 0.986 0.045 ;
      RECT 0.936 0.495 0.986 0.513 ;
      RECT 0.936 0.297 0.954 0.513 ;
      RECT 0.936 0.297 0.986 0.315 ;
      RECT 0.801 0.126 0.819 0.203 ;
      RECT 0.767 0.126 0.819 0.144 ;
      RECT 0.767 0.396 0.819 0.414 ;
      RECT 0.801 0.337 0.819 0.414 ;
      RECT 0.666 0.225 0.77 0.243 ;
      RECT 0.666 0.027 0.684 0.243 ;
      RECT 0.558 0.122 0.684 0.14 ;
      RECT 0.666 0.027 0.716 0.045 ;
      RECT 0.666 0.495 0.716 0.513 ;
      RECT 0.666 0.297 0.684 0.513 ;
      RECT 0.558 0.4 0.684 0.418 ;
      RECT 0.666 0.297 0.77 0.315 ;
      RECT 0.504 0.225 0.558 0.243 ;
      RECT 0.504 0.081 0.522 0.243 ;
      RECT 0.504 0.081 0.638 0.099 ;
      RECT 0.531 0.045 0.549 0.099 ;
      RECT 0.531 0.441 0.549 0.495 ;
      RECT 0.504 0.441 0.638 0.459 ;
      RECT 0.504 0.297 0.522 0.459 ;
      RECT 0.504 0.297 0.558 0.315 ;
      RECT 0.396 0.224 0.446 0.242 ;
      RECT 0.396 0.027 0.414 0.242 ;
      RECT 0.234 0.153 0.414 0.171 ;
      RECT 0.288 0.117 0.306 0.171 ;
      RECT 0.234 0.117 0.252 0.171 ;
      RECT 0.396 0.027 0.5 0.045 ;
      RECT 0.396 0.495 0.5 0.513 ;
      RECT 0.396 0.298 0.414 0.513 ;
      RECT 0.288 0.369 0.306 0.423 ;
      RECT 0.234 0.369 0.252 0.423 ;
      RECT 0.234 0.369 0.414 0.387 ;
      RECT 0.396 0.298 0.446 0.316 ;
      RECT 0.18 0.225 0.284 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.342 0.027 0.36 0.119 ;
      RECT 0.18 0.027 0.36 0.045 ;
      RECT 0.18 0.495 0.36 0.513 ;
      RECT 0.342 0.421 0.36 0.513 ;
      RECT 0.18 0.297 0.198 0.513 ;
      RECT 0.18 0.297 0.284 0.315 ;
      RECT 2.124 0.09 2.142 0.167 ;
      RECT 2.124 0.373 2.142 0.45 ;
      RECT 1.8 0.101 1.818 0.167 ;
      RECT 1.8 0.373 1.818 0.439 ;
      RECT 1.638 0.165 1.656 0.203 ;
      RECT 1.638 0.337 1.656 0.375 ;
      RECT 1.53 0.106 1.548 0.167 ;
      RECT 1.53 0.373 1.548 0.434 ;
      RECT 1.276 0.106 1.294 0.167 ;
      RECT 1.276 0.373 1.294 0.434 ;
      RECT 0.974 0.106 0.992 0.167 ;
      RECT 0.974 0.373 0.992 0.434 ;
      RECT 0.72 0.106 0.738 0.167 ;
      RECT 0.72 0.373 0.738 0.434 ;
      RECT 0.612 0.165 0.63 0.203 ;
      RECT 0.612 0.337 0.63 0.375 ;
      RECT 0.45 0.101 0.468 0.167 ;
      RECT 0.45 0.373 0.468 0.439 ;
      RECT 0.126 0.09 0.144 0.167 ;
      RECT 0.126 0.373 0.144 0.45 ;
    LAYER M2 ;
      RECT 2.011 0.144 2.147 0.162 ;
      RECT 2.011 0.378 2.147 0.396 ;
      RECT 1.153 0.144 1.823 0.162 ;
      RECT 1.153 0.378 1.823 0.396 ;
      RECT 1.309 0.18 1.661 0.198 ;
      RECT 1.309 0.342 1.661 0.36 ;
      RECT 0.445 0.144 1.115 0.162 ;
      RECT 0.445 0.378 1.115 0.396 ;
      RECT 0.607 0.18 0.959 0.198 ;
      RECT 0.607 0.342 0.959 0.36 ;
      RECT 0.121 0.144 0.257 0.162 ;
      RECT 0.121 0.378 0.257 0.396 ;
    LAYER V1 ;
      RECT 2.124 0.144 2.142 0.162 ;
      RECT 2.124 0.378 2.142 0.396 ;
      RECT 2.016 0.144 2.034 0.162 ;
      RECT 2.016 0.378 2.034 0.396 ;
      RECT 1.8 0.144 1.818 0.162 ;
      RECT 1.8 0.378 1.818 0.396 ;
      RECT 1.638 0.18 1.656 0.198 ;
      RECT 1.638 0.342 1.656 0.36 ;
      RECT 1.53 0.144 1.548 0.162 ;
      RECT 1.53 0.378 1.548 0.396 ;
      RECT 1.449 0.18 1.467 0.198 ;
      RECT 1.449 0.342 1.467 0.36 ;
      RECT 1.314 0.18 1.332 0.198 ;
      RECT 1.314 0.342 1.332 0.36 ;
      RECT 1.276 0.144 1.294 0.162 ;
      RECT 1.276 0.378 1.294 0.396 ;
      RECT 1.158 0.144 1.176 0.162 ;
      RECT 1.158 0.378 1.176 0.396 ;
      RECT 1.092 0.144 1.11 0.162 ;
      RECT 1.092 0.378 1.11 0.396 ;
      RECT 0.974 0.144 0.992 0.162 ;
      RECT 0.974 0.378 0.992 0.396 ;
      RECT 0.936 0.18 0.954 0.198 ;
      RECT 0.936 0.342 0.954 0.36 ;
      RECT 0.801 0.18 0.819 0.198 ;
      RECT 0.801 0.342 0.819 0.36 ;
      RECT 0.72 0.144 0.738 0.162 ;
      RECT 0.72 0.378 0.738 0.396 ;
      RECT 0.612 0.18 0.63 0.198 ;
      RECT 0.612 0.342 0.63 0.36 ;
      RECT 0.45 0.144 0.468 0.162 ;
      RECT 0.45 0.378 0.468 0.396 ;
      RECT 0.234 0.144 0.252 0.162 ;
      RECT 0.234 0.378 0.252 0.396 ;
      RECT 0.126 0.144 0.144 0.162 ;
      RECT 0.126 0.378 0.144 0.396 ;
  END
END DFFHQNH2V2Xx2_ASAP7_75t_L

MACRO DFFHQNH2V2Xx2_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNH2V2Xx2_ASAP7_75t_R 0 0 ;
  SIZE 2.268 BY 0.54 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t_pg ;
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.126 1.424 0.144 ;
        RECT 1.368 0.225 1.405 0.243 ;
        RECT 1.368 0.027 1.405 0.045 ;
        RECT 1.368 0.027 1.386 0.243 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.396 1.424 0.414 ;
        RECT 1.368 0.495 1.405 0.513 ;
        RECT 1.368 0.297 1.405 0.315 ;
        RECT 1.368 0.297 1.386 0.513 ;
    END
  END D1
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.863 0.225 0.9 0.243 ;
        RECT 0.882 0.027 0.9 0.243 ;
        RECT 0.844 0.126 0.9 0.144 ;
        RECT 0.863 0.027 0.9 0.045 ;
    END
  END D2
  PIN D3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.863 0.495 0.9 0.513 ;
        RECT 0.882 0.297 0.9 0.513 ;
        RECT 0.844 0.396 0.9 0.414 ;
        RECT 0.863 0.297 0.9 0.315 ;
    END
  END D3
  PIN QN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.146 0.216 2.251 0.234 ;
        RECT 2.233 0.036 2.251 0.234 ;
        RECT 2.146 0.036 2.251 0.054 ;
    END
  END QN0
  PIN QN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.146 0.486 2.251 0.504 ;
        RECT 2.233 0.306 2.251 0.504 ;
        RECT 2.146 0.306 2.251 0.324 ;
    END
  END QN1
  PIN QN2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.017 0.216 0.122 0.234 ;
        RECT 0.017 0.036 0.122 0.054 ;
        RECT 0.017 0.036 0.035 0.234 ;
    END
  END QN2
  PIN QN3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.017 0.486 0.122 0.504 ;
        RECT 0.017 0.306 0.122 0.324 ;
        RECT 0.017 0.306 0.035 0.504 ;
    END
  END QN3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 2.268 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 2.268 0.009 ;
        RECT 0 0.531 2.268 0.549 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 1.012 0.07 1.256 0.088 ;
        RECT 1.012 0.452 1.256 0.47 ;
      LAYER M3 ;
        RECT 1.071 0.05 1.089 0.492 ;
      LAYER M1 ;
        RECT 1.233 0.164 1.251 0.236 ;
        RECT 1.206 0.07 1.251 0.106 ;
        RECT 1.233 0.034 1.251 0.106 ;
        RECT 1.206 0.164 1.251 0.2 ;
        RECT 1.206 0.07 1.224 0.2 ;
        RECT 1.233 0.434 1.251 0.506 ;
        RECT 1.206 0.34 1.251 0.376 ;
        RECT 1.233 0.304 1.251 0.376 ;
        RECT 1.206 0.434 1.251 0.47 ;
        RECT 1.206 0.34 1.224 0.47 ;
        RECT 1.017 0.164 1.062 0.2 ;
        RECT 1.044 0.07 1.062 0.2 ;
        RECT 1.017 0.07 1.062 0.106 ;
        RECT 1.017 0.164 1.035 0.236 ;
        RECT 1.017 0.034 1.035 0.106 ;
        RECT 1.017 0.434 1.062 0.47 ;
        RECT 1.044 0.34 1.062 0.47 ;
        RECT 1.017 0.34 1.062 0.376 ;
        RECT 1.017 0.434 1.035 0.506 ;
        RECT 1.017 0.304 1.035 0.376 ;
      LAYER V2 ;
        RECT 1.071 0.452 1.089 0.47 ;
        RECT 1.071 0.07 1.089 0.088 ;
      LAYER V1 ;
        RECT 1.017 0.452 1.035 0.47 ;
        RECT 1.017 0.07 1.035 0.088 ;
        RECT 1.233 0.452 1.251 0.47 ;
        RECT 1.233 0.07 1.251 0.088 ;
    END
  END CLK
  OBS
    LAYER M1 ;
      RECT 1.984 0.225 2.088 0.243 ;
      RECT 2.07 0.027 2.088 0.243 ;
      RECT 1.908 0.027 1.926 0.119 ;
      RECT 1.908 0.027 2.088 0.045 ;
      RECT 1.908 0.495 2.088 0.513 ;
      RECT 2.07 0.297 2.088 0.513 ;
      RECT 1.908 0.421 1.926 0.513 ;
      RECT 1.984 0.297 2.088 0.315 ;
      RECT 1.822 0.224 1.872 0.242 ;
      RECT 1.854 0.027 1.872 0.242 ;
      RECT 1.854 0.153 2.034 0.171 ;
      RECT 2.016 0.117 2.034 0.171 ;
      RECT 1.962 0.117 1.98 0.171 ;
      RECT 1.768 0.027 1.872 0.045 ;
      RECT 1.768 0.495 1.872 0.513 ;
      RECT 1.854 0.298 1.872 0.513 ;
      RECT 2.016 0.369 2.034 0.423 ;
      RECT 1.962 0.369 1.98 0.423 ;
      RECT 1.854 0.369 2.034 0.387 ;
      RECT 1.822 0.298 1.872 0.316 ;
      RECT 1.71 0.225 1.764 0.243 ;
      RECT 1.746 0.081 1.764 0.243 ;
      RECT 1.63 0.081 1.764 0.099 ;
      RECT 1.719 0.045 1.737 0.099 ;
      RECT 1.719 0.441 1.737 0.495 ;
      RECT 1.63 0.441 1.764 0.459 ;
      RECT 1.746 0.297 1.764 0.459 ;
      RECT 1.71 0.297 1.764 0.315 ;
      RECT 1.498 0.225 1.602 0.243 ;
      RECT 1.584 0.027 1.602 0.243 ;
      RECT 1.584 0.122 1.71 0.14 ;
      RECT 1.552 0.027 1.602 0.045 ;
      RECT 1.552 0.495 1.602 0.513 ;
      RECT 1.584 0.297 1.602 0.513 ;
      RECT 1.584 0.4 1.71 0.418 ;
      RECT 1.498 0.297 1.602 0.315 ;
      RECT 1.449 0.126 1.467 0.203 ;
      RECT 1.449 0.126 1.501 0.144 ;
      RECT 1.449 0.396 1.501 0.414 ;
      RECT 1.449 0.337 1.467 0.414 ;
      RECT 1.282 0.225 1.332 0.243 ;
      RECT 1.314 0.027 1.332 0.243 ;
      RECT 1.282 0.027 1.332 0.045 ;
      RECT 1.282 0.495 1.332 0.513 ;
      RECT 1.314 0.297 1.332 0.513 ;
      RECT 1.282 0.297 1.332 0.315 ;
      RECT 1.143 0.225 1.202 0.243 ;
      RECT 1.143 0.027 1.161 0.243 ;
      RECT 1.143 0.144 1.181 0.162 ;
      RECT 1.143 0.027 1.202 0.045 ;
      RECT 1.143 0.495 1.202 0.513 ;
      RECT 1.143 0.297 1.161 0.513 ;
      RECT 1.143 0.378 1.181 0.396 ;
      RECT 1.143 0.297 1.202 0.315 ;
      RECT 1.066 0.225 1.125 0.243 ;
      RECT 1.107 0.027 1.125 0.243 ;
      RECT 1.087 0.144 1.125 0.162 ;
      RECT 1.066 0.027 1.125 0.045 ;
      RECT 1.066 0.495 1.125 0.513 ;
      RECT 1.107 0.297 1.125 0.513 ;
      RECT 1.087 0.378 1.125 0.396 ;
      RECT 1.066 0.297 1.125 0.315 ;
      RECT 0.936 0.225 0.986 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.936 0.027 0.986 0.045 ;
      RECT 0.936 0.495 0.986 0.513 ;
      RECT 0.936 0.297 0.954 0.513 ;
      RECT 0.936 0.297 0.986 0.315 ;
      RECT 0.801 0.126 0.819 0.203 ;
      RECT 0.767 0.126 0.819 0.144 ;
      RECT 0.767 0.396 0.819 0.414 ;
      RECT 0.801 0.337 0.819 0.414 ;
      RECT 0.666 0.225 0.77 0.243 ;
      RECT 0.666 0.027 0.684 0.243 ;
      RECT 0.558 0.122 0.684 0.14 ;
      RECT 0.666 0.027 0.716 0.045 ;
      RECT 0.666 0.495 0.716 0.513 ;
      RECT 0.666 0.297 0.684 0.513 ;
      RECT 0.558 0.4 0.684 0.418 ;
      RECT 0.666 0.297 0.77 0.315 ;
      RECT 0.504 0.225 0.558 0.243 ;
      RECT 0.504 0.081 0.522 0.243 ;
      RECT 0.504 0.081 0.638 0.099 ;
      RECT 0.531 0.045 0.549 0.099 ;
      RECT 0.531 0.441 0.549 0.495 ;
      RECT 0.504 0.441 0.638 0.459 ;
      RECT 0.504 0.297 0.522 0.459 ;
      RECT 0.504 0.297 0.558 0.315 ;
      RECT 0.396 0.224 0.446 0.242 ;
      RECT 0.396 0.027 0.414 0.242 ;
      RECT 0.234 0.153 0.414 0.171 ;
      RECT 0.288 0.117 0.306 0.171 ;
      RECT 0.234 0.117 0.252 0.171 ;
      RECT 0.396 0.027 0.5 0.045 ;
      RECT 0.396 0.495 0.5 0.513 ;
      RECT 0.396 0.298 0.414 0.513 ;
      RECT 0.288 0.369 0.306 0.423 ;
      RECT 0.234 0.369 0.252 0.423 ;
      RECT 0.234 0.369 0.414 0.387 ;
      RECT 0.396 0.298 0.446 0.316 ;
      RECT 0.18 0.225 0.284 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.342 0.027 0.36 0.119 ;
      RECT 0.18 0.027 0.36 0.045 ;
      RECT 0.18 0.495 0.36 0.513 ;
      RECT 0.342 0.421 0.36 0.513 ;
      RECT 0.18 0.297 0.198 0.513 ;
      RECT 0.18 0.297 0.284 0.315 ;
      RECT 2.124 0.09 2.142 0.167 ;
      RECT 2.124 0.373 2.142 0.45 ;
      RECT 1.8 0.101 1.818 0.167 ;
      RECT 1.8 0.373 1.818 0.439 ;
      RECT 1.638 0.165 1.656 0.203 ;
      RECT 1.638 0.337 1.656 0.375 ;
      RECT 1.53 0.106 1.548 0.167 ;
      RECT 1.53 0.373 1.548 0.434 ;
      RECT 1.276 0.106 1.294 0.167 ;
      RECT 1.276 0.373 1.294 0.434 ;
      RECT 0.974 0.106 0.992 0.167 ;
      RECT 0.974 0.373 0.992 0.434 ;
      RECT 0.72 0.106 0.738 0.167 ;
      RECT 0.72 0.373 0.738 0.434 ;
      RECT 0.612 0.165 0.63 0.203 ;
      RECT 0.612 0.337 0.63 0.375 ;
      RECT 0.45 0.101 0.468 0.167 ;
      RECT 0.45 0.373 0.468 0.439 ;
      RECT 0.126 0.09 0.144 0.167 ;
      RECT 0.126 0.373 0.144 0.45 ;
    LAYER M2 ;
      RECT 2.011 0.144 2.147 0.162 ;
      RECT 2.011 0.378 2.147 0.396 ;
      RECT 1.153 0.144 1.823 0.162 ;
      RECT 1.153 0.378 1.823 0.396 ;
      RECT 1.309 0.18 1.661 0.198 ;
      RECT 1.309 0.342 1.661 0.36 ;
      RECT 0.445 0.144 1.115 0.162 ;
      RECT 0.445 0.378 1.115 0.396 ;
      RECT 0.607 0.18 0.959 0.198 ;
      RECT 0.607 0.342 0.959 0.36 ;
      RECT 0.121 0.144 0.257 0.162 ;
      RECT 0.121 0.378 0.257 0.396 ;
    LAYER V1 ;
      RECT 2.124 0.144 2.142 0.162 ;
      RECT 2.124 0.378 2.142 0.396 ;
      RECT 2.016 0.144 2.034 0.162 ;
      RECT 2.016 0.378 2.034 0.396 ;
      RECT 1.8 0.144 1.818 0.162 ;
      RECT 1.8 0.378 1.818 0.396 ;
      RECT 1.638 0.18 1.656 0.198 ;
      RECT 1.638 0.342 1.656 0.36 ;
      RECT 1.53 0.144 1.548 0.162 ;
      RECT 1.53 0.378 1.548 0.396 ;
      RECT 1.449 0.18 1.467 0.198 ;
      RECT 1.449 0.342 1.467 0.36 ;
      RECT 1.314 0.18 1.332 0.198 ;
      RECT 1.314 0.342 1.332 0.36 ;
      RECT 1.276 0.144 1.294 0.162 ;
      RECT 1.276 0.378 1.294 0.396 ;
      RECT 1.158 0.144 1.176 0.162 ;
      RECT 1.158 0.378 1.176 0.396 ;
      RECT 1.092 0.144 1.11 0.162 ;
      RECT 1.092 0.378 1.11 0.396 ;
      RECT 0.974 0.144 0.992 0.162 ;
      RECT 0.974 0.378 0.992 0.396 ;
      RECT 0.936 0.18 0.954 0.198 ;
      RECT 0.936 0.342 0.954 0.36 ;
      RECT 0.801 0.18 0.819 0.198 ;
      RECT 0.801 0.342 0.819 0.36 ;
      RECT 0.72 0.144 0.738 0.162 ;
      RECT 0.72 0.378 0.738 0.396 ;
      RECT 0.612 0.18 0.63 0.198 ;
      RECT 0.612 0.342 0.63 0.36 ;
      RECT 0.45 0.144 0.468 0.162 ;
      RECT 0.45 0.378 0.468 0.396 ;
      RECT 0.234 0.144 0.252 0.162 ;
      RECT 0.234 0.378 0.252 0.396 ;
      RECT 0.126 0.144 0.144 0.162 ;
      RECT 0.126 0.378 0.144 0.396 ;
  END
END DFFHQNH2V2Xx2_ASAP7_75t_R

MACRO DFFHQNH2V2Xx2_ASAP7_75t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNH2V2Xx2_ASAP7_75t_SL 0 0 ;
  SIZE 2.268 BY 0.54 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t_pg ;
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.126 1.424 0.144 ;
        RECT 1.368 0.225 1.405 0.243 ;
        RECT 1.368 0.027 1.405 0.045 ;
        RECT 1.368 0.027 1.386 0.243 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.396 1.424 0.414 ;
        RECT 1.368 0.495 1.405 0.513 ;
        RECT 1.368 0.297 1.405 0.315 ;
        RECT 1.368 0.297 1.386 0.513 ;
    END
  END D1
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.863 0.225 0.9 0.243 ;
        RECT 0.882 0.027 0.9 0.243 ;
        RECT 0.844 0.126 0.9 0.144 ;
        RECT 0.863 0.027 0.9 0.045 ;
    END
  END D2
  PIN D3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.863 0.495 0.9 0.513 ;
        RECT 0.882 0.297 0.9 0.513 ;
        RECT 0.844 0.396 0.9 0.414 ;
        RECT 0.863 0.297 0.9 0.315 ;
    END
  END D3
  PIN QN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.146 0.216 2.251 0.234 ;
        RECT 2.233 0.036 2.251 0.234 ;
        RECT 2.146 0.036 2.251 0.054 ;
    END
  END QN0
  PIN QN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.146 0.486 2.251 0.504 ;
        RECT 2.233 0.306 2.251 0.504 ;
        RECT 2.146 0.306 2.251 0.324 ;
    END
  END QN1
  PIN QN2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.017 0.216 0.122 0.234 ;
        RECT 0.017 0.036 0.122 0.054 ;
        RECT 0.017 0.036 0.035 0.234 ;
    END
  END QN2
  PIN QN3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.017 0.486 0.122 0.504 ;
        RECT 0.017 0.306 0.122 0.324 ;
        RECT 0.017 0.306 0.035 0.504 ;
    END
  END QN3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 2.268 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 2.268 0.009 ;
        RECT 0 0.531 2.268 0.549 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 1.012 0.07 1.256 0.088 ;
        RECT 1.012 0.452 1.256 0.47 ;
      LAYER M3 ;
        RECT 1.071 0.05 1.089 0.492 ;
      LAYER M1 ;
        RECT 1.233 0.164 1.251 0.236 ;
        RECT 1.206 0.07 1.251 0.106 ;
        RECT 1.233 0.034 1.251 0.106 ;
        RECT 1.206 0.164 1.251 0.2 ;
        RECT 1.206 0.07 1.224 0.2 ;
        RECT 1.233 0.434 1.251 0.506 ;
        RECT 1.206 0.34 1.251 0.376 ;
        RECT 1.233 0.304 1.251 0.376 ;
        RECT 1.206 0.434 1.251 0.47 ;
        RECT 1.206 0.34 1.224 0.47 ;
        RECT 1.017 0.164 1.062 0.2 ;
        RECT 1.044 0.07 1.062 0.2 ;
        RECT 1.017 0.07 1.062 0.106 ;
        RECT 1.017 0.164 1.035 0.236 ;
        RECT 1.017 0.034 1.035 0.106 ;
        RECT 1.017 0.434 1.062 0.47 ;
        RECT 1.044 0.34 1.062 0.47 ;
        RECT 1.017 0.34 1.062 0.376 ;
        RECT 1.017 0.434 1.035 0.506 ;
        RECT 1.017 0.304 1.035 0.376 ;
      LAYER V2 ;
        RECT 1.071 0.452 1.089 0.47 ;
        RECT 1.071 0.07 1.089 0.088 ;
      LAYER V1 ;
        RECT 1.017 0.452 1.035 0.47 ;
        RECT 1.017 0.07 1.035 0.088 ;
        RECT 1.233 0.452 1.251 0.47 ;
        RECT 1.233 0.07 1.251 0.088 ;
    END
  END CLK
  OBS
    LAYER M1 ;
      RECT 1.984 0.225 2.088 0.243 ;
      RECT 2.07 0.027 2.088 0.243 ;
      RECT 1.908 0.027 1.926 0.119 ;
      RECT 1.908 0.027 2.088 0.045 ;
      RECT 1.908 0.495 2.088 0.513 ;
      RECT 2.07 0.297 2.088 0.513 ;
      RECT 1.908 0.421 1.926 0.513 ;
      RECT 1.984 0.297 2.088 0.315 ;
      RECT 1.822 0.224 1.872 0.242 ;
      RECT 1.854 0.027 1.872 0.242 ;
      RECT 1.854 0.153 2.034 0.171 ;
      RECT 2.016 0.117 2.034 0.171 ;
      RECT 1.962 0.117 1.98 0.171 ;
      RECT 1.768 0.027 1.872 0.045 ;
      RECT 1.768 0.495 1.872 0.513 ;
      RECT 1.854 0.298 1.872 0.513 ;
      RECT 2.016 0.369 2.034 0.423 ;
      RECT 1.962 0.369 1.98 0.423 ;
      RECT 1.854 0.369 2.034 0.387 ;
      RECT 1.822 0.298 1.872 0.316 ;
      RECT 1.71 0.225 1.764 0.243 ;
      RECT 1.746 0.081 1.764 0.243 ;
      RECT 1.63 0.081 1.764 0.099 ;
      RECT 1.719 0.045 1.737 0.099 ;
      RECT 1.719 0.441 1.737 0.495 ;
      RECT 1.63 0.441 1.764 0.459 ;
      RECT 1.746 0.297 1.764 0.459 ;
      RECT 1.71 0.297 1.764 0.315 ;
      RECT 1.498 0.225 1.602 0.243 ;
      RECT 1.584 0.027 1.602 0.243 ;
      RECT 1.584 0.122 1.71 0.14 ;
      RECT 1.552 0.027 1.602 0.045 ;
      RECT 1.552 0.495 1.602 0.513 ;
      RECT 1.584 0.297 1.602 0.513 ;
      RECT 1.584 0.4 1.71 0.418 ;
      RECT 1.498 0.297 1.602 0.315 ;
      RECT 1.449 0.126 1.467 0.203 ;
      RECT 1.449 0.126 1.501 0.144 ;
      RECT 1.449 0.396 1.501 0.414 ;
      RECT 1.449 0.337 1.467 0.414 ;
      RECT 1.282 0.225 1.332 0.243 ;
      RECT 1.314 0.027 1.332 0.243 ;
      RECT 1.282 0.027 1.332 0.045 ;
      RECT 1.282 0.495 1.332 0.513 ;
      RECT 1.314 0.297 1.332 0.513 ;
      RECT 1.282 0.297 1.332 0.315 ;
      RECT 1.143 0.225 1.202 0.243 ;
      RECT 1.143 0.027 1.161 0.243 ;
      RECT 1.143 0.144 1.181 0.162 ;
      RECT 1.143 0.027 1.202 0.045 ;
      RECT 1.143 0.495 1.202 0.513 ;
      RECT 1.143 0.297 1.161 0.513 ;
      RECT 1.143 0.378 1.181 0.396 ;
      RECT 1.143 0.297 1.202 0.315 ;
      RECT 1.066 0.225 1.125 0.243 ;
      RECT 1.107 0.027 1.125 0.243 ;
      RECT 1.087 0.144 1.125 0.162 ;
      RECT 1.066 0.027 1.125 0.045 ;
      RECT 1.066 0.495 1.125 0.513 ;
      RECT 1.107 0.297 1.125 0.513 ;
      RECT 1.087 0.378 1.125 0.396 ;
      RECT 1.066 0.297 1.125 0.315 ;
      RECT 0.936 0.225 0.986 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.936 0.027 0.986 0.045 ;
      RECT 0.936 0.495 0.986 0.513 ;
      RECT 0.936 0.297 0.954 0.513 ;
      RECT 0.936 0.297 0.986 0.315 ;
      RECT 0.801 0.126 0.819 0.203 ;
      RECT 0.767 0.126 0.819 0.144 ;
      RECT 0.767 0.396 0.819 0.414 ;
      RECT 0.801 0.337 0.819 0.414 ;
      RECT 0.666 0.225 0.77 0.243 ;
      RECT 0.666 0.027 0.684 0.243 ;
      RECT 0.558 0.122 0.684 0.14 ;
      RECT 0.666 0.027 0.716 0.045 ;
      RECT 0.666 0.495 0.716 0.513 ;
      RECT 0.666 0.297 0.684 0.513 ;
      RECT 0.558 0.4 0.684 0.418 ;
      RECT 0.666 0.297 0.77 0.315 ;
      RECT 0.504 0.225 0.558 0.243 ;
      RECT 0.504 0.081 0.522 0.243 ;
      RECT 0.504 0.081 0.638 0.099 ;
      RECT 0.531 0.045 0.549 0.099 ;
      RECT 0.531 0.441 0.549 0.495 ;
      RECT 0.504 0.441 0.638 0.459 ;
      RECT 0.504 0.297 0.522 0.459 ;
      RECT 0.504 0.297 0.558 0.315 ;
      RECT 0.396 0.224 0.446 0.242 ;
      RECT 0.396 0.027 0.414 0.242 ;
      RECT 0.234 0.153 0.414 0.171 ;
      RECT 0.288 0.117 0.306 0.171 ;
      RECT 0.234 0.117 0.252 0.171 ;
      RECT 0.396 0.027 0.5 0.045 ;
      RECT 0.396 0.495 0.5 0.513 ;
      RECT 0.396 0.298 0.414 0.513 ;
      RECT 0.288 0.369 0.306 0.423 ;
      RECT 0.234 0.369 0.252 0.423 ;
      RECT 0.234 0.369 0.414 0.387 ;
      RECT 0.396 0.298 0.446 0.316 ;
      RECT 0.18 0.225 0.284 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.342 0.027 0.36 0.119 ;
      RECT 0.18 0.027 0.36 0.045 ;
      RECT 0.18 0.495 0.36 0.513 ;
      RECT 0.342 0.421 0.36 0.513 ;
      RECT 0.18 0.297 0.198 0.513 ;
      RECT 0.18 0.297 0.284 0.315 ;
      RECT 2.124 0.09 2.142 0.167 ;
      RECT 2.124 0.373 2.142 0.45 ;
      RECT 1.8 0.101 1.818 0.167 ;
      RECT 1.8 0.373 1.818 0.439 ;
      RECT 1.638 0.165 1.656 0.203 ;
      RECT 1.638 0.337 1.656 0.375 ;
      RECT 1.53 0.106 1.548 0.167 ;
      RECT 1.53 0.373 1.548 0.434 ;
      RECT 1.276 0.106 1.294 0.167 ;
      RECT 1.276 0.373 1.294 0.434 ;
      RECT 0.974 0.106 0.992 0.167 ;
      RECT 0.974 0.373 0.992 0.434 ;
      RECT 0.72 0.106 0.738 0.167 ;
      RECT 0.72 0.373 0.738 0.434 ;
      RECT 0.612 0.165 0.63 0.203 ;
      RECT 0.612 0.337 0.63 0.375 ;
      RECT 0.45 0.101 0.468 0.167 ;
      RECT 0.45 0.373 0.468 0.439 ;
      RECT 0.126 0.09 0.144 0.167 ;
      RECT 0.126 0.373 0.144 0.45 ;
    LAYER M2 ;
      RECT 2.011 0.144 2.147 0.162 ;
      RECT 2.011 0.378 2.147 0.396 ;
      RECT 1.153 0.144 1.823 0.162 ;
      RECT 1.153 0.378 1.823 0.396 ;
      RECT 1.309 0.18 1.661 0.198 ;
      RECT 1.309 0.342 1.661 0.36 ;
      RECT 0.445 0.144 1.115 0.162 ;
      RECT 0.445 0.378 1.115 0.396 ;
      RECT 0.607 0.18 0.959 0.198 ;
      RECT 0.607 0.342 0.959 0.36 ;
      RECT 0.121 0.144 0.257 0.162 ;
      RECT 0.121 0.378 0.257 0.396 ;
    LAYER V1 ;
      RECT 2.124 0.144 2.142 0.162 ;
      RECT 2.124 0.378 2.142 0.396 ;
      RECT 2.016 0.144 2.034 0.162 ;
      RECT 2.016 0.378 2.034 0.396 ;
      RECT 1.8 0.144 1.818 0.162 ;
      RECT 1.8 0.378 1.818 0.396 ;
      RECT 1.638 0.18 1.656 0.198 ;
      RECT 1.638 0.342 1.656 0.36 ;
      RECT 1.53 0.144 1.548 0.162 ;
      RECT 1.53 0.378 1.548 0.396 ;
      RECT 1.449 0.18 1.467 0.198 ;
      RECT 1.449 0.342 1.467 0.36 ;
      RECT 1.314 0.18 1.332 0.198 ;
      RECT 1.314 0.342 1.332 0.36 ;
      RECT 1.276 0.144 1.294 0.162 ;
      RECT 1.276 0.378 1.294 0.396 ;
      RECT 1.158 0.144 1.176 0.162 ;
      RECT 1.158 0.378 1.176 0.396 ;
      RECT 1.092 0.144 1.11 0.162 ;
      RECT 1.092 0.378 1.11 0.396 ;
      RECT 0.974 0.144 0.992 0.162 ;
      RECT 0.974 0.378 0.992 0.396 ;
      RECT 0.936 0.18 0.954 0.198 ;
      RECT 0.936 0.342 0.954 0.36 ;
      RECT 0.801 0.18 0.819 0.198 ;
      RECT 0.801 0.342 0.819 0.36 ;
      RECT 0.72 0.144 0.738 0.162 ;
      RECT 0.72 0.378 0.738 0.396 ;
      RECT 0.612 0.18 0.63 0.198 ;
      RECT 0.612 0.342 0.63 0.36 ;
      RECT 0.45 0.144 0.468 0.162 ;
      RECT 0.45 0.378 0.468 0.396 ;
      RECT 0.234 0.144 0.252 0.162 ;
      RECT 0.234 0.378 0.252 0.396 ;
      RECT 0.126 0.144 0.144 0.162 ;
      RECT 0.126 0.378 0.144 0.396 ;
  END
END DFFHQNH2V2Xx2_ASAP7_75t_SL

MACRO DFFHQNH2V2Xx3_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNH2V2Xx3_ASAP7_75t_L 0 0 ;
  SIZE 2.376 BY 0.54 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t_pg ;
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.422 0.126 1.478 0.144 ;
        RECT 1.422 0.225 1.459 0.243 ;
        RECT 1.422 0.027 1.459 0.045 ;
        RECT 1.422 0.027 1.44 0.243 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.422 0.396 1.478 0.414 ;
        RECT 1.422 0.495 1.459 0.513 ;
        RECT 1.422 0.297 1.459 0.315 ;
        RECT 1.422 0.297 1.44 0.513 ;
    END
  END D1
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.917 0.225 0.954 0.243 ;
        RECT 0.936 0.027 0.954 0.243 ;
        RECT 0.898 0.126 0.954 0.144 ;
        RECT 0.917 0.027 0.954 0.045 ;
    END
  END D2
  PIN D3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.917 0.495 0.954 0.513 ;
        RECT 0.936 0.297 0.954 0.513 ;
        RECT 0.898 0.396 0.954 0.414 ;
        RECT 0.917 0.297 0.954 0.315 ;
    END
  END D3
  PIN QN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2 0.225 2.359 0.243 ;
        RECT 2.341 0.027 2.359 0.243 ;
        RECT 2.2 0.027 2.359 0.045 ;
    END
  END QN0
  PIN QN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2 0.495 2.359 0.513 ;
        RECT 2.341 0.297 2.359 0.513 ;
        RECT 2.2 0.297 2.359 0.315 ;
    END
  END QN1
  PIN QN2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.017 0.225 0.176 0.243 ;
        RECT 0.017 0.027 0.176 0.045 ;
        RECT 0.017 0.027 0.035 0.243 ;
    END
  END QN2
  PIN QN3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.017 0.495 0.176 0.513 ;
        RECT 0.017 0.297 0.176 0.315 ;
        RECT 0.017 0.297 0.035 0.513 ;
    END
  END QN3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 2.376 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 2.376 0.009 ;
        RECT 0 0.531 2.376 0.549 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 1.066 0.07 1.31 0.088 ;
        RECT 1.066 0.452 1.31 0.47 ;
      LAYER M3 ;
        RECT 1.125 0.05 1.143 0.492 ;
      LAYER M1 ;
        RECT 1.287 0.164 1.305 0.236 ;
        RECT 1.26 0.07 1.305 0.106 ;
        RECT 1.287 0.034 1.305 0.106 ;
        RECT 1.26 0.164 1.305 0.2 ;
        RECT 1.26 0.07 1.278 0.2 ;
        RECT 1.287 0.434 1.305 0.506 ;
        RECT 1.26 0.34 1.305 0.376 ;
        RECT 1.287 0.304 1.305 0.376 ;
        RECT 1.26 0.434 1.305 0.47 ;
        RECT 1.26 0.34 1.278 0.47 ;
        RECT 1.071 0.164 1.116 0.2 ;
        RECT 1.098 0.07 1.116 0.2 ;
        RECT 1.071 0.07 1.116 0.106 ;
        RECT 1.071 0.164 1.089 0.236 ;
        RECT 1.071 0.034 1.089 0.106 ;
        RECT 1.071 0.434 1.116 0.47 ;
        RECT 1.098 0.34 1.116 0.47 ;
        RECT 1.071 0.34 1.116 0.376 ;
        RECT 1.071 0.434 1.089 0.506 ;
        RECT 1.071 0.304 1.089 0.376 ;
      LAYER V2 ;
        RECT 1.125 0.452 1.143 0.47 ;
        RECT 1.125 0.07 1.143 0.088 ;
      LAYER V1 ;
        RECT 1.071 0.452 1.089 0.47 ;
        RECT 1.071 0.07 1.089 0.088 ;
        RECT 1.287 0.452 1.305 0.47 ;
        RECT 1.287 0.07 1.305 0.088 ;
    END
  END CLK
  OBS
    LAYER M1 ;
      RECT 2.038 0.225 2.142 0.243 ;
      RECT 2.124 0.027 2.142 0.243 ;
      RECT 1.962 0.027 1.98 0.119 ;
      RECT 1.962 0.027 2.142 0.045 ;
      RECT 1.962 0.495 2.142 0.513 ;
      RECT 2.124 0.297 2.142 0.513 ;
      RECT 1.962 0.421 1.98 0.513 ;
      RECT 2.038 0.297 2.142 0.315 ;
      RECT 1.876 0.224 1.926 0.242 ;
      RECT 1.908 0.027 1.926 0.242 ;
      RECT 1.908 0.153 2.088 0.171 ;
      RECT 2.07 0.117 2.088 0.171 ;
      RECT 2.016 0.117 2.034 0.171 ;
      RECT 1.822 0.027 1.926 0.045 ;
      RECT 1.822 0.495 1.926 0.513 ;
      RECT 1.908 0.298 1.926 0.513 ;
      RECT 2.07 0.369 2.088 0.423 ;
      RECT 2.016 0.369 2.034 0.423 ;
      RECT 1.908 0.369 2.088 0.387 ;
      RECT 1.876 0.298 1.926 0.316 ;
      RECT 1.764 0.225 1.818 0.243 ;
      RECT 1.8 0.081 1.818 0.243 ;
      RECT 1.684 0.081 1.818 0.099 ;
      RECT 1.773 0.045 1.791 0.099 ;
      RECT 1.773 0.441 1.791 0.495 ;
      RECT 1.684 0.441 1.818 0.459 ;
      RECT 1.8 0.297 1.818 0.459 ;
      RECT 1.764 0.297 1.818 0.315 ;
      RECT 1.552 0.225 1.656 0.243 ;
      RECT 1.638 0.027 1.656 0.243 ;
      RECT 1.638 0.122 1.764 0.14 ;
      RECT 1.606 0.027 1.656 0.045 ;
      RECT 1.606 0.495 1.656 0.513 ;
      RECT 1.638 0.297 1.656 0.513 ;
      RECT 1.638 0.4 1.764 0.418 ;
      RECT 1.552 0.297 1.656 0.315 ;
      RECT 1.503 0.126 1.521 0.203 ;
      RECT 1.503 0.126 1.555 0.144 ;
      RECT 1.503 0.396 1.555 0.414 ;
      RECT 1.503 0.337 1.521 0.414 ;
      RECT 1.336 0.225 1.386 0.243 ;
      RECT 1.368 0.027 1.386 0.243 ;
      RECT 1.336 0.027 1.386 0.045 ;
      RECT 1.336 0.495 1.386 0.513 ;
      RECT 1.368 0.297 1.386 0.513 ;
      RECT 1.336 0.297 1.386 0.315 ;
      RECT 1.197 0.225 1.256 0.243 ;
      RECT 1.197 0.027 1.215 0.243 ;
      RECT 1.197 0.144 1.235 0.162 ;
      RECT 1.197 0.027 1.256 0.045 ;
      RECT 1.197 0.495 1.256 0.513 ;
      RECT 1.197 0.297 1.215 0.513 ;
      RECT 1.197 0.378 1.235 0.396 ;
      RECT 1.197 0.297 1.256 0.315 ;
      RECT 1.12 0.225 1.179 0.243 ;
      RECT 1.161 0.027 1.179 0.243 ;
      RECT 1.141 0.144 1.179 0.162 ;
      RECT 1.12 0.027 1.179 0.045 ;
      RECT 1.12 0.495 1.179 0.513 ;
      RECT 1.161 0.297 1.179 0.513 ;
      RECT 1.141 0.378 1.179 0.396 ;
      RECT 1.12 0.297 1.179 0.315 ;
      RECT 0.99 0.225 1.04 0.243 ;
      RECT 0.99 0.027 1.008 0.243 ;
      RECT 0.99 0.027 1.04 0.045 ;
      RECT 0.99 0.495 1.04 0.513 ;
      RECT 0.99 0.297 1.008 0.513 ;
      RECT 0.99 0.297 1.04 0.315 ;
      RECT 0.855 0.126 0.873 0.203 ;
      RECT 0.821 0.126 0.873 0.144 ;
      RECT 0.821 0.396 0.873 0.414 ;
      RECT 0.855 0.337 0.873 0.414 ;
      RECT 0.72 0.225 0.824 0.243 ;
      RECT 0.72 0.027 0.738 0.243 ;
      RECT 0.612 0.122 0.738 0.14 ;
      RECT 0.72 0.027 0.77 0.045 ;
      RECT 0.72 0.495 0.77 0.513 ;
      RECT 0.72 0.297 0.738 0.513 ;
      RECT 0.612 0.4 0.738 0.418 ;
      RECT 0.72 0.297 0.824 0.315 ;
      RECT 0.558 0.225 0.612 0.243 ;
      RECT 0.558 0.081 0.576 0.243 ;
      RECT 0.558 0.081 0.692 0.099 ;
      RECT 0.585 0.045 0.603 0.099 ;
      RECT 0.585 0.441 0.603 0.495 ;
      RECT 0.558 0.441 0.692 0.459 ;
      RECT 0.558 0.297 0.576 0.459 ;
      RECT 0.558 0.297 0.612 0.315 ;
      RECT 0.45 0.224 0.5 0.242 ;
      RECT 0.45 0.027 0.468 0.242 ;
      RECT 0.288 0.153 0.468 0.171 ;
      RECT 0.342 0.117 0.36 0.171 ;
      RECT 0.288 0.117 0.306 0.171 ;
      RECT 0.45 0.027 0.554 0.045 ;
      RECT 0.45 0.495 0.554 0.513 ;
      RECT 0.45 0.298 0.468 0.513 ;
      RECT 0.342 0.369 0.36 0.423 ;
      RECT 0.288 0.369 0.306 0.423 ;
      RECT 0.288 0.369 0.468 0.387 ;
      RECT 0.45 0.298 0.5 0.316 ;
      RECT 0.234 0.225 0.338 0.243 ;
      RECT 0.234 0.027 0.252 0.243 ;
      RECT 0.396 0.027 0.414 0.119 ;
      RECT 0.234 0.027 0.414 0.045 ;
      RECT 0.234 0.495 0.414 0.513 ;
      RECT 0.396 0.421 0.414 0.513 ;
      RECT 0.234 0.297 0.252 0.513 ;
      RECT 0.234 0.297 0.338 0.315 ;
      RECT 2.178 0.122 2.196 0.167 ;
      RECT 2.178 0.373 2.196 0.418 ;
      RECT 1.854 0.101 1.872 0.167 ;
      RECT 1.854 0.373 1.872 0.439 ;
      RECT 1.692 0.165 1.71 0.203 ;
      RECT 1.692 0.337 1.71 0.375 ;
      RECT 1.584 0.106 1.602 0.167 ;
      RECT 1.584 0.373 1.602 0.434 ;
      RECT 1.33 0.106 1.348 0.167 ;
      RECT 1.33 0.373 1.348 0.434 ;
      RECT 1.028 0.106 1.046 0.167 ;
      RECT 1.028 0.373 1.046 0.434 ;
      RECT 0.774 0.106 0.792 0.167 ;
      RECT 0.774 0.373 0.792 0.434 ;
      RECT 0.666 0.165 0.684 0.203 ;
      RECT 0.666 0.337 0.684 0.375 ;
      RECT 0.504 0.101 0.522 0.167 ;
      RECT 0.504 0.373 0.522 0.439 ;
      RECT 0.18 0.122 0.198 0.167 ;
      RECT 0.18 0.373 0.198 0.418 ;
    LAYER M2 ;
      RECT 2.065 0.144 2.201 0.162 ;
      RECT 2.065 0.378 2.201 0.396 ;
      RECT 1.207 0.144 1.877 0.162 ;
      RECT 1.207 0.378 1.877 0.396 ;
      RECT 1.363 0.18 1.715 0.198 ;
      RECT 1.363 0.342 1.715 0.36 ;
      RECT 0.499 0.144 1.169 0.162 ;
      RECT 0.499 0.378 1.169 0.396 ;
      RECT 0.661 0.18 1.013 0.198 ;
      RECT 0.661 0.342 1.013 0.36 ;
      RECT 0.175 0.144 0.311 0.162 ;
      RECT 0.175 0.378 0.311 0.396 ;
    LAYER V1 ;
      RECT 2.178 0.144 2.196 0.162 ;
      RECT 2.178 0.378 2.196 0.396 ;
      RECT 2.07 0.144 2.088 0.162 ;
      RECT 2.07 0.378 2.088 0.396 ;
      RECT 1.854 0.144 1.872 0.162 ;
      RECT 1.854 0.378 1.872 0.396 ;
      RECT 1.692 0.18 1.71 0.198 ;
      RECT 1.692 0.342 1.71 0.36 ;
      RECT 1.584 0.144 1.602 0.162 ;
      RECT 1.584 0.378 1.602 0.396 ;
      RECT 1.503 0.18 1.521 0.198 ;
      RECT 1.503 0.342 1.521 0.36 ;
      RECT 1.368 0.18 1.386 0.198 ;
      RECT 1.368 0.342 1.386 0.36 ;
      RECT 1.33 0.144 1.348 0.162 ;
      RECT 1.33 0.378 1.348 0.396 ;
      RECT 1.212 0.144 1.23 0.162 ;
      RECT 1.212 0.378 1.23 0.396 ;
      RECT 1.146 0.144 1.164 0.162 ;
      RECT 1.146 0.378 1.164 0.396 ;
      RECT 1.028 0.144 1.046 0.162 ;
      RECT 1.028 0.378 1.046 0.396 ;
      RECT 0.99 0.18 1.008 0.198 ;
      RECT 0.99 0.342 1.008 0.36 ;
      RECT 0.855 0.18 0.873 0.198 ;
      RECT 0.855 0.342 0.873 0.36 ;
      RECT 0.774 0.144 0.792 0.162 ;
      RECT 0.774 0.378 0.792 0.396 ;
      RECT 0.666 0.18 0.684 0.198 ;
      RECT 0.666 0.342 0.684 0.36 ;
      RECT 0.504 0.144 0.522 0.162 ;
      RECT 0.504 0.378 0.522 0.396 ;
      RECT 0.288 0.144 0.306 0.162 ;
      RECT 0.288 0.378 0.306 0.396 ;
      RECT 0.18 0.144 0.198 0.162 ;
      RECT 0.18 0.378 0.198 0.396 ;
  END
END DFFHQNH2V2Xx3_ASAP7_75t_L

MACRO DFFHQNH2V2Xx3_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNH2V2Xx3_ASAP7_75t_R 0 0 ;
  SIZE 2.376 BY 0.54 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t_pg ;
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.422 0.126 1.478 0.144 ;
        RECT 1.422 0.225 1.459 0.243 ;
        RECT 1.422 0.027 1.459 0.045 ;
        RECT 1.422 0.027 1.44 0.243 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.422 0.396 1.478 0.414 ;
        RECT 1.422 0.495 1.459 0.513 ;
        RECT 1.422 0.297 1.459 0.315 ;
        RECT 1.422 0.297 1.44 0.513 ;
    END
  END D1
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.917 0.225 0.954 0.243 ;
        RECT 0.936 0.027 0.954 0.243 ;
        RECT 0.898 0.126 0.954 0.144 ;
        RECT 0.917 0.027 0.954 0.045 ;
    END
  END D2
  PIN D3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.917 0.495 0.954 0.513 ;
        RECT 0.936 0.297 0.954 0.513 ;
        RECT 0.898 0.396 0.954 0.414 ;
        RECT 0.917 0.297 0.954 0.315 ;
    END
  END D3
  PIN QN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2 0.225 2.359 0.243 ;
        RECT 2.341 0.027 2.359 0.243 ;
        RECT 2.2 0.027 2.359 0.045 ;
    END
  END QN0
  PIN QN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2 0.495 2.359 0.513 ;
        RECT 2.341 0.297 2.359 0.513 ;
        RECT 2.2 0.297 2.359 0.315 ;
    END
  END QN1
  PIN QN2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.017 0.225 0.176 0.243 ;
        RECT 0.017 0.027 0.176 0.045 ;
        RECT 0.017 0.027 0.035 0.243 ;
    END
  END QN2
  PIN QN3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.017 0.495 0.176 0.513 ;
        RECT 0.017 0.297 0.176 0.315 ;
        RECT 0.017 0.297 0.035 0.513 ;
    END
  END QN3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 2.376 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 2.376 0.009 ;
        RECT 0 0.531 2.376 0.549 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 1.066 0.07 1.31 0.088 ;
        RECT 1.066 0.452 1.31 0.47 ;
      LAYER M3 ;
        RECT 1.125 0.05 1.143 0.492 ;
      LAYER M1 ;
        RECT 1.287 0.164 1.305 0.236 ;
        RECT 1.26 0.07 1.305 0.106 ;
        RECT 1.287 0.034 1.305 0.106 ;
        RECT 1.26 0.164 1.305 0.2 ;
        RECT 1.26 0.07 1.278 0.2 ;
        RECT 1.287 0.434 1.305 0.506 ;
        RECT 1.26 0.34 1.305 0.376 ;
        RECT 1.287 0.304 1.305 0.376 ;
        RECT 1.26 0.434 1.305 0.47 ;
        RECT 1.26 0.34 1.278 0.47 ;
        RECT 1.071 0.164 1.116 0.2 ;
        RECT 1.098 0.07 1.116 0.2 ;
        RECT 1.071 0.07 1.116 0.106 ;
        RECT 1.071 0.164 1.089 0.236 ;
        RECT 1.071 0.034 1.089 0.106 ;
        RECT 1.071 0.434 1.116 0.47 ;
        RECT 1.098 0.34 1.116 0.47 ;
        RECT 1.071 0.34 1.116 0.376 ;
        RECT 1.071 0.434 1.089 0.506 ;
        RECT 1.071 0.304 1.089 0.376 ;
      LAYER V2 ;
        RECT 1.125 0.452 1.143 0.47 ;
        RECT 1.125 0.07 1.143 0.088 ;
      LAYER V1 ;
        RECT 1.071 0.452 1.089 0.47 ;
        RECT 1.071 0.07 1.089 0.088 ;
        RECT 1.287 0.452 1.305 0.47 ;
        RECT 1.287 0.07 1.305 0.088 ;
    END
  END CLK
  OBS
    LAYER M1 ;
      RECT 2.038 0.225 2.142 0.243 ;
      RECT 2.124 0.027 2.142 0.243 ;
      RECT 1.962 0.027 1.98 0.119 ;
      RECT 1.962 0.027 2.142 0.045 ;
      RECT 1.962 0.495 2.142 0.513 ;
      RECT 2.124 0.297 2.142 0.513 ;
      RECT 1.962 0.421 1.98 0.513 ;
      RECT 2.038 0.297 2.142 0.315 ;
      RECT 1.876 0.224 1.926 0.242 ;
      RECT 1.908 0.027 1.926 0.242 ;
      RECT 1.908 0.153 2.088 0.171 ;
      RECT 2.07 0.117 2.088 0.171 ;
      RECT 2.016 0.117 2.034 0.171 ;
      RECT 1.822 0.027 1.926 0.045 ;
      RECT 1.822 0.495 1.926 0.513 ;
      RECT 1.908 0.298 1.926 0.513 ;
      RECT 2.07 0.369 2.088 0.423 ;
      RECT 2.016 0.369 2.034 0.423 ;
      RECT 1.908 0.369 2.088 0.387 ;
      RECT 1.876 0.298 1.926 0.316 ;
      RECT 1.764 0.225 1.818 0.243 ;
      RECT 1.8 0.081 1.818 0.243 ;
      RECT 1.684 0.081 1.818 0.099 ;
      RECT 1.773 0.045 1.791 0.099 ;
      RECT 1.773 0.441 1.791 0.495 ;
      RECT 1.684 0.441 1.818 0.459 ;
      RECT 1.8 0.297 1.818 0.459 ;
      RECT 1.764 0.297 1.818 0.315 ;
      RECT 1.552 0.225 1.656 0.243 ;
      RECT 1.638 0.027 1.656 0.243 ;
      RECT 1.638 0.122 1.764 0.14 ;
      RECT 1.606 0.027 1.656 0.045 ;
      RECT 1.606 0.495 1.656 0.513 ;
      RECT 1.638 0.297 1.656 0.513 ;
      RECT 1.638 0.4 1.764 0.418 ;
      RECT 1.552 0.297 1.656 0.315 ;
      RECT 1.503 0.126 1.521 0.203 ;
      RECT 1.503 0.126 1.555 0.144 ;
      RECT 1.503 0.396 1.555 0.414 ;
      RECT 1.503 0.337 1.521 0.414 ;
      RECT 1.336 0.225 1.386 0.243 ;
      RECT 1.368 0.027 1.386 0.243 ;
      RECT 1.336 0.027 1.386 0.045 ;
      RECT 1.336 0.495 1.386 0.513 ;
      RECT 1.368 0.297 1.386 0.513 ;
      RECT 1.336 0.297 1.386 0.315 ;
      RECT 1.197 0.225 1.256 0.243 ;
      RECT 1.197 0.027 1.215 0.243 ;
      RECT 1.197 0.144 1.235 0.162 ;
      RECT 1.197 0.027 1.256 0.045 ;
      RECT 1.197 0.495 1.256 0.513 ;
      RECT 1.197 0.297 1.215 0.513 ;
      RECT 1.197 0.378 1.235 0.396 ;
      RECT 1.197 0.297 1.256 0.315 ;
      RECT 1.12 0.225 1.179 0.243 ;
      RECT 1.161 0.027 1.179 0.243 ;
      RECT 1.141 0.144 1.179 0.162 ;
      RECT 1.12 0.027 1.179 0.045 ;
      RECT 1.12 0.495 1.179 0.513 ;
      RECT 1.161 0.297 1.179 0.513 ;
      RECT 1.141 0.378 1.179 0.396 ;
      RECT 1.12 0.297 1.179 0.315 ;
      RECT 0.99 0.225 1.04 0.243 ;
      RECT 0.99 0.027 1.008 0.243 ;
      RECT 0.99 0.027 1.04 0.045 ;
      RECT 0.99 0.495 1.04 0.513 ;
      RECT 0.99 0.297 1.008 0.513 ;
      RECT 0.99 0.297 1.04 0.315 ;
      RECT 0.855 0.126 0.873 0.203 ;
      RECT 0.821 0.126 0.873 0.144 ;
      RECT 0.821 0.396 0.873 0.414 ;
      RECT 0.855 0.337 0.873 0.414 ;
      RECT 0.72 0.225 0.824 0.243 ;
      RECT 0.72 0.027 0.738 0.243 ;
      RECT 0.612 0.122 0.738 0.14 ;
      RECT 0.72 0.027 0.77 0.045 ;
      RECT 0.72 0.495 0.77 0.513 ;
      RECT 0.72 0.297 0.738 0.513 ;
      RECT 0.612 0.4 0.738 0.418 ;
      RECT 0.72 0.297 0.824 0.315 ;
      RECT 0.558 0.225 0.612 0.243 ;
      RECT 0.558 0.081 0.576 0.243 ;
      RECT 0.558 0.081 0.692 0.099 ;
      RECT 0.585 0.045 0.603 0.099 ;
      RECT 0.585 0.441 0.603 0.495 ;
      RECT 0.558 0.441 0.692 0.459 ;
      RECT 0.558 0.297 0.576 0.459 ;
      RECT 0.558 0.297 0.612 0.315 ;
      RECT 0.45 0.224 0.5 0.242 ;
      RECT 0.45 0.027 0.468 0.242 ;
      RECT 0.288 0.153 0.468 0.171 ;
      RECT 0.342 0.117 0.36 0.171 ;
      RECT 0.288 0.117 0.306 0.171 ;
      RECT 0.45 0.027 0.554 0.045 ;
      RECT 0.45 0.495 0.554 0.513 ;
      RECT 0.45 0.298 0.468 0.513 ;
      RECT 0.342 0.369 0.36 0.423 ;
      RECT 0.288 0.369 0.306 0.423 ;
      RECT 0.288 0.369 0.468 0.387 ;
      RECT 0.45 0.298 0.5 0.316 ;
      RECT 0.234 0.225 0.338 0.243 ;
      RECT 0.234 0.027 0.252 0.243 ;
      RECT 0.396 0.027 0.414 0.119 ;
      RECT 0.234 0.027 0.414 0.045 ;
      RECT 0.234 0.495 0.414 0.513 ;
      RECT 0.396 0.421 0.414 0.513 ;
      RECT 0.234 0.297 0.252 0.513 ;
      RECT 0.234 0.297 0.338 0.315 ;
      RECT 2.178 0.122 2.196 0.167 ;
      RECT 2.178 0.373 2.196 0.418 ;
      RECT 1.854 0.101 1.872 0.167 ;
      RECT 1.854 0.373 1.872 0.439 ;
      RECT 1.692 0.165 1.71 0.203 ;
      RECT 1.692 0.337 1.71 0.375 ;
      RECT 1.584 0.106 1.602 0.167 ;
      RECT 1.584 0.373 1.602 0.434 ;
      RECT 1.33 0.106 1.348 0.167 ;
      RECT 1.33 0.373 1.348 0.434 ;
      RECT 1.028 0.106 1.046 0.167 ;
      RECT 1.028 0.373 1.046 0.434 ;
      RECT 0.774 0.106 0.792 0.167 ;
      RECT 0.774 0.373 0.792 0.434 ;
      RECT 0.666 0.165 0.684 0.203 ;
      RECT 0.666 0.337 0.684 0.375 ;
      RECT 0.504 0.101 0.522 0.167 ;
      RECT 0.504 0.373 0.522 0.439 ;
      RECT 0.18 0.122 0.198 0.167 ;
      RECT 0.18 0.373 0.198 0.418 ;
    LAYER M2 ;
      RECT 2.065 0.144 2.201 0.162 ;
      RECT 2.065 0.378 2.201 0.396 ;
      RECT 1.207 0.144 1.877 0.162 ;
      RECT 1.207 0.378 1.877 0.396 ;
      RECT 1.363 0.18 1.715 0.198 ;
      RECT 1.363 0.342 1.715 0.36 ;
      RECT 0.499 0.144 1.169 0.162 ;
      RECT 0.499 0.378 1.169 0.396 ;
      RECT 0.661 0.18 1.013 0.198 ;
      RECT 0.661 0.342 1.013 0.36 ;
      RECT 0.175 0.144 0.311 0.162 ;
      RECT 0.175 0.378 0.311 0.396 ;
    LAYER V1 ;
      RECT 2.178 0.144 2.196 0.162 ;
      RECT 2.178 0.378 2.196 0.396 ;
      RECT 2.07 0.144 2.088 0.162 ;
      RECT 2.07 0.378 2.088 0.396 ;
      RECT 1.854 0.144 1.872 0.162 ;
      RECT 1.854 0.378 1.872 0.396 ;
      RECT 1.692 0.18 1.71 0.198 ;
      RECT 1.692 0.342 1.71 0.36 ;
      RECT 1.584 0.144 1.602 0.162 ;
      RECT 1.584 0.378 1.602 0.396 ;
      RECT 1.503 0.18 1.521 0.198 ;
      RECT 1.503 0.342 1.521 0.36 ;
      RECT 1.368 0.18 1.386 0.198 ;
      RECT 1.368 0.342 1.386 0.36 ;
      RECT 1.33 0.144 1.348 0.162 ;
      RECT 1.33 0.378 1.348 0.396 ;
      RECT 1.212 0.144 1.23 0.162 ;
      RECT 1.212 0.378 1.23 0.396 ;
      RECT 1.146 0.144 1.164 0.162 ;
      RECT 1.146 0.378 1.164 0.396 ;
      RECT 1.028 0.144 1.046 0.162 ;
      RECT 1.028 0.378 1.046 0.396 ;
      RECT 0.99 0.18 1.008 0.198 ;
      RECT 0.99 0.342 1.008 0.36 ;
      RECT 0.855 0.18 0.873 0.198 ;
      RECT 0.855 0.342 0.873 0.36 ;
      RECT 0.774 0.144 0.792 0.162 ;
      RECT 0.774 0.378 0.792 0.396 ;
      RECT 0.666 0.18 0.684 0.198 ;
      RECT 0.666 0.342 0.684 0.36 ;
      RECT 0.504 0.144 0.522 0.162 ;
      RECT 0.504 0.378 0.522 0.396 ;
      RECT 0.288 0.144 0.306 0.162 ;
      RECT 0.288 0.378 0.306 0.396 ;
      RECT 0.18 0.144 0.198 0.162 ;
      RECT 0.18 0.378 0.198 0.396 ;
  END
END DFFHQNH2V2Xx3_ASAP7_75t_R

MACRO DFFHQNH2V2Xx3_ASAP7_75t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNH2V2Xx3_ASAP7_75t_SL 0 0 ;
  SIZE 2.376 BY 0.54 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t_pg ;
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.422 0.126 1.478 0.144 ;
        RECT 1.422 0.225 1.459 0.243 ;
        RECT 1.422 0.027 1.459 0.045 ;
        RECT 1.422 0.027 1.44 0.243 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.422 0.396 1.478 0.414 ;
        RECT 1.422 0.495 1.459 0.513 ;
        RECT 1.422 0.297 1.459 0.315 ;
        RECT 1.422 0.297 1.44 0.513 ;
    END
  END D1
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.917 0.225 0.954 0.243 ;
        RECT 0.936 0.027 0.954 0.243 ;
        RECT 0.898 0.126 0.954 0.144 ;
        RECT 0.917 0.027 0.954 0.045 ;
    END
  END D2
  PIN D3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.917 0.495 0.954 0.513 ;
        RECT 0.936 0.297 0.954 0.513 ;
        RECT 0.898 0.396 0.954 0.414 ;
        RECT 0.917 0.297 0.954 0.315 ;
    END
  END D3
  PIN QN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2 0.225 2.359 0.243 ;
        RECT 2.341 0.027 2.359 0.243 ;
        RECT 2.2 0.027 2.359 0.045 ;
    END
  END QN0
  PIN QN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2 0.495 2.359 0.513 ;
        RECT 2.341 0.297 2.359 0.513 ;
        RECT 2.2 0.297 2.359 0.315 ;
    END
  END QN1
  PIN QN2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.017 0.225 0.176 0.243 ;
        RECT 0.017 0.027 0.176 0.045 ;
        RECT 0.017 0.027 0.035 0.243 ;
    END
  END QN2
  PIN QN3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.017 0.495 0.176 0.513 ;
        RECT 0.017 0.297 0.176 0.315 ;
        RECT 0.017 0.297 0.035 0.513 ;
    END
  END QN3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 2.376 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 2.376 0.009 ;
        RECT 0 0.531 2.376 0.549 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 1.066 0.07 1.31 0.088 ;
        RECT 1.066 0.452 1.31 0.47 ;
      LAYER M3 ;
        RECT 1.125 0.05 1.143 0.492 ;
      LAYER M1 ;
        RECT 1.287 0.164 1.305 0.236 ;
        RECT 1.26 0.07 1.305 0.106 ;
        RECT 1.287 0.034 1.305 0.106 ;
        RECT 1.26 0.164 1.305 0.2 ;
        RECT 1.26 0.07 1.278 0.2 ;
        RECT 1.287 0.434 1.305 0.506 ;
        RECT 1.26 0.34 1.305 0.376 ;
        RECT 1.287 0.304 1.305 0.376 ;
        RECT 1.26 0.434 1.305 0.47 ;
        RECT 1.26 0.34 1.278 0.47 ;
        RECT 1.071 0.164 1.116 0.2 ;
        RECT 1.098 0.07 1.116 0.2 ;
        RECT 1.071 0.07 1.116 0.106 ;
        RECT 1.071 0.164 1.089 0.236 ;
        RECT 1.071 0.034 1.089 0.106 ;
        RECT 1.071 0.434 1.116 0.47 ;
        RECT 1.098 0.34 1.116 0.47 ;
        RECT 1.071 0.34 1.116 0.376 ;
        RECT 1.071 0.434 1.089 0.506 ;
        RECT 1.071 0.304 1.089 0.376 ;
      LAYER V2 ;
        RECT 1.125 0.452 1.143 0.47 ;
        RECT 1.125 0.07 1.143 0.088 ;
      LAYER V1 ;
        RECT 1.071 0.452 1.089 0.47 ;
        RECT 1.071 0.07 1.089 0.088 ;
        RECT 1.287 0.452 1.305 0.47 ;
        RECT 1.287 0.07 1.305 0.088 ;
    END
  END CLK
  OBS
    LAYER M1 ;
      RECT 2.038 0.225 2.142 0.243 ;
      RECT 2.124 0.027 2.142 0.243 ;
      RECT 1.962 0.027 1.98 0.119 ;
      RECT 1.962 0.027 2.142 0.045 ;
      RECT 1.962 0.495 2.142 0.513 ;
      RECT 2.124 0.297 2.142 0.513 ;
      RECT 1.962 0.421 1.98 0.513 ;
      RECT 2.038 0.297 2.142 0.315 ;
      RECT 1.876 0.224 1.926 0.242 ;
      RECT 1.908 0.027 1.926 0.242 ;
      RECT 1.908 0.153 2.088 0.171 ;
      RECT 2.07 0.117 2.088 0.171 ;
      RECT 2.016 0.117 2.034 0.171 ;
      RECT 1.822 0.027 1.926 0.045 ;
      RECT 1.822 0.495 1.926 0.513 ;
      RECT 1.908 0.298 1.926 0.513 ;
      RECT 2.07 0.369 2.088 0.423 ;
      RECT 2.016 0.369 2.034 0.423 ;
      RECT 1.908 0.369 2.088 0.387 ;
      RECT 1.876 0.298 1.926 0.316 ;
      RECT 1.764 0.225 1.818 0.243 ;
      RECT 1.8 0.081 1.818 0.243 ;
      RECT 1.684 0.081 1.818 0.099 ;
      RECT 1.773 0.045 1.791 0.099 ;
      RECT 1.773 0.441 1.791 0.495 ;
      RECT 1.684 0.441 1.818 0.459 ;
      RECT 1.8 0.297 1.818 0.459 ;
      RECT 1.764 0.297 1.818 0.315 ;
      RECT 1.552 0.225 1.656 0.243 ;
      RECT 1.638 0.027 1.656 0.243 ;
      RECT 1.638 0.122 1.764 0.14 ;
      RECT 1.606 0.027 1.656 0.045 ;
      RECT 1.606 0.495 1.656 0.513 ;
      RECT 1.638 0.297 1.656 0.513 ;
      RECT 1.638 0.4 1.764 0.418 ;
      RECT 1.552 0.297 1.656 0.315 ;
      RECT 1.503 0.126 1.521 0.203 ;
      RECT 1.503 0.126 1.555 0.144 ;
      RECT 1.503 0.396 1.555 0.414 ;
      RECT 1.503 0.337 1.521 0.414 ;
      RECT 1.336 0.225 1.386 0.243 ;
      RECT 1.368 0.027 1.386 0.243 ;
      RECT 1.336 0.027 1.386 0.045 ;
      RECT 1.336 0.495 1.386 0.513 ;
      RECT 1.368 0.297 1.386 0.513 ;
      RECT 1.336 0.297 1.386 0.315 ;
      RECT 1.197 0.225 1.256 0.243 ;
      RECT 1.197 0.027 1.215 0.243 ;
      RECT 1.197 0.144 1.235 0.162 ;
      RECT 1.197 0.027 1.256 0.045 ;
      RECT 1.197 0.495 1.256 0.513 ;
      RECT 1.197 0.297 1.215 0.513 ;
      RECT 1.197 0.378 1.235 0.396 ;
      RECT 1.197 0.297 1.256 0.315 ;
      RECT 1.12 0.225 1.179 0.243 ;
      RECT 1.161 0.027 1.179 0.243 ;
      RECT 1.141 0.144 1.179 0.162 ;
      RECT 1.12 0.027 1.179 0.045 ;
      RECT 1.12 0.495 1.179 0.513 ;
      RECT 1.161 0.297 1.179 0.513 ;
      RECT 1.141 0.378 1.179 0.396 ;
      RECT 1.12 0.297 1.179 0.315 ;
      RECT 0.99 0.225 1.04 0.243 ;
      RECT 0.99 0.027 1.008 0.243 ;
      RECT 0.99 0.027 1.04 0.045 ;
      RECT 0.99 0.495 1.04 0.513 ;
      RECT 0.99 0.297 1.008 0.513 ;
      RECT 0.99 0.297 1.04 0.315 ;
      RECT 0.855 0.126 0.873 0.203 ;
      RECT 0.821 0.126 0.873 0.144 ;
      RECT 0.821 0.396 0.873 0.414 ;
      RECT 0.855 0.337 0.873 0.414 ;
      RECT 0.72 0.225 0.824 0.243 ;
      RECT 0.72 0.027 0.738 0.243 ;
      RECT 0.612 0.122 0.738 0.14 ;
      RECT 0.72 0.027 0.77 0.045 ;
      RECT 0.72 0.495 0.77 0.513 ;
      RECT 0.72 0.297 0.738 0.513 ;
      RECT 0.612 0.4 0.738 0.418 ;
      RECT 0.72 0.297 0.824 0.315 ;
      RECT 0.558 0.225 0.612 0.243 ;
      RECT 0.558 0.081 0.576 0.243 ;
      RECT 0.558 0.081 0.692 0.099 ;
      RECT 0.585 0.045 0.603 0.099 ;
      RECT 0.585 0.441 0.603 0.495 ;
      RECT 0.558 0.441 0.692 0.459 ;
      RECT 0.558 0.297 0.576 0.459 ;
      RECT 0.558 0.297 0.612 0.315 ;
      RECT 0.45 0.224 0.5 0.242 ;
      RECT 0.45 0.027 0.468 0.242 ;
      RECT 0.288 0.153 0.468 0.171 ;
      RECT 0.342 0.117 0.36 0.171 ;
      RECT 0.288 0.117 0.306 0.171 ;
      RECT 0.45 0.027 0.554 0.045 ;
      RECT 0.45 0.495 0.554 0.513 ;
      RECT 0.45 0.298 0.468 0.513 ;
      RECT 0.342 0.369 0.36 0.423 ;
      RECT 0.288 0.369 0.306 0.423 ;
      RECT 0.288 0.369 0.468 0.387 ;
      RECT 0.45 0.298 0.5 0.316 ;
      RECT 0.234 0.225 0.338 0.243 ;
      RECT 0.234 0.027 0.252 0.243 ;
      RECT 0.396 0.027 0.414 0.119 ;
      RECT 0.234 0.027 0.414 0.045 ;
      RECT 0.234 0.495 0.414 0.513 ;
      RECT 0.396 0.421 0.414 0.513 ;
      RECT 0.234 0.297 0.252 0.513 ;
      RECT 0.234 0.297 0.338 0.315 ;
      RECT 2.178 0.122 2.196 0.167 ;
      RECT 2.178 0.373 2.196 0.418 ;
      RECT 1.854 0.101 1.872 0.167 ;
      RECT 1.854 0.373 1.872 0.439 ;
      RECT 1.692 0.165 1.71 0.203 ;
      RECT 1.692 0.337 1.71 0.375 ;
      RECT 1.584 0.106 1.602 0.167 ;
      RECT 1.584 0.373 1.602 0.434 ;
      RECT 1.33 0.106 1.348 0.167 ;
      RECT 1.33 0.373 1.348 0.434 ;
      RECT 1.028 0.106 1.046 0.167 ;
      RECT 1.028 0.373 1.046 0.434 ;
      RECT 0.774 0.106 0.792 0.167 ;
      RECT 0.774 0.373 0.792 0.434 ;
      RECT 0.666 0.165 0.684 0.203 ;
      RECT 0.666 0.337 0.684 0.375 ;
      RECT 0.504 0.101 0.522 0.167 ;
      RECT 0.504 0.373 0.522 0.439 ;
      RECT 0.18 0.122 0.198 0.167 ;
      RECT 0.18 0.373 0.198 0.418 ;
    LAYER M2 ;
      RECT 2.065 0.144 2.201 0.162 ;
      RECT 2.065 0.378 2.201 0.396 ;
      RECT 1.207 0.144 1.877 0.162 ;
      RECT 1.207 0.378 1.877 0.396 ;
      RECT 1.363 0.18 1.715 0.198 ;
      RECT 1.363 0.342 1.715 0.36 ;
      RECT 0.499 0.144 1.169 0.162 ;
      RECT 0.499 0.378 1.169 0.396 ;
      RECT 0.661 0.18 1.013 0.198 ;
      RECT 0.661 0.342 1.013 0.36 ;
      RECT 0.175 0.144 0.311 0.162 ;
      RECT 0.175 0.378 0.311 0.396 ;
    LAYER V1 ;
      RECT 2.178 0.144 2.196 0.162 ;
      RECT 2.178 0.378 2.196 0.396 ;
      RECT 2.07 0.144 2.088 0.162 ;
      RECT 2.07 0.378 2.088 0.396 ;
      RECT 1.854 0.144 1.872 0.162 ;
      RECT 1.854 0.378 1.872 0.396 ;
      RECT 1.692 0.18 1.71 0.198 ;
      RECT 1.692 0.342 1.71 0.36 ;
      RECT 1.584 0.144 1.602 0.162 ;
      RECT 1.584 0.378 1.602 0.396 ;
      RECT 1.503 0.18 1.521 0.198 ;
      RECT 1.503 0.342 1.521 0.36 ;
      RECT 1.368 0.18 1.386 0.198 ;
      RECT 1.368 0.342 1.386 0.36 ;
      RECT 1.33 0.144 1.348 0.162 ;
      RECT 1.33 0.378 1.348 0.396 ;
      RECT 1.212 0.144 1.23 0.162 ;
      RECT 1.212 0.378 1.23 0.396 ;
      RECT 1.146 0.144 1.164 0.162 ;
      RECT 1.146 0.378 1.164 0.396 ;
      RECT 1.028 0.144 1.046 0.162 ;
      RECT 1.028 0.378 1.046 0.396 ;
      RECT 0.99 0.18 1.008 0.198 ;
      RECT 0.99 0.342 1.008 0.36 ;
      RECT 0.855 0.18 0.873 0.198 ;
      RECT 0.855 0.342 0.873 0.36 ;
      RECT 0.774 0.144 0.792 0.162 ;
      RECT 0.774 0.378 0.792 0.396 ;
      RECT 0.666 0.18 0.684 0.198 ;
      RECT 0.666 0.342 0.684 0.36 ;
      RECT 0.504 0.144 0.522 0.162 ;
      RECT 0.504 0.378 0.522 0.396 ;
      RECT 0.288 0.144 0.306 0.162 ;
      RECT 0.288 0.378 0.306 0.396 ;
      RECT 0.18 0.144 0.198 0.162 ;
      RECT 0.18 0.378 0.198 0.396 ;
  END
END DFFHQNH2V2Xx3_ASAP7_75t_SL

END LIBRARY
