../../../../test/Nangate45/Nangate45_stdcell.lef