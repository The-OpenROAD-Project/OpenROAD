VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO DFF
  ORIGIN 0 0 ;
  SIZE 1.0 BY 0.1 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
  END VSS
  PIN CP
    DIRECTION INPUT ;
    USE SIGNAL ;
  END CP
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
  END SI
  PIN VBB
    DIRECTION INOUT ;
    USE GROUND ;
  END VBB
  PIN VPP
    DIRECTION INOUT ;
    USE POWER ;
  END VPP
END DFF

MACRO MBFF2
  ORIGIN 0 0 ;
  SIZE 1.0 BY 0.1 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
  END VSS
  PIN CP
    DIRECTION INPUT ;
    USE SIGNAL ;
  END CP
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
  END D1
  PIN Q0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END Q0
  PIN Q1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END Q1
  PIN VBB
    DIRECTION INOUT ;
    USE GROUND ;
  END VBB
  PIN VPP
    DIRECTION INOUT ;
    USE POWER ;
  END VPP
END MBFF2

MACRO MBFF2CLPS
  ORIGIN 0 0 ;
  SIZE 1.0 BY 0.1 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
  END VSS
  PIN CP
    DIRECTION INPUT ;
    USE SIGNAL ;
  END CP
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
  END D1
  PIN Q0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END Q0
  PIN Q1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END Q1
  PIN CLEAR
    DIRECTION INPUT ;
    USE SIGNAL ;
  END CLEAR
  PIN PRESET
    DIRECTION INPUT ;
    USE SIGNAL ;
  END PRESET
  PIN VBB
    DIRECTION INOUT ;
    USE GROUND ;
  END VBB
  PIN VPP
    DIRECTION INOUT ;
    USE POWER ;
  END VPP
END MBFF2CLPS

MACRO MBFF2SE
  ORIGIN 0 0 ;
  SIZE 1.0 BY 0.1 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
  END VSS
  PIN CP
    DIRECTION INPUT ;
    USE SIGNAL ;
  END CP
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
  END D1
  PIN Q0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END Q0
  PIN Q1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END Q1
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
  END SI
  PIN VBB
    DIRECTION INOUT ;
    USE GROUND ;
  END VBB
  PIN VPP
    DIRECTION INOUT ;
    USE POWER ;
  END VPP
END MBFF2SE

MACRO MBFF2SECLPS
  ORIGIN 0 0 ;
  SIZE 1.0 BY 0.1 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
  END VSS
  PIN CP
    DIRECTION INPUT ;
    USE SIGNAL ;
  END CP
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
  END D1
  PIN Q0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END Q0
  PIN Q1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END Q1
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
  END SI
  PIN CLEAR
    DIRECTION INPUT ;
    USE SIGNAL ;
  END CLEAR
  PIN PRESET
    DIRECTION INPUT ;
    USE SIGNAL ;
  END PRESET
  PIN VBB
    DIRECTION INOUT ;
    USE GROUND ;
  END VBB
  PIN VPP
    DIRECTION INOUT ;
    USE POWER ;
  END VPP
END MBFF2SECLPS

MACRO INV
  ORIGIN 0 0 ;
  SIZE 0.1 BY 0.1 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
  END A
  PIN Z
    DIRECTION INPUT ;
    USE SIGNAL ;
  END Z
  PIN VBB
    DIRECTION INOUT ;
    USE GROUND ;
  END VBB
  PIN VPP
    DIRECTION INOUT ;
    USE POWER ;
  END VPP
END INV

END LIBRARY
