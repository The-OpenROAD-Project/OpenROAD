module MockArray (clock,
    io_lsbs_0,
    io_lsbs_1,
    io_lsbs_10,
    io_lsbs_11,
    io_lsbs_12,
    io_lsbs_13,
    io_lsbs_14,
    io_lsbs_15,
    io_lsbs_2,
    io_lsbs_3,
    io_lsbs_4,
    io_lsbs_5,
    io_lsbs_6,
    io_lsbs_7,
    io_lsbs_8,
    io_lsbs_9,
    reset,
    io_ins_down_0,
    io_ins_down_1,
    io_ins_down_2,
    io_ins_down_3,
    io_ins_left_0,
    io_ins_left_1,
    io_ins_left_2,
    io_ins_left_3,
    io_ins_right_0,
    io_ins_right_1,
    io_ins_right_2,
    io_ins_right_3,
    io_ins_up_0,
    io_ins_up_1,
    io_ins_up_2,
    io_ins_up_3,
    io_outs_down_0,
    io_outs_down_1,
    io_outs_down_2,
    io_outs_down_3,
    io_outs_left_0,
    io_outs_left_1,
    io_outs_left_2,
    io_outs_left_3,
    io_outs_right_0,
    io_outs_right_1,
    io_outs_right_2,
    io_outs_right_3,
    io_outs_up_0,
    io_outs_up_1,
    io_outs_up_2,
    io_outs_up_3);
 input clock;
 output io_lsbs_0;
 output io_lsbs_1;
 output io_lsbs_10;
 output io_lsbs_11;
 output io_lsbs_12;
 output io_lsbs_13;
 output io_lsbs_14;
 output io_lsbs_15;
 output io_lsbs_2;
 output io_lsbs_3;
 output io_lsbs_4;
 output io_lsbs_5;
 output io_lsbs_6;
 output io_lsbs_7;
 output io_lsbs_8;
 output io_lsbs_9;
 input reset;
 input [63:0] io_ins_down_0;
 input [63:0] io_ins_down_1;
 input [63:0] io_ins_down_2;
 input [63:0] io_ins_down_3;
 input [63:0] io_ins_left_0;
 input [63:0] io_ins_left_1;
 input [63:0] io_ins_left_2;
 input [63:0] io_ins_left_3;
 input [63:0] io_ins_right_0;
 input [63:0] io_ins_right_1;
 input [63:0] io_ins_right_2;
 input [63:0] io_ins_right_3;
 input [63:0] io_ins_up_0;
 input [63:0] io_ins_up_1;
 input [63:0] io_ins_up_2;
 input [63:0] io_ins_up_3;
 output [63:0] io_outs_down_0;
 output [63:0] io_outs_down_1;
 output [63:0] io_outs_down_2;
 output [63:0] io_outs_down_3;
 output [63:0] io_outs_left_0;
 output [63:0] io_outs_left_1;
 output [63:0] io_outs_left_2;
 output [63:0] io_outs_left_3;
 output [63:0] io_outs_right_0;
 output [63:0] io_outs_right_1;
 output [63:0] io_outs_right_2;
 output [63:0] io_outs_right_3;
 output [63:0] io_outs_up_0;
 output [63:0] io_outs_up_1;
 output [63:0] io_outs_up_2;
 output [63:0] io_outs_up_3;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _ces_0_0_io_lsbOuts_1;
 wire _ces_0_0_io_lsbOuts_2;
 wire _ces_0_0_io_lsbOuts_3;
 wire \_ces_0_0_io_outs_right[0] ;
 wire \_ces_0_0_io_outs_right[10] ;
 wire \_ces_0_0_io_outs_right[11] ;
 wire \_ces_0_0_io_outs_right[12] ;
 wire \_ces_0_0_io_outs_right[13] ;
 wire \_ces_0_0_io_outs_right[14] ;
 wire \_ces_0_0_io_outs_right[15] ;
 wire \_ces_0_0_io_outs_right[16] ;
 wire \_ces_0_0_io_outs_right[17] ;
 wire \_ces_0_0_io_outs_right[18] ;
 wire \_ces_0_0_io_outs_right[19] ;
 wire \_ces_0_0_io_outs_right[1] ;
 wire \_ces_0_0_io_outs_right[20] ;
 wire \_ces_0_0_io_outs_right[21] ;
 wire \_ces_0_0_io_outs_right[22] ;
 wire \_ces_0_0_io_outs_right[23] ;
 wire \_ces_0_0_io_outs_right[24] ;
 wire \_ces_0_0_io_outs_right[25] ;
 wire \_ces_0_0_io_outs_right[26] ;
 wire \_ces_0_0_io_outs_right[27] ;
 wire \_ces_0_0_io_outs_right[28] ;
 wire \_ces_0_0_io_outs_right[29] ;
 wire \_ces_0_0_io_outs_right[2] ;
 wire \_ces_0_0_io_outs_right[30] ;
 wire \_ces_0_0_io_outs_right[31] ;
 wire \_ces_0_0_io_outs_right[32] ;
 wire \_ces_0_0_io_outs_right[33] ;
 wire \_ces_0_0_io_outs_right[34] ;
 wire \_ces_0_0_io_outs_right[35] ;
 wire \_ces_0_0_io_outs_right[36] ;
 wire \_ces_0_0_io_outs_right[37] ;
 wire \_ces_0_0_io_outs_right[38] ;
 wire \_ces_0_0_io_outs_right[39] ;
 wire \_ces_0_0_io_outs_right[3] ;
 wire \_ces_0_0_io_outs_right[40] ;
 wire \_ces_0_0_io_outs_right[41] ;
 wire \_ces_0_0_io_outs_right[42] ;
 wire \_ces_0_0_io_outs_right[43] ;
 wire \_ces_0_0_io_outs_right[44] ;
 wire \_ces_0_0_io_outs_right[45] ;
 wire \_ces_0_0_io_outs_right[46] ;
 wire \_ces_0_0_io_outs_right[47] ;
 wire \_ces_0_0_io_outs_right[48] ;
 wire \_ces_0_0_io_outs_right[49] ;
 wire \_ces_0_0_io_outs_right[4] ;
 wire \_ces_0_0_io_outs_right[50] ;
 wire \_ces_0_0_io_outs_right[51] ;
 wire \_ces_0_0_io_outs_right[52] ;
 wire \_ces_0_0_io_outs_right[53] ;
 wire \_ces_0_0_io_outs_right[54] ;
 wire \_ces_0_0_io_outs_right[55] ;
 wire \_ces_0_0_io_outs_right[56] ;
 wire \_ces_0_0_io_outs_right[57] ;
 wire \_ces_0_0_io_outs_right[58] ;
 wire \_ces_0_0_io_outs_right[59] ;
 wire \_ces_0_0_io_outs_right[5] ;
 wire \_ces_0_0_io_outs_right[60] ;
 wire \_ces_0_0_io_outs_right[61] ;
 wire \_ces_0_0_io_outs_right[62] ;
 wire \_ces_0_0_io_outs_right[63] ;
 wire \_ces_0_0_io_outs_right[6] ;
 wire \_ces_0_0_io_outs_right[7] ;
 wire \_ces_0_0_io_outs_right[8] ;
 wire \_ces_0_0_io_outs_right[9] ;
 wire \_ces_0_0_io_outs_up[0] ;
 wire \_ces_0_0_io_outs_up[10] ;
 wire \_ces_0_0_io_outs_up[11] ;
 wire \_ces_0_0_io_outs_up[12] ;
 wire \_ces_0_0_io_outs_up[13] ;
 wire \_ces_0_0_io_outs_up[14] ;
 wire \_ces_0_0_io_outs_up[15] ;
 wire \_ces_0_0_io_outs_up[16] ;
 wire \_ces_0_0_io_outs_up[17] ;
 wire \_ces_0_0_io_outs_up[18] ;
 wire \_ces_0_0_io_outs_up[19] ;
 wire \_ces_0_0_io_outs_up[1] ;
 wire \_ces_0_0_io_outs_up[20] ;
 wire \_ces_0_0_io_outs_up[21] ;
 wire \_ces_0_0_io_outs_up[22] ;
 wire \_ces_0_0_io_outs_up[23] ;
 wire \_ces_0_0_io_outs_up[24] ;
 wire \_ces_0_0_io_outs_up[25] ;
 wire \_ces_0_0_io_outs_up[26] ;
 wire \_ces_0_0_io_outs_up[27] ;
 wire \_ces_0_0_io_outs_up[28] ;
 wire \_ces_0_0_io_outs_up[29] ;
 wire \_ces_0_0_io_outs_up[2] ;
 wire \_ces_0_0_io_outs_up[30] ;
 wire \_ces_0_0_io_outs_up[31] ;
 wire \_ces_0_0_io_outs_up[32] ;
 wire \_ces_0_0_io_outs_up[33] ;
 wire \_ces_0_0_io_outs_up[34] ;
 wire \_ces_0_0_io_outs_up[35] ;
 wire \_ces_0_0_io_outs_up[36] ;
 wire \_ces_0_0_io_outs_up[37] ;
 wire \_ces_0_0_io_outs_up[38] ;
 wire \_ces_0_0_io_outs_up[39] ;
 wire \_ces_0_0_io_outs_up[3] ;
 wire \_ces_0_0_io_outs_up[40] ;
 wire \_ces_0_0_io_outs_up[41] ;
 wire \_ces_0_0_io_outs_up[42] ;
 wire \_ces_0_0_io_outs_up[43] ;
 wire \_ces_0_0_io_outs_up[44] ;
 wire \_ces_0_0_io_outs_up[45] ;
 wire \_ces_0_0_io_outs_up[46] ;
 wire \_ces_0_0_io_outs_up[47] ;
 wire \_ces_0_0_io_outs_up[48] ;
 wire \_ces_0_0_io_outs_up[49] ;
 wire \_ces_0_0_io_outs_up[4] ;
 wire \_ces_0_0_io_outs_up[50] ;
 wire \_ces_0_0_io_outs_up[51] ;
 wire \_ces_0_0_io_outs_up[52] ;
 wire \_ces_0_0_io_outs_up[53] ;
 wire \_ces_0_0_io_outs_up[54] ;
 wire \_ces_0_0_io_outs_up[55] ;
 wire \_ces_0_0_io_outs_up[56] ;
 wire \_ces_0_0_io_outs_up[57] ;
 wire \_ces_0_0_io_outs_up[58] ;
 wire \_ces_0_0_io_outs_up[59] ;
 wire \_ces_0_0_io_outs_up[5] ;
 wire \_ces_0_0_io_outs_up[60] ;
 wire \_ces_0_0_io_outs_up[61] ;
 wire \_ces_0_0_io_outs_up[62] ;
 wire \_ces_0_0_io_outs_up[63] ;
 wire \_ces_0_0_io_outs_up[6] ;
 wire \_ces_0_0_io_outs_up[7] ;
 wire \_ces_0_0_io_outs_up[8] ;
 wire \_ces_0_0_io_outs_up[9] ;
 wire _ces_0_1_io_lsbOuts_1;
 wire _ces_0_1_io_lsbOuts_2;
 wire _ces_0_1_io_lsbOuts_3;
 wire \_ces_0_1_io_outs_left[0] ;
 wire \_ces_0_1_io_outs_left[10] ;
 wire \_ces_0_1_io_outs_left[11] ;
 wire \_ces_0_1_io_outs_left[12] ;
 wire \_ces_0_1_io_outs_left[13] ;
 wire \_ces_0_1_io_outs_left[14] ;
 wire \_ces_0_1_io_outs_left[15] ;
 wire \_ces_0_1_io_outs_left[16] ;
 wire \_ces_0_1_io_outs_left[17] ;
 wire \_ces_0_1_io_outs_left[18] ;
 wire \_ces_0_1_io_outs_left[19] ;
 wire \_ces_0_1_io_outs_left[1] ;
 wire \_ces_0_1_io_outs_left[20] ;
 wire \_ces_0_1_io_outs_left[21] ;
 wire \_ces_0_1_io_outs_left[22] ;
 wire \_ces_0_1_io_outs_left[23] ;
 wire \_ces_0_1_io_outs_left[24] ;
 wire \_ces_0_1_io_outs_left[25] ;
 wire \_ces_0_1_io_outs_left[26] ;
 wire \_ces_0_1_io_outs_left[27] ;
 wire \_ces_0_1_io_outs_left[28] ;
 wire \_ces_0_1_io_outs_left[29] ;
 wire \_ces_0_1_io_outs_left[2] ;
 wire \_ces_0_1_io_outs_left[30] ;
 wire \_ces_0_1_io_outs_left[31] ;
 wire \_ces_0_1_io_outs_left[32] ;
 wire \_ces_0_1_io_outs_left[33] ;
 wire \_ces_0_1_io_outs_left[34] ;
 wire \_ces_0_1_io_outs_left[35] ;
 wire \_ces_0_1_io_outs_left[36] ;
 wire \_ces_0_1_io_outs_left[37] ;
 wire \_ces_0_1_io_outs_left[38] ;
 wire \_ces_0_1_io_outs_left[39] ;
 wire \_ces_0_1_io_outs_left[3] ;
 wire \_ces_0_1_io_outs_left[40] ;
 wire \_ces_0_1_io_outs_left[41] ;
 wire \_ces_0_1_io_outs_left[42] ;
 wire \_ces_0_1_io_outs_left[43] ;
 wire \_ces_0_1_io_outs_left[44] ;
 wire \_ces_0_1_io_outs_left[45] ;
 wire \_ces_0_1_io_outs_left[46] ;
 wire \_ces_0_1_io_outs_left[47] ;
 wire \_ces_0_1_io_outs_left[48] ;
 wire \_ces_0_1_io_outs_left[49] ;
 wire \_ces_0_1_io_outs_left[4] ;
 wire \_ces_0_1_io_outs_left[50] ;
 wire \_ces_0_1_io_outs_left[51] ;
 wire \_ces_0_1_io_outs_left[52] ;
 wire \_ces_0_1_io_outs_left[53] ;
 wire \_ces_0_1_io_outs_left[54] ;
 wire \_ces_0_1_io_outs_left[55] ;
 wire \_ces_0_1_io_outs_left[56] ;
 wire \_ces_0_1_io_outs_left[57] ;
 wire \_ces_0_1_io_outs_left[58] ;
 wire \_ces_0_1_io_outs_left[59] ;
 wire \_ces_0_1_io_outs_left[5] ;
 wire \_ces_0_1_io_outs_left[60] ;
 wire \_ces_0_1_io_outs_left[61] ;
 wire \_ces_0_1_io_outs_left[62] ;
 wire \_ces_0_1_io_outs_left[63] ;
 wire \_ces_0_1_io_outs_left[6] ;
 wire \_ces_0_1_io_outs_left[7] ;
 wire \_ces_0_1_io_outs_left[8] ;
 wire \_ces_0_1_io_outs_left[9] ;
 wire \_ces_0_1_io_outs_right[0] ;
 wire \_ces_0_1_io_outs_right[10] ;
 wire \_ces_0_1_io_outs_right[11] ;
 wire \_ces_0_1_io_outs_right[12] ;
 wire \_ces_0_1_io_outs_right[13] ;
 wire \_ces_0_1_io_outs_right[14] ;
 wire \_ces_0_1_io_outs_right[15] ;
 wire \_ces_0_1_io_outs_right[16] ;
 wire \_ces_0_1_io_outs_right[17] ;
 wire \_ces_0_1_io_outs_right[18] ;
 wire \_ces_0_1_io_outs_right[19] ;
 wire \_ces_0_1_io_outs_right[1] ;
 wire \_ces_0_1_io_outs_right[20] ;
 wire \_ces_0_1_io_outs_right[21] ;
 wire \_ces_0_1_io_outs_right[22] ;
 wire \_ces_0_1_io_outs_right[23] ;
 wire \_ces_0_1_io_outs_right[24] ;
 wire \_ces_0_1_io_outs_right[25] ;
 wire \_ces_0_1_io_outs_right[26] ;
 wire \_ces_0_1_io_outs_right[27] ;
 wire \_ces_0_1_io_outs_right[28] ;
 wire \_ces_0_1_io_outs_right[29] ;
 wire \_ces_0_1_io_outs_right[2] ;
 wire \_ces_0_1_io_outs_right[30] ;
 wire \_ces_0_1_io_outs_right[31] ;
 wire \_ces_0_1_io_outs_right[32] ;
 wire \_ces_0_1_io_outs_right[33] ;
 wire \_ces_0_1_io_outs_right[34] ;
 wire \_ces_0_1_io_outs_right[35] ;
 wire \_ces_0_1_io_outs_right[36] ;
 wire \_ces_0_1_io_outs_right[37] ;
 wire \_ces_0_1_io_outs_right[38] ;
 wire \_ces_0_1_io_outs_right[39] ;
 wire \_ces_0_1_io_outs_right[3] ;
 wire \_ces_0_1_io_outs_right[40] ;
 wire \_ces_0_1_io_outs_right[41] ;
 wire \_ces_0_1_io_outs_right[42] ;
 wire \_ces_0_1_io_outs_right[43] ;
 wire \_ces_0_1_io_outs_right[44] ;
 wire \_ces_0_1_io_outs_right[45] ;
 wire \_ces_0_1_io_outs_right[46] ;
 wire \_ces_0_1_io_outs_right[47] ;
 wire \_ces_0_1_io_outs_right[48] ;
 wire \_ces_0_1_io_outs_right[49] ;
 wire \_ces_0_1_io_outs_right[4] ;
 wire \_ces_0_1_io_outs_right[50] ;
 wire \_ces_0_1_io_outs_right[51] ;
 wire \_ces_0_1_io_outs_right[52] ;
 wire \_ces_0_1_io_outs_right[53] ;
 wire \_ces_0_1_io_outs_right[54] ;
 wire \_ces_0_1_io_outs_right[55] ;
 wire \_ces_0_1_io_outs_right[56] ;
 wire \_ces_0_1_io_outs_right[57] ;
 wire \_ces_0_1_io_outs_right[58] ;
 wire \_ces_0_1_io_outs_right[59] ;
 wire \_ces_0_1_io_outs_right[5] ;
 wire \_ces_0_1_io_outs_right[60] ;
 wire \_ces_0_1_io_outs_right[61] ;
 wire \_ces_0_1_io_outs_right[62] ;
 wire \_ces_0_1_io_outs_right[63] ;
 wire \_ces_0_1_io_outs_right[6] ;
 wire \_ces_0_1_io_outs_right[7] ;
 wire \_ces_0_1_io_outs_right[8] ;
 wire \_ces_0_1_io_outs_right[9] ;
 wire \_ces_0_1_io_outs_up[0] ;
 wire \_ces_0_1_io_outs_up[10] ;
 wire \_ces_0_1_io_outs_up[11] ;
 wire \_ces_0_1_io_outs_up[12] ;
 wire \_ces_0_1_io_outs_up[13] ;
 wire \_ces_0_1_io_outs_up[14] ;
 wire \_ces_0_1_io_outs_up[15] ;
 wire \_ces_0_1_io_outs_up[16] ;
 wire \_ces_0_1_io_outs_up[17] ;
 wire \_ces_0_1_io_outs_up[18] ;
 wire \_ces_0_1_io_outs_up[19] ;
 wire \_ces_0_1_io_outs_up[1] ;
 wire \_ces_0_1_io_outs_up[20] ;
 wire \_ces_0_1_io_outs_up[21] ;
 wire \_ces_0_1_io_outs_up[22] ;
 wire \_ces_0_1_io_outs_up[23] ;
 wire \_ces_0_1_io_outs_up[24] ;
 wire \_ces_0_1_io_outs_up[25] ;
 wire \_ces_0_1_io_outs_up[26] ;
 wire \_ces_0_1_io_outs_up[27] ;
 wire \_ces_0_1_io_outs_up[28] ;
 wire \_ces_0_1_io_outs_up[29] ;
 wire \_ces_0_1_io_outs_up[2] ;
 wire \_ces_0_1_io_outs_up[30] ;
 wire \_ces_0_1_io_outs_up[31] ;
 wire \_ces_0_1_io_outs_up[32] ;
 wire \_ces_0_1_io_outs_up[33] ;
 wire \_ces_0_1_io_outs_up[34] ;
 wire \_ces_0_1_io_outs_up[35] ;
 wire \_ces_0_1_io_outs_up[36] ;
 wire \_ces_0_1_io_outs_up[37] ;
 wire \_ces_0_1_io_outs_up[38] ;
 wire \_ces_0_1_io_outs_up[39] ;
 wire \_ces_0_1_io_outs_up[3] ;
 wire \_ces_0_1_io_outs_up[40] ;
 wire \_ces_0_1_io_outs_up[41] ;
 wire \_ces_0_1_io_outs_up[42] ;
 wire \_ces_0_1_io_outs_up[43] ;
 wire \_ces_0_1_io_outs_up[44] ;
 wire \_ces_0_1_io_outs_up[45] ;
 wire \_ces_0_1_io_outs_up[46] ;
 wire \_ces_0_1_io_outs_up[47] ;
 wire \_ces_0_1_io_outs_up[48] ;
 wire \_ces_0_1_io_outs_up[49] ;
 wire \_ces_0_1_io_outs_up[4] ;
 wire \_ces_0_1_io_outs_up[50] ;
 wire \_ces_0_1_io_outs_up[51] ;
 wire \_ces_0_1_io_outs_up[52] ;
 wire \_ces_0_1_io_outs_up[53] ;
 wire \_ces_0_1_io_outs_up[54] ;
 wire \_ces_0_1_io_outs_up[55] ;
 wire \_ces_0_1_io_outs_up[56] ;
 wire \_ces_0_1_io_outs_up[57] ;
 wire \_ces_0_1_io_outs_up[58] ;
 wire \_ces_0_1_io_outs_up[59] ;
 wire \_ces_0_1_io_outs_up[5] ;
 wire \_ces_0_1_io_outs_up[60] ;
 wire \_ces_0_1_io_outs_up[61] ;
 wire \_ces_0_1_io_outs_up[62] ;
 wire \_ces_0_1_io_outs_up[63] ;
 wire \_ces_0_1_io_outs_up[6] ;
 wire \_ces_0_1_io_outs_up[7] ;
 wire \_ces_0_1_io_outs_up[8] ;
 wire \_ces_0_1_io_outs_up[9] ;
 wire _ces_0_2_io_lsbOuts_1;
 wire _ces_0_2_io_lsbOuts_2;
 wire _ces_0_2_io_lsbOuts_3;
 wire \_ces_0_2_io_outs_left[0] ;
 wire \_ces_0_2_io_outs_left[10] ;
 wire \_ces_0_2_io_outs_left[11] ;
 wire \_ces_0_2_io_outs_left[12] ;
 wire \_ces_0_2_io_outs_left[13] ;
 wire \_ces_0_2_io_outs_left[14] ;
 wire \_ces_0_2_io_outs_left[15] ;
 wire \_ces_0_2_io_outs_left[16] ;
 wire \_ces_0_2_io_outs_left[17] ;
 wire \_ces_0_2_io_outs_left[18] ;
 wire \_ces_0_2_io_outs_left[19] ;
 wire \_ces_0_2_io_outs_left[1] ;
 wire \_ces_0_2_io_outs_left[20] ;
 wire \_ces_0_2_io_outs_left[21] ;
 wire \_ces_0_2_io_outs_left[22] ;
 wire \_ces_0_2_io_outs_left[23] ;
 wire \_ces_0_2_io_outs_left[24] ;
 wire \_ces_0_2_io_outs_left[25] ;
 wire \_ces_0_2_io_outs_left[26] ;
 wire \_ces_0_2_io_outs_left[27] ;
 wire \_ces_0_2_io_outs_left[28] ;
 wire \_ces_0_2_io_outs_left[29] ;
 wire \_ces_0_2_io_outs_left[2] ;
 wire \_ces_0_2_io_outs_left[30] ;
 wire \_ces_0_2_io_outs_left[31] ;
 wire \_ces_0_2_io_outs_left[32] ;
 wire \_ces_0_2_io_outs_left[33] ;
 wire \_ces_0_2_io_outs_left[34] ;
 wire \_ces_0_2_io_outs_left[35] ;
 wire \_ces_0_2_io_outs_left[36] ;
 wire \_ces_0_2_io_outs_left[37] ;
 wire \_ces_0_2_io_outs_left[38] ;
 wire \_ces_0_2_io_outs_left[39] ;
 wire \_ces_0_2_io_outs_left[3] ;
 wire \_ces_0_2_io_outs_left[40] ;
 wire \_ces_0_2_io_outs_left[41] ;
 wire \_ces_0_2_io_outs_left[42] ;
 wire \_ces_0_2_io_outs_left[43] ;
 wire \_ces_0_2_io_outs_left[44] ;
 wire \_ces_0_2_io_outs_left[45] ;
 wire \_ces_0_2_io_outs_left[46] ;
 wire \_ces_0_2_io_outs_left[47] ;
 wire \_ces_0_2_io_outs_left[48] ;
 wire \_ces_0_2_io_outs_left[49] ;
 wire \_ces_0_2_io_outs_left[4] ;
 wire \_ces_0_2_io_outs_left[50] ;
 wire \_ces_0_2_io_outs_left[51] ;
 wire \_ces_0_2_io_outs_left[52] ;
 wire \_ces_0_2_io_outs_left[53] ;
 wire \_ces_0_2_io_outs_left[54] ;
 wire \_ces_0_2_io_outs_left[55] ;
 wire \_ces_0_2_io_outs_left[56] ;
 wire \_ces_0_2_io_outs_left[57] ;
 wire \_ces_0_2_io_outs_left[58] ;
 wire \_ces_0_2_io_outs_left[59] ;
 wire \_ces_0_2_io_outs_left[5] ;
 wire \_ces_0_2_io_outs_left[60] ;
 wire \_ces_0_2_io_outs_left[61] ;
 wire \_ces_0_2_io_outs_left[62] ;
 wire \_ces_0_2_io_outs_left[63] ;
 wire \_ces_0_2_io_outs_left[6] ;
 wire \_ces_0_2_io_outs_left[7] ;
 wire \_ces_0_2_io_outs_left[8] ;
 wire \_ces_0_2_io_outs_left[9] ;
 wire \_ces_0_2_io_outs_right[0] ;
 wire \_ces_0_2_io_outs_right[10] ;
 wire \_ces_0_2_io_outs_right[11] ;
 wire \_ces_0_2_io_outs_right[12] ;
 wire \_ces_0_2_io_outs_right[13] ;
 wire \_ces_0_2_io_outs_right[14] ;
 wire \_ces_0_2_io_outs_right[15] ;
 wire \_ces_0_2_io_outs_right[16] ;
 wire \_ces_0_2_io_outs_right[17] ;
 wire \_ces_0_2_io_outs_right[18] ;
 wire \_ces_0_2_io_outs_right[19] ;
 wire \_ces_0_2_io_outs_right[1] ;
 wire \_ces_0_2_io_outs_right[20] ;
 wire \_ces_0_2_io_outs_right[21] ;
 wire \_ces_0_2_io_outs_right[22] ;
 wire \_ces_0_2_io_outs_right[23] ;
 wire \_ces_0_2_io_outs_right[24] ;
 wire \_ces_0_2_io_outs_right[25] ;
 wire \_ces_0_2_io_outs_right[26] ;
 wire \_ces_0_2_io_outs_right[27] ;
 wire \_ces_0_2_io_outs_right[28] ;
 wire \_ces_0_2_io_outs_right[29] ;
 wire \_ces_0_2_io_outs_right[2] ;
 wire \_ces_0_2_io_outs_right[30] ;
 wire \_ces_0_2_io_outs_right[31] ;
 wire \_ces_0_2_io_outs_right[32] ;
 wire \_ces_0_2_io_outs_right[33] ;
 wire \_ces_0_2_io_outs_right[34] ;
 wire \_ces_0_2_io_outs_right[35] ;
 wire \_ces_0_2_io_outs_right[36] ;
 wire \_ces_0_2_io_outs_right[37] ;
 wire \_ces_0_2_io_outs_right[38] ;
 wire \_ces_0_2_io_outs_right[39] ;
 wire \_ces_0_2_io_outs_right[3] ;
 wire \_ces_0_2_io_outs_right[40] ;
 wire \_ces_0_2_io_outs_right[41] ;
 wire \_ces_0_2_io_outs_right[42] ;
 wire \_ces_0_2_io_outs_right[43] ;
 wire \_ces_0_2_io_outs_right[44] ;
 wire \_ces_0_2_io_outs_right[45] ;
 wire \_ces_0_2_io_outs_right[46] ;
 wire \_ces_0_2_io_outs_right[47] ;
 wire \_ces_0_2_io_outs_right[48] ;
 wire \_ces_0_2_io_outs_right[49] ;
 wire \_ces_0_2_io_outs_right[4] ;
 wire \_ces_0_2_io_outs_right[50] ;
 wire \_ces_0_2_io_outs_right[51] ;
 wire \_ces_0_2_io_outs_right[52] ;
 wire \_ces_0_2_io_outs_right[53] ;
 wire \_ces_0_2_io_outs_right[54] ;
 wire \_ces_0_2_io_outs_right[55] ;
 wire \_ces_0_2_io_outs_right[56] ;
 wire \_ces_0_2_io_outs_right[57] ;
 wire \_ces_0_2_io_outs_right[58] ;
 wire \_ces_0_2_io_outs_right[59] ;
 wire \_ces_0_2_io_outs_right[5] ;
 wire \_ces_0_2_io_outs_right[60] ;
 wire \_ces_0_2_io_outs_right[61] ;
 wire \_ces_0_2_io_outs_right[62] ;
 wire \_ces_0_2_io_outs_right[63] ;
 wire \_ces_0_2_io_outs_right[6] ;
 wire \_ces_0_2_io_outs_right[7] ;
 wire \_ces_0_2_io_outs_right[8] ;
 wire \_ces_0_2_io_outs_right[9] ;
 wire \_ces_0_2_io_outs_up[0] ;
 wire \_ces_0_2_io_outs_up[10] ;
 wire \_ces_0_2_io_outs_up[11] ;
 wire \_ces_0_2_io_outs_up[12] ;
 wire \_ces_0_2_io_outs_up[13] ;
 wire \_ces_0_2_io_outs_up[14] ;
 wire \_ces_0_2_io_outs_up[15] ;
 wire \_ces_0_2_io_outs_up[16] ;
 wire \_ces_0_2_io_outs_up[17] ;
 wire \_ces_0_2_io_outs_up[18] ;
 wire \_ces_0_2_io_outs_up[19] ;
 wire \_ces_0_2_io_outs_up[1] ;
 wire \_ces_0_2_io_outs_up[20] ;
 wire \_ces_0_2_io_outs_up[21] ;
 wire \_ces_0_2_io_outs_up[22] ;
 wire \_ces_0_2_io_outs_up[23] ;
 wire \_ces_0_2_io_outs_up[24] ;
 wire \_ces_0_2_io_outs_up[25] ;
 wire \_ces_0_2_io_outs_up[26] ;
 wire \_ces_0_2_io_outs_up[27] ;
 wire \_ces_0_2_io_outs_up[28] ;
 wire \_ces_0_2_io_outs_up[29] ;
 wire \_ces_0_2_io_outs_up[2] ;
 wire \_ces_0_2_io_outs_up[30] ;
 wire \_ces_0_2_io_outs_up[31] ;
 wire \_ces_0_2_io_outs_up[32] ;
 wire \_ces_0_2_io_outs_up[33] ;
 wire \_ces_0_2_io_outs_up[34] ;
 wire \_ces_0_2_io_outs_up[35] ;
 wire \_ces_0_2_io_outs_up[36] ;
 wire \_ces_0_2_io_outs_up[37] ;
 wire \_ces_0_2_io_outs_up[38] ;
 wire \_ces_0_2_io_outs_up[39] ;
 wire \_ces_0_2_io_outs_up[3] ;
 wire \_ces_0_2_io_outs_up[40] ;
 wire \_ces_0_2_io_outs_up[41] ;
 wire \_ces_0_2_io_outs_up[42] ;
 wire \_ces_0_2_io_outs_up[43] ;
 wire \_ces_0_2_io_outs_up[44] ;
 wire \_ces_0_2_io_outs_up[45] ;
 wire \_ces_0_2_io_outs_up[46] ;
 wire \_ces_0_2_io_outs_up[47] ;
 wire \_ces_0_2_io_outs_up[48] ;
 wire \_ces_0_2_io_outs_up[49] ;
 wire \_ces_0_2_io_outs_up[4] ;
 wire \_ces_0_2_io_outs_up[50] ;
 wire \_ces_0_2_io_outs_up[51] ;
 wire \_ces_0_2_io_outs_up[52] ;
 wire \_ces_0_2_io_outs_up[53] ;
 wire \_ces_0_2_io_outs_up[54] ;
 wire \_ces_0_2_io_outs_up[55] ;
 wire \_ces_0_2_io_outs_up[56] ;
 wire \_ces_0_2_io_outs_up[57] ;
 wire \_ces_0_2_io_outs_up[58] ;
 wire \_ces_0_2_io_outs_up[59] ;
 wire \_ces_0_2_io_outs_up[5] ;
 wire \_ces_0_2_io_outs_up[60] ;
 wire \_ces_0_2_io_outs_up[61] ;
 wire \_ces_0_2_io_outs_up[62] ;
 wire \_ces_0_2_io_outs_up[63] ;
 wire \_ces_0_2_io_outs_up[6] ;
 wire \_ces_0_2_io_outs_up[7] ;
 wire \_ces_0_2_io_outs_up[8] ;
 wire \_ces_0_2_io_outs_up[9] ;
 wire _ces_0_3_io_lsbOuts_0;
 wire _ces_0_3_io_lsbOuts_1;
 wire _ces_0_3_io_lsbOuts_2;
 wire _ces_0_3_io_lsbOuts_3;
 wire \_ces_0_3_io_outs_left[0] ;
 wire \_ces_0_3_io_outs_left[10] ;
 wire \_ces_0_3_io_outs_left[11] ;
 wire \_ces_0_3_io_outs_left[12] ;
 wire \_ces_0_3_io_outs_left[13] ;
 wire \_ces_0_3_io_outs_left[14] ;
 wire \_ces_0_3_io_outs_left[15] ;
 wire \_ces_0_3_io_outs_left[16] ;
 wire \_ces_0_3_io_outs_left[17] ;
 wire \_ces_0_3_io_outs_left[18] ;
 wire \_ces_0_3_io_outs_left[19] ;
 wire \_ces_0_3_io_outs_left[1] ;
 wire \_ces_0_3_io_outs_left[20] ;
 wire \_ces_0_3_io_outs_left[21] ;
 wire \_ces_0_3_io_outs_left[22] ;
 wire \_ces_0_3_io_outs_left[23] ;
 wire \_ces_0_3_io_outs_left[24] ;
 wire \_ces_0_3_io_outs_left[25] ;
 wire \_ces_0_3_io_outs_left[26] ;
 wire \_ces_0_3_io_outs_left[27] ;
 wire \_ces_0_3_io_outs_left[28] ;
 wire \_ces_0_3_io_outs_left[29] ;
 wire \_ces_0_3_io_outs_left[2] ;
 wire \_ces_0_3_io_outs_left[30] ;
 wire \_ces_0_3_io_outs_left[31] ;
 wire \_ces_0_3_io_outs_left[32] ;
 wire \_ces_0_3_io_outs_left[33] ;
 wire \_ces_0_3_io_outs_left[34] ;
 wire \_ces_0_3_io_outs_left[35] ;
 wire \_ces_0_3_io_outs_left[36] ;
 wire \_ces_0_3_io_outs_left[37] ;
 wire \_ces_0_3_io_outs_left[38] ;
 wire \_ces_0_3_io_outs_left[39] ;
 wire \_ces_0_3_io_outs_left[3] ;
 wire \_ces_0_3_io_outs_left[40] ;
 wire \_ces_0_3_io_outs_left[41] ;
 wire \_ces_0_3_io_outs_left[42] ;
 wire \_ces_0_3_io_outs_left[43] ;
 wire \_ces_0_3_io_outs_left[44] ;
 wire \_ces_0_3_io_outs_left[45] ;
 wire \_ces_0_3_io_outs_left[46] ;
 wire \_ces_0_3_io_outs_left[47] ;
 wire \_ces_0_3_io_outs_left[48] ;
 wire \_ces_0_3_io_outs_left[49] ;
 wire \_ces_0_3_io_outs_left[4] ;
 wire \_ces_0_3_io_outs_left[50] ;
 wire \_ces_0_3_io_outs_left[51] ;
 wire \_ces_0_3_io_outs_left[52] ;
 wire \_ces_0_3_io_outs_left[53] ;
 wire \_ces_0_3_io_outs_left[54] ;
 wire \_ces_0_3_io_outs_left[55] ;
 wire \_ces_0_3_io_outs_left[56] ;
 wire \_ces_0_3_io_outs_left[57] ;
 wire \_ces_0_3_io_outs_left[58] ;
 wire \_ces_0_3_io_outs_left[59] ;
 wire \_ces_0_3_io_outs_left[5] ;
 wire \_ces_0_3_io_outs_left[60] ;
 wire \_ces_0_3_io_outs_left[61] ;
 wire \_ces_0_3_io_outs_left[62] ;
 wire \_ces_0_3_io_outs_left[63] ;
 wire \_ces_0_3_io_outs_left[6] ;
 wire \_ces_0_3_io_outs_left[7] ;
 wire \_ces_0_3_io_outs_left[8] ;
 wire \_ces_0_3_io_outs_left[9] ;
 wire \_ces_0_3_io_outs_up[0] ;
 wire \_ces_0_3_io_outs_up[10] ;
 wire \_ces_0_3_io_outs_up[11] ;
 wire \_ces_0_3_io_outs_up[12] ;
 wire \_ces_0_3_io_outs_up[13] ;
 wire \_ces_0_3_io_outs_up[14] ;
 wire \_ces_0_3_io_outs_up[15] ;
 wire \_ces_0_3_io_outs_up[16] ;
 wire \_ces_0_3_io_outs_up[17] ;
 wire \_ces_0_3_io_outs_up[18] ;
 wire \_ces_0_3_io_outs_up[19] ;
 wire \_ces_0_3_io_outs_up[1] ;
 wire \_ces_0_3_io_outs_up[20] ;
 wire \_ces_0_3_io_outs_up[21] ;
 wire \_ces_0_3_io_outs_up[22] ;
 wire \_ces_0_3_io_outs_up[23] ;
 wire \_ces_0_3_io_outs_up[24] ;
 wire \_ces_0_3_io_outs_up[25] ;
 wire \_ces_0_3_io_outs_up[26] ;
 wire \_ces_0_3_io_outs_up[27] ;
 wire \_ces_0_3_io_outs_up[28] ;
 wire \_ces_0_3_io_outs_up[29] ;
 wire \_ces_0_3_io_outs_up[2] ;
 wire \_ces_0_3_io_outs_up[30] ;
 wire \_ces_0_3_io_outs_up[31] ;
 wire \_ces_0_3_io_outs_up[32] ;
 wire \_ces_0_3_io_outs_up[33] ;
 wire \_ces_0_3_io_outs_up[34] ;
 wire \_ces_0_3_io_outs_up[35] ;
 wire \_ces_0_3_io_outs_up[36] ;
 wire \_ces_0_3_io_outs_up[37] ;
 wire \_ces_0_3_io_outs_up[38] ;
 wire \_ces_0_3_io_outs_up[39] ;
 wire \_ces_0_3_io_outs_up[3] ;
 wire \_ces_0_3_io_outs_up[40] ;
 wire \_ces_0_3_io_outs_up[41] ;
 wire \_ces_0_3_io_outs_up[42] ;
 wire \_ces_0_3_io_outs_up[43] ;
 wire \_ces_0_3_io_outs_up[44] ;
 wire \_ces_0_3_io_outs_up[45] ;
 wire \_ces_0_3_io_outs_up[46] ;
 wire \_ces_0_3_io_outs_up[47] ;
 wire \_ces_0_3_io_outs_up[48] ;
 wire \_ces_0_3_io_outs_up[49] ;
 wire \_ces_0_3_io_outs_up[4] ;
 wire \_ces_0_3_io_outs_up[50] ;
 wire \_ces_0_3_io_outs_up[51] ;
 wire \_ces_0_3_io_outs_up[52] ;
 wire \_ces_0_3_io_outs_up[53] ;
 wire \_ces_0_3_io_outs_up[54] ;
 wire \_ces_0_3_io_outs_up[55] ;
 wire \_ces_0_3_io_outs_up[56] ;
 wire \_ces_0_3_io_outs_up[57] ;
 wire \_ces_0_3_io_outs_up[58] ;
 wire \_ces_0_3_io_outs_up[59] ;
 wire \_ces_0_3_io_outs_up[5] ;
 wire \_ces_0_3_io_outs_up[60] ;
 wire \_ces_0_3_io_outs_up[61] ;
 wire \_ces_0_3_io_outs_up[62] ;
 wire \_ces_0_3_io_outs_up[63] ;
 wire \_ces_0_3_io_outs_up[6] ;
 wire \_ces_0_3_io_outs_up[7] ;
 wire \_ces_0_3_io_outs_up[8] ;
 wire \_ces_0_3_io_outs_up[9] ;
 wire _ces_1_0_io_lsbOuts_1;
 wire _ces_1_0_io_lsbOuts_2;
 wire _ces_1_0_io_lsbOuts_3;
 wire \_ces_1_0_io_outs_down[0] ;
 wire \_ces_1_0_io_outs_down[10] ;
 wire \_ces_1_0_io_outs_down[11] ;
 wire \_ces_1_0_io_outs_down[12] ;
 wire \_ces_1_0_io_outs_down[13] ;
 wire \_ces_1_0_io_outs_down[14] ;
 wire \_ces_1_0_io_outs_down[15] ;
 wire \_ces_1_0_io_outs_down[16] ;
 wire \_ces_1_0_io_outs_down[17] ;
 wire \_ces_1_0_io_outs_down[18] ;
 wire \_ces_1_0_io_outs_down[19] ;
 wire \_ces_1_0_io_outs_down[1] ;
 wire \_ces_1_0_io_outs_down[20] ;
 wire \_ces_1_0_io_outs_down[21] ;
 wire \_ces_1_0_io_outs_down[22] ;
 wire \_ces_1_0_io_outs_down[23] ;
 wire \_ces_1_0_io_outs_down[24] ;
 wire \_ces_1_0_io_outs_down[25] ;
 wire \_ces_1_0_io_outs_down[26] ;
 wire \_ces_1_0_io_outs_down[27] ;
 wire \_ces_1_0_io_outs_down[28] ;
 wire \_ces_1_0_io_outs_down[29] ;
 wire \_ces_1_0_io_outs_down[2] ;
 wire \_ces_1_0_io_outs_down[30] ;
 wire \_ces_1_0_io_outs_down[31] ;
 wire \_ces_1_0_io_outs_down[32] ;
 wire \_ces_1_0_io_outs_down[33] ;
 wire \_ces_1_0_io_outs_down[34] ;
 wire \_ces_1_0_io_outs_down[35] ;
 wire \_ces_1_0_io_outs_down[36] ;
 wire \_ces_1_0_io_outs_down[37] ;
 wire \_ces_1_0_io_outs_down[38] ;
 wire \_ces_1_0_io_outs_down[39] ;
 wire \_ces_1_0_io_outs_down[3] ;
 wire \_ces_1_0_io_outs_down[40] ;
 wire \_ces_1_0_io_outs_down[41] ;
 wire \_ces_1_0_io_outs_down[42] ;
 wire \_ces_1_0_io_outs_down[43] ;
 wire \_ces_1_0_io_outs_down[44] ;
 wire \_ces_1_0_io_outs_down[45] ;
 wire \_ces_1_0_io_outs_down[46] ;
 wire \_ces_1_0_io_outs_down[47] ;
 wire \_ces_1_0_io_outs_down[48] ;
 wire \_ces_1_0_io_outs_down[49] ;
 wire \_ces_1_0_io_outs_down[4] ;
 wire \_ces_1_0_io_outs_down[50] ;
 wire \_ces_1_0_io_outs_down[51] ;
 wire \_ces_1_0_io_outs_down[52] ;
 wire \_ces_1_0_io_outs_down[53] ;
 wire \_ces_1_0_io_outs_down[54] ;
 wire \_ces_1_0_io_outs_down[55] ;
 wire \_ces_1_0_io_outs_down[56] ;
 wire \_ces_1_0_io_outs_down[57] ;
 wire \_ces_1_0_io_outs_down[58] ;
 wire \_ces_1_0_io_outs_down[59] ;
 wire \_ces_1_0_io_outs_down[5] ;
 wire \_ces_1_0_io_outs_down[60] ;
 wire \_ces_1_0_io_outs_down[61] ;
 wire \_ces_1_0_io_outs_down[62] ;
 wire \_ces_1_0_io_outs_down[63] ;
 wire \_ces_1_0_io_outs_down[6] ;
 wire \_ces_1_0_io_outs_down[7] ;
 wire \_ces_1_0_io_outs_down[8] ;
 wire \_ces_1_0_io_outs_down[9] ;
 wire \_ces_1_0_io_outs_right[0] ;
 wire \_ces_1_0_io_outs_right[10] ;
 wire \_ces_1_0_io_outs_right[11] ;
 wire \_ces_1_0_io_outs_right[12] ;
 wire \_ces_1_0_io_outs_right[13] ;
 wire \_ces_1_0_io_outs_right[14] ;
 wire \_ces_1_0_io_outs_right[15] ;
 wire \_ces_1_0_io_outs_right[16] ;
 wire \_ces_1_0_io_outs_right[17] ;
 wire \_ces_1_0_io_outs_right[18] ;
 wire \_ces_1_0_io_outs_right[19] ;
 wire \_ces_1_0_io_outs_right[1] ;
 wire \_ces_1_0_io_outs_right[20] ;
 wire \_ces_1_0_io_outs_right[21] ;
 wire \_ces_1_0_io_outs_right[22] ;
 wire \_ces_1_0_io_outs_right[23] ;
 wire \_ces_1_0_io_outs_right[24] ;
 wire \_ces_1_0_io_outs_right[25] ;
 wire \_ces_1_0_io_outs_right[26] ;
 wire \_ces_1_0_io_outs_right[27] ;
 wire \_ces_1_0_io_outs_right[28] ;
 wire \_ces_1_0_io_outs_right[29] ;
 wire \_ces_1_0_io_outs_right[2] ;
 wire \_ces_1_0_io_outs_right[30] ;
 wire \_ces_1_0_io_outs_right[31] ;
 wire \_ces_1_0_io_outs_right[32] ;
 wire \_ces_1_0_io_outs_right[33] ;
 wire \_ces_1_0_io_outs_right[34] ;
 wire \_ces_1_0_io_outs_right[35] ;
 wire \_ces_1_0_io_outs_right[36] ;
 wire \_ces_1_0_io_outs_right[37] ;
 wire \_ces_1_0_io_outs_right[38] ;
 wire \_ces_1_0_io_outs_right[39] ;
 wire \_ces_1_0_io_outs_right[3] ;
 wire \_ces_1_0_io_outs_right[40] ;
 wire \_ces_1_0_io_outs_right[41] ;
 wire \_ces_1_0_io_outs_right[42] ;
 wire \_ces_1_0_io_outs_right[43] ;
 wire \_ces_1_0_io_outs_right[44] ;
 wire \_ces_1_0_io_outs_right[45] ;
 wire \_ces_1_0_io_outs_right[46] ;
 wire \_ces_1_0_io_outs_right[47] ;
 wire \_ces_1_0_io_outs_right[48] ;
 wire \_ces_1_0_io_outs_right[49] ;
 wire \_ces_1_0_io_outs_right[4] ;
 wire \_ces_1_0_io_outs_right[50] ;
 wire \_ces_1_0_io_outs_right[51] ;
 wire \_ces_1_0_io_outs_right[52] ;
 wire \_ces_1_0_io_outs_right[53] ;
 wire \_ces_1_0_io_outs_right[54] ;
 wire \_ces_1_0_io_outs_right[55] ;
 wire \_ces_1_0_io_outs_right[56] ;
 wire \_ces_1_0_io_outs_right[57] ;
 wire \_ces_1_0_io_outs_right[58] ;
 wire \_ces_1_0_io_outs_right[59] ;
 wire \_ces_1_0_io_outs_right[5] ;
 wire \_ces_1_0_io_outs_right[60] ;
 wire \_ces_1_0_io_outs_right[61] ;
 wire \_ces_1_0_io_outs_right[62] ;
 wire \_ces_1_0_io_outs_right[63] ;
 wire \_ces_1_0_io_outs_right[6] ;
 wire \_ces_1_0_io_outs_right[7] ;
 wire \_ces_1_0_io_outs_right[8] ;
 wire \_ces_1_0_io_outs_right[9] ;
 wire \_ces_1_0_io_outs_up[0] ;
 wire \_ces_1_0_io_outs_up[10] ;
 wire \_ces_1_0_io_outs_up[11] ;
 wire \_ces_1_0_io_outs_up[12] ;
 wire \_ces_1_0_io_outs_up[13] ;
 wire \_ces_1_0_io_outs_up[14] ;
 wire \_ces_1_0_io_outs_up[15] ;
 wire \_ces_1_0_io_outs_up[16] ;
 wire \_ces_1_0_io_outs_up[17] ;
 wire \_ces_1_0_io_outs_up[18] ;
 wire \_ces_1_0_io_outs_up[19] ;
 wire \_ces_1_0_io_outs_up[1] ;
 wire \_ces_1_0_io_outs_up[20] ;
 wire \_ces_1_0_io_outs_up[21] ;
 wire \_ces_1_0_io_outs_up[22] ;
 wire \_ces_1_0_io_outs_up[23] ;
 wire \_ces_1_0_io_outs_up[24] ;
 wire \_ces_1_0_io_outs_up[25] ;
 wire \_ces_1_0_io_outs_up[26] ;
 wire \_ces_1_0_io_outs_up[27] ;
 wire \_ces_1_0_io_outs_up[28] ;
 wire \_ces_1_0_io_outs_up[29] ;
 wire \_ces_1_0_io_outs_up[2] ;
 wire \_ces_1_0_io_outs_up[30] ;
 wire \_ces_1_0_io_outs_up[31] ;
 wire \_ces_1_0_io_outs_up[32] ;
 wire \_ces_1_0_io_outs_up[33] ;
 wire \_ces_1_0_io_outs_up[34] ;
 wire \_ces_1_0_io_outs_up[35] ;
 wire \_ces_1_0_io_outs_up[36] ;
 wire \_ces_1_0_io_outs_up[37] ;
 wire \_ces_1_0_io_outs_up[38] ;
 wire \_ces_1_0_io_outs_up[39] ;
 wire \_ces_1_0_io_outs_up[3] ;
 wire \_ces_1_0_io_outs_up[40] ;
 wire \_ces_1_0_io_outs_up[41] ;
 wire \_ces_1_0_io_outs_up[42] ;
 wire \_ces_1_0_io_outs_up[43] ;
 wire \_ces_1_0_io_outs_up[44] ;
 wire \_ces_1_0_io_outs_up[45] ;
 wire \_ces_1_0_io_outs_up[46] ;
 wire \_ces_1_0_io_outs_up[47] ;
 wire \_ces_1_0_io_outs_up[48] ;
 wire \_ces_1_0_io_outs_up[49] ;
 wire \_ces_1_0_io_outs_up[4] ;
 wire \_ces_1_0_io_outs_up[50] ;
 wire \_ces_1_0_io_outs_up[51] ;
 wire \_ces_1_0_io_outs_up[52] ;
 wire \_ces_1_0_io_outs_up[53] ;
 wire \_ces_1_0_io_outs_up[54] ;
 wire \_ces_1_0_io_outs_up[55] ;
 wire \_ces_1_0_io_outs_up[56] ;
 wire \_ces_1_0_io_outs_up[57] ;
 wire \_ces_1_0_io_outs_up[58] ;
 wire \_ces_1_0_io_outs_up[59] ;
 wire \_ces_1_0_io_outs_up[5] ;
 wire \_ces_1_0_io_outs_up[60] ;
 wire \_ces_1_0_io_outs_up[61] ;
 wire \_ces_1_0_io_outs_up[62] ;
 wire \_ces_1_0_io_outs_up[63] ;
 wire \_ces_1_0_io_outs_up[6] ;
 wire \_ces_1_0_io_outs_up[7] ;
 wire \_ces_1_0_io_outs_up[8] ;
 wire \_ces_1_0_io_outs_up[9] ;
 wire _ces_1_1_io_lsbOuts_1;
 wire _ces_1_1_io_lsbOuts_2;
 wire _ces_1_1_io_lsbOuts_3;
 wire \_ces_1_1_io_outs_down[0] ;
 wire \_ces_1_1_io_outs_down[10] ;
 wire \_ces_1_1_io_outs_down[11] ;
 wire \_ces_1_1_io_outs_down[12] ;
 wire \_ces_1_1_io_outs_down[13] ;
 wire \_ces_1_1_io_outs_down[14] ;
 wire \_ces_1_1_io_outs_down[15] ;
 wire \_ces_1_1_io_outs_down[16] ;
 wire \_ces_1_1_io_outs_down[17] ;
 wire \_ces_1_1_io_outs_down[18] ;
 wire \_ces_1_1_io_outs_down[19] ;
 wire \_ces_1_1_io_outs_down[1] ;
 wire \_ces_1_1_io_outs_down[20] ;
 wire \_ces_1_1_io_outs_down[21] ;
 wire \_ces_1_1_io_outs_down[22] ;
 wire \_ces_1_1_io_outs_down[23] ;
 wire \_ces_1_1_io_outs_down[24] ;
 wire \_ces_1_1_io_outs_down[25] ;
 wire \_ces_1_1_io_outs_down[26] ;
 wire \_ces_1_1_io_outs_down[27] ;
 wire \_ces_1_1_io_outs_down[28] ;
 wire \_ces_1_1_io_outs_down[29] ;
 wire \_ces_1_1_io_outs_down[2] ;
 wire \_ces_1_1_io_outs_down[30] ;
 wire \_ces_1_1_io_outs_down[31] ;
 wire \_ces_1_1_io_outs_down[32] ;
 wire \_ces_1_1_io_outs_down[33] ;
 wire \_ces_1_1_io_outs_down[34] ;
 wire \_ces_1_1_io_outs_down[35] ;
 wire \_ces_1_1_io_outs_down[36] ;
 wire \_ces_1_1_io_outs_down[37] ;
 wire \_ces_1_1_io_outs_down[38] ;
 wire \_ces_1_1_io_outs_down[39] ;
 wire \_ces_1_1_io_outs_down[3] ;
 wire \_ces_1_1_io_outs_down[40] ;
 wire \_ces_1_1_io_outs_down[41] ;
 wire \_ces_1_1_io_outs_down[42] ;
 wire \_ces_1_1_io_outs_down[43] ;
 wire \_ces_1_1_io_outs_down[44] ;
 wire \_ces_1_1_io_outs_down[45] ;
 wire \_ces_1_1_io_outs_down[46] ;
 wire \_ces_1_1_io_outs_down[47] ;
 wire \_ces_1_1_io_outs_down[48] ;
 wire \_ces_1_1_io_outs_down[49] ;
 wire \_ces_1_1_io_outs_down[4] ;
 wire \_ces_1_1_io_outs_down[50] ;
 wire \_ces_1_1_io_outs_down[51] ;
 wire \_ces_1_1_io_outs_down[52] ;
 wire \_ces_1_1_io_outs_down[53] ;
 wire \_ces_1_1_io_outs_down[54] ;
 wire \_ces_1_1_io_outs_down[55] ;
 wire \_ces_1_1_io_outs_down[56] ;
 wire \_ces_1_1_io_outs_down[57] ;
 wire \_ces_1_1_io_outs_down[58] ;
 wire \_ces_1_1_io_outs_down[59] ;
 wire \_ces_1_1_io_outs_down[5] ;
 wire \_ces_1_1_io_outs_down[60] ;
 wire \_ces_1_1_io_outs_down[61] ;
 wire \_ces_1_1_io_outs_down[62] ;
 wire \_ces_1_1_io_outs_down[63] ;
 wire \_ces_1_1_io_outs_down[6] ;
 wire \_ces_1_1_io_outs_down[7] ;
 wire \_ces_1_1_io_outs_down[8] ;
 wire \_ces_1_1_io_outs_down[9] ;
 wire \_ces_1_1_io_outs_left[0] ;
 wire \_ces_1_1_io_outs_left[10] ;
 wire \_ces_1_1_io_outs_left[11] ;
 wire \_ces_1_1_io_outs_left[12] ;
 wire \_ces_1_1_io_outs_left[13] ;
 wire \_ces_1_1_io_outs_left[14] ;
 wire \_ces_1_1_io_outs_left[15] ;
 wire \_ces_1_1_io_outs_left[16] ;
 wire \_ces_1_1_io_outs_left[17] ;
 wire \_ces_1_1_io_outs_left[18] ;
 wire \_ces_1_1_io_outs_left[19] ;
 wire \_ces_1_1_io_outs_left[1] ;
 wire \_ces_1_1_io_outs_left[20] ;
 wire \_ces_1_1_io_outs_left[21] ;
 wire \_ces_1_1_io_outs_left[22] ;
 wire \_ces_1_1_io_outs_left[23] ;
 wire \_ces_1_1_io_outs_left[24] ;
 wire \_ces_1_1_io_outs_left[25] ;
 wire \_ces_1_1_io_outs_left[26] ;
 wire \_ces_1_1_io_outs_left[27] ;
 wire \_ces_1_1_io_outs_left[28] ;
 wire \_ces_1_1_io_outs_left[29] ;
 wire \_ces_1_1_io_outs_left[2] ;
 wire \_ces_1_1_io_outs_left[30] ;
 wire \_ces_1_1_io_outs_left[31] ;
 wire \_ces_1_1_io_outs_left[32] ;
 wire \_ces_1_1_io_outs_left[33] ;
 wire \_ces_1_1_io_outs_left[34] ;
 wire \_ces_1_1_io_outs_left[35] ;
 wire \_ces_1_1_io_outs_left[36] ;
 wire \_ces_1_1_io_outs_left[37] ;
 wire \_ces_1_1_io_outs_left[38] ;
 wire \_ces_1_1_io_outs_left[39] ;
 wire \_ces_1_1_io_outs_left[3] ;
 wire \_ces_1_1_io_outs_left[40] ;
 wire \_ces_1_1_io_outs_left[41] ;
 wire \_ces_1_1_io_outs_left[42] ;
 wire \_ces_1_1_io_outs_left[43] ;
 wire \_ces_1_1_io_outs_left[44] ;
 wire \_ces_1_1_io_outs_left[45] ;
 wire \_ces_1_1_io_outs_left[46] ;
 wire \_ces_1_1_io_outs_left[47] ;
 wire \_ces_1_1_io_outs_left[48] ;
 wire \_ces_1_1_io_outs_left[49] ;
 wire \_ces_1_1_io_outs_left[4] ;
 wire \_ces_1_1_io_outs_left[50] ;
 wire \_ces_1_1_io_outs_left[51] ;
 wire \_ces_1_1_io_outs_left[52] ;
 wire \_ces_1_1_io_outs_left[53] ;
 wire \_ces_1_1_io_outs_left[54] ;
 wire \_ces_1_1_io_outs_left[55] ;
 wire \_ces_1_1_io_outs_left[56] ;
 wire \_ces_1_1_io_outs_left[57] ;
 wire \_ces_1_1_io_outs_left[58] ;
 wire \_ces_1_1_io_outs_left[59] ;
 wire \_ces_1_1_io_outs_left[5] ;
 wire \_ces_1_1_io_outs_left[60] ;
 wire \_ces_1_1_io_outs_left[61] ;
 wire \_ces_1_1_io_outs_left[62] ;
 wire \_ces_1_1_io_outs_left[63] ;
 wire \_ces_1_1_io_outs_left[6] ;
 wire \_ces_1_1_io_outs_left[7] ;
 wire \_ces_1_1_io_outs_left[8] ;
 wire \_ces_1_1_io_outs_left[9] ;
 wire \_ces_1_1_io_outs_right[0] ;
 wire \_ces_1_1_io_outs_right[10] ;
 wire \_ces_1_1_io_outs_right[11] ;
 wire \_ces_1_1_io_outs_right[12] ;
 wire \_ces_1_1_io_outs_right[13] ;
 wire \_ces_1_1_io_outs_right[14] ;
 wire \_ces_1_1_io_outs_right[15] ;
 wire \_ces_1_1_io_outs_right[16] ;
 wire \_ces_1_1_io_outs_right[17] ;
 wire \_ces_1_1_io_outs_right[18] ;
 wire \_ces_1_1_io_outs_right[19] ;
 wire \_ces_1_1_io_outs_right[1] ;
 wire \_ces_1_1_io_outs_right[20] ;
 wire \_ces_1_1_io_outs_right[21] ;
 wire \_ces_1_1_io_outs_right[22] ;
 wire \_ces_1_1_io_outs_right[23] ;
 wire \_ces_1_1_io_outs_right[24] ;
 wire \_ces_1_1_io_outs_right[25] ;
 wire \_ces_1_1_io_outs_right[26] ;
 wire \_ces_1_1_io_outs_right[27] ;
 wire \_ces_1_1_io_outs_right[28] ;
 wire \_ces_1_1_io_outs_right[29] ;
 wire \_ces_1_1_io_outs_right[2] ;
 wire \_ces_1_1_io_outs_right[30] ;
 wire \_ces_1_1_io_outs_right[31] ;
 wire \_ces_1_1_io_outs_right[32] ;
 wire \_ces_1_1_io_outs_right[33] ;
 wire \_ces_1_1_io_outs_right[34] ;
 wire \_ces_1_1_io_outs_right[35] ;
 wire \_ces_1_1_io_outs_right[36] ;
 wire \_ces_1_1_io_outs_right[37] ;
 wire \_ces_1_1_io_outs_right[38] ;
 wire \_ces_1_1_io_outs_right[39] ;
 wire \_ces_1_1_io_outs_right[3] ;
 wire \_ces_1_1_io_outs_right[40] ;
 wire \_ces_1_1_io_outs_right[41] ;
 wire \_ces_1_1_io_outs_right[42] ;
 wire \_ces_1_1_io_outs_right[43] ;
 wire \_ces_1_1_io_outs_right[44] ;
 wire \_ces_1_1_io_outs_right[45] ;
 wire \_ces_1_1_io_outs_right[46] ;
 wire \_ces_1_1_io_outs_right[47] ;
 wire \_ces_1_1_io_outs_right[48] ;
 wire \_ces_1_1_io_outs_right[49] ;
 wire \_ces_1_1_io_outs_right[4] ;
 wire \_ces_1_1_io_outs_right[50] ;
 wire \_ces_1_1_io_outs_right[51] ;
 wire \_ces_1_1_io_outs_right[52] ;
 wire \_ces_1_1_io_outs_right[53] ;
 wire \_ces_1_1_io_outs_right[54] ;
 wire \_ces_1_1_io_outs_right[55] ;
 wire \_ces_1_1_io_outs_right[56] ;
 wire \_ces_1_1_io_outs_right[57] ;
 wire \_ces_1_1_io_outs_right[58] ;
 wire \_ces_1_1_io_outs_right[59] ;
 wire \_ces_1_1_io_outs_right[5] ;
 wire \_ces_1_1_io_outs_right[60] ;
 wire \_ces_1_1_io_outs_right[61] ;
 wire \_ces_1_1_io_outs_right[62] ;
 wire \_ces_1_1_io_outs_right[63] ;
 wire \_ces_1_1_io_outs_right[6] ;
 wire \_ces_1_1_io_outs_right[7] ;
 wire \_ces_1_1_io_outs_right[8] ;
 wire \_ces_1_1_io_outs_right[9] ;
 wire \_ces_1_1_io_outs_up[0] ;
 wire \_ces_1_1_io_outs_up[10] ;
 wire \_ces_1_1_io_outs_up[11] ;
 wire \_ces_1_1_io_outs_up[12] ;
 wire \_ces_1_1_io_outs_up[13] ;
 wire \_ces_1_1_io_outs_up[14] ;
 wire \_ces_1_1_io_outs_up[15] ;
 wire \_ces_1_1_io_outs_up[16] ;
 wire \_ces_1_1_io_outs_up[17] ;
 wire \_ces_1_1_io_outs_up[18] ;
 wire \_ces_1_1_io_outs_up[19] ;
 wire \_ces_1_1_io_outs_up[1] ;
 wire \_ces_1_1_io_outs_up[20] ;
 wire \_ces_1_1_io_outs_up[21] ;
 wire \_ces_1_1_io_outs_up[22] ;
 wire \_ces_1_1_io_outs_up[23] ;
 wire \_ces_1_1_io_outs_up[24] ;
 wire \_ces_1_1_io_outs_up[25] ;
 wire \_ces_1_1_io_outs_up[26] ;
 wire \_ces_1_1_io_outs_up[27] ;
 wire \_ces_1_1_io_outs_up[28] ;
 wire \_ces_1_1_io_outs_up[29] ;
 wire \_ces_1_1_io_outs_up[2] ;
 wire \_ces_1_1_io_outs_up[30] ;
 wire \_ces_1_1_io_outs_up[31] ;
 wire \_ces_1_1_io_outs_up[32] ;
 wire \_ces_1_1_io_outs_up[33] ;
 wire \_ces_1_1_io_outs_up[34] ;
 wire \_ces_1_1_io_outs_up[35] ;
 wire \_ces_1_1_io_outs_up[36] ;
 wire \_ces_1_1_io_outs_up[37] ;
 wire \_ces_1_1_io_outs_up[38] ;
 wire \_ces_1_1_io_outs_up[39] ;
 wire \_ces_1_1_io_outs_up[3] ;
 wire \_ces_1_1_io_outs_up[40] ;
 wire \_ces_1_1_io_outs_up[41] ;
 wire \_ces_1_1_io_outs_up[42] ;
 wire \_ces_1_1_io_outs_up[43] ;
 wire \_ces_1_1_io_outs_up[44] ;
 wire \_ces_1_1_io_outs_up[45] ;
 wire \_ces_1_1_io_outs_up[46] ;
 wire \_ces_1_1_io_outs_up[47] ;
 wire \_ces_1_1_io_outs_up[48] ;
 wire \_ces_1_1_io_outs_up[49] ;
 wire \_ces_1_1_io_outs_up[4] ;
 wire \_ces_1_1_io_outs_up[50] ;
 wire \_ces_1_1_io_outs_up[51] ;
 wire \_ces_1_1_io_outs_up[52] ;
 wire \_ces_1_1_io_outs_up[53] ;
 wire \_ces_1_1_io_outs_up[54] ;
 wire \_ces_1_1_io_outs_up[55] ;
 wire \_ces_1_1_io_outs_up[56] ;
 wire \_ces_1_1_io_outs_up[57] ;
 wire \_ces_1_1_io_outs_up[58] ;
 wire \_ces_1_1_io_outs_up[59] ;
 wire \_ces_1_1_io_outs_up[5] ;
 wire \_ces_1_1_io_outs_up[60] ;
 wire \_ces_1_1_io_outs_up[61] ;
 wire \_ces_1_1_io_outs_up[62] ;
 wire \_ces_1_1_io_outs_up[63] ;
 wire \_ces_1_1_io_outs_up[6] ;
 wire \_ces_1_1_io_outs_up[7] ;
 wire \_ces_1_1_io_outs_up[8] ;
 wire \_ces_1_1_io_outs_up[9] ;
 wire _ces_1_2_io_lsbOuts_1;
 wire _ces_1_2_io_lsbOuts_2;
 wire _ces_1_2_io_lsbOuts_3;
 wire \_ces_1_2_io_outs_down[0] ;
 wire \_ces_1_2_io_outs_down[10] ;
 wire \_ces_1_2_io_outs_down[11] ;
 wire \_ces_1_2_io_outs_down[12] ;
 wire \_ces_1_2_io_outs_down[13] ;
 wire \_ces_1_2_io_outs_down[14] ;
 wire \_ces_1_2_io_outs_down[15] ;
 wire \_ces_1_2_io_outs_down[16] ;
 wire \_ces_1_2_io_outs_down[17] ;
 wire \_ces_1_2_io_outs_down[18] ;
 wire \_ces_1_2_io_outs_down[19] ;
 wire \_ces_1_2_io_outs_down[1] ;
 wire \_ces_1_2_io_outs_down[20] ;
 wire \_ces_1_2_io_outs_down[21] ;
 wire \_ces_1_2_io_outs_down[22] ;
 wire \_ces_1_2_io_outs_down[23] ;
 wire \_ces_1_2_io_outs_down[24] ;
 wire \_ces_1_2_io_outs_down[25] ;
 wire \_ces_1_2_io_outs_down[26] ;
 wire \_ces_1_2_io_outs_down[27] ;
 wire \_ces_1_2_io_outs_down[28] ;
 wire \_ces_1_2_io_outs_down[29] ;
 wire \_ces_1_2_io_outs_down[2] ;
 wire \_ces_1_2_io_outs_down[30] ;
 wire \_ces_1_2_io_outs_down[31] ;
 wire \_ces_1_2_io_outs_down[32] ;
 wire \_ces_1_2_io_outs_down[33] ;
 wire \_ces_1_2_io_outs_down[34] ;
 wire \_ces_1_2_io_outs_down[35] ;
 wire \_ces_1_2_io_outs_down[36] ;
 wire \_ces_1_2_io_outs_down[37] ;
 wire \_ces_1_2_io_outs_down[38] ;
 wire \_ces_1_2_io_outs_down[39] ;
 wire \_ces_1_2_io_outs_down[3] ;
 wire \_ces_1_2_io_outs_down[40] ;
 wire \_ces_1_2_io_outs_down[41] ;
 wire \_ces_1_2_io_outs_down[42] ;
 wire \_ces_1_2_io_outs_down[43] ;
 wire \_ces_1_2_io_outs_down[44] ;
 wire \_ces_1_2_io_outs_down[45] ;
 wire \_ces_1_2_io_outs_down[46] ;
 wire \_ces_1_2_io_outs_down[47] ;
 wire \_ces_1_2_io_outs_down[48] ;
 wire \_ces_1_2_io_outs_down[49] ;
 wire \_ces_1_2_io_outs_down[4] ;
 wire \_ces_1_2_io_outs_down[50] ;
 wire \_ces_1_2_io_outs_down[51] ;
 wire \_ces_1_2_io_outs_down[52] ;
 wire \_ces_1_2_io_outs_down[53] ;
 wire \_ces_1_2_io_outs_down[54] ;
 wire \_ces_1_2_io_outs_down[55] ;
 wire \_ces_1_2_io_outs_down[56] ;
 wire \_ces_1_2_io_outs_down[57] ;
 wire \_ces_1_2_io_outs_down[58] ;
 wire \_ces_1_2_io_outs_down[59] ;
 wire \_ces_1_2_io_outs_down[5] ;
 wire \_ces_1_2_io_outs_down[60] ;
 wire \_ces_1_2_io_outs_down[61] ;
 wire \_ces_1_2_io_outs_down[62] ;
 wire \_ces_1_2_io_outs_down[63] ;
 wire \_ces_1_2_io_outs_down[6] ;
 wire \_ces_1_2_io_outs_down[7] ;
 wire \_ces_1_2_io_outs_down[8] ;
 wire \_ces_1_2_io_outs_down[9] ;
 wire \_ces_1_2_io_outs_left[0] ;
 wire \_ces_1_2_io_outs_left[10] ;
 wire \_ces_1_2_io_outs_left[11] ;
 wire \_ces_1_2_io_outs_left[12] ;
 wire \_ces_1_2_io_outs_left[13] ;
 wire \_ces_1_2_io_outs_left[14] ;
 wire \_ces_1_2_io_outs_left[15] ;
 wire \_ces_1_2_io_outs_left[16] ;
 wire \_ces_1_2_io_outs_left[17] ;
 wire \_ces_1_2_io_outs_left[18] ;
 wire \_ces_1_2_io_outs_left[19] ;
 wire \_ces_1_2_io_outs_left[1] ;
 wire \_ces_1_2_io_outs_left[20] ;
 wire \_ces_1_2_io_outs_left[21] ;
 wire \_ces_1_2_io_outs_left[22] ;
 wire \_ces_1_2_io_outs_left[23] ;
 wire \_ces_1_2_io_outs_left[24] ;
 wire \_ces_1_2_io_outs_left[25] ;
 wire \_ces_1_2_io_outs_left[26] ;
 wire \_ces_1_2_io_outs_left[27] ;
 wire \_ces_1_2_io_outs_left[28] ;
 wire \_ces_1_2_io_outs_left[29] ;
 wire \_ces_1_2_io_outs_left[2] ;
 wire \_ces_1_2_io_outs_left[30] ;
 wire \_ces_1_2_io_outs_left[31] ;
 wire \_ces_1_2_io_outs_left[32] ;
 wire \_ces_1_2_io_outs_left[33] ;
 wire \_ces_1_2_io_outs_left[34] ;
 wire \_ces_1_2_io_outs_left[35] ;
 wire \_ces_1_2_io_outs_left[36] ;
 wire \_ces_1_2_io_outs_left[37] ;
 wire \_ces_1_2_io_outs_left[38] ;
 wire \_ces_1_2_io_outs_left[39] ;
 wire \_ces_1_2_io_outs_left[3] ;
 wire \_ces_1_2_io_outs_left[40] ;
 wire \_ces_1_2_io_outs_left[41] ;
 wire \_ces_1_2_io_outs_left[42] ;
 wire \_ces_1_2_io_outs_left[43] ;
 wire \_ces_1_2_io_outs_left[44] ;
 wire \_ces_1_2_io_outs_left[45] ;
 wire \_ces_1_2_io_outs_left[46] ;
 wire \_ces_1_2_io_outs_left[47] ;
 wire \_ces_1_2_io_outs_left[48] ;
 wire \_ces_1_2_io_outs_left[49] ;
 wire \_ces_1_2_io_outs_left[4] ;
 wire \_ces_1_2_io_outs_left[50] ;
 wire \_ces_1_2_io_outs_left[51] ;
 wire \_ces_1_2_io_outs_left[52] ;
 wire \_ces_1_2_io_outs_left[53] ;
 wire \_ces_1_2_io_outs_left[54] ;
 wire \_ces_1_2_io_outs_left[55] ;
 wire \_ces_1_2_io_outs_left[56] ;
 wire \_ces_1_2_io_outs_left[57] ;
 wire \_ces_1_2_io_outs_left[58] ;
 wire \_ces_1_2_io_outs_left[59] ;
 wire \_ces_1_2_io_outs_left[5] ;
 wire \_ces_1_2_io_outs_left[60] ;
 wire \_ces_1_2_io_outs_left[61] ;
 wire \_ces_1_2_io_outs_left[62] ;
 wire \_ces_1_2_io_outs_left[63] ;
 wire \_ces_1_2_io_outs_left[6] ;
 wire \_ces_1_2_io_outs_left[7] ;
 wire \_ces_1_2_io_outs_left[8] ;
 wire \_ces_1_2_io_outs_left[9] ;
 wire \_ces_1_2_io_outs_right[0] ;
 wire \_ces_1_2_io_outs_right[10] ;
 wire \_ces_1_2_io_outs_right[11] ;
 wire \_ces_1_2_io_outs_right[12] ;
 wire \_ces_1_2_io_outs_right[13] ;
 wire \_ces_1_2_io_outs_right[14] ;
 wire \_ces_1_2_io_outs_right[15] ;
 wire \_ces_1_2_io_outs_right[16] ;
 wire \_ces_1_2_io_outs_right[17] ;
 wire \_ces_1_2_io_outs_right[18] ;
 wire \_ces_1_2_io_outs_right[19] ;
 wire \_ces_1_2_io_outs_right[1] ;
 wire \_ces_1_2_io_outs_right[20] ;
 wire \_ces_1_2_io_outs_right[21] ;
 wire \_ces_1_2_io_outs_right[22] ;
 wire \_ces_1_2_io_outs_right[23] ;
 wire \_ces_1_2_io_outs_right[24] ;
 wire \_ces_1_2_io_outs_right[25] ;
 wire \_ces_1_2_io_outs_right[26] ;
 wire \_ces_1_2_io_outs_right[27] ;
 wire \_ces_1_2_io_outs_right[28] ;
 wire \_ces_1_2_io_outs_right[29] ;
 wire \_ces_1_2_io_outs_right[2] ;
 wire \_ces_1_2_io_outs_right[30] ;
 wire \_ces_1_2_io_outs_right[31] ;
 wire \_ces_1_2_io_outs_right[32] ;
 wire \_ces_1_2_io_outs_right[33] ;
 wire \_ces_1_2_io_outs_right[34] ;
 wire \_ces_1_2_io_outs_right[35] ;
 wire \_ces_1_2_io_outs_right[36] ;
 wire \_ces_1_2_io_outs_right[37] ;
 wire \_ces_1_2_io_outs_right[38] ;
 wire \_ces_1_2_io_outs_right[39] ;
 wire \_ces_1_2_io_outs_right[3] ;
 wire \_ces_1_2_io_outs_right[40] ;
 wire \_ces_1_2_io_outs_right[41] ;
 wire \_ces_1_2_io_outs_right[42] ;
 wire \_ces_1_2_io_outs_right[43] ;
 wire \_ces_1_2_io_outs_right[44] ;
 wire \_ces_1_2_io_outs_right[45] ;
 wire \_ces_1_2_io_outs_right[46] ;
 wire \_ces_1_2_io_outs_right[47] ;
 wire \_ces_1_2_io_outs_right[48] ;
 wire \_ces_1_2_io_outs_right[49] ;
 wire \_ces_1_2_io_outs_right[4] ;
 wire \_ces_1_2_io_outs_right[50] ;
 wire \_ces_1_2_io_outs_right[51] ;
 wire \_ces_1_2_io_outs_right[52] ;
 wire \_ces_1_2_io_outs_right[53] ;
 wire \_ces_1_2_io_outs_right[54] ;
 wire \_ces_1_2_io_outs_right[55] ;
 wire \_ces_1_2_io_outs_right[56] ;
 wire \_ces_1_2_io_outs_right[57] ;
 wire \_ces_1_2_io_outs_right[58] ;
 wire \_ces_1_2_io_outs_right[59] ;
 wire \_ces_1_2_io_outs_right[5] ;
 wire \_ces_1_2_io_outs_right[60] ;
 wire \_ces_1_2_io_outs_right[61] ;
 wire \_ces_1_2_io_outs_right[62] ;
 wire \_ces_1_2_io_outs_right[63] ;
 wire \_ces_1_2_io_outs_right[6] ;
 wire \_ces_1_2_io_outs_right[7] ;
 wire \_ces_1_2_io_outs_right[8] ;
 wire \_ces_1_2_io_outs_right[9] ;
 wire \_ces_1_2_io_outs_up[0] ;
 wire \_ces_1_2_io_outs_up[10] ;
 wire \_ces_1_2_io_outs_up[11] ;
 wire \_ces_1_2_io_outs_up[12] ;
 wire \_ces_1_2_io_outs_up[13] ;
 wire \_ces_1_2_io_outs_up[14] ;
 wire \_ces_1_2_io_outs_up[15] ;
 wire \_ces_1_2_io_outs_up[16] ;
 wire \_ces_1_2_io_outs_up[17] ;
 wire \_ces_1_2_io_outs_up[18] ;
 wire \_ces_1_2_io_outs_up[19] ;
 wire \_ces_1_2_io_outs_up[1] ;
 wire \_ces_1_2_io_outs_up[20] ;
 wire \_ces_1_2_io_outs_up[21] ;
 wire \_ces_1_2_io_outs_up[22] ;
 wire \_ces_1_2_io_outs_up[23] ;
 wire \_ces_1_2_io_outs_up[24] ;
 wire \_ces_1_2_io_outs_up[25] ;
 wire \_ces_1_2_io_outs_up[26] ;
 wire \_ces_1_2_io_outs_up[27] ;
 wire \_ces_1_2_io_outs_up[28] ;
 wire \_ces_1_2_io_outs_up[29] ;
 wire \_ces_1_2_io_outs_up[2] ;
 wire \_ces_1_2_io_outs_up[30] ;
 wire \_ces_1_2_io_outs_up[31] ;
 wire \_ces_1_2_io_outs_up[32] ;
 wire \_ces_1_2_io_outs_up[33] ;
 wire \_ces_1_2_io_outs_up[34] ;
 wire \_ces_1_2_io_outs_up[35] ;
 wire \_ces_1_2_io_outs_up[36] ;
 wire \_ces_1_2_io_outs_up[37] ;
 wire \_ces_1_2_io_outs_up[38] ;
 wire \_ces_1_2_io_outs_up[39] ;
 wire \_ces_1_2_io_outs_up[3] ;
 wire \_ces_1_2_io_outs_up[40] ;
 wire \_ces_1_2_io_outs_up[41] ;
 wire \_ces_1_2_io_outs_up[42] ;
 wire \_ces_1_2_io_outs_up[43] ;
 wire \_ces_1_2_io_outs_up[44] ;
 wire \_ces_1_2_io_outs_up[45] ;
 wire \_ces_1_2_io_outs_up[46] ;
 wire \_ces_1_2_io_outs_up[47] ;
 wire \_ces_1_2_io_outs_up[48] ;
 wire \_ces_1_2_io_outs_up[49] ;
 wire \_ces_1_2_io_outs_up[4] ;
 wire \_ces_1_2_io_outs_up[50] ;
 wire \_ces_1_2_io_outs_up[51] ;
 wire \_ces_1_2_io_outs_up[52] ;
 wire \_ces_1_2_io_outs_up[53] ;
 wire \_ces_1_2_io_outs_up[54] ;
 wire \_ces_1_2_io_outs_up[55] ;
 wire \_ces_1_2_io_outs_up[56] ;
 wire \_ces_1_2_io_outs_up[57] ;
 wire \_ces_1_2_io_outs_up[58] ;
 wire \_ces_1_2_io_outs_up[59] ;
 wire \_ces_1_2_io_outs_up[5] ;
 wire \_ces_1_2_io_outs_up[60] ;
 wire \_ces_1_2_io_outs_up[61] ;
 wire \_ces_1_2_io_outs_up[62] ;
 wire \_ces_1_2_io_outs_up[63] ;
 wire \_ces_1_2_io_outs_up[6] ;
 wire \_ces_1_2_io_outs_up[7] ;
 wire \_ces_1_2_io_outs_up[8] ;
 wire \_ces_1_2_io_outs_up[9] ;
 wire _ces_1_3_io_lsbOuts_0;
 wire _ces_1_3_io_lsbOuts_1;
 wire _ces_1_3_io_lsbOuts_2;
 wire _ces_1_3_io_lsbOuts_3;
 wire \_ces_1_3_io_outs_down[0] ;
 wire \_ces_1_3_io_outs_down[10] ;
 wire \_ces_1_3_io_outs_down[11] ;
 wire \_ces_1_3_io_outs_down[12] ;
 wire \_ces_1_3_io_outs_down[13] ;
 wire \_ces_1_3_io_outs_down[14] ;
 wire \_ces_1_3_io_outs_down[15] ;
 wire \_ces_1_3_io_outs_down[16] ;
 wire \_ces_1_3_io_outs_down[17] ;
 wire \_ces_1_3_io_outs_down[18] ;
 wire \_ces_1_3_io_outs_down[19] ;
 wire \_ces_1_3_io_outs_down[1] ;
 wire \_ces_1_3_io_outs_down[20] ;
 wire \_ces_1_3_io_outs_down[21] ;
 wire \_ces_1_3_io_outs_down[22] ;
 wire \_ces_1_3_io_outs_down[23] ;
 wire \_ces_1_3_io_outs_down[24] ;
 wire \_ces_1_3_io_outs_down[25] ;
 wire \_ces_1_3_io_outs_down[26] ;
 wire \_ces_1_3_io_outs_down[27] ;
 wire \_ces_1_3_io_outs_down[28] ;
 wire \_ces_1_3_io_outs_down[29] ;
 wire \_ces_1_3_io_outs_down[2] ;
 wire \_ces_1_3_io_outs_down[30] ;
 wire \_ces_1_3_io_outs_down[31] ;
 wire \_ces_1_3_io_outs_down[32] ;
 wire \_ces_1_3_io_outs_down[33] ;
 wire \_ces_1_3_io_outs_down[34] ;
 wire \_ces_1_3_io_outs_down[35] ;
 wire \_ces_1_3_io_outs_down[36] ;
 wire \_ces_1_3_io_outs_down[37] ;
 wire \_ces_1_3_io_outs_down[38] ;
 wire \_ces_1_3_io_outs_down[39] ;
 wire \_ces_1_3_io_outs_down[3] ;
 wire \_ces_1_3_io_outs_down[40] ;
 wire \_ces_1_3_io_outs_down[41] ;
 wire \_ces_1_3_io_outs_down[42] ;
 wire \_ces_1_3_io_outs_down[43] ;
 wire \_ces_1_3_io_outs_down[44] ;
 wire \_ces_1_3_io_outs_down[45] ;
 wire \_ces_1_3_io_outs_down[46] ;
 wire \_ces_1_3_io_outs_down[47] ;
 wire \_ces_1_3_io_outs_down[48] ;
 wire \_ces_1_3_io_outs_down[49] ;
 wire \_ces_1_3_io_outs_down[4] ;
 wire \_ces_1_3_io_outs_down[50] ;
 wire \_ces_1_3_io_outs_down[51] ;
 wire \_ces_1_3_io_outs_down[52] ;
 wire \_ces_1_3_io_outs_down[53] ;
 wire \_ces_1_3_io_outs_down[54] ;
 wire \_ces_1_3_io_outs_down[55] ;
 wire \_ces_1_3_io_outs_down[56] ;
 wire \_ces_1_3_io_outs_down[57] ;
 wire \_ces_1_3_io_outs_down[58] ;
 wire \_ces_1_3_io_outs_down[59] ;
 wire \_ces_1_3_io_outs_down[5] ;
 wire \_ces_1_3_io_outs_down[60] ;
 wire \_ces_1_3_io_outs_down[61] ;
 wire \_ces_1_3_io_outs_down[62] ;
 wire \_ces_1_3_io_outs_down[63] ;
 wire \_ces_1_3_io_outs_down[6] ;
 wire \_ces_1_3_io_outs_down[7] ;
 wire \_ces_1_3_io_outs_down[8] ;
 wire \_ces_1_3_io_outs_down[9] ;
 wire \_ces_1_3_io_outs_left[0] ;
 wire \_ces_1_3_io_outs_left[10] ;
 wire \_ces_1_3_io_outs_left[11] ;
 wire \_ces_1_3_io_outs_left[12] ;
 wire \_ces_1_3_io_outs_left[13] ;
 wire \_ces_1_3_io_outs_left[14] ;
 wire \_ces_1_3_io_outs_left[15] ;
 wire \_ces_1_3_io_outs_left[16] ;
 wire \_ces_1_3_io_outs_left[17] ;
 wire \_ces_1_3_io_outs_left[18] ;
 wire \_ces_1_3_io_outs_left[19] ;
 wire \_ces_1_3_io_outs_left[1] ;
 wire \_ces_1_3_io_outs_left[20] ;
 wire \_ces_1_3_io_outs_left[21] ;
 wire \_ces_1_3_io_outs_left[22] ;
 wire \_ces_1_3_io_outs_left[23] ;
 wire \_ces_1_3_io_outs_left[24] ;
 wire \_ces_1_3_io_outs_left[25] ;
 wire \_ces_1_3_io_outs_left[26] ;
 wire \_ces_1_3_io_outs_left[27] ;
 wire \_ces_1_3_io_outs_left[28] ;
 wire \_ces_1_3_io_outs_left[29] ;
 wire \_ces_1_3_io_outs_left[2] ;
 wire \_ces_1_3_io_outs_left[30] ;
 wire \_ces_1_3_io_outs_left[31] ;
 wire \_ces_1_3_io_outs_left[32] ;
 wire \_ces_1_3_io_outs_left[33] ;
 wire \_ces_1_3_io_outs_left[34] ;
 wire \_ces_1_3_io_outs_left[35] ;
 wire \_ces_1_3_io_outs_left[36] ;
 wire \_ces_1_3_io_outs_left[37] ;
 wire \_ces_1_3_io_outs_left[38] ;
 wire \_ces_1_3_io_outs_left[39] ;
 wire \_ces_1_3_io_outs_left[3] ;
 wire \_ces_1_3_io_outs_left[40] ;
 wire \_ces_1_3_io_outs_left[41] ;
 wire \_ces_1_3_io_outs_left[42] ;
 wire \_ces_1_3_io_outs_left[43] ;
 wire \_ces_1_3_io_outs_left[44] ;
 wire \_ces_1_3_io_outs_left[45] ;
 wire \_ces_1_3_io_outs_left[46] ;
 wire \_ces_1_3_io_outs_left[47] ;
 wire \_ces_1_3_io_outs_left[48] ;
 wire \_ces_1_3_io_outs_left[49] ;
 wire \_ces_1_3_io_outs_left[4] ;
 wire \_ces_1_3_io_outs_left[50] ;
 wire \_ces_1_3_io_outs_left[51] ;
 wire \_ces_1_3_io_outs_left[52] ;
 wire \_ces_1_3_io_outs_left[53] ;
 wire \_ces_1_3_io_outs_left[54] ;
 wire \_ces_1_3_io_outs_left[55] ;
 wire \_ces_1_3_io_outs_left[56] ;
 wire \_ces_1_3_io_outs_left[57] ;
 wire \_ces_1_3_io_outs_left[58] ;
 wire \_ces_1_3_io_outs_left[59] ;
 wire \_ces_1_3_io_outs_left[5] ;
 wire \_ces_1_3_io_outs_left[60] ;
 wire \_ces_1_3_io_outs_left[61] ;
 wire \_ces_1_3_io_outs_left[62] ;
 wire \_ces_1_3_io_outs_left[63] ;
 wire \_ces_1_3_io_outs_left[6] ;
 wire \_ces_1_3_io_outs_left[7] ;
 wire \_ces_1_3_io_outs_left[8] ;
 wire \_ces_1_3_io_outs_left[9] ;
 wire \_ces_1_3_io_outs_up[0] ;
 wire \_ces_1_3_io_outs_up[10] ;
 wire \_ces_1_3_io_outs_up[11] ;
 wire \_ces_1_3_io_outs_up[12] ;
 wire \_ces_1_3_io_outs_up[13] ;
 wire \_ces_1_3_io_outs_up[14] ;
 wire \_ces_1_3_io_outs_up[15] ;
 wire \_ces_1_3_io_outs_up[16] ;
 wire \_ces_1_3_io_outs_up[17] ;
 wire \_ces_1_3_io_outs_up[18] ;
 wire \_ces_1_3_io_outs_up[19] ;
 wire \_ces_1_3_io_outs_up[1] ;
 wire \_ces_1_3_io_outs_up[20] ;
 wire \_ces_1_3_io_outs_up[21] ;
 wire \_ces_1_3_io_outs_up[22] ;
 wire \_ces_1_3_io_outs_up[23] ;
 wire \_ces_1_3_io_outs_up[24] ;
 wire \_ces_1_3_io_outs_up[25] ;
 wire \_ces_1_3_io_outs_up[26] ;
 wire \_ces_1_3_io_outs_up[27] ;
 wire \_ces_1_3_io_outs_up[28] ;
 wire \_ces_1_3_io_outs_up[29] ;
 wire \_ces_1_3_io_outs_up[2] ;
 wire \_ces_1_3_io_outs_up[30] ;
 wire \_ces_1_3_io_outs_up[31] ;
 wire \_ces_1_3_io_outs_up[32] ;
 wire \_ces_1_3_io_outs_up[33] ;
 wire \_ces_1_3_io_outs_up[34] ;
 wire \_ces_1_3_io_outs_up[35] ;
 wire \_ces_1_3_io_outs_up[36] ;
 wire \_ces_1_3_io_outs_up[37] ;
 wire \_ces_1_3_io_outs_up[38] ;
 wire \_ces_1_3_io_outs_up[39] ;
 wire \_ces_1_3_io_outs_up[3] ;
 wire \_ces_1_3_io_outs_up[40] ;
 wire \_ces_1_3_io_outs_up[41] ;
 wire \_ces_1_3_io_outs_up[42] ;
 wire \_ces_1_3_io_outs_up[43] ;
 wire \_ces_1_3_io_outs_up[44] ;
 wire \_ces_1_3_io_outs_up[45] ;
 wire \_ces_1_3_io_outs_up[46] ;
 wire \_ces_1_3_io_outs_up[47] ;
 wire \_ces_1_3_io_outs_up[48] ;
 wire \_ces_1_3_io_outs_up[49] ;
 wire \_ces_1_3_io_outs_up[4] ;
 wire \_ces_1_3_io_outs_up[50] ;
 wire \_ces_1_3_io_outs_up[51] ;
 wire \_ces_1_3_io_outs_up[52] ;
 wire \_ces_1_3_io_outs_up[53] ;
 wire \_ces_1_3_io_outs_up[54] ;
 wire \_ces_1_3_io_outs_up[55] ;
 wire \_ces_1_3_io_outs_up[56] ;
 wire \_ces_1_3_io_outs_up[57] ;
 wire \_ces_1_3_io_outs_up[58] ;
 wire \_ces_1_3_io_outs_up[59] ;
 wire \_ces_1_3_io_outs_up[5] ;
 wire \_ces_1_3_io_outs_up[60] ;
 wire \_ces_1_3_io_outs_up[61] ;
 wire \_ces_1_3_io_outs_up[62] ;
 wire \_ces_1_3_io_outs_up[63] ;
 wire \_ces_1_3_io_outs_up[6] ;
 wire \_ces_1_3_io_outs_up[7] ;
 wire \_ces_1_3_io_outs_up[8] ;
 wire \_ces_1_3_io_outs_up[9] ;
 wire _ces_2_0_io_lsbOuts_1;
 wire _ces_2_0_io_lsbOuts_2;
 wire _ces_2_0_io_lsbOuts_3;
 wire \_ces_2_0_io_outs_down[0] ;
 wire \_ces_2_0_io_outs_down[10] ;
 wire \_ces_2_0_io_outs_down[11] ;
 wire \_ces_2_0_io_outs_down[12] ;
 wire \_ces_2_0_io_outs_down[13] ;
 wire \_ces_2_0_io_outs_down[14] ;
 wire \_ces_2_0_io_outs_down[15] ;
 wire \_ces_2_0_io_outs_down[16] ;
 wire \_ces_2_0_io_outs_down[17] ;
 wire \_ces_2_0_io_outs_down[18] ;
 wire \_ces_2_0_io_outs_down[19] ;
 wire \_ces_2_0_io_outs_down[1] ;
 wire \_ces_2_0_io_outs_down[20] ;
 wire \_ces_2_0_io_outs_down[21] ;
 wire \_ces_2_0_io_outs_down[22] ;
 wire \_ces_2_0_io_outs_down[23] ;
 wire \_ces_2_0_io_outs_down[24] ;
 wire \_ces_2_0_io_outs_down[25] ;
 wire \_ces_2_0_io_outs_down[26] ;
 wire \_ces_2_0_io_outs_down[27] ;
 wire \_ces_2_0_io_outs_down[28] ;
 wire \_ces_2_0_io_outs_down[29] ;
 wire \_ces_2_0_io_outs_down[2] ;
 wire \_ces_2_0_io_outs_down[30] ;
 wire \_ces_2_0_io_outs_down[31] ;
 wire \_ces_2_0_io_outs_down[32] ;
 wire \_ces_2_0_io_outs_down[33] ;
 wire \_ces_2_0_io_outs_down[34] ;
 wire \_ces_2_0_io_outs_down[35] ;
 wire \_ces_2_0_io_outs_down[36] ;
 wire \_ces_2_0_io_outs_down[37] ;
 wire \_ces_2_0_io_outs_down[38] ;
 wire \_ces_2_0_io_outs_down[39] ;
 wire \_ces_2_0_io_outs_down[3] ;
 wire \_ces_2_0_io_outs_down[40] ;
 wire \_ces_2_0_io_outs_down[41] ;
 wire \_ces_2_0_io_outs_down[42] ;
 wire \_ces_2_0_io_outs_down[43] ;
 wire \_ces_2_0_io_outs_down[44] ;
 wire \_ces_2_0_io_outs_down[45] ;
 wire \_ces_2_0_io_outs_down[46] ;
 wire \_ces_2_0_io_outs_down[47] ;
 wire \_ces_2_0_io_outs_down[48] ;
 wire \_ces_2_0_io_outs_down[49] ;
 wire \_ces_2_0_io_outs_down[4] ;
 wire \_ces_2_0_io_outs_down[50] ;
 wire \_ces_2_0_io_outs_down[51] ;
 wire \_ces_2_0_io_outs_down[52] ;
 wire \_ces_2_0_io_outs_down[53] ;
 wire \_ces_2_0_io_outs_down[54] ;
 wire \_ces_2_0_io_outs_down[55] ;
 wire \_ces_2_0_io_outs_down[56] ;
 wire \_ces_2_0_io_outs_down[57] ;
 wire \_ces_2_0_io_outs_down[58] ;
 wire \_ces_2_0_io_outs_down[59] ;
 wire \_ces_2_0_io_outs_down[5] ;
 wire \_ces_2_0_io_outs_down[60] ;
 wire \_ces_2_0_io_outs_down[61] ;
 wire \_ces_2_0_io_outs_down[62] ;
 wire \_ces_2_0_io_outs_down[63] ;
 wire \_ces_2_0_io_outs_down[6] ;
 wire \_ces_2_0_io_outs_down[7] ;
 wire \_ces_2_0_io_outs_down[8] ;
 wire \_ces_2_0_io_outs_down[9] ;
 wire \_ces_2_0_io_outs_right[0] ;
 wire \_ces_2_0_io_outs_right[10] ;
 wire \_ces_2_0_io_outs_right[11] ;
 wire \_ces_2_0_io_outs_right[12] ;
 wire \_ces_2_0_io_outs_right[13] ;
 wire \_ces_2_0_io_outs_right[14] ;
 wire \_ces_2_0_io_outs_right[15] ;
 wire \_ces_2_0_io_outs_right[16] ;
 wire \_ces_2_0_io_outs_right[17] ;
 wire \_ces_2_0_io_outs_right[18] ;
 wire \_ces_2_0_io_outs_right[19] ;
 wire \_ces_2_0_io_outs_right[1] ;
 wire \_ces_2_0_io_outs_right[20] ;
 wire \_ces_2_0_io_outs_right[21] ;
 wire \_ces_2_0_io_outs_right[22] ;
 wire \_ces_2_0_io_outs_right[23] ;
 wire \_ces_2_0_io_outs_right[24] ;
 wire \_ces_2_0_io_outs_right[25] ;
 wire \_ces_2_0_io_outs_right[26] ;
 wire \_ces_2_0_io_outs_right[27] ;
 wire \_ces_2_0_io_outs_right[28] ;
 wire \_ces_2_0_io_outs_right[29] ;
 wire \_ces_2_0_io_outs_right[2] ;
 wire \_ces_2_0_io_outs_right[30] ;
 wire \_ces_2_0_io_outs_right[31] ;
 wire \_ces_2_0_io_outs_right[32] ;
 wire \_ces_2_0_io_outs_right[33] ;
 wire \_ces_2_0_io_outs_right[34] ;
 wire \_ces_2_0_io_outs_right[35] ;
 wire \_ces_2_0_io_outs_right[36] ;
 wire \_ces_2_0_io_outs_right[37] ;
 wire \_ces_2_0_io_outs_right[38] ;
 wire \_ces_2_0_io_outs_right[39] ;
 wire \_ces_2_0_io_outs_right[3] ;
 wire \_ces_2_0_io_outs_right[40] ;
 wire \_ces_2_0_io_outs_right[41] ;
 wire \_ces_2_0_io_outs_right[42] ;
 wire \_ces_2_0_io_outs_right[43] ;
 wire \_ces_2_0_io_outs_right[44] ;
 wire \_ces_2_0_io_outs_right[45] ;
 wire \_ces_2_0_io_outs_right[46] ;
 wire \_ces_2_0_io_outs_right[47] ;
 wire \_ces_2_0_io_outs_right[48] ;
 wire \_ces_2_0_io_outs_right[49] ;
 wire \_ces_2_0_io_outs_right[4] ;
 wire \_ces_2_0_io_outs_right[50] ;
 wire \_ces_2_0_io_outs_right[51] ;
 wire \_ces_2_0_io_outs_right[52] ;
 wire \_ces_2_0_io_outs_right[53] ;
 wire \_ces_2_0_io_outs_right[54] ;
 wire \_ces_2_0_io_outs_right[55] ;
 wire \_ces_2_0_io_outs_right[56] ;
 wire \_ces_2_0_io_outs_right[57] ;
 wire \_ces_2_0_io_outs_right[58] ;
 wire \_ces_2_0_io_outs_right[59] ;
 wire \_ces_2_0_io_outs_right[5] ;
 wire \_ces_2_0_io_outs_right[60] ;
 wire \_ces_2_0_io_outs_right[61] ;
 wire \_ces_2_0_io_outs_right[62] ;
 wire \_ces_2_0_io_outs_right[63] ;
 wire \_ces_2_0_io_outs_right[6] ;
 wire \_ces_2_0_io_outs_right[7] ;
 wire \_ces_2_0_io_outs_right[8] ;
 wire \_ces_2_0_io_outs_right[9] ;
 wire \_ces_2_0_io_outs_up[0] ;
 wire \_ces_2_0_io_outs_up[10] ;
 wire \_ces_2_0_io_outs_up[11] ;
 wire \_ces_2_0_io_outs_up[12] ;
 wire \_ces_2_0_io_outs_up[13] ;
 wire \_ces_2_0_io_outs_up[14] ;
 wire \_ces_2_0_io_outs_up[15] ;
 wire \_ces_2_0_io_outs_up[16] ;
 wire \_ces_2_0_io_outs_up[17] ;
 wire \_ces_2_0_io_outs_up[18] ;
 wire \_ces_2_0_io_outs_up[19] ;
 wire \_ces_2_0_io_outs_up[1] ;
 wire \_ces_2_0_io_outs_up[20] ;
 wire \_ces_2_0_io_outs_up[21] ;
 wire \_ces_2_0_io_outs_up[22] ;
 wire \_ces_2_0_io_outs_up[23] ;
 wire \_ces_2_0_io_outs_up[24] ;
 wire \_ces_2_0_io_outs_up[25] ;
 wire \_ces_2_0_io_outs_up[26] ;
 wire \_ces_2_0_io_outs_up[27] ;
 wire \_ces_2_0_io_outs_up[28] ;
 wire \_ces_2_0_io_outs_up[29] ;
 wire \_ces_2_0_io_outs_up[2] ;
 wire \_ces_2_0_io_outs_up[30] ;
 wire \_ces_2_0_io_outs_up[31] ;
 wire \_ces_2_0_io_outs_up[32] ;
 wire \_ces_2_0_io_outs_up[33] ;
 wire \_ces_2_0_io_outs_up[34] ;
 wire \_ces_2_0_io_outs_up[35] ;
 wire \_ces_2_0_io_outs_up[36] ;
 wire \_ces_2_0_io_outs_up[37] ;
 wire \_ces_2_0_io_outs_up[38] ;
 wire \_ces_2_0_io_outs_up[39] ;
 wire \_ces_2_0_io_outs_up[3] ;
 wire \_ces_2_0_io_outs_up[40] ;
 wire \_ces_2_0_io_outs_up[41] ;
 wire \_ces_2_0_io_outs_up[42] ;
 wire \_ces_2_0_io_outs_up[43] ;
 wire \_ces_2_0_io_outs_up[44] ;
 wire \_ces_2_0_io_outs_up[45] ;
 wire \_ces_2_0_io_outs_up[46] ;
 wire \_ces_2_0_io_outs_up[47] ;
 wire \_ces_2_0_io_outs_up[48] ;
 wire \_ces_2_0_io_outs_up[49] ;
 wire \_ces_2_0_io_outs_up[4] ;
 wire \_ces_2_0_io_outs_up[50] ;
 wire \_ces_2_0_io_outs_up[51] ;
 wire \_ces_2_0_io_outs_up[52] ;
 wire \_ces_2_0_io_outs_up[53] ;
 wire \_ces_2_0_io_outs_up[54] ;
 wire \_ces_2_0_io_outs_up[55] ;
 wire \_ces_2_0_io_outs_up[56] ;
 wire \_ces_2_0_io_outs_up[57] ;
 wire \_ces_2_0_io_outs_up[58] ;
 wire \_ces_2_0_io_outs_up[59] ;
 wire \_ces_2_0_io_outs_up[5] ;
 wire \_ces_2_0_io_outs_up[60] ;
 wire \_ces_2_0_io_outs_up[61] ;
 wire \_ces_2_0_io_outs_up[62] ;
 wire \_ces_2_0_io_outs_up[63] ;
 wire \_ces_2_0_io_outs_up[6] ;
 wire \_ces_2_0_io_outs_up[7] ;
 wire \_ces_2_0_io_outs_up[8] ;
 wire \_ces_2_0_io_outs_up[9] ;
 wire _ces_2_1_io_lsbOuts_1;
 wire _ces_2_1_io_lsbOuts_2;
 wire _ces_2_1_io_lsbOuts_3;
 wire \_ces_2_1_io_outs_down[0] ;
 wire \_ces_2_1_io_outs_down[10] ;
 wire \_ces_2_1_io_outs_down[11] ;
 wire \_ces_2_1_io_outs_down[12] ;
 wire \_ces_2_1_io_outs_down[13] ;
 wire \_ces_2_1_io_outs_down[14] ;
 wire \_ces_2_1_io_outs_down[15] ;
 wire \_ces_2_1_io_outs_down[16] ;
 wire \_ces_2_1_io_outs_down[17] ;
 wire \_ces_2_1_io_outs_down[18] ;
 wire \_ces_2_1_io_outs_down[19] ;
 wire \_ces_2_1_io_outs_down[1] ;
 wire \_ces_2_1_io_outs_down[20] ;
 wire \_ces_2_1_io_outs_down[21] ;
 wire \_ces_2_1_io_outs_down[22] ;
 wire \_ces_2_1_io_outs_down[23] ;
 wire \_ces_2_1_io_outs_down[24] ;
 wire \_ces_2_1_io_outs_down[25] ;
 wire \_ces_2_1_io_outs_down[26] ;
 wire \_ces_2_1_io_outs_down[27] ;
 wire \_ces_2_1_io_outs_down[28] ;
 wire \_ces_2_1_io_outs_down[29] ;
 wire \_ces_2_1_io_outs_down[2] ;
 wire \_ces_2_1_io_outs_down[30] ;
 wire \_ces_2_1_io_outs_down[31] ;
 wire \_ces_2_1_io_outs_down[32] ;
 wire \_ces_2_1_io_outs_down[33] ;
 wire \_ces_2_1_io_outs_down[34] ;
 wire \_ces_2_1_io_outs_down[35] ;
 wire \_ces_2_1_io_outs_down[36] ;
 wire \_ces_2_1_io_outs_down[37] ;
 wire \_ces_2_1_io_outs_down[38] ;
 wire \_ces_2_1_io_outs_down[39] ;
 wire \_ces_2_1_io_outs_down[3] ;
 wire \_ces_2_1_io_outs_down[40] ;
 wire \_ces_2_1_io_outs_down[41] ;
 wire \_ces_2_1_io_outs_down[42] ;
 wire \_ces_2_1_io_outs_down[43] ;
 wire \_ces_2_1_io_outs_down[44] ;
 wire \_ces_2_1_io_outs_down[45] ;
 wire \_ces_2_1_io_outs_down[46] ;
 wire \_ces_2_1_io_outs_down[47] ;
 wire \_ces_2_1_io_outs_down[48] ;
 wire \_ces_2_1_io_outs_down[49] ;
 wire \_ces_2_1_io_outs_down[4] ;
 wire \_ces_2_1_io_outs_down[50] ;
 wire \_ces_2_1_io_outs_down[51] ;
 wire \_ces_2_1_io_outs_down[52] ;
 wire \_ces_2_1_io_outs_down[53] ;
 wire \_ces_2_1_io_outs_down[54] ;
 wire \_ces_2_1_io_outs_down[55] ;
 wire \_ces_2_1_io_outs_down[56] ;
 wire \_ces_2_1_io_outs_down[57] ;
 wire \_ces_2_1_io_outs_down[58] ;
 wire \_ces_2_1_io_outs_down[59] ;
 wire \_ces_2_1_io_outs_down[5] ;
 wire \_ces_2_1_io_outs_down[60] ;
 wire \_ces_2_1_io_outs_down[61] ;
 wire \_ces_2_1_io_outs_down[62] ;
 wire \_ces_2_1_io_outs_down[63] ;
 wire \_ces_2_1_io_outs_down[6] ;
 wire \_ces_2_1_io_outs_down[7] ;
 wire \_ces_2_1_io_outs_down[8] ;
 wire \_ces_2_1_io_outs_down[9] ;
 wire \_ces_2_1_io_outs_left[0] ;
 wire \_ces_2_1_io_outs_left[10] ;
 wire \_ces_2_1_io_outs_left[11] ;
 wire \_ces_2_1_io_outs_left[12] ;
 wire \_ces_2_1_io_outs_left[13] ;
 wire \_ces_2_1_io_outs_left[14] ;
 wire \_ces_2_1_io_outs_left[15] ;
 wire \_ces_2_1_io_outs_left[16] ;
 wire \_ces_2_1_io_outs_left[17] ;
 wire \_ces_2_1_io_outs_left[18] ;
 wire \_ces_2_1_io_outs_left[19] ;
 wire \_ces_2_1_io_outs_left[1] ;
 wire \_ces_2_1_io_outs_left[20] ;
 wire \_ces_2_1_io_outs_left[21] ;
 wire \_ces_2_1_io_outs_left[22] ;
 wire \_ces_2_1_io_outs_left[23] ;
 wire \_ces_2_1_io_outs_left[24] ;
 wire \_ces_2_1_io_outs_left[25] ;
 wire \_ces_2_1_io_outs_left[26] ;
 wire \_ces_2_1_io_outs_left[27] ;
 wire \_ces_2_1_io_outs_left[28] ;
 wire \_ces_2_1_io_outs_left[29] ;
 wire \_ces_2_1_io_outs_left[2] ;
 wire \_ces_2_1_io_outs_left[30] ;
 wire \_ces_2_1_io_outs_left[31] ;
 wire \_ces_2_1_io_outs_left[32] ;
 wire \_ces_2_1_io_outs_left[33] ;
 wire \_ces_2_1_io_outs_left[34] ;
 wire \_ces_2_1_io_outs_left[35] ;
 wire \_ces_2_1_io_outs_left[36] ;
 wire \_ces_2_1_io_outs_left[37] ;
 wire \_ces_2_1_io_outs_left[38] ;
 wire \_ces_2_1_io_outs_left[39] ;
 wire \_ces_2_1_io_outs_left[3] ;
 wire \_ces_2_1_io_outs_left[40] ;
 wire \_ces_2_1_io_outs_left[41] ;
 wire \_ces_2_1_io_outs_left[42] ;
 wire \_ces_2_1_io_outs_left[43] ;
 wire \_ces_2_1_io_outs_left[44] ;
 wire \_ces_2_1_io_outs_left[45] ;
 wire \_ces_2_1_io_outs_left[46] ;
 wire \_ces_2_1_io_outs_left[47] ;
 wire \_ces_2_1_io_outs_left[48] ;
 wire \_ces_2_1_io_outs_left[49] ;
 wire \_ces_2_1_io_outs_left[4] ;
 wire \_ces_2_1_io_outs_left[50] ;
 wire \_ces_2_1_io_outs_left[51] ;
 wire \_ces_2_1_io_outs_left[52] ;
 wire \_ces_2_1_io_outs_left[53] ;
 wire \_ces_2_1_io_outs_left[54] ;
 wire \_ces_2_1_io_outs_left[55] ;
 wire \_ces_2_1_io_outs_left[56] ;
 wire \_ces_2_1_io_outs_left[57] ;
 wire \_ces_2_1_io_outs_left[58] ;
 wire \_ces_2_1_io_outs_left[59] ;
 wire \_ces_2_1_io_outs_left[5] ;
 wire \_ces_2_1_io_outs_left[60] ;
 wire \_ces_2_1_io_outs_left[61] ;
 wire \_ces_2_1_io_outs_left[62] ;
 wire \_ces_2_1_io_outs_left[63] ;
 wire \_ces_2_1_io_outs_left[6] ;
 wire \_ces_2_1_io_outs_left[7] ;
 wire \_ces_2_1_io_outs_left[8] ;
 wire \_ces_2_1_io_outs_left[9] ;
 wire \_ces_2_1_io_outs_right[0] ;
 wire \_ces_2_1_io_outs_right[10] ;
 wire \_ces_2_1_io_outs_right[11] ;
 wire \_ces_2_1_io_outs_right[12] ;
 wire \_ces_2_1_io_outs_right[13] ;
 wire \_ces_2_1_io_outs_right[14] ;
 wire \_ces_2_1_io_outs_right[15] ;
 wire \_ces_2_1_io_outs_right[16] ;
 wire \_ces_2_1_io_outs_right[17] ;
 wire \_ces_2_1_io_outs_right[18] ;
 wire \_ces_2_1_io_outs_right[19] ;
 wire \_ces_2_1_io_outs_right[1] ;
 wire \_ces_2_1_io_outs_right[20] ;
 wire \_ces_2_1_io_outs_right[21] ;
 wire \_ces_2_1_io_outs_right[22] ;
 wire \_ces_2_1_io_outs_right[23] ;
 wire \_ces_2_1_io_outs_right[24] ;
 wire \_ces_2_1_io_outs_right[25] ;
 wire \_ces_2_1_io_outs_right[26] ;
 wire \_ces_2_1_io_outs_right[27] ;
 wire \_ces_2_1_io_outs_right[28] ;
 wire \_ces_2_1_io_outs_right[29] ;
 wire \_ces_2_1_io_outs_right[2] ;
 wire \_ces_2_1_io_outs_right[30] ;
 wire \_ces_2_1_io_outs_right[31] ;
 wire \_ces_2_1_io_outs_right[32] ;
 wire \_ces_2_1_io_outs_right[33] ;
 wire \_ces_2_1_io_outs_right[34] ;
 wire \_ces_2_1_io_outs_right[35] ;
 wire \_ces_2_1_io_outs_right[36] ;
 wire \_ces_2_1_io_outs_right[37] ;
 wire \_ces_2_1_io_outs_right[38] ;
 wire \_ces_2_1_io_outs_right[39] ;
 wire \_ces_2_1_io_outs_right[3] ;
 wire \_ces_2_1_io_outs_right[40] ;
 wire \_ces_2_1_io_outs_right[41] ;
 wire \_ces_2_1_io_outs_right[42] ;
 wire \_ces_2_1_io_outs_right[43] ;
 wire \_ces_2_1_io_outs_right[44] ;
 wire \_ces_2_1_io_outs_right[45] ;
 wire \_ces_2_1_io_outs_right[46] ;
 wire \_ces_2_1_io_outs_right[47] ;
 wire \_ces_2_1_io_outs_right[48] ;
 wire \_ces_2_1_io_outs_right[49] ;
 wire \_ces_2_1_io_outs_right[4] ;
 wire \_ces_2_1_io_outs_right[50] ;
 wire \_ces_2_1_io_outs_right[51] ;
 wire \_ces_2_1_io_outs_right[52] ;
 wire \_ces_2_1_io_outs_right[53] ;
 wire \_ces_2_1_io_outs_right[54] ;
 wire \_ces_2_1_io_outs_right[55] ;
 wire \_ces_2_1_io_outs_right[56] ;
 wire \_ces_2_1_io_outs_right[57] ;
 wire \_ces_2_1_io_outs_right[58] ;
 wire \_ces_2_1_io_outs_right[59] ;
 wire \_ces_2_1_io_outs_right[5] ;
 wire \_ces_2_1_io_outs_right[60] ;
 wire \_ces_2_1_io_outs_right[61] ;
 wire \_ces_2_1_io_outs_right[62] ;
 wire \_ces_2_1_io_outs_right[63] ;
 wire \_ces_2_1_io_outs_right[6] ;
 wire \_ces_2_1_io_outs_right[7] ;
 wire \_ces_2_1_io_outs_right[8] ;
 wire \_ces_2_1_io_outs_right[9] ;
 wire \_ces_2_1_io_outs_up[0] ;
 wire \_ces_2_1_io_outs_up[10] ;
 wire \_ces_2_1_io_outs_up[11] ;
 wire \_ces_2_1_io_outs_up[12] ;
 wire \_ces_2_1_io_outs_up[13] ;
 wire \_ces_2_1_io_outs_up[14] ;
 wire \_ces_2_1_io_outs_up[15] ;
 wire \_ces_2_1_io_outs_up[16] ;
 wire \_ces_2_1_io_outs_up[17] ;
 wire \_ces_2_1_io_outs_up[18] ;
 wire \_ces_2_1_io_outs_up[19] ;
 wire \_ces_2_1_io_outs_up[1] ;
 wire \_ces_2_1_io_outs_up[20] ;
 wire \_ces_2_1_io_outs_up[21] ;
 wire \_ces_2_1_io_outs_up[22] ;
 wire \_ces_2_1_io_outs_up[23] ;
 wire \_ces_2_1_io_outs_up[24] ;
 wire \_ces_2_1_io_outs_up[25] ;
 wire \_ces_2_1_io_outs_up[26] ;
 wire \_ces_2_1_io_outs_up[27] ;
 wire \_ces_2_1_io_outs_up[28] ;
 wire \_ces_2_1_io_outs_up[29] ;
 wire \_ces_2_1_io_outs_up[2] ;
 wire \_ces_2_1_io_outs_up[30] ;
 wire \_ces_2_1_io_outs_up[31] ;
 wire \_ces_2_1_io_outs_up[32] ;
 wire \_ces_2_1_io_outs_up[33] ;
 wire \_ces_2_1_io_outs_up[34] ;
 wire \_ces_2_1_io_outs_up[35] ;
 wire \_ces_2_1_io_outs_up[36] ;
 wire \_ces_2_1_io_outs_up[37] ;
 wire \_ces_2_1_io_outs_up[38] ;
 wire \_ces_2_1_io_outs_up[39] ;
 wire \_ces_2_1_io_outs_up[3] ;
 wire \_ces_2_1_io_outs_up[40] ;
 wire \_ces_2_1_io_outs_up[41] ;
 wire \_ces_2_1_io_outs_up[42] ;
 wire \_ces_2_1_io_outs_up[43] ;
 wire \_ces_2_1_io_outs_up[44] ;
 wire \_ces_2_1_io_outs_up[45] ;
 wire \_ces_2_1_io_outs_up[46] ;
 wire \_ces_2_1_io_outs_up[47] ;
 wire \_ces_2_1_io_outs_up[48] ;
 wire \_ces_2_1_io_outs_up[49] ;
 wire \_ces_2_1_io_outs_up[4] ;
 wire \_ces_2_1_io_outs_up[50] ;
 wire \_ces_2_1_io_outs_up[51] ;
 wire \_ces_2_1_io_outs_up[52] ;
 wire \_ces_2_1_io_outs_up[53] ;
 wire \_ces_2_1_io_outs_up[54] ;
 wire \_ces_2_1_io_outs_up[55] ;
 wire \_ces_2_1_io_outs_up[56] ;
 wire \_ces_2_1_io_outs_up[57] ;
 wire \_ces_2_1_io_outs_up[58] ;
 wire \_ces_2_1_io_outs_up[59] ;
 wire \_ces_2_1_io_outs_up[5] ;
 wire \_ces_2_1_io_outs_up[60] ;
 wire \_ces_2_1_io_outs_up[61] ;
 wire \_ces_2_1_io_outs_up[62] ;
 wire \_ces_2_1_io_outs_up[63] ;
 wire \_ces_2_1_io_outs_up[6] ;
 wire \_ces_2_1_io_outs_up[7] ;
 wire \_ces_2_1_io_outs_up[8] ;
 wire \_ces_2_1_io_outs_up[9] ;
 wire _ces_2_2_io_lsbOuts_1;
 wire _ces_2_2_io_lsbOuts_2;
 wire _ces_2_2_io_lsbOuts_3;
 wire \_ces_2_2_io_outs_down[0] ;
 wire \_ces_2_2_io_outs_down[10] ;
 wire \_ces_2_2_io_outs_down[11] ;
 wire \_ces_2_2_io_outs_down[12] ;
 wire \_ces_2_2_io_outs_down[13] ;
 wire \_ces_2_2_io_outs_down[14] ;
 wire \_ces_2_2_io_outs_down[15] ;
 wire \_ces_2_2_io_outs_down[16] ;
 wire \_ces_2_2_io_outs_down[17] ;
 wire \_ces_2_2_io_outs_down[18] ;
 wire \_ces_2_2_io_outs_down[19] ;
 wire \_ces_2_2_io_outs_down[1] ;
 wire \_ces_2_2_io_outs_down[20] ;
 wire \_ces_2_2_io_outs_down[21] ;
 wire \_ces_2_2_io_outs_down[22] ;
 wire \_ces_2_2_io_outs_down[23] ;
 wire \_ces_2_2_io_outs_down[24] ;
 wire \_ces_2_2_io_outs_down[25] ;
 wire \_ces_2_2_io_outs_down[26] ;
 wire \_ces_2_2_io_outs_down[27] ;
 wire \_ces_2_2_io_outs_down[28] ;
 wire \_ces_2_2_io_outs_down[29] ;
 wire \_ces_2_2_io_outs_down[2] ;
 wire \_ces_2_2_io_outs_down[30] ;
 wire \_ces_2_2_io_outs_down[31] ;
 wire \_ces_2_2_io_outs_down[32] ;
 wire \_ces_2_2_io_outs_down[33] ;
 wire \_ces_2_2_io_outs_down[34] ;
 wire \_ces_2_2_io_outs_down[35] ;
 wire \_ces_2_2_io_outs_down[36] ;
 wire \_ces_2_2_io_outs_down[37] ;
 wire \_ces_2_2_io_outs_down[38] ;
 wire \_ces_2_2_io_outs_down[39] ;
 wire \_ces_2_2_io_outs_down[3] ;
 wire \_ces_2_2_io_outs_down[40] ;
 wire \_ces_2_2_io_outs_down[41] ;
 wire \_ces_2_2_io_outs_down[42] ;
 wire \_ces_2_2_io_outs_down[43] ;
 wire \_ces_2_2_io_outs_down[44] ;
 wire \_ces_2_2_io_outs_down[45] ;
 wire \_ces_2_2_io_outs_down[46] ;
 wire \_ces_2_2_io_outs_down[47] ;
 wire \_ces_2_2_io_outs_down[48] ;
 wire \_ces_2_2_io_outs_down[49] ;
 wire \_ces_2_2_io_outs_down[4] ;
 wire \_ces_2_2_io_outs_down[50] ;
 wire \_ces_2_2_io_outs_down[51] ;
 wire \_ces_2_2_io_outs_down[52] ;
 wire \_ces_2_2_io_outs_down[53] ;
 wire \_ces_2_2_io_outs_down[54] ;
 wire \_ces_2_2_io_outs_down[55] ;
 wire \_ces_2_2_io_outs_down[56] ;
 wire \_ces_2_2_io_outs_down[57] ;
 wire \_ces_2_2_io_outs_down[58] ;
 wire \_ces_2_2_io_outs_down[59] ;
 wire \_ces_2_2_io_outs_down[5] ;
 wire \_ces_2_2_io_outs_down[60] ;
 wire \_ces_2_2_io_outs_down[61] ;
 wire \_ces_2_2_io_outs_down[62] ;
 wire \_ces_2_2_io_outs_down[63] ;
 wire \_ces_2_2_io_outs_down[6] ;
 wire \_ces_2_2_io_outs_down[7] ;
 wire \_ces_2_2_io_outs_down[8] ;
 wire \_ces_2_2_io_outs_down[9] ;
 wire \_ces_2_2_io_outs_left[0] ;
 wire \_ces_2_2_io_outs_left[10] ;
 wire \_ces_2_2_io_outs_left[11] ;
 wire \_ces_2_2_io_outs_left[12] ;
 wire \_ces_2_2_io_outs_left[13] ;
 wire \_ces_2_2_io_outs_left[14] ;
 wire \_ces_2_2_io_outs_left[15] ;
 wire \_ces_2_2_io_outs_left[16] ;
 wire \_ces_2_2_io_outs_left[17] ;
 wire \_ces_2_2_io_outs_left[18] ;
 wire \_ces_2_2_io_outs_left[19] ;
 wire \_ces_2_2_io_outs_left[1] ;
 wire \_ces_2_2_io_outs_left[20] ;
 wire \_ces_2_2_io_outs_left[21] ;
 wire \_ces_2_2_io_outs_left[22] ;
 wire \_ces_2_2_io_outs_left[23] ;
 wire \_ces_2_2_io_outs_left[24] ;
 wire \_ces_2_2_io_outs_left[25] ;
 wire \_ces_2_2_io_outs_left[26] ;
 wire \_ces_2_2_io_outs_left[27] ;
 wire \_ces_2_2_io_outs_left[28] ;
 wire \_ces_2_2_io_outs_left[29] ;
 wire \_ces_2_2_io_outs_left[2] ;
 wire \_ces_2_2_io_outs_left[30] ;
 wire \_ces_2_2_io_outs_left[31] ;
 wire \_ces_2_2_io_outs_left[32] ;
 wire \_ces_2_2_io_outs_left[33] ;
 wire \_ces_2_2_io_outs_left[34] ;
 wire \_ces_2_2_io_outs_left[35] ;
 wire \_ces_2_2_io_outs_left[36] ;
 wire \_ces_2_2_io_outs_left[37] ;
 wire \_ces_2_2_io_outs_left[38] ;
 wire \_ces_2_2_io_outs_left[39] ;
 wire \_ces_2_2_io_outs_left[3] ;
 wire \_ces_2_2_io_outs_left[40] ;
 wire \_ces_2_2_io_outs_left[41] ;
 wire \_ces_2_2_io_outs_left[42] ;
 wire \_ces_2_2_io_outs_left[43] ;
 wire \_ces_2_2_io_outs_left[44] ;
 wire \_ces_2_2_io_outs_left[45] ;
 wire \_ces_2_2_io_outs_left[46] ;
 wire \_ces_2_2_io_outs_left[47] ;
 wire \_ces_2_2_io_outs_left[48] ;
 wire \_ces_2_2_io_outs_left[49] ;
 wire \_ces_2_2_io_outs_left[4] ;
 wire \_ces_2_2_io_outs_left[50] ;
 wire \_ces_2_2_io_outs_left[51] ;
 wire \_ces_2_2_io_outs_left[52] ;
 wire \_ces_2_2_io_outs_left[53] ;
 wire \_ces_2_2_io_outs_left[54] ;
 wire \_ces_2_2_io_outs_left[55] ;
 wire \_ces_2_2_io_outs_left[56] ;
 wire \_ces_2_2_io_outs_left[57] ;
 wire \_ces_2_2_io_outs_left[58] ;
 wire \_ces_2_2_io_outs_left[59] ;
 wire \_ces_2_2_io_outs_left[5] ;
 wire \_ces_2_2_io_outs_left[60] ;
 wire \_ces_2_2_io_outs_left[61] ;
 wire \_ces_2_2_io_outs_left[62] ;
 wire \_ces_2_2_io_outs_left[63] ;
 wire \_ces_2_2_io_outs_left[6] ;
 wire \_ces_2_2_io_outs_left[7] ;
 wire \_ces_2_2_io_outs_left[8] ;
 wire \_ces_2_2_io_outs_left[9] ;
 wire \_ces_2_2_io_outs_right[0] ;
 wire \_ces_2_2_io_outs_right[10] ;
 wire \_ces_2_2_io_outs_right[11] ;
 wire \_ces_2_2_io_outs_right[12] ;
 wire \_ces_2_2_io_outs_right[13] ;
 wire \_ces_2_2_io_outs_right[14] ;
 wire \_ces_2_2_io_outs_right[15] ;
 wire \_ces_2_2_io_outs_right[16] ;
 wire \_ces_2_2_io_outs_right[17] ;
 wire \_ces_2_2_io_outs_right[18] ;
 wire \_ces_2_2_io_outs_right[19] ;
 wire \_ces_2_2_io_outs_right[1] ;
 wire \_ces_2_2_io_outs_right[20] ;
 wire \_ces_2_2_io_outs_right[21] ;
 wire \_ces_2_2_io_outs_right[22] ;
 wire \_ces_2_2_io_outs_right[23] ;
 wire \_ces_2_2_io_outs_right[24] ;
 wire \_ces_2_2_io_outs_right[25] ;
 wire \_ces_2_2_io_outs_right[26] ;
 wire \_ces_2_2_io_outs_right[27] ;
 wire \_ces_2_2_io_outs_right[28] ;
 wire \_ces_2_2_io_outs_right[29] ;
 wire \_ces_2_2_io_outs_right[2] ;
 wire \_ces_2_2_io_outs_right[30] ;
 wire \_ces_2_2_io_outs_right[31] ;
 wire \_ces_2_2_io_outs_right[32] ;
 wire \_ces_2_2_io_outs_right[33] ;
 wire \_ces_2_2_io_outs_right[34] ;
 wire \_ces_2_2_io_outs_right[35] ;
 wire \_ces_2_2_io_outs_right[36] ;
 wire \_ces_2_2_io_outs_right[37] ;
 wire \_ces_2_2_io_outs_right[38] ;
 wire \_ces_2_2_io_outs_right[39] ;
 wire \_ces_2_2_io_outs_right[3] ;
 wire \_ces_2_2_io_outs_right[40] ;
 wire \_ces_2_2_io_outs_right[41] ;
 wire \_ces_2_2_io_outs_right[42] ;
 wire \_ces_2_2_io_outs_right[43] ;
 wire \_ces_2_2_io_outs_right[44] ;
 wire \_ces_2_2_io_outs_right[45] ;
 wire \_ces_2_2_io_outs_right[46] ;
 wire \_ces_2_2_io_outs_right[47] ;
 wire \_ces_2_2_io_outs_right[48] ;
 wire \_ces_2_2_io_outs_right[49] ;
 wire \_ces_2_2_io_outs_right[4] ;
 wire \_ces_2_2_io_outs_right[50] ;
 wire \_ces_2_2_io_outs_right[51] ;
 wire \_ces_2_2_io_outs_right[52] ;
 wire \_ces_2_2_io_outs_right[53] ;
 wire \_ces_2_2_io_outs_right[54] ;
 wire \_ces_2_2_io_outs_right[55] ;
 wire \_ces_2_2_io_outs_right[56] ;
 wire \_ces_2_2_io_outs_right[57] ;
 wire \_ces_2_2_io_outs_right[58] ;
 wire \_ces_2_2_io_outs_right[59] ;
 wire \_ces_2_2_io_outs_right[5] ;
 wire \_ces_2_2_io_outs_right[60] ;
 wire \_ces_2_2_io_outs_right[61] ;
 wire \_ces_2_2_io_outs_right[62] ;
 wire \_ces_2_2_io_outs_right[63] ;
 wire \_ces_2_2_io_outs_right[6] ;
 wire \_ces_2_2_io_outs_right[7] ;
 wire \_ces_2_2_io_outs_right[8] ;
 wire \_ces_2_2_io_outs_right[9] ;
 wire \_ces_2_2_io_outs_up[0] ;
 wire \_ces_2_2_io_outs_up[10] ;
 wire \_ces_2_2_io_outs_up[11] ;
 wire \_ces_2_2_io_outs_up[12] ;
 wire \_ces_2_2_io_outs_up[13] ;
 wire \_ces_2_2_io_outs_up[14] ;
 wire \_ces_2_2_io_outs_up[15] ;
 wire \_ces_2_2_io_outs_up[16] ;
 wire \_ces_2_2_io_outs_up[17] ;
 wire \_ces_2_2_io_outs_up[18] ;
 wire \_ces_2_2_io_outs_up[19] ;
 wire \_ces_2_2_io_outs_up[1] ;
 wire \_ces_2_2_io_outs_up[20] ;
 wire \_ces_2_2_io_outs_up[21] ;
 wire \_ces_2_2_io_outs_up[22] ;
 wire \_ces_2_2_io_outs_up[23] ;
 wire \_ces_2_2_io_outs_up[24] ;
 wire \_ces_2_2_io_outs_up[25] ;
 wire \_ces_2_2_io_outs_up[26] ;
 wire \_ces_2_2_io_outs_up[27] ;
 wire \_ces_2_2_io_outs_up[28] ;
 wire \_ces_2_2_io_outs_up[29] ;
 wire \_ces_2_2_io_outs_up[2] ;
 wire \_ces_2_2_io_outs_up[30] ;
 wire \_ces_2_2_io_outs_up[31] ;
 wire \_ces_2_2_io_outs_up[32] ;
 wire \_ces_2_2_io_outs_up[33] ;
 wire \_ces_2_2_io_outs_up[34] ;
 wire \_ces_2_2_io_outs_up[35] ;
 wire \_ces_2_2_io_outs_up[36] ;
 wire \_ces_2_2_io_outs_up[37] ;
 wire \_ces_2_2_io_outs_up[38] ;
 wire \_ces_2_2_io_outs_up[39] ;
 wire \_ces_2_2_io_outs_up[3] ;
 wire \_ces_2_2_io_outs_up[40] ;
 wire \_ces_2_2_io_outs_up[41] ;
 wire \_ces_2_2_io_outs_up[42] ;
 wire \_ces_2_2_io_outs_up[43] ;
 wire \_ces_2_2_io_outs_up[44] ;
 wire \_ces_2_2_io_outs_up[45] ;
 wire \_ces_2_2_io_outs_up[46] ;
 wire \_ces_2_2_io_outs_up[47] ;
 wire \_ces_2_2_io_outs_up[48] ;
 wire \_ces_2_2_io_outs_up[49] ;
 wire \_ces_2_2_io_outs_up[4] ;
 wire \_ces_2_2_io_outs_up[50] ;
 wire \_ces_2_2_io_outs_up[51] ;
 wire \_ces_2_2_io_outs_up[52] ;
 wire \_ces_2_2_io_outs_up[53] ;
 wire \_ces_2_2_io_outs_up[54] ;
 wire \_ces_2_2_io_outs_up[55] ;
 wire \_ces_2_2_io_outs_up[56] ;
 wire \_ces_2_2_io_outs_up[57] ;
 wire \_ces_2_2_io_outs_up[58] ;
 wire \_ces_2_2_io_outs_up[59] ;
 wire \_ces_2_2_io_outs_up[5] ;
 wire \_ces_2_2_io_outs_up[60] ;
 wire \_ces_2_2_io_outs_up[61] ;
 wire \_ces_2_2_io_outs_up[62] ;
 wire \_ces_2_2_io_outs_up[63] ;
 wire \_ces_2_2_io_outs_up[6] ;
 wire \_ces_2_2_io_outs_up[7] ;
 wire \_ces_2_2_io_outs_up[8] ;
 wire \_ces_2_2_io_outs_up[9] ;
 wire _ces_2_3_io_lsbOuts_0;
 wire _ces_2_3_io_lsbOuts_1;
 wire _ces_2_3_io_lsbOuts_2;
 wire _ces_2_3_io_lsbOuts_3;
 wire \_ces_2_3_io_outs_down[0] ;
 wire \_ces_2_3_io_outs_down[10] ;
 wire \_ces_2_3_io_outs_down[11] ;
 wire \_ces_2_3_io_outs_down[12] ;
 wire \_ces_2_3_io_outs_down[13] ;
 wire \_ces_2_3_io_outs_down[14] ;
 wire \_ces_2_3_io_outs_down[15] ;
 wire \_ces_2_3_io_outs_down[16] ;
 wire \_ces_2_3_io_outs_down[17] ;
 wire \_ces_2_3_io_outs_down[18] ;
 wire \_ces_2_3_io_outs_down[19] ;
 wire \_ces_2_3_io_outs_down[1] ;
 wire \_ces_2_3_io_outs_down[20] ;
 wire \_ces_2_3_io_outs_down[21] ;
 wire \_ces_2_3_io_outs_down[22] ;
 wire \_ces_2_3_io_outs_down[23] ;
 wire \_ces_2_3_io_outs_down[24] ;
 wire \_ces_2_3_io_outs_down[25] ;
 wire \_ces_2_3_io_outs_down[26] ;
 wire \_ces_2_3_io_outs_down[27] ;
 wire \_ces_2_3_io_outs_down[28] ;
 wire \_ces_2_3_io_outs_down[29] ;
 wire \_ces_2_3_io_outs_down[2] ;
 wire \_ces_2_3_io_outs_down[30] ;
 wire \_ces_2_3_io_outs_down[31] ;
 wire \_ces_2_3_io_outs_down[32] ;
 wire \_ces_2_3_io_outs_down[33] ;
 wire \_ces_2_3_io_outs_down[34] ;
 wire \_ces_2_3_io_outs_down[35] ;
 wire \_ces_2_3_io_outs_down[36] ;
 wire \_ces_2_3_io_outs_down[37] ;
 wire \_ces_2_3_io_outs_down[38] ;
 wire \_ces_2_3_io_outs_down[39] ;
 wire \_ces_2_3_io_outs_down[3] ;
 wire \_ces_2_3_io_outs_down[40] ;
 wire \_ces_2_3_io_outs_down[41] ;
 wire \_ces_2_3_io_outs_down[42] ;
 wire \_ces_2_3_io_outs_down[43] ;
 wire \_ces_2_3_io_outs_down[44] ;
 wire \_ces_2_3_io_outs_down[45] ;
 wire \_ces_2_3_io_outs_down[46] ;
 wire \_ces_2_3_io_outs_down[47] ;
 wire \_ces_2_3_io_outs_down[48] ;
 wire \_ces_2_3_io_outs_down[49] ;
 wire \_ces_2_3_io_outs_down[4] ;
 wire \_ces_2_3_io_outs_down[50] ;
 wire \_ces_2_3_io_outs_down[51] ;
 wire \_ces_2_3_io_outs_down[52] ;
 wire \_ces_2_3_io_outs_down[53] ;
 wire \_ces_2_3_io_outs_down[54] ;
 wire \_ces_2_3_io_outs_down[55] ;
 wire \_ces_2_3_io_outs_down[56] ;
 wire \_ces_2_3_io_outs_down[57] ;
 wire \_ces_2_3_io_outs_down[58] ;
 wire \_ces_2_3_io_outs_down[59] ;
 wire \_ces_2_3_io_outs_down[5] ;
 wire \_ces_2_3_io_outs_down[60] ;
 wire \_ces_2_3_io_outs_down[61] ;
 wire \_ces_2_3_io_outs_down[62] ;
 wire \_ces_2_3_io_outs_down[63] ;
 wire \_ces_2_3_io_outs_down[6] ;
 wire \_ces_2_3_io_outs_down[7] ;
 wire \_ces_2_3_io_outs_down[8] ;
 wire \_ces_2_3_io_outs_down[9] ;
 wire \_ces_2_3_io_outs_left[0] ;
 wire \_ces_2_3_io_outs_left[10] ;
 wire \_ces_2_3_io_outs_left[11] ;
 wire \_ces_2_3_io_outs_left[12] ;
 wire \_ces_2_3_io_outs_left[13] ;
 wire \_ces_2_3_io_outs_left[14] ;
 wire \_ces_2_3_io_outs_left[15] ;
 wire \_ces_2_3_io_outs_left[16] ;
 wire \_ces_2_3_io_outs_left[17] ;
 wire \_ces_2_3_io_outs_left[18] ;
 wire \_ces_2_3_io_outs_left[19] ;
 wire \_ces_2_3_io_outs_left[1] ;
 wire \_ces_2_3_io_outs_left[20] ;
 wire \_ces_2_3_io_outs_left[21] ;
 wire \_ces_2_3_io_outs_left[22] ;
 wire \_ces_2_3_io_outs_left[23] ;
 wire \_ces_2_3_io_outs_left[24] ;
 wire \_ces_2_3_io_outs_left[25] ;
 wire \_ces_2_3_io_outs_left[26] ;
 wire \_ces_2_3_io_outs_left[27] ;
 wire \_ces_2_3_io_outs_left[28] ;
 wire \_ces_2_3_io_outs_left[29] ;
 wire \_ces_2_3_io_outs_left[2] ;
 wire \_ces_2_3_io_outs_left[30] ;
 wire \_ces_2_3_io_outs_left[31] ;
 wire \_ces_2_3_io_outs_left[32] ;
 wire \_ces_2_3_io_outs_left[33] ;
 wire \_ces_2_3_io_outs_left[34] ;
 wire \_ces_2_3_io_outs_left[35] ;
 wire \_ces_2_3_io_outs_left[36] ;
 wire \_ces_2_3_io_outs_left[37] ;
 wire \_ces_2_3_io_outs_left[38] ;
 wire \_ces_2_3_io_outs_left[39] ;
 wire \_ces_2_3_io_outs_left[3] ;
 wire \_ces_2_3_io_outs_left[40] ;
 wire \_ces_2_3_io_outs_left[41] ;
 wire \_ces_2_3_io_outs_left[42] ;
 wire \_ces_2_3_io_outs_left[43] ;
 wire \_ces_2_3_io_outs_left[44] ;
 wire \_ces_2_3_io_outs_left[45] ;
 wire \_ces_2_3_io_outs_left[46] ;
 wire \_ces_2_3_io_outs_left[47] ;
 wire \_ces_2_3_io_outs_left[48] ;
 wire \_ces_2_3_io_outs_left[49] ;
 wire \_ces_2_3_io_outs_left[4] ;
 wire \_ces_2_3_io_outs_left[50] ;
 wire \_ces_2_3_io_outs_left[51] ;
 wire \_ces_2_3_io_outs_left[52] ;
 wire \_ces_2_3_io_outs_left[53] ;
 wire \_ces_2_3_io_outs_left[54] ;
 wire \_ces_2_3_io_outs_left[55] ;
 wire \_ces_2_3_io_outs_left[56] ;
 wire \_ces_2_3_io_outs_left[57] ;
 wire \_ces_2_3_io_outs_left[58] ;
 wire \_ces_2_3_io_outs_left[59] ;
 wire \_ces_2_3_io_outs_left[5] ;
 wire \_ces_2_3_io_outs_left[60] ;
 wire \_ces_2_3_io_outs_left[61] ;
 wire \_ces_2_3_io_outs_left[62] ;
 wire \_ces_2_3_io_outs_left[63] ;
 wire \_ces_2_3_io_outs_left[6] ;
 wire \_ces_2_3_io_outs_left[7] ;
 wire \_ces_2_3_io_outs_left[8] ;
 wire \_ces_2_3_io_outs_left[9] ;
 wire \_ces_2_3_io_outs_up[0] ;
 wire \_ces_2_3_io_outs_up[10] ;
 wire \_ces_2_3_io_outs_up[11] ;
 wire \_ces_2_3_io_outs_up[12] ;
 wire \_ces_2_3_io_outs_up[13] ;
 wire \_ces_2_3_io_outs_up[14] ;
 wire \_ces_2_3_io_outs_up[15] ;
 wire \_ces_2_3_io_outs_up[16] ;
 wire \_ces_2_3_io_outs_up[17] ;
 wire \_ces_2_3_io_outs_up[18] ;
 wire \_ces_2_3_io_outs_up[19] ;
 wire \_ces_2_3_io_outs_up[1] ;
 wire \_ces_2_3_io_outs_up[20] ;
 wire \_ces_2_3_io_outs_up[21] ;
 wire \_ces_2_3_io_outs_up[22] ;
 wire \_ces_2_3_io_outs_up[23] ;
 wire \_ces_2_3_io_outs_up[24] ;
 wire \_ces_2_3_io_outs_up[25] ;
 wire \_ces_2_3_io_outs_up[26] ;
 wire \_ces_2_3_io_outs_up[27] ;
 wire \_ces_2_3_io_outs_up[28] ;
 wire \_ces_2_3_io_outs_up[29] ;
 wire \_ces_2_3_io_outs_up[2] ;
 wire \_ces_2_3_io_outs_up[30] ;
 wire \_ces_2_3_io_outs_up[31] ;
 wire \_ces_2_3_io_outs_up[32] ;
 wire \_ces_2_3_io_outs_up[33] ;
 wire \_ces_2_3_io_outs_up[34] ;
 wire \_ces_2_3_io_outs_up[35] ;
 wire \_ces_2_3_io_outs_up[36] ;
 wire \_ces_2_3_io_outs_up[37] ;
 wire \_ces_2_3_io_outs_up[38] ;
 wire \_ces_2_3_io_outs_up[39] ;
 wire \_ces_2_3_io_outs_up[3] ;
 wire \_ces_2_3_io_outs_up[40] ;
 wire \_ces_2_3_io_outs_up[41] ;
 wire \_ces_2_3_io_outs_up[42] ;
 wire \_ces_2_3_io_outs_up[43] ;
 wire \_ces_2_3_io_outs_up[44] ;
 wire \_ces_2_3_io_outs_up[45] ;
 wire \_ces_2_3_io_outs_up[46] ;
 wire \_ces_2_3_io_outs_up[47] ;
 wire \_ces_2_3_io_outs_up[48] ;
 wire \_ces_2_3_io_outs_up[49] ;
 wire \_ces_2_3_io_outs_up[4] ;
 wire \_ces_2_3_io_outs_up[50] ;
 wire \_ces_2_3_io_outs_up[51] ;
 wire \_ces_2_3_io_outs_up[52] ;
 wire \_ces_2_3_io_outs_up[53] ;
 wire \_ces_2_3_io_outs_up[54] ;
 wire \_ces_2_3_io_outs_up[55] ;
 wire \_ces_2_3_io_outs_up[56] ;
 wire \_ces_2_3_io_outs_up[57] ;
 wire \_ces_2_3_io_outs_up[58] ;
 wire \_ces_2_3_io_outs_up[59] ;
 wire \_ces_2_3_io_outs_up[5] ;
 wire \_ces_2_3_io_outs_up[60] ;
 wire \_ces_2_3_io_outs_up[61] ;
 wire \_ces_2_3_io_outs_up[62] ;
 wire \_ces_2_3_io_outs_up[63] ;
 wire \_ces_2_3_io_outs_up[6] ;
 wire \_ces_2_3_io_outs_up[7] ;
 wire \_ces_2_3_io_outs_up[8] ;
 wire \_ces_2_3_io_outs_up[9] ;
 wire _ces_3_0_io_lsbOuts_1;
 wire _ces_3_0_io_lsbOuts_2;
 wire _ces_3_0_io_lsbOuts_3;
 wire \_ces_3_0_io_outs_down[0] ;
 wire \_ces_3_0_io_outs_down[10] ;
 wire \_ces_3_0_io_outs_down[11] ;
 wire \_ces_3_0_io_outs_down[12] ;
 wire \_ces_3_0_io_outs_down[13] ;
 wire \_ces_3_0_io_outs_down[14] ;
 wire \_ces_3_0_io_outs_down[15] ;
 wire \_ces_3_0_io_outs_down[16] ;
 wire \_ces_3_0_io_outs_down[17] ;
 wire \_ces_3_0_io_outs_down[18] ;
 wire \_ces_3_0_io_outs_down[19] ;
 wire \_ces_3_0_io_outs_down[1] ;
 wire \_ces_3_0_io_outs_down[20] ;
 wire \_ces_3_0_io_outs_down[21] ;
 wire \_ces_3_0_io_outs_down[22] ;
 wire \_ces_3_0_io_outs_down[23] ;
 wire \_ces_3_0_io_outs_down[24] ;
 wire \_ces_3_0_io_outs_down[25] ;
 wire \_ces_3_0_io_outs_down[26] ;
 wire \_ces_3_0_io_outs_down[27] ;
 wire \_ces_3_0_io_outs_down[28] ;
 wire \_ces_3_0_io_outs_down[29] ;
 wire \_ces_3_0_io_outs_down[2] ;
 wire \_ces_3_0_io_outs_down[30] ;
 wire \_ces_3_0_io_outs_down[31] ;
 wire \_ces_3_0_io_outs_down[32] ;
 wire \_ces_3_0_io_outs_down[33] ;
 wire \_ces_3_0_io_outs_down[34] ;
 wire \_ces_3_0_io_outs_down[35] ;
 wire \_ces_3_0_io_outs_down[36] ;
 wire \_ces_3_0_io_outs_down[37] ;
 wire \_ces_3_0_io_outs_down[38] ;
 wire \_ces_3_0_io_outs_down[39] ;
 wire \_ces_3_0_io_outs_down[3] ;
 wire \_ces_3_0_io_outs_down[40] ;
 wire \_ces_3_0_io_outs_down[41] ;
 wire \_ces_3_0_io_outs_down[42] ;
 wire \_ces_3_0_io_outs_down[43] ;
 wire \_ces_3_0_io_outs_down[44] ;
 wire \_ces_3_0_io_outs_down[45] ;
 wire \_ces_3_0_io_outs_down[46] ;
 wire \_ces_3_0_io_outs_down[47] ;
 wire \_ces_3_0_io_outs_down[48] ;
 wire \_ces_3_0_io_outs_down[49] ;
 wire \_ces_3_0_io_outs_down[4] ;
 wire \_ces_3_0_io_outs_down[50] ;
 wire \_ces_3_0_io_outs_down[51] ;
 wire \_ces_3_0_io_outs_down[52] ;
 wire \_ces_3_0_io_outs_down[53] ;
 wire \_ces_3_0_io_outs_down[54] ;
 wire \_ces_3_0_io_outs_down[55] ;
 wire \_ces_3_0_io_outs_down[56] ;
 wire \_ces_3_0_io_outs_down[57] ;
 wire \_ces_3_0_io_outs_down[58] ;
 wire \_ces_3_0_io_outs_down[59] ;
 wire \_ces_3_0_io_outs_down[5] ;
 wire \_ces_3_0_io_outs_down[60] ;
 wire \_ces_3_0_io_outs_down[61] ;
 wire \_ces_3_0_io_outs_down[62] ;
 wire \_ces_3_0_io_outs_down[63] ;
 wire \_ces_3_0_io_outs_down[6] ;
 wire \_ces_3_0_io_outs_down[7] ;
 wire \_ces_3_0_io_outs_down[8] ;
 wire \_ces_3_0_io_outs_down[9] ;
 wire \_ces_3_0_io_outs_right[0] ;
 wire \_ces_3_0_io_outs_right[10] ;
 wire \_ces_3_0_io_outs_right[11] ;
 wire \_ces_3_0_io_outs_right[12] ;
 wire \_ces_3_0_io_outs_right[13] ;
 wire \_ces_3_0_io_outs_right[14] ;
 wire \_ces_3_0_io_outs_right[15] ;
 wire \_ces_3_0_io_outs_right[16] ;
 wire \_ces_3_0_io_outs_right[17] ;
 wire \_ces_3_0_io_outs_right[18] ;
 wire \_ces_3_0_io_outs_right[19] ;
 wire \_ces_3_0_io_outs_right[1] ;
 wire \_ces_3_0_io_outs_right[20] ;
 wire \_ces_3_0_io_outs_right[21] ;
 wire \_ces_3_0_io_outs_right[22] ;
 wire \_ces_3_0_io_outs_right[23] ;
 wire \_ces_3_0_io_outs_right[24] ;
 wire \_ces_3_0_io_outs_right[25] ;
 wire \_ces_3_0_io_outs_right[26] ;
 wire \_ces_3_0_io_outs_right[27] ;
 wire \_ces_3_0_io_outs_right[28] ;
 wire \_ces_3_0_io_outs_right[29] ;
 wire \_ces_3_0_io_outs_right[2] ;
 wire \_ces_3_0_io_outs_right[30] ;
 wire \_ces_3_0_io_outs_right[31] ;
 wire \_ces_3_0_io_outs_right[32] ;
 wire \_ces_3_0_io_outs_right[33] ;
 wire \_ces_3_0_io_outs_right[34] ;
 wire \_ces_3_0_io_outs_right[35] ;
 wire \_ces_3_0_io_outs_right[36] ;
 wire \_ces_3_0_io_outs_right[37] ;
 wire \_ces_3_0_io_outs_right[38] ;
 wire \_ces_3_0_io_outs_right[39] ;
 wire \_ces_3_0_io_outs_right[3] ;
 wire \_ces_3_0_io_outs_right[40] ;
 wire \_ces_3_0_io_outs_right[41] ;
 wire \_ces_3_0_io_outs_right[42] ;
 wire \_ces_3_0_io_outs_right[43] ;
 wire \_ces_3_0_io_outs_right[44] ;
 wire \_ces_3_0_io_outs_right[45] ;
 wire \_ces_3_0_io_outs_right[46] ;
 wire \_ces_3_0_io_outs_right[47] ;
 wire \_ces_3_0_io_outs_right[48] ;
 wire \_ces_3_0_io_outs_right[49] ;
 wire \_ces_3_0_io_outs_right[4] ;
 wire \_ces_3_0_io_outs_right[50] ;
 wire \_ces_3_0_io_outs_right[51] ;
 wire \_ces_3_0_io_outs_right[52] ;
 wire \_ces_3_0_io_outs_right[53] ;
 wire \_ces_3_0_io_outs_right[54] ;
 wire \_ces_3_0_io_outs_right[55] ;
 wire \_ces_3_0_io_outs_right[56] ;
 wire \_ces_3_0_io_outs_right[57] ;
 wire \_ces_3_0_io_outs_right[58] ;
 wire \_ces_3_0_io_outs_right[59] ;
 wire \_ces_3_0_io_outs_right[5] ;
 wire \_ces_3_0_io_outs_right[60] ;
 wire \_ces_3_0_io_outs_right[61] ;
 wire \_ces_3_0_io_outs_right[62] ;
 wire \_ces_3_0_io_outs_right[63] ;
 wire \_ces_3_0_io_outs_right[6] ;
 wire \_ces_3_0_io_outs_right[7] ;
 wire \_ces_3_0_io_outs_right[8] ;
 wire \_ces_3_0_io_outs_right[9] ;
 wire _ces_3_1_io_lsbOuts_1;
 wire _ces_3_1_io_lsbOuts_2;
 wire _ces_3_1_io_lsbOuts_3;
 wire \_ces_3_1_io_outs_down[0] ;
 wire \_ces_3_1_io_outs_down[10] ;
 wire \_ces_3_1_io_outs_down[11] ;
 wire \_ces_3_1_io_outs_down[12] ;
 wire \_ces_3_1_io_outs_down[13] ;
 wire \_ces_3_1_io_outs_down[14] ;
 wire \_ces_3_1_io_outs_down[15] ;
 wire \_ces_3_1_io_outs_down[16] ;
 wire \_ces_3_1_io_outs_down[17] ;
 wire \_ces_3_1_io_outs_down[18] ;
 wire \_ces_3_1_io_outs_down[19] ;
 wire \_ces_3_1_io_outs_down[1] ;
 wire \_ces_3_1_io_outs_down[20] ;
 wire \_ces_3_1_io_outs_down[21] ;
 wire \_ces_3_1_io_outs_down[22] ;
 wire \_ces_3_1_io_outs_down[23] ;
 wire \_ces_3_1_io_outs_down[24] ;
 wire \_ces_3_1_io_outs_down[25] ;
 wire \_ces_3_1_io_outs_down[26] ;
 wire \_ces_3_1_io_outs_down[27] ;
 wire \_ces_3_1_io_outs_down[28] ;
 wire \_ces_3_1_io_outs_down[29] ;
 wire \_ces_3_1_io_outs_down[2] ;
 wire \_ces_3_1_io_outs_down[30] ;
 wire \_ces_3_1_io_outs_down[31] ;
 wire \_ces_3_1_io_outs_down[32] ;
 wire \_ces_3_1_io_outs_down[33] ;
 wire \_ces_3_1_io_outs_down[34] ;
 wire \_ces_3_1_io_outs_down[35] ;
 wire \_ces_3_1_io_outs_down[36] ;
 wire \_ces_3_1_io_outs_down[37] ;
 wire \_ces_3_1_io_outs_down[38] ;
 wire \_ces_3_1_io_outs_down[39] ;
 wire \_ces_3_1_io_outs_down[3] ;
 wire \_ces_3_1_io_outs_down[40] ;
 wire \_ces_3_1_io_outs_down[41] ;
 wire \_ces_3_1_io_outs_down[42] ;
 wire \_ces_3_1_io_outs_down[43] ;
 wire \_ces_3_1_io_outs_down[44] ;
 wire \_ces_3_1_io_outs_down[45] ;
 wire \_ces_3_1_io_outs_down[46] ;
 wire \_ces_3_1_io_outs_down[47] ;
 wire \_ces_3_1_io_outs_down[48] ;
 wire \_ces_3_1_io_outs_down[49] ;
 wire \_ces_3_1_io_outs_down[4] ;
 wire \_ces_3_1_io_outs_down[50] ;
 wire \_ces_3_1_io_outs_down[51] ;
 wire \_ces_3_1_io_outs_down[52] ;
 wire \_ces_3_1_io_outs_down[53] ;
 wire \_ces_3_1_io_outs_down[54] ;
 wire \_ces_3_1_io_outs_down[55] ;
 wire \_ces_3_1_io_outs_down[56] ;
 wire \_ces_3_1_io_outs_down[57] ;
 wire \_ces_3_1_io_outs_down[58] ;
 wire \_ces_3_1_io_outs_down[59] ;
 wire \_ces_3_1_io_outs_down[5] ;
 wire \_ces_3_1_io_outs_down[60] ;
 wire \_ces_3_1_io_outs_down[61] ;
 wire \_ces_3_1_io_outs_down[62] ;
 wire \_ces_3_1_io_outs_down[63] ;
 wire \_ces_3_1_io_outs_down[6] ;
 wire \_ces_3_1_io_outs_down[7] ;
 wire \_ces_3_1_io_outs_down[8] ;
 wire \_ces_3_1_io_outs_down[9] ;
 wire \_ces_3_1_io_outs_left[0] ;
 wire \_ces_3_1_io_outs_left[10] ;
 wire \_ces_3_1_io_outs_left[11] ;
 wire \_ces_3_1_io_outs_left[12] ;
 wire \_ces_3_1_io_outs_left[13] ;
 wire \_ces_3_1_io_outs_left[14] ;
 wire \_ces_3_1_io_outs_left[15] ;
 wire \_ces_3_1_io_outs_left[16] ;
 wire \_ces_3_1_io_outs_left[17] ;
 wire \_ces_3_1_io_outs_left[18] ;
 wire \_ces_3_1_io_outs_left[19] ;
 wire \_ces_3_1_io_outs_left[1] ;
 wire \_ces_3_1_io_outs_left[20] ;
 wire \_ces_3_1_io_outs_left[21] ;
 wire \_ces_3_1_io_outs_left[22] ;
 wire \_ces_3_1_io_outs_left[23] ;
 wire \_ces_3_1_io_outs_left[24] ;
 wire \_ces_3_1_io_outs_left[25] ;
 wire \_ces_3_1_io_outs_left[26] ;
 wire \_ces_3_1_io_outs_left[27] ;
 wire \_ces_3_1_io_outs_left[28] ;
 wire \_ces_3_1_io_outs_left[29] ;
 wire \_ces_3_1_io_outs_left[2] ;
 wire \_ces_3_1_io_outs_left[30] ;
 wire \_ces_3_1_io_outs_left[31] ;
 wire \_ces_3_1_io_outs_left[32] ;
 wire \_ces_3_1_io_outs_left[33] ;
 wire \_ces_3_1_io_outs_left[34] ;
 wire \_ces_3_1_io_outs_left[35] ;
 wire \_ces_3_1_io_outs_left[36] ;
 wire \_ces_3_1_io_outs_left[37] ;
 wire \_ces_3_1_io_outs_left[38] ;
 wire \_ces_3_1_io_outs_left[39] ;
 wire \_ces_3_1_io_outs_left[3] ;
 wire \_ces_3_1_io_outs_left[40] ;
 wire \_ces_3_1_io_outs_left[41] ;
 wire \_ces_3_1_io_outs_left[42] ;
 wire \_ces_3_1_io_outs_left[43] ;
 wire \_ces_3_1_io_outs_left[44] ;
 wire \_ces_3_1_io_outs_left[45] ;
 wire \_ces_3_1_io_outs_left[46] ;
 wire \_ces_3_1_io_outs_left[47] ;
 wire \_ces_3_1_io_outs_left[48] ;
 wire \_ces_3_1_io_outs_left[49] ;
 wire \_ces_3_1_io_outs_left[4] ;
 wire \_ces_3_1_io_outs_left[50] ;
 wire \_ces_3_1_io_outs_left[51] ;
 wire \_ces_3_1_io_outs_left[52] ;
 wire \_ces_3_1_io_outs_left[53] ;
 wire \_ces_3_1_io_outs_left[54] ;
 wire \_ces_3_1_io_outs_left[55] ;
 wire \_ces_3_1_io_outs_left[56] ;
 wire \_ces_3_1_io_outs_left[57] ;
 wire \_ces_3_1_io_outs_left[58] ;
 wire \_ces_3_1_io_outs_left[59] ;
 wire \_ces_3_1_io_outs_left[5] ;
 wire \_ces_3_1_io_outs_left[60] ;
 wire \_ces_3_1_io_outs_left[61] ;
 wire \_ces_3_1_io_outs_left[62] ;
 wire \_ces_3_1_io_outs_left[63] ;
 wire \_ces_3_1_io_outs_left[6] ;
 wire \_ces_3_1_io_outs_left[7] ;
 wire \_ces_3_1_io_outs_left[8] ;
 wire \_ces_3_1_io_outs_left[9] ;
 wire \_ces_3_1_io_outs_right[0] ;
 wire \_ces_3_1_io_outs_right[10] ;
 wire \_ces_3_1_io_outs_right[11] ;
 wire \_ces_3_1_io_outs_right[12] ;
 wire \_ces_3_1_io_outs_right[13] ;
 wire \_ces_3_1_io_outs_right[14] ;
 wire \_ces_3_1_io_outs_right[15] ;
 wire \_ces_3_1_io_outs_right[16] ;
 wire \_ces_3_1_io_outs_right[17] ;
 wire \_ces_3_1_io_outs_right[18] ;
 wire \_ces_3_1_io_outs_right[19] ;
 wire \_ces_3_1_io_outs_right[1] ;
 wire \_ces_3_1_io_outs_right[20] ;
 wire \_ces_3_1_io_outs_right[21] ;
 wire \_ces_3_1_io_outs_right[22] ;
 wire \_ces_3_1_io_outs_right[23] ;
 wire \_ces_3_1_io_outs_right[24] ;
 wire \_ces_3_1_io_outs_right[25] ;
 wire \_ces_3_1_io_outs_right[26] ;
 wire \_ces_3_1_io_outs_right[27] ;
 wire \_ces_3_1_io_outs_right[28] ;
 wire \_ces_3_1_io_outs_right[29] ;
 wire \_ces_3_1_io_outs_right[2] ;
 wire \_ces_3_1_io_outs_right[30] ;
 wire \_ces_3_1_io_outs_right[31] ;
 wire \_ces_3_1_io_outs_right[32] ;
 wire \_ces_3_1_io_outs_right[33] ;
 wire \_ces_3_1_io_outs_right[34] ;
 wire \_ces_3_1_io_outs_right[35] ;
 wire \_ces_3_1_io_outs_right[36] ;
 wire \_ces_3_1_io_outs_right[37] ;
 wire \_ces_3_1_io_outs_right[38] ;
 wire \_ces_3_1_io_outs_right[39] ;
 wire \_ces_3_1_io_outs_right[3] ;
 wire \_ces_3_1_io_outs_right[40] ;
 wire \_ces_3_1_io_outs_right[41] ;
 wire \_ces_3_1_io_outs_right[42] ;
 wire \_ces_3_1_io_outs_right[43] ;
 wire \_ces_3_1_io_outs_right[44] ;
 wire \_ces_3_1_io_outs_right[45] ;
 wire \_ces_3_1_io_outs_right[46] ;
 wire \_ces_3_1_io_outs_right[47] ;
 wire \_ces_3_1_io_outs_right[48] ;
 wire \_ces_3_1_io_outs_right[49] ;
 wire \_ces_3_1_io_outs_right[4] ;
 wire \_ces_3_1_io_outs_right[50] ;
 wire \_ces_3_1_io_outs_right[51] ;
 wire \_ces_3_1_io_outs_right[52] ;
 wire \_ces_3_1_io_outs_right[53] ;
 wire \_ces_3_1_io_outs_right[54] ;
 wire \_ces_3_1_io_outs_right[55] ;
 wire \_ces_3_1_io_outs_right[56] ;
 wire \_ces_3_1_io_outs_right[57] ;
 wire \_ces_3_1_io_outs_right[58] ;
 wire \_ces_3_1_io_outs_right[59] ;
 wire \_ces_3_1_io_outs_right[5] ;
 wire \_ces_3_1_io_outs_right[60] ;
 wire \_ces_3_1_io_outs_right[61] ;
 wire \_ces_3_1_io_outs_right[62] ;
 wire \_ces_3_1_io_outs_right[63] ;
 wire \_ces_3_1_io_outs_right[6] ;
 wire \_ces_3_1_io_outs_right[7] ;
 wire \_ces_3_1_io_outs_right[8] ;
 wire \_ces_3_1_io_outs_right[9] ;
 wire _ces_3_2_io_lsbOuts_1;
 wire _ces_3_2_io_lsbOuts_2;
 wire _ces_3_2_io_lsbOuts_3;
 wire \_ces_3_2_io_outs_down[0] ;
 wire \_ces_3_2_io_outs_down[10] ;
 wire \_ces_3_2_io_outs_down[11] ;
 wire \_ces_3_2_io_outs_down[12] ;
 wire \_ces_3_2_io_outs_down[13] ;
 wire \_ces_3_2_io_outs_down[14] ;
 wire \_ces_3_2_io_outs_down[15] ;
 wire \_ces_3_2_io_outs_down[16] ;
 wire \_ces_3_2_io_outs_down[17] ;
 wire \_ces_3_2_io_outs_down[18] ;
 wire \_ces_3_2_io_outs_down[19] ;
 wire \_ces_3_2_io_outs_down[1] ;
 wire \_ces_3_2_io_outs_down[20] ;
 wire \_ces_3_2_io_outs_down[21] ;
 wire \_ces_3_2_io_outs_down[22] ;
 wire \_ces_3_2_io_outs_down[23] ;
 wire \_ces_3_2_io_outs_down[24] ;
 wire \_ces_3_2_io_outs_down[25] ;
 wire \_ces_3_2_io_outs_down[26] ;
 wire \_ces_3_2_io_outs_down[27] ;
 wire \_ces_3_2_io_outs_down[28] ;
 wire \_ces_3_2_io_outs_down[29] ;
 wire \_ces_3_2_io_outs_down[2] ;
 wire \_ces_3_2_io_outs_down[30] ;
 wire \_ces_3_2_io_outs_down[31] ;
 wire \_ces_3_2_io_outs_down[32] ;
 wire \_ces_3_2_io_outs_down[33] ;
 wire \_ces_3_2_io_outs_down[34] ;
 wire \_ces_3_2_io_outs_down[35] ;
 wire \_ces_3_2_io_outs_down[36] ;
 wire \_ces_3_2_io_outs_down[37] ;
 wire \_ces_3_2_io_outs_down[38] ;
 wire \_ces_3_2_io_outs_down[39] ;
 wire \_ces_3_2_io_outs_down[3] ;
 wire \_ces_3_2_io_outs_down[40] ;
 wire \_ces_3_2_io_outs_down[41] ;
 wire \_ces_3_2_io_outs_down[42] ;
 wire \_ces_3_2_io_outs_down[43] ;
 wire \_ces_3_2_io_outs_down[44] ;
 wire \_ces_3_2_io_outs_down[45] ;
 wire \_ces_3_2_io_outs_down[46] ;
 wire \_ces_3_2_io_outs_down[47] ;
 wire \_ces_3_2_io_outs_down[48] ;
 wire \_ces_3_2_io_outs_down[49] ;
 wire \_ces_3_2_io_outs_down[4] ;
 wire \_ces_3_2_io_outs_down[50] ;
 wire \_ces_3_2_io_outs_down[51] ;
 wire \_ces_3_2_io_outs_down[52] ;
 wire \_ces_3_2_io_outs_down[53] ;
 wire \_ces_3_2_io_outs_down[54] ;
 wire \_ces_3_2_io_outs_down[55] ;
 wire \_ces_3_2_io_outs_down[56] ;
 wire \_ces_3_2_io_outs_down[57] ;
 wire \_ces_3_2_io_outs_down[58] ;
 wire \_ces_3_2_io_outs_down[59] ;
 wire \_ces_3_2_io_outs_down[5] ;
 wire \_ces_3_2_io_outs_down[60] ;
 wire \_ces_3_2_io_outs_down[61] ;
 wire \_ces_3_2_io_outs_down[62] ;
 wire \_ces_3_2_io_outs_down[63] ;
 wire \_ces_3_2_io_outs_down[6] ;
 wire \_ces_3_2_io_outs_down[7] ;
 wire \_ces_3_2_io_outs_down[8] ;
 wire \_ces_3_2_io_outs_down[9] ;
 wire \_ces_3_2_io_outs_left[0] ;
 wire \_ces_3_2_io_outs_left[10] ;
 wire \_ces_3_2_io_outs_left[11] ;
 wire \_ces_3_2_io_outs_left[12] ;
 wire \_ces_3_2_io_outs_left[13] ;
 wire \_ces_3_2_io_outs_left[14] ;
 wire \_ces_3_2_io_outs_left[15] ;
 wire \_ces_3_2_io_outs_left[16] ;
 wire \_ces_3_2_io_outs_left[17] ;
 wire \_ces_3_2_io_outs_left[18] ;
 wire \_ces_3_2_io_outs_left[19] ;
 wire \_ces_3_2_io_outs_left[1] ;
 wire \_ces_3_2_io_outs_left[20] ;
 wire \_ces_3_2_io_outs_left[21] ;
 wire \_ces_3_2_io_outs_left[22] ;
 wire \_ces_3_2_io_outs_left[23] ;
 wire \_ces_3_2_io_outs_left[24] ;
 wire \_ces_3_2_io_outs_left[25] ;
 wire \_ces_3_2_io_outs_left[26] ;
 wire \_ces_3_2_io_outs_left[27] ;
 wire \_ces_3_2_io_outs_left[28] ;
 wire \_ces_3_2_io_outs_left[29] ;
 wire \_ces_3_2_io_outs_left[2] ;
 wire \_ces_3_2_io_outs_left[30] ;
 wire \_ces_3_2_io_outs_left[31] ;
 wire \_ces_3_2_io_outs_left[32] ;
 wire \_ces_3_2_io_outs_left[33] ;
 wire \_ces_3_2_io_outs_left[34] ;
 wire \_ces_3_2_io_outs_left[35] ;
 wire \_ces_3_2_io_outs_left[36] ;
 wire \_ces_3_2_io_outs_left[37] ;
 wire \_ces_3_2_io_outs_left[38] ;
 wire \_ces_3_2_io_outs_left[39] ;
 wire \_ces_3_2_io_outs_left[3] ;
 wire \_ces_3_2_io_outs_left[40] ;
 wire \_ces_3_2_io_outs_left[41] ;
 wire \_ces_3_2_io_outs_left[42] ;
 wire \_ces_3_2_io_outs_left[43] ;
 wire \_ces_3_2_io_outs_left[44] ;
 wire \_ces_3_2_io_outs_left[45] ;
 wire \_ces_3_2_io_outs_left[46] ;
 wire \_ces_3_2_io_outs_left[47] ;
 wire \_ces_3_2_io_outs_left[48] ;
 wire \_ces_3_2_io_outs_left[49] ;
 wire \_ces_3_2_io_outs_left[4] ;
 wire \_ces_3_2_io_outs_left[50] ;
 wire \_ces_3_2_io_outs_left[51] ;
 wire \_ces_3_2_io_outs_left[52] ;
 wire \_ces_3_2_io_outs_left[53] ;
 wire \_ces_3_2_io_outs_left[54] ;
 wire \_ces_3_2_io_outs_left[55] ;
 wire \_ces_3_2_io_outs_left[56] ;
 wire \_ces_3_2_io_outs_left[57] ;
 wire \_ces_3_2_io_outs_left[58] ;
 wire \_ces_3_2_io_outs_left[59] ;
 wire \_ces_3_2_io_outs_left[5] ;
 wire \_ces_3_2_io_outs_left[60] ;
 wire \_ces_3_2_io_outs_left[61] ;
 wire \_ces_3_2_io_outs_left[62] ;
 wire \_ces_3_2_io_outs_left[63] ;
 wire \_ces_3_2_io_outs_left[6] ;
 wire \_ces_3_2_io_outs_left[7] ;
 wire \_ces_3_2_io_outs_left[8] ;
 wire \_ces_3_2_io_outs_left[9] ;
 wire \_ces_3_2_io_outs_right[0] ;
 wire \_ces_3_2_io_outs_right[10] ;
 wire \_ces_3_2_io_outs_right[11] ;
 wire \_ces_3_2_io_outs_right[12] ;
 wire \_ces_3_2_io_outs_right[13] ;
 wire \_ces_3_2_io_outs_right[14] ;
 wire \_ces_3_2_io_outs_right[15] ;
 wire \_ces_3_2_io_outs_right[16] ;
 wire \_ces_3_2_io_outs_right[17] ;
 wire \_ces_3_2_io_outs_right[18] ;
 wire \_ces_3_2_io_outs_right[19] ;
 wire \_ces_3_2_io_outs_right[1] ;
 wire \_ces_3_2_io_outs_right[20] ;
 wire \_ces_3_2_io_outs_right[21] ;
 wire \_ces_3_2_io_outs_right[22] ;
 wire \_ces_3_2_io_outs_right[23] ;
 wire \_ces_3_2_io_outs_right[24] ;
 wire \_ces_3_2_io_outs_right[25] ;
 wire \_ces_3_2_io_outs_right[26] ;
 wire \_ces_3_2_io_outs_right[27] ;
 wire \_ces_3_2_io_outs_right[28] ;
 wire \_ces_3_2_io_outs_right[29] ;
 wire \_ces_3_2_io_outs_right[2] ;
 wire \_ces_3_2_io_outs_right[30] ;
 wire \_ces_3_2_io_outs_right[31] ;
 wire \_ces_3_2_io_outs_right[32] ;
 wire \_ces_3_2_io_outs_right[33] ;
 wire \_ces_3_2_io_outs_right[34] ;
 wire \_ces_3_2_io_outs_right[35] ;
 wire \_ces_3_2_io_outs_right[36] ;
 wire \_ces_3_2_io_outs_right[37] ;
 wire \_ces_3_2_io_outs_right[38] ;
 wire \_ces_3_2_io_outs_right[39] ;
 wire \_ces_3_2_io_outs_right[3] ;
 wire \_ces_3_2_io_outs_right[40] ;
 wire \_ces_3_2_io_outs_right[41] ;
 wire \_ces_3_2_io_outs_right[42] ;
 wire \_ces_3_2_io_outs_right[43] ;
 wire \_ces_3_2_io_outs_right[44] ;
 wire \_ces_3_2_io_outs_right[45] ;
 wire \_ces_3_2_io_outs_right[46] ;
 wire \_ces_3_2_io_outs_right[47] ;
 wire \_ces_3_2_io_outs_right[48] ;
 wire \_ces_3_2_io_outs_right[49] ;
 wire \_ces_3_2_io_outs_right[4] ;
 wire \_ces_3_2_io_outs_right[50] ;
 wire \_ces_3_2_io_outs_right[51] ;
 wire \_ces_3_2_io_outs_right[52] ;
 wire \_ces_3_2_io_outs_right[53] ;
 wire \_ces_3_2_io_outs_right[54] ;
 wire \_ces_3_2_io_outs_right[55] ;
 wire \_ces_3_2_io_outs_right[56] ;
 wire \_ces_3_2_io_outs_right[57] ;
 wire \_ces_3_2_io_outs_right[58] ;
 wire \_ces_3_2_io_outs_right[59] ;
 wire \_ces_3_2_io_outs_right[5] ;
 wire \_ces_3_2_io_outs_right[60] ;
 wire \_ces_3_2_io_outs_right[61] ;
 wire \_ces_3_2_io_outs_right[62] ;
 wire \_ces_3_2_io_outs_right[63] ;
 wire \_ces_3_2_io_outs_right[6] ;
 wire \_ces_3_2_io_outs_right[7] ;
 wire \_ces_3_2_io_outs_right[8] ;
 wire \_ces_3_2_io_outs_right[9] ;
 wire _ces_3_3_io_lsbOuts_0;
 wire _ces_3_3_io_lsbOuts_1;
 wire _ces_3_3_io_lsbOuts_2;
 wire _ces_3_3_io_lsbOuts_3;
 wire \_ces_3_3_io_outs_down[0] ;
 wire \_ces_3_3_io_outs_down[10] ;
 wire \_ces_3_3_io_outs_down[11] ;
 wire \_ces_3_3_io_outs_down[12] ;
 wire \_ces_3_3_io_outs_down[13] ;
 wire \_ces_3_3_io_outs_down[14] ;
 wire \_ces_3_3_io_outs_down[15] ;
 wire \_ces_3_3_io_outs_down[16] ;
 wire \_ces_3_3_io_outs_down[17] ;
 wire \_ces_3_3_io_outs_down[18] ;
 wire \_ces_3_3_io_outs_down[19] ;
 wire \_ces_3_3_io_outs_down[1] ;
 wire \_ces_3_3_io_outs_down[20] ;
 wire \_ces_3_3_io_outs_down[21] ;
 wire \_ces_3_3_io_outs_down[22] ;
 wire \_ces_3_3_io_outs_down[23] ;
 wire \_ces_3_3_io_outs_down[24] ;
 wire \_ces_3_3_io_outs_down[25] ;
 wire \_ces_3_3_io_outs_down[26] ;
 wire \_ces_3_3_io_outs_down[27] ;
 wire \_ces_3_3_io_outs_down[28] ;
 wire \_ces_3_3_io_outs_down[29] ;
 wire \_ces_3_3_io_outs_down[2] ;
 wire \_ces_3_3_io_outs_down[30] ;
 wire \_ces_3_3_io_outs_down[31] ;
 wire \_ces_3_3_io_outs_down[32] ;
 wire \_ces_3_3_io_outs_down[33] ;
 wire \_ces_3_3_io_outs_down[34] ;
 wire \_ces_3_3_io_outs_down[35] ;
 wire \_ces_3_3_io_outs_down[36] ;
 wire \_ces_3_3_io_outs_down[37] ;
 wire \_ces_3_3_io_outs_down[38] ;
 wire \_ces_3_3_io_outs_down[39] ;
 wire \_ces_3_3_io_outs_down[3] ;
 wire \_ces_3_3_io_outs_down[40] ;
 wire \_ces_3_3_io_outs_down[41] ;
 wire \_ces_3_3_io_outs_down[42] ;
 wire \_ces_3_3_io_outs_down[43] ;
 wire \_ces_3_3_io_outs_down[44] ;
 wire \_ces_3_3_io_outs_down[45] ;
 wire \_ces_3_3_io_outs_down[46] ;
 wire \_ces_3_3_io_outs_down[47] ;
 wire \_ces_3_3_io_outs_down[48] ;
 wire \_ces_3_3_io_outs_down[49] ;
 wire \_ces_3_3_io_outs_down[4] ;
 wire \_ces_3_3_io_outs_down[50] ;
 wire \_ces_3_3_io_outs_down[51] ;
 wire \_ces_3_3_io_outs_down[52] ;
 wire \_ces_3_3_io_outs_down[53] ;
 wire \_ces_3_3_io_outs_down[54] ;
 wire \_ces_3_3_io_outs_down[55] ;
 wire \_ces_3_3_io_outs_down[56] ;
 wire \_ces_3_3_io_outs_down[57] ;
 wire \_ces_3_3_io_outs_down[58] ;
 wire \_ces_3_3_io_outs_down[59] ;
 wire \_ces_3_3_io_outs_down[5] ;
 wire \_ces_3_3_io_outs_down[60] ;
 wire \_ces_3_3_io_outs_down[61] ;
 wire \_ces_3_3_io_outs_down[62] ;
 wire \_ces_3_3_io_outs_down[63] ;
 wire \_ces_3_3_io_outs_down[6] ;
 wire \_ces_3_3_io_outs_down[7] ;
 wire \_ces_3_3_io_outs_down[8] ;
 wire \_ces_3_3_io_outs_down[9] ;
 wire \_ces_3_3_io_outs_left[0] ;
 wire \_ces_3_3_io_outs_left[10] ;
 wire \_ces_3_3_io_outs_left[11] ;
 wire \_ces_3_3_io_outs_left[12] ;
 wire \_ces_3_3_io_outs_left[13] ;
 wire \_ces_3_3_io_outs_left[14] ;
 wire \_ces_3_3_io_outs_left[15] ;
 wire \_ces_3_3_io_outs_left[16] ;
 wire \_ces_3_3_io_outs_left[17] ;
 wire \_ces_3_3_io_outs_left[18] ;
 wire \_ces_3_3_io_outs_left[19] ;
 wire \_ces_3_3_io_outs_left[1] ;
 wire \_ces_3_3_io_outs_left[20] ;
 wire \_ces_3_3_io_outs_left[21] ;
 wire \_ces_3_3_io_outs_left[22] ;
 wire \_ces_3_3_io_outs_left[23] ;
 wire \_ces_3_3_io_outs_left[24] ;
 wire \_ces_3_3_io_outs_left[25] ;
 wire \_ces_3_3_io_outs_left[26] ;
 wire \_ces_3_3_io_outs_left[27] ;
 wire \_ces_3_3_io_outs_left[28] ;
 wire \_ces_3_3_io_outs_left[29] ;
 wire \_ces_3_3_io_outs_left[2] ;
 wire \_ces_3_3_io_outs_left[30] ;
 wire \_ces_3_3_io_outs_left[31] ;
 wire \_ces_3_3_io_outs_left[32] ;
 wire \_ces_3_3_io_outs_left[33] ;
 wire \_ces_3_3_io_outs_left[34] ;
 wire \_ces_3_3_io_outs_left[35] ;
 wire \_ces_3_3_io_outs_left[36] ;
 wire \_ces_3_3_io_outs_left[37] ;
 wire \_ces_3_3_io_outs_left[38] ;
 wire \_ces_3_3_io_outs_left[39] ;
 wire \_ces_3_3_io_outs_left[3] ;
 wire \_ces_3_3_io_outs_left[40] ;
 wire \_ces_3_3_io_outs_left[41] ;
 wire \_ces_3_3_io_outs_left[42] ;
 wire \_ces_3_3_io_outs_left[43] ;
 wire \_ces_3_3_io_outs_left[44] ;
 wire \_ces_3_3_io_outs_left[45] ;
 wire \_ces_3_3_io_outs_left[46] ;
 wire \_ces_3_3_io_outs_left[47] ;
 wire \_ces_3_3_io_outs_left[48] ;
 wire \_ces_3_3_io_outs_left[49] ;
 wire \_ces_3_3_io_outs_left[4] ;
 wire \_ces_3_3_io_outs_left[50] ;
 wire \_ces_3_3_io_outs_left[51] ;
 wire \_ces_3_3_io_outs_left[52] ;
 wire \_ces_3_3_io_outs_left[53] ;
 wire \_ces_3_3_io_outs_left[54] ;
 wire \_ces_3_3_io_outs_left[55] ;
 wire \_ces_3_3_io_outs_left[56] ;
 wire \_ces_3_3_io_outs_left[57] ;
 wire \_ces_3_3_io_outs_left[58] ;
 wire \_ces_3_3_io_outs_left[59] ;
 wire \_ces_3_3_io_outs_left[5] ;
 wire \_ces_3_3_io_outs_left[60] ;
 wire \_ces_3_3_io_outs_left[61] ;
 wire \_ces_3_3_io_outs_left[62] ;
 wire \_ces_3_3_io_outs_left[63] ;
 wire \_ces_3_3_io_outs_left[6] ;
 wire \_ces_3_3_io_outs_left[7] ;
 wire \_ces_3_3_io_outs_left[8] ;
 wire \_ces_3_3_io_outs_left[9] ;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire clock_regs;
 wire clknet_leaf_0_clock;
 wire clknet_leaf_1_clock;
 wire clknet_leaf_2_clock;
 wire clknet_leaf_3_clock;
 wire clknet_0_clock;
 wire clknet_1_0__leaf_clock;
 wire clknet_1_1__leaf_clock;
 wire clknet_0_clock_regs;
 wire clknet_1_0__leaf_clock_regs;
 wire clknet_1_1__leaf_clock_regs;
 wire delaynet_0_clock;
 wire delaynet_1_clock;
 wire delaynet_2_clock;
 wire delaynet_3_clock;
 wire delaynet_4_clock;
 wire delaynet_5_clock;

 BUFx24_ASAP7_75t_R delaybuf_5_clock (.A(delaynet_4_clock),
    .Y(delaynet_5_clock));
 BUFx24_ASAP7_75t_R delaybuf_4_clock (.A(delaynet_3_clock),
    .Y(delaynet_4_clock));
 BUFx24_ASAP7_75t_R delaybuf_3_clock (.A(delaynet_2_clock),
    .Y(delaynet_3_clock));
 BUFx24_ASAP7_75t_R delaybuf_2_clock (.A(delaynet_1_clock),
    .Y(delaynet_2_clock));
 BUFx24_ASAP7_75t_R delaybuf_1_clock (.A(delaynet_0_clock),
    .Y(delaynet_1_clock));
 BUFx24_ASAP7_75t_R delaybuf_0_clock (.A(clock),
    .Y(delaynet_0_clock));
 BUFx24_ASAP7_75t_R clkbuf_1_1__f_clock_regs (.A(clknet_0_clock_regs),
    .Y(clknet_1_1__leaf_clock_regs));
 BUFx24_ASAP7_75t_R clkbuf_1_0__f_clock_regs (.A(clknet_0_clock_regs),
    .Y(clknet_1_0__leaf_clock_regs));
 BUFx24_ASAP7_75t_R clkbuf_0_clock_regs (.A(clock_regs),
    .Y(clknet_0_clock_regs));
 BUFx24_ASAP7_75t_R clkbuf_1_1__f_clock (.A(clknet_0_clock),
    .Y(clknet_1_1__leaf_clock));
 BUFx24_ASAP7_75t_R clkbuf_1_0__f_clock (.A(clknet_0_clock),
    .Y(clknet_1_0__leaf_clock));
 BUFx24_ASAP7_75t_R clkbuf_0_clock (.A(clock),
    .Y(clknet_0_clock));
 BUFx24_ASAP7_75t_R clkbuf_leaf_3_clock (.A(clknet_1_0__leaf_clock),
    .Y(clknet_leaf_3_clock));
 BUFx24_ASAP7_75t_R clkbuf_leaf_2_clock (.A(clknet_1_0__leaf_clock),
    .Y(clknet_leaf_2_clock));
 BUFx24_ASAP7_75t_R clkbuf_leaf_1_clock (.A(clknet_1_1__leaf_clock),
    .Y(clknet_leaf_1_clock));
 BUFx24_ASAP7_75t_R clkbuf_leaf_0_clock (.A(clknet_1_1__leaf_clock),
    .Y(clknet_leaf_0_clock));
 BUFx24_ASAP7_75t_R clkbuf_regs_0_clock (.A(delaynet_5_clock),
    .Y(clock_regs));
 BUFx2_ASAP7_75t_R output2076 (.A(net2075),
    .Y(io_outs_up_3[9]));
 BUFx2_ASAP7_75t_R output2075 (.A(net2074),
    .Y(io_outs_up_3[8]));
 BUFx2_ASAP7_75t_R output2074 (.A(net2073),
    .Y(io_outs_up_3[7]));
 BUFx2_ASAP7_75t_R output2073 (.A(net2072),
    .Y(io_outs_up_3[6]));
 BUFx2_ASAP7_75t_R output2072 (.A(net2071),
    .Y(io_outs_up_3[63]));
 BUFx2_ASAP7_75t_R output2071 (.A(net2070),
    .Y(io_outs_up_3[62]));
 BUFx2_ASAP7_75t_R output2070 (.A(net2069),
    .Y(io_outs_up_3[61]));
 BUFx2_ASAP7_75t_R output2069 (.A(net2068),
    .Y(io_outs_up_3[60]));
 BUFx2_ASAP7_75t_R output2068 (.A(net2067),
    .Y(io_outs_up_3[5]));
 BUFx2_ASAP7_75t_R output2067 (.A(net2066),
    .Y(io_outs_up_3[59]));
 BUFx2_ASAP7_75t_R output2066 (.A(net2065),
    .Y(io_outs_up_3[58]));
 BUFx2_ASAP7_75t_R output2065 (.A(net2064),
    .Y(io_outs_up_3[57]));
 BUFx2_ASAP7_75t_R output2064 (.A(net2063),
    .Y(io_outs_up_3[56]));
 BUFx2_ASAP7_75t_R output2063 (.A(net2062),
    .Y(io_outs_up_3[55]));
 BUFx2_ASAP7_75t_R output2062 (.A(net2061),
    .Y(io_outs_up_3[54]));
 BUFx2_ASAP7_75t_R output2061 (.A(net2060),
    .Y(io_outs_up_3[53]));
 BUFx2_ASAP7_75t_R output2060 (.A(net2059),
    .Y(io_outs_up_3[52]));
 BUFx2_ASAP7_75t_R output2059 (.A(net2058),
    .Y(io_outs_up_3[51]));
 BUFx2_ASAP7_75t_R output2058 (.A(net2057),
    .Y(io_outs_up_3[50]));
 BUFx2_ASAP7_75t_R output2057 (.A(net2056),
    .Y(io_outs_up_3[4]));
 BUFx2_ASAP7_75t_R output2056 (.A(net2055),
    .Y(io_outs_up_3[49]));
 BUFx2_ASAP7_75t_R output2055 (.A(net2054),
    .Y(io_outs_up_3[48]));
 BUFx2_ASAP7_75t_R output2054 (.A(net2053),
    .Y(io_outs_up_3[47]));
 BUFx2_ASAP7_75t_R output2053 (.A(net2052),
    .Y(io_outs_up_3[46]));
 BUFx2_ASAP7_75t_R output2052 (.A(net2051),
    .Y(io_outs_up_3[45]));
 BUFx2_ASAP7_75t_R output2051 (.A(net2050),
    .Y(io_outs_up_3[44]));
 BUFx2_ASAP7_75t_R output2050 (.A(net2049),
    .Y(io_outs_up_3[43]));
 BUFx2_ASAP7_75t_R output2049 (.A(net2048),
    .Y(io_outs_up_3[42]));
 BUFx2_ASAP7_75t_R output2048 (.A(net2047),
    .Y(io_outs_up_3[41]));
 BUFx2_ASAP7_75t_R output2047 (.A(net2046),
    .Y(io_outs_up_3[40]));
 BUFx2_ASAP7_75t_R output2046 (.A(net2045),
    .Y(io_outs_up_3[3]));
 BUFx2_ASAP7_75t_R output2045 (.A(net2044),
    .Y(io_outs_up_3[39]));
 BUFx2_ASAP7_75t_R output2044 (.A(net2043),
    .Y(io_outs_up_3[38]));
 BUFx2_ASAP7_75t_R output2043 (.A(net2042),
    .Y(io_outs_up_3[37]));
 BUFx2_ASAP7_75t_R output2042 (.A(net2041),
    .Y(io_outs_up_3[36]));
 BUFx2_ASAP7_75t_R output2041 (.A(net2040),
    .Y(io_outs_up_3[35]));
 BUFx2_ASAP7_75t_R output2040 (.A(net2039),
    .Y(io_outs_up_3[34]));
 BUFx2_ASAP7_75t_R output2039 (.A(net2038),
    .Y(io_outs_up_3[33]));
 BUFx2_ASAP7_75t_R output2038 (.A(net2037),
    .Y(io_outs_up_3[32]));
 BUFx2_ASAP7_75t_R output2037 (.A(net2036),
    .Y(io_outs_up_3[31]));
 BUFx2_ASAP7_75t_R output2036 (.A(net2035),
    .Y(io_outs_up_3[30]));
 BUFx2_ASAP7_75t_R output2035 (.A(net2034),
    .Y(io_outs_up_3[2]));
 BUFx2_ASAP7_75t_R output2034 (.A(net2033),
    .Y(io_outs_up_3[29]));
 BUFx2_ASAP7_75t_R output2033 (.A(net2032),
    .Y(io_outs_up_3[28]));
 BUFx2_ASAP7_75t_R output2032 (.A(net2031),
    .Y(io_outs_up_3[27]));
 BUFx2_ASAP7_75t_R output2031 (.A(net2030),
    .Y(io_outs_up_3[26]));
 BUFx2_ASAP7_75t_R output2030 (.A(net2029),
    .Y(io_outs_up_3[25]));
 BUFx2_ASAP7_75t_R output2029 (.A(net2028),
    .Y(io_outs_up_3[24]));
 BUFx2_ASAP7_75t_R output2028 (.A(net2027),
    .Y(io_outs_up_3[23]));
 BUFx2_ASAP7_75t_R output2027 (.A(net2026),
    .Y(io_outs_up_3[22]));
 BUFx2_ASAP7_75t_R output2026 (.A(net2025),
    .Y(io_outs_up_3[21]));
 BUFx2_ASAP7_75t_R output2025 (.A(net2024),
    .Y(io_outs_up_3[20]));
 BUFx2_ASAP7_75t_R output2024 (.A(net2023),
    .Y(io_outs_up_3[1]));
 BUFx2_ASAP7_75t_R output2023 (.A(net2022),
    .Y(io_outs_up_3[19]));
 BUFx2_ASAP7_75t_R output2022 (.A(net2021),
    .Y(io_outs_up_3[18]));
 BUFx2_ASAP7_75t_R output2021 (.A(net2020),
    .Y(io_outs_up_3[17]));
 BUFx2_ASAP7_75t_R output2020 (.A(net2019),
    .Y(io_outs_up_3[16]));
 BUFx2_ASAP7_75t_R output2019 (.A(net2018),
    .Y(io_outs_up_3[15]));
 BUFx2_ASAP7_75t_R output2018 (.A(net2017),
    .Y(io_outs_up_3[14]));
 BUFx2_ASAP7_75t_R output2017 (.A(net2016),
    .Y(io_outs_up_3[13]));
 BUFx2_ASAP7_75t_R output2016 (.A(net2015),
    .Y(io_outs_up_3[12]));
 BUFx2_ASAP7_75t_R output2015 (.A(net2014),
    .Y(io_outs_up_3[11]));
 BUFx2_ASAP7_75t_R output2014 (.A(net2013),
    .Y(io_outs_up_3[10]));
 BUFx2_ASAP7_75t_R output2013 (.A(net2012),
    .Y(io_outs_up_3[0]));
 BUFx2_ASAP7_75t_R output2012 (.A(net2011),
    .Y(io_outs_up_2[9]));
 BUFx2_ASAP7_75t_R output2011 (.A(net2010),
    .Y(io_outs_up_2[8]));
 BUFx2_ASAP7_75t_R output2010 (.A(net2009),
    .Y(io_outs_up_2[7]));
 BUFx2_ASAP7_75t_R output2009 (.A(net2008),
    .Y(io_outs_up_2[6]));
 BUFx2_ASAP7_75t_R output2008 (.A(net2007),
    .Y(io_outs_up_2[63]));
 BUFx2_ASAP7_75t_R output2007 (.A(net2006),
    .Y(io_outs_up_2[62]));
 BUFx2_ASAP7_75t_R output2006 (.A(net2005),
    .Y(io_outs_up_2[61]));
 BUFx2_ASAP7_75t_R output2005 (.A(net2004),
    .Y(io_outs_up_2[60]));
 BUFx2_ASAP7_75t_R output2004 (.A(net2003),
    .Y(io_outs_up_2[5]));
 BUFx2_ASAP7_75t_R output2003 (.A(net2002),
    .Y(io_outs_up_2[59]));
 BUFx2_ASAP7_75t_R output2002 (.A(net2001),
    .Y(io_outs_up_2[58]));
 BUFx2_ASAP7_75t_R output2001 (.A(net2000),
    .Y(io_outs_up_2[57]));
 BUFx2_ASAP7_75t_R output2000 (.A(net1999),
    .Y(io_outs_up_2[56]));
 BUFx2_ASAP7_75t_R output1999 (.A(net1998),
    .Y(io_outs_up_2[55]));
 BUFx2_ASAP7_75t_R output1998 (.A(net1997),
    .Y(io_outs_up_2[54]));
 BUFx2_ASAP7_75t_R output1997 (.A(net1996),
    .Y(io_outs_up_2[53]));
 BUFx2_ASAP7_75t_R output1996 (.A(net1995),
    .Y(io_outs_up_2[52]));
 BUFx2_ASAP7_75t_R output1995 (.A(net1994),
    .Y(io_outs_up_2[51]));
 BUFx2_ASAP7_75t_R output1994 (.A(net1993),
    .Y(io_outs_up_2[50]));
 BUFx2_ASAP7_75t_R output1993 (.A(net1992),
    .Y(io_outs_up_2[4]));
 BUFx2_ASAP7_75t_R output1992 (.A(net1991),
    .Y(io_outs_up_2[49]));
 BUFx2_ASAP7_75t_R output1991 (.A(net1990),
    .Y(io_outs_up_2[48]));
 BUFx2_ASAP7_75t_R output1990 (.A(net1989),
    .Y(io_outs_up_2[47]));
 BUFx2_ASAP7_75t_R output1989 (.A(net1988),
    .Y(io_outs_up_2[46]));
 BUFx2_ASAP7_75t_R output1988 (.A(net1987),
    .Y(io_outs_up_2[45]));
 BUFx2_ASAP7_75t_R output1987 (.A(net1986),
    .Y(io_outs_up_2[44]));
 BUFx2_ASAP7_75t_R output1986 (.A(net1985),
    .Y(io_outs_up_2[43]));
 BUFx2_ASAP7_75t_R output1985 (.A(net1984),
    .Y(io_outs_up_2[42]));
 BUFx2_ASAP7_75t_R output1984 (.A(net1983),
    .Y(io_outs_up_2[41]));
 BUFx2_ASAP7_75t_R output1983 (.A(net1982),
    .Y(io_outs_up_2[40]));
 BUFx2_ASAP7_75t_R output1982 (.A(net1981),
    .Y(io_outs_up_2[3]));
 BUFx2_ASAP7_75t_R output1981 (.A(net1980),
    .Y(io_outs_up_2[39]));
 BUFx2_ASAP7_75t_R output1980 (.A(net1979),
    .Y(io_outs_up_2[38]));
 BUFx2_ASAP7_75t_R output1979 (.A(net1978),
    .Y(io_outs_up_2[37]));
 BUFx2_ASAP7_75t_R output1978 (.A(net1977),
    .Y(io_outs_up_2[36]));
 BUFx2_ASAP7_75t_R output1977 (.A(net1976),
    .Y(io_outs_up_2[35]));
 BUFx2_ASAP7_75t_R output1976 (.A(net1975),
    .Y(io_outs_up_2[34]));
 BUFx2_ASAP7_75t_R output1975 (.A(net1974),
    .Y(io_outs_up_2[33]));
 BUFx2_ASAP7_75t_R output1974 (.A(net1973),
    .Y(io_outs_up_2[32]));
 BUFx2_ASAP7_75t_R output1973 (.A(net1972),
    .Y(io_outs_up_2[31]));
 BUFx2_ASAP7_75t_R output1972 (.A(net1971),
    .Y(io_outs_up_2[30]));
 BUFx2_ASAP7_75t_R output1971 (.A(net1970),
    .Y(io_outs_up_2[2]));
 BUFx2_ASAP7_75t_R output1970 (.A(net1969),
    .Y(io_outs_up_2[29]));
 BUFx2_ASAP7_75t_R output1969 (.A(net1968),
    .Y(io_outs_up_2[28]));
 BUFx2_ASAP7_75t_R output1968 (.A(net1967),
    .Y(io_outs_up_2[27]));
 BUFx2_ASAP7_75t_R output1967 (.A(net1966),
    .Y(io_outs_up_2[26]));
 BUFx2_ASAP7_75t_R output1966 (.A(net1965),
    .Y(io_outs_up_2[25]));
 BUFx2_ASAP7_75t_R output1965 (.A(net1964),
    .Y(io_outs_up_2[24]));
 BUFx2_ASAP7_75t_R output1964 (.A(net1963),
    .Y(io_outs_up_2[23]));
 BUFx2_ASAP7_75t_R output1963 (.A(net1962),
    .Y(io_outs_up_2[22]));
 BUFx2_ASAP7_75t_R output1962 (.A(net1961),
    .Y(io_outs_up_2[21]));
 BUFx2_ASAP7_75t_R output1961 (.A(net1960),
    .Y(io_outs_up_2[20]));
 BUFx2_ASAP7_75t_R output1960 (.A(net1959),
    .Y(io_outs_up_2[1]));
 BUFx2_ASAP7_75t_R output1959 (.A(net1958),
    .Y(io_outs_up_2[19]));
 BUFx2_ASAP7_75t_R output1958 (.A(net1957),
    .Y(io_outs_up_2[18]));
 BUFx2_ASAP7_75t_R output1957 (.A(net1956),
    .Y(io_outs_up_2[17]));
 BUFx2_ASAP7_75t_R output1956 (.A(net1955),
    .Y(io_outs_up_2[16]));
 BUFx2_ASAP7_75t_R output1955 (.A(net1954),
    .Y(io_outs_up_2[15]));
 BUFx2_ASAP7_75t_R output1954 (.A(net1953),
    .Y(io_outs_up_2[14]));
 BUFx2_ASAP7_75t_R output1953 (.A(net1952),
    .Y(io_outs_up_2[13]));
 BUFx2_ASAP7_75t_R output1952 (.A(net1951),
    .Y(io_outs_up_2[12]));
 BUFx2_ASAP7_75t_R output1951 (.A(net1950),
    .Y(io_outs_up_2[11]));
 BUFx2_ASAP7_75t_R output1950 (.A(net1949),
    .Y(io_outs_up_2[10]));
 BUFx2_ASAP7_75t_R output1949 (.A(net1948),
    .Y(io_outs_up_2[0]));
 BUFx2_ASAP7_75t_R output1948 (.A(net1947),
    .Y(io_outs_up_1[9]));
 BUFx2_ASAP7_75t_R output1947 (.A(net1946),
    .Y(io_outs_up_1[8]));
 BUFx2_ASAP7_75t_R output1946 (.A(net1945),
    .Y(io_outs_up_1[7]));
 BUFx2_ASAP7_75t_R output1945 (.A(net1944),
    .Y(io_outs_up_1[6]));
 BUFx2_ASAP7_75t_R output1944 (.A(net1943),
    .Y(io_outs_up_1[63]));
 BUFx2_ASAP7_75t_R output1943 (.A(net1942),
    .Y(io_outs_up_1[62]));
 BUFx2_ASAP7_75t_R output1942 (.A(net1941),
    .Y(io_outs_up_1[61]));
 BUFx2_ASAP7_75t_R output1941 (.A(net1940),
    .Y(io_outs_up_1[60]));
 BUFx2_ASAP7_75t_R output1940 (.A(net1939),
    .Y(io_outs_up_1[5]));
 BUFx2_ASAP7_75t_R output1939 (.A(net1938),
    .Y(io_outs_up_1[59]));
 BUFx2_ASAP7_75t_R output1938 (.A(net1937),
    .Y(io_outs_up_1[58]));
 BUFx2_ASAP7_75t_R output1937 (.A(net1936),
    .Y(io_outs_up_1[57]));
 BUFx2_ASAP7_75t_R output1936 (.A(net1935),
    .Y(io_outs_up_1[56]));
 BUFx2_ASAP7_75t_R output1935 (.A(net1934),
    .Y(io_outs_up_1[55]));
 BUFx2_ASAP7_75t_R output1934 (.A(net1933),
    .Y(io_outs_up_1[54]));
 BUFx2_ASAP7_75t_R output1933 (.A(net1932),
    .Y(io_outs_up_1[53]));
 BUFx2_ASAP7_75t_R output1932 (.A(net1931),
    .Y(io_outs_up_1[52]));
 BUFx2_ASAP7_75t_R output1931 (.A(net1930),
    .Y(io_outs_up_1[51]));
 BUFx2_ASAP7_75t_R output1930 (.A(net1929),
    .Y(io_outs_up_1[50]));
 BUFx2_ASAP7_75t_R output1929 (.A(net1928),
    .Y(io_outs_up_1[4]));
 BUFx2_ASAP7_75t_R output1928 (.A(net1927),
    .Y(io_outs_up_1[49]));
 BUFx2_ASAP7_75t_R output1927 (.A(net1926),
    .Y(io_outs_up_1[48]));
 BUFx2_ASAP7_75t_R output1926 (.A(net1925),
    .Y(io_outs_up_1[47]));
 BUFx2_ASAP7_75t_R output1925 (.A(net1924),
    .Y(io_outs_up_1[46]));
 BUFx2_ASAP7_75t_R output1924 (.A(net1923),
    .Y(io_outs_up_1[45]));
 BUFx2_ASAP7_75t_R output1923 (.A(net1922),
    .Y(io_outs_up_1[44]));
 BUFx2_ASAP7_75t_R output1922 (.A(net1921),
    .Y(io_outs_up_1[43]));
 BUFx2_ASAP7_75t_R output1921 (.A(net1920),
    .Y(io_outs_up_1[42]));
 BUFx2_ASAP7_75t_R output1920 (.A(net1919),
    .Y(io_outs_up_1[41]));
 BUFx2_ASAP7_75t_R output1919 (.A(net1918),
    .Y(io_outs_up_1[40]));
 BUFx2_ASAP7_75t_R output1918 (.A(net1917),
    .Y(io_outs_up_1[3]));
 BUFx2_ASAP7_75t_R output1917 (.A(net1916),
    .Y(io_outs_up_1[39]));
 BUFx2_ASAP7_75t_R output1916 (.A(net1915),
    .Y(io_outs_up_1[38]));
 BUFx2_ASAP7_75t_R output1915 (.A(net1914),
    .Y(io_outs_up_1[37]));
 BUFx2_ASAP7_75t_R output1914 (.A(net1913),
    .Y(io_outs_up_1[36]));
 BUFx2_ASAP7_75t_R output1913 (.A(net1912),
    .Y(io_outs_up_1[35]));
 BUFx2_ASAP7_75t_R output1912 (.A(net1911),
    .Y(io_outs_up_1[34]));
 BUFx2_ASAP7_75t_R output1911 (.A(net1910),
    .Y(io_outs_up_1[33]));
 BUFx2_ASAP7_75t_R output1910 (.A(net1909),
    .Y(io_outs_up_1[32]));
 BUFx2_ASAP7_75t_R output1909 (.A(net1908),
    .Y(io_outs_up_1[31]));
 BUFx2_ASAP7_75t_R output1908 (.A(net1907),
    .Y(io_outs_up_1[30]));
 BUFx2_ASAP7_75t_R output1907 (.A(net1906),
    .Y(io_outs_up_1[2]));
 BUFx2_ASAP7_75t_R output1906 (.A(net1905),
    .Y(io_outs_up_1[29]));
 BUFx2_ASAP7_75t_R output1905 (.A(net1904),
    .Y(io_outs_up_1[28]));
 BUFx2_ASAP7_75t_R output1904 (.A(net1903),
    .Y(io_outs_up_1[27]));
 BUFx2_ASAP7_75t_R output1903 (.A(net1902),
    .Y(io_outs_up_1[26]));
 BUFx2_ASAP7_75t_R output1902 (.A(net1901),
    .Y(io_outs_up_1[25]));
 BUFx2_ASAP7_75t_R output1901 (.A(net1900),
    .Y(io_outs_up_1[24]));
 BUFx2_ASAP7_75t_R output1900 (.A(net1899),
    .Y(io_outs_up_1[23]));
 BUFx2_ASAP7_75t_R output1899 (.A(net1898),
    .Y(io_outs_up_1[22]));
 BUFx2_ASAP7_75t_R output1898 (.A(net1897),
    .Y(io_outs_up_1[21]));
 BUFx2_ASAP7_75t_R output1897 (.A(net1896),
    .Y(io_outs_up_1[20]));
 BUFx2_ASAP7_75t_R output1896 (.A(net1895),
    .Y(io_outs_up_1[1]));
 BUFx2_ASAP7_75t_R output1895 (.A(net1894),
    .Y(io_outs_up_1[19]));
 BUFx2_ASAP7_75t_R output1894 (.A(net1893),
    .Y(io_outs_up_1[18]));
 BUFx2_ASAP7_75t_R output1893 (.A(net1892),
    .Y(io_outs_up_1[17]));
 BUFx2_ASAP7_75t_R output1892 (.A(net1891),
    .Y(io_outs_up_1[16]));
 BUFx2_ASAP7_75t_R output1891 (.A(net1890),
    .Y(io_outs_up_1[15]));
 BUFx2_ASAP7_75t_R output1890 (.A(net1889),
    .Y(io_outs_up_1[14]));
 BUFx2_ASAP7_75t_R output1889 (.A(net1888),
    .Y(io_outs_up_1[13]));
 BUFx2_ASAP7_75t_R output1888 (.A(net1887),
    .Y(io_outs_up_1[12]));
 BUFx2_ASAP7_75t_R output1887 (.A(net1886),
    .Y(io_outs_up_1[11]));
 BUFx2_ASAP7_75t_R output1886 (.A(net1885),
    .Y(io_outs_up_1[10]));
 BUFx2_ASAP7_75t_R output1885 (.A(net1884),
    .Y(io_outs_up_1[0]));
 BUFx2_ASAP7_75t_R output1884 (.A(net1883),
    .Y(io_outs_up_0[9]));
 BUFx2_ASAP7_75t_R output1883 (.A(net1882),
    .Y(io_outs_up_0[8]));
 BUFx2_ASAP7_75t_R output1882 (.A(net1881),
    .Y(io_outs_up_0[7]));
 BUFx2_ASAP7_75t_R output1881 (.A(net1880),
    .Y(io_outs_up_0[6]));
 BUFx2_ASAP7_75t_R output1880 (.A(net1879),
    .Y(io_outs_up_0[63]));
 BUFx2_ASAP7_75t_R output1879 (.A(net1878),
    .Y(io_outs_up_0[62]));
 BUFx2_ASAP7_75t_R output1878 (.A(net1877),
    .Y(io_outs_up_0[61]));
 BUFx2_ASAP7_75t_R output1877 (.A(net1876),
    .Y(io_outs_up_0[60]));
 BUFx2_ASAP7_75t_R output1876 (.A(net1875),
    .Y(io_outs_up_0[5]));
 BUFx2_ASAP7_75t_R output1875 (.A(net1874),
    .Y(io_outs_up_0[59]));
 BUFx2_ASAP7_75t_R output1874 (.A(net1873),
    .Y(io_outs_up_0[58]));
 BUFx2_ASAP7_75t_R output1873 (.A(net1872),
    .Y(io_outs_up_0[57]));
 BUFx2_ASAP7_75t_R output1872 (.A(net1871),
    .Y(io_outs_up_0[56]));
 BUFx2_ASAP7_75t_R output1871 (.A(net1870),
    .Y(io_outs_up_0[55]));
 BUFx2_ASAP7_75t_R output1870 (.A(net1869),
    .Y(io_outs_up_0[54]));
 BUFx2_ASAP7_75t_R output1869 (.A(net1868),
    .Y(io_outs_up_0[53]));
 BUFx2_ASAP7_75t_R output1868 (.A(net1867),
    .Y(io_outs_up_0[52]));
 BUFx2_ASAP7_75t_R output1867 (.A(net1866),
    .Y(io_outs_up_0[51]));
 BUFx2_ASAP7_75t_R output1866 (.A(net1865),
    .Y(io_outs_up_0[50]));
 BUFx2_ASAP7_75t_R output1865 (.A(net1864),
    .Y(io_outs_up_0[4]));
 BUFx2_ASAP7_75t_R output1864 (.A(net1863),
    .Y(io_outs_up_0[49]));
 BUFx2_ASAP7_75t_R output1863 (.A(net1862),
    .Y(io_outs_up_0[48]));
 BUFx2_ASAP7_75t_R output1862 (.A(net1861),
    .Y(io_outs_up_0[47]));
 BUFx2_ASAP7_75t_R output1861 (.A(net1860),
    .Y(io_outs_up_0[46]));
 BUFx2_ASAP7_75t_R output1860 (.A(net1859),
    .Y(io_outs_up_0[45]));
 BUFx2_ASAP7_75t_R output1859 (.A(net1858),
    .Y(io_outs_up_0[44]));
 BUFx2_ASAP7_75t_R output1858 (.A(net1857),
    .Y(io_outs_up_0[43]));
 BUFx2_ASAP7_75t_R output1857 (.A(net1856),
    .Y(io_outs_up_0[42]));
 BUFx2_ASAP7_75t_R output1856 (.A(net1855),
    .Y(io_outs_up_0[41]));
 BUFx2_ASAP7_75t_R output1855 (.A(net1854),
    .Y(io_outs_up_0[40]));
 BUFx2_ASAP7_75t_R output1854 (.A(net1853),
    .Y(io_outs_up_0[3]));
 BUFx2_ASAP7_75t_R output1853 (.A(net1852),
    .Y(io_outs_up_0[39]));
 BUFx2_ASAP7_75t_R output1852 (.A(net1851),
    .Y(io_outs_up_0[38]));
 BUFx2_ASAP7_75t_R output1851 (.A(net1850),
    .Y(io_outs_up_0[37]));
 BUFx2_ASAP7_75t_R output1850 (.A(net1849),
    .Y(io_outs_up_0[36]));
 BUFx2_ASAP7_75t_R output1849 (.A(net1848),
    .Y(io_outs_up_0[35]));
 BUFx2_ASAP7_75t_R output1848 (.A(net1847),
    .Y(io_outs_up_0[34]));
 BUFx2_ASAP7_75t_R output1847 (.A(net1846),
    .Y(io_outs_up_0[33]));
 BUFx2_ASAP7_75t_R output1846 (.A(net1845),
    .Y(io_outs_up_0[32]));
 BUFx2_ASAP7_75t_R output1845 (.A(net1844),
    .Y(io_outs_up_0[31]));
 BUFx2_ASAP7_75t_R output1844 (.A(net1843),
    .Y(io_outs_up_0[30]));
 BUFx2_ASAP7_75t_R output1843 (.A(net1842),
    .Y(io_outs_up_0[2]));
 BUFx2_ASAP7_75t_R output1842 (.A(net1841),
    .Y(io_outs_up_0[29]));
 BUFx2_ASAP7_75t_R output1841 (.A(net1840),
    .Y(io_outs_up_0[28]));
 BUFx2_ASAP7_75t_R output1840 (.A(net1839),
    .Y(io_outs_up_0[27]));
 BUFx2_ASAP7_75t_R output1839 (.A(net1838),
    .Y(io_outs_up_0[26]));
 BUFx2_ASAP7_75t_R output1838 (.A(net1837),
    .Y(io_outs_up_0[25]));
 BUFx2_ASAP7_75t_R output1837 (.A(net1836),
    .Y(io_outs_up_0[24]));
 BUFx2_ASAP7_75t_R output1836 (.A(net1835),
    .Y(io_outs_up_0[23]));
 BUFx2_ASAP7_75t_R output1835 (.A(net1834),
    .Y(io_outs_up_0[22]));
 BUFx2_ASAP7_75t_R output1834 (.A(net1833),
    .Y(io_outs_up_0[21]));
 BUFx2_ASAP7_75t_R output1833 (.A(net1832),
    .Y(io_outs_up_0[20]));
 BUFx2_ASAP7_75t_R output1832 (.A(net1831),
    .Y(io_outs_up_0[1]));
 BUFx2_ASAP7_75t_R output1831 (.A(net1830),
    .Y(io_outs_up_0[19]));
 BUFx2_ASAP7_75t_R output1830 (.A(net1829),
    .Y(io_outs_up_0[18]));
 BUFx2_ASAP7_75t_R output1829 (.A(net1828),
    .Y(io_outs_up_0[17]));
 BUFx2_ASAP7_75t_R output1828 (.A(net1827),
    .Y(io_outs_up_0[16]));
 BUFx2_ASAP7_75t_R output1827 (.A(net1826),
    .Y(io_outs_up_0[15]));
 BUFx2_ASAP7_75t_R output1826 (.A(net1825),
    .Y(io_outs_up_0[14]));
 BUFx2_ASAP7_75t_R output1825 (.A(net1824),
    .Y(io_outs_up_0[13]));
 BUFx2_ASAP7_75t_R output1824 (.A(net1823),
    .Y(io_outs_up_0[12]));
 BUFx2_ASAP7_75t_R output1823 (.A(net1822),
    .Y(io_outs_up_0[11]));
 BUFx2_ASAP7_75t_R output1822 (.A(net1821),
    .Y(io_outs_up_0[10]));
 BUFx2_ASAP7_75t_R output1821 (.A(net1820),
    .Y(io_outs_up_0[0]));
 BUFx2_ASAP7_75t_R output1820 (.A(net1819),
    .Y(io_outs_right_3[9]));
 BUFx2_ASAP7_75t_R output1819 (.A(net1818),
    .Y(io_outs_right_3[8]));
 BUFx2_ASAP7_75t_R output1818 (.A(net1817),
    .Y(io_outs_right_3[7]));
 BUFx2_ASAP7_75t_R output1817 (.A(net1816),
    .Y(io_outs_right_3[6]));
 BUFx2_ASAP7_75t_R output1816 (.A(net1815),
    .Y(io_outs_right_3[63]));
 BUFx2_ASAP7_75t_R output1815 (.A(net1814),
    .Y(io_outs_right_3[62]));
 BUFx2_ASAP7_75t_R output1814 (.A(net1813),
    .Y(io_outs_right_3[61]));
 BUFx2_ASAP7_75t_R output1813 (.A(net1812),
    .Y(io_outs_right_3[60]));
 BUFx2_ASAP7_75t_R output1812 (.A(net1811),
    .Y(io_outs_right_3[5]));
 BUFx2_ASAP7_75t_R output1811 (.A(net1810),
    .Y(io_outs_right_3[59]));
 BUFx2_ASAP7_75t_R output1810 (.A(net1809),
    .Y(io_outs_right_3[58]));
 BUFx2_ASAP7_75t_R output1809 (.A(net1808),
    .Y(io_outs_right_3[57]));
 BUFx2_ASAP7_75t_R output1808 (.A(net1807),
    .Y(io_outs_right_3[56]));
 BUFx2_ASAP7_75t_R output1807 (.A(net1806),
    .Y(io_outs_right_3[55]));
 BUFx2_ASAP7_75t_R output1806 (.A(net1805),
    .Y(io_outs_right_3[54]));
 BUFx2_ASAP7_75t_R output1805 (.A(net1804),
    .Y(io_outs_right_3[53]));
 BUFx2_ASAP7_75t_R output1804 (.A(net1803),
    .Y(io_outs_right_3[52]));
 BUFx2_ASAP7_75t_R output1803 (.A(net1802),
    .Y(io_outs_right_3[51]));
 BUFx2_ASAP7_75t_R output1802 (.A(net1801),
    .Y(io_outs_right_3[50]));
 BUFx2_ASAP7_75t_R output1801 (.A(net1800),
    .Y(io_outs_right_3[4]));
 BUFx2_ASAP7_75t_R output1800 (.A(net1799),
    .Y(io_outs_right_3[49]));
 BUFx2_ASAP7_75t_R output1799 (.A(net1798),
    .Y(io_outs_right_3[48]));
 BUFx2_ASAP7_75t_R output1798 (.A(net1797),
    .Y(io_outs_right_3[47]));
 BUFx2_ASAP7_75t_R output1797 (.A(net1796),
    .Y(io_outs_right_3[46]));
 BUFx2_ASAP7_75t_R output1796 (.A(net1795),
    .Y(io_outs_right_3[45]));
 BUFx2_ASAP7_75t_R output1795 (.A(net1794),
    .Y(io_outs_right_3[44]));
 BUFx2_ASAP7_75t_R output1794 (.A(net1793),
    .Y(io_outs_right_3[43]));
 BUFx2_ASAP7_75t_R output1793 (.A(net1792),
    .Y(io_outs_right_3[42]));
 BUFx2_ASAP7_75t_R output1792 (.A(net1791),
    .Y(io_outs_right_3[41]));
 BUFx2_ASAP7_75t_R output1791 (.A(net1790),
    .Y(io_outs_right_3[40]));
 BUFx2_ASAP7_75t_R output1790 (.A(net1789),
    .Y(io_outs_right_3[3]));
 BUFx2_ASAP7_75t_R output1789 (.A(net1788),
    .Y(io_outs_right_3[39]));
 BUFx2_ASAP7_75t_R output1788 (.A(net1787),
    .Y(io_outs_right_3[38]));
 BUFx2_ASAP7_75t_R output1787 (.A(net1786),
    .Y(io_outs_right_3[37]));
 BUFx2_ASAP7_75t_R output1786 (.A(net1785),
    .Y(io_outs_right_3[36]));
 BUFx2_ASAP7_75t_R output1785 (.A(net1784),
    .Y(io_outs_right_3[35]));
 BUFx2_ASAP7_75t_R output1784 (.A(net1783),
    .Y(io_outs_right_3[34]));
 BUFx2_ASAP7_75t_R output1783 (.A(net1782),
    .Y(io_outs_right_3[33]));
 BUFx2_ASAP7_75t_R output1782 (.A(net1781),
    .Y(io_outs_right_3[32]));
 BUFx2_ASAP7_75t_R output1781 (.A(net1780),
    .Y(io_outs_right_3[31]));
 BUFx2_ASAP7_75t_R output1780 (.A(net1779),
    .Y(io_outs_right_3[30]));
 BUFx2_ASAP7_75t_R output1779 (.A(net1778),
    .Y(io_outs_right_3[2]));
 BUFx2_ASAP7_75t_R output1778 (.A(net1777),
    .Y(io_outs_right_3[29]));
 BUFx2_ASAP7_75t_R output1777 (.A(net1776),
    .Y(io_outs_right_3[28]));
 BUFx2_ASAP7_75t_R output1776 (.A(net1775),
    .Y(io_outs_right_3[27]));
 BUFx2_ASAP7_75t_R output1775 (.A(net1774),
    .Y(io_outs_right_3[26]));
 BUFx2_ASAP7_75t_R output1774 (.A(net1773),
    .Y(io_outs_right_3[25]));
 BUFx2_ASAP7_75t_R output1773 (.A(net1772),
    .Y(io_outs_right_3[24]));
 BUFx2_ASAP7_75t_R output1772 (.A(net1771),
    .Y(io_outs_right_3[23]));
 BUFx2_ASAP7_75t_R output1771 (.A(net1770),
    .Y(io_outs_right_3[22]));
 BUFx2_ASAP7_75t_R output1770 (.A(net1769),
    .Y(io_outs_right_3[21]));
 BUFx2_ASAP7_75t_R output1769 (.A(net1768),
    .Y(io_outs_right_3[20]));
 BUFx2_ASAP7_75t_R output1768 (.A(net1767),
    .Y(io_outs_right_3[1]));
 BUFx2_ASAP7_75t_R output1767 (.A(net1766),
    .Y(io_outs_right_3[19]));
 BUFx2_ASAP7_75t_R output1766 (.A(net1765),
    .Y(io_outs_right_3[18]));
 BUFx2_ASAP7_75t_R output1765 (.A(net1764),
    .Y(io_outs_right_3[17]));
 BUFx2_ASAP7_75t_R output1764 (.A(net1763),
    .Y(io_outs_right_3[16]));
 BUFx2_ASAP7_75t_R output1763 (.A(net1762),
    .Y(io_outs_right_3[15]));
 BUFx2_ASAP7_75t_R output1762 (.A(net1761),
    .Y(io_outs_right_3[14]));
 BUFx2_ASAP7_75t_R output1761 (.A(net1760),
    .Y(io_outs_right_3[13]));
 BUFx2_ASAP7_75t_R output1760 (.A(net1759),
    .Y(io_outs_right_3[12]));
 BUFx2_ASAP7_75t_R output1759 (.A(net1758),
    .Y(io_outs_right_3[11]));
 BUFx2_ASAP7_75t_R output1758 (.A(net1757),
    .Y(io_outs_right_3[10]));
 BUFx2_ASAP7_75t_R output1757 (.A(net1756),
    .Y(io_outs_right_3[0]));
 BUFx2_ASAP7_75t_R output1756 (.A(net1755),
    .Y(io_outs_right_2[9]));
 BUFx2_ASAP7_75t_R output1755 (.A(net1754),
    .Y(io_outs_right_2[8]));
 BUFx2_ASAP7_75t_R output1754 (.A(net1753),
    .Y(io_outs_right_2[7]));
 BUFx2_ASAP7_75t_R output1753 (.A(net1752),
    .Y(io_outs_right_2[6]));
 BUFx2_ASAP7_75t_R output1752 (.A(net1751),
    .Y(io_outs_right_2[63]));
 BUFx2_ASAP7_75t_R output1751 (.A(net1750),
    .Y(io_outs_right_2[62]));
 BUFx2_ASAP7_75t_R output1750 (.A(net1749),
    .Y(io_outs_right_2[61]));
 BUFx2_ASAP7_75t_R output1749 (.A(net1748),
    .Y(io_outs_right_2[60]));
 BUFx2_ASAP7_75t_R output1748 (.A(net1747),
    .Y(io_outs_right_2[5]));
 BUFx2_ASAP7_75t_R output1747 (.A(net1746),
    .Y(io_outs_right_2[59]));
 BUFx2_ASAP7_75t_R output1746 (.A(net1745),
    .Y(io_outs_right_2[58]));
 BUFx2_ASAP7_75t_R output1745 (.A(net1744),
    .Y(io_outs_right_2[57]));
 BUFx2_ASAP7_75t_R output1744 (.A(net1743),
    .Y(io_outs_right_2[56]));
 BUFx2_ASAP7_75t_R output1743 (.A(net1742),
    .Y(io_outs_right_2[55]));
 BUFx2_ASAP7_75t_R output1742 (.A(net1741),
    .Y(io_outs_right_2[54]));
 BUFx2_ASAP7_75t_R output1741 (.A(net1740),
    .Y(io_outs_right_2[53]));
 BUFx2_ASAP7_75t_R output1740 (.A(net1739),
    .Y(io_outs_right_2[52]));
 BUFx2_ASAP7_75t_R output1739 (.A(net1738),
    .Y(io_outs_right_2[51]));
 BUFx2_ASAP7_75t_R output1738 (.A(net1737),
    .Y(io_outs_right_2[50]));
 BUFx2_ASAP7_75t_R output1737 (.A(net1736),
    .Y(io_outs_right_2[4]));
 BUFx2_ASAP7_75t_R output1736 (.A(net1735),
    .Y(io_outs_right_2[49]));
 BUFx2_ASAP7_75t_R output1735 (.A(net1734),
    .Y(io_outs_right_2[48]));
 BUFx2_ASAP7_75t_R output1734 (.A(net1733),
    .Y(io_outs_right_2[47]));
 BUFx2_ASAP7_75t_R output1733 (.A(net1732),
    .Y(io_outs_right_2[46]));
 BUFx2_ASAP7_75t_R output1732 (.A(net1731),
    .Y(io_outs_right_2[45]));
 BUFx2_ASAP7_75t_R output1731 (.A(net1730),
    .Y(io_outs_right_2[44]));
 BUFx2_ASAP7_75t_R output1730 (.A(net1729),
    .Y(io_outs_right_2[43]));
 BUFx2_ASAP7_75t_R output1729 (.A(net1728),
    .Y(io_outs_right_2[42]));
 BUFx2_ASAP7_75t_R output1728 (.A(net1727),
    .Y(io_outs_right_2[41]));
 BUFx2_ASAP7_75t_R output1727 (.A(net1726),
    .Y(io_outs_right_2[40]));
 BUFx2_ASAP7_75t_R output1726 (.A(net1725),
    .Y(io_outs_right_2[3]));
 BUFx2_ASAP7_75t_R output1725 (.A(net1724),
    .Y(io_outs_right_2[39]));
 BUFx2_ASAP7_75t_R output1724 (.A(net1723),
    .Y(io_outs_right_2[38]));
 BUFx2_ASAP7_75t_R output1723 (.A(net1722),
    .Y(io_outs_right_2[37]));
 BUFx2_ASAP7_75t_R output1722 (.A(net1721),
    .Y(io_outs_right_2[36]));
 BUFx2_ASAP7_75t_R output1721 (.A(net1720),
    .Y(io_outs_right_2[35]));
 BUFx2_ASAP7_75t_R output1720 (.A(net1719),
    .Y(io_outs_right_2[34]));
 BUFx2_ASAP7_75t_R output1719 (.A(net1718),
    .Y(io_outs_right_2[33]));
 BUFx2_ASAP7_75t_R output1718 (.A(net1717),
    .Y(io_outs_right_2[32]));
 BUFx2_ASAP7_75t_R output1717 (.A(net1716),
    .Y(io_outs_right_2[31]));
 BUFx2_ASAP7_75t_R output1716 (.A(net1715),
    .Y(io_outs_right_2[30]));
 BUFx2_ASAP7_75t_R output1715 (.A(net1714),
    .Y(io_outs_right_2[2]));
 BUFx2_ASAP7_75t_R output1714 (.A(net1713),
    .Y(io_outs_right_2[29]));
 BUFx2_ASAP7_75t_R output1713 (.A(net1712),
    .Y(io_outs_right_2[28]));
 BUFx2_ASAP7_75t_R output1712 (.A(net1711),
    .Y(io_outs_right_2[27]));
 BUFx2_ASAP7_75t_R output1711 (.A(net1710),
    .Y(io_outs_right_2[26]));
 BUFx2_ASAP7_75t_R output1710 (.A(net1709),
    .Y(io_outs_right_2[25]));
 BUFx2_ASAP7_75t_R output1709 (.A(net1708),
    .Y(io_outs_right_2[24]));
 BUFx2_ASAP7_75t_R output1708 (.A(net1707),
    .Y(io_outs_right_2[23]));
 BUFx2_ASAP7_75t_R output1707 (.A(net1706),
    .Y(io_outs_right_2[22]));
 BUFx2_ASAP7_75t_R output1706 (.A(net1705),
    .Y(io_outs_right_2[21]));
 BUFx2_ASAP7_75t_R output1705 (.A(net1704),
    .Y(io_outs_right_2[20]));
 BUFx2_ASAP7_75t_R output1704 (.A(net1703),
    .Y(io_outs_right_2[1]));
 BUFx2_ASAP7_75t_R output1703 (.A(net1702),
    .Y(io_outs_right_2[19]));
 BUFx2_ASAP7_75t_R output1702 (.A(net1701),
    .Y(io_outs_right_2[18]));
 BUFx2_ASAP7_75t_R output1701 (.A(net1700),
    .Y(io_outs_right_2[17]));
 BUFx2_ASAP7_75t_R output1700 (.A(net1699),
    .Y(io_outs_right_2[16]));
 BUFx2_ASAP7_75t_R output1699 (.A(net1698),
    .Y(io_outs_right_2[15]));
 BUFx2_ASAP7_75t_R output1698 (.A(net1697),
    .Y(io_outs_right_2[14]));
 BUFx2_ASAP7_75t_R output1697 (.A(net1696),
    .Y(io_outs_right_2[13]));
 BUFx2_ASAP7_75t_R output1696 (.A(net1695),
    .Y(io_outs_right_2[12]));
 BUFx2_ASAP7_75t_R output1695 (.A(net1694),
    .Y(io_outs_right_2[11]));
 BUFx2_ASAP7_75t_R output1694 (.A(net1693),
    .Y(io_outs_right_2[10]));
 BUFx2_ASAP7_75t_R output1693 (.A(net1692),
    .Y(io_outs_right_2[0]));
 BUFx2_ASAP7_75t_R output1692 (.A(net1691),
    .Y(io_outs_right_1[9]));
 BUFx2_ASAP7_75t_R output1691 (.A(net1690),
    .Y(io_outs_right_1[8]));
 BUFx2_ASAP7_75t_R output1690 (.A(net1689),
    .Y(io_outs_right_1[7]));
 BUFx2_ASAP7_75t_R output1689 (.A(net1688),
    .Y(io_outs_right_1[6]));
 BUFx2_ASAP7_75t_R output1688 (.A(net1687),
    .Y(io_outs_right_1[63]));
 BUFx2_ASAP7_75t_R output1687 (.A(net1686),
    .Y(io_outs_right_1[62]));
 BUFx2_ASAP7_75t_R output1686 (.A(net1685),
    .Y(io_outs_right_1[61]));
 BUFx2_ASAP7_75t_R output1685 (.A(net1684),
    .Y(io_outs_right_1[60]));
 BUFx2_ASAP7_75t_R output1684 (.A(net1683),
    .Y(io_outs_right_1[5]));
 BUFx2_ASAP7_75t_R output1683 (.A(net1682),
    .Y(io_outs_right_1[59]));
 BUFx2_ASAP7_75t_R output1682 (.A(net1681),
    .Y(io_outs_right_1[58]));
 BUFx2_ASAP7_75t_R output1681 (.A(net1680),
    .Y(io_outs_right_1[57]));
 BUFx2_ASAP7_75t_R output1680 (.A(net1679),
    .Y(io_outs_right_1[56]));
 BUFx2_ASAP7_75t_R output1679 (.A(net1678),
    .Y(io_outs_right_1[55]));
 BUFx2_ASAP7_75t_R output1678 (.A(net1677),
    .Y(io_outs_right_1[54]));
 BUFx2_ASAP7_75t_R output1677 (.A(net1676),
    .Y(io_outs_right_1[53]));
 BUFx2_ASAP7_75t_R output1676 (.A(net1675),
    .Y(io_outs_right_1[52]));
 BUFx2_ASAP7_75t_R output1675 (.A(net1674),
    .Y(io_outs_right_1[51]));
 BUFx2_ASAP7_75t_R output1674 (.A(net1673),
    .Y(io_outs_right_1[50]));
 BUFx2_ASAP7_75t_R output1673 (.A(net1672),
    .Y(io_outs_right_1[4]));
 BUFx2_ASAP7_75t_R output1672 (.A(net1671),
    .Y(io_outs_right_1[49]));
 BUFx2_ASAP7_75t_R output1671 (.A(net1670),
    .Y(io_outs_right_1[48]));
 BUFx2_ASAP7_75t_R output1670 (.A(net1669),
    .Y(io_outs_right_1[47]));
 BUFx2_ASAP7_75t_R output1669 (.A(net1668),
    .Y(io_outs_right_1[46]));
 BUFx2_ASAP7_75t_R output1668 (.A(net1667),
    .Y(io_outs_right_1[45]));
 BUFx2_ASAP7_75t_R output1667 (.A(net1666),
    .Y(io_outs_right_1[44]));
 BUFx2_ASAP7_75t_R output1666 (.A(net1665),
    .Y(io_outs_right_1[43]));
 BUFx2_ASAP7_75t_R output1665 (.A(net1664),
    .Y(io_outs_right_1[42]));
 BUFx2_ASAP7_75t_R output1664 (.A(net1663),
    .Y(io_outs_right_1[41]));
 BUFx2_ASAP7_75t_R output1663 (.A(net1662),
    .Y(io_outs_right_1[40]));
 BUFx2_ASAP7_75t_R output1662 (.A(net1661),
    .Y(io_outs_right_1[3]));
 BUFx2_ASAP7_75t_R output1661 (.A(net1660),
    .Y(io_outs_right_1[39]));
 BUFx2_ASAP7_75t_R output1660 (.A(net1659),
    .Y(io_outs_right_1[38]));
 BUFx2_ASAP7_75t_R output1659 (.A(net1658),
    .Y(io_outs_right_1[37]));
 BUFx2_ASAP7_75t_R output1658 (.A(net1657),
    .Y(io_outs_right_1[36]));
 BUFx2_ASAP7_75t_R output1657 (.A(net1656),
    .Y(io_outs_right_1[35]));
 BUFx2_ASAP7_75t_R output1656 (.A(net1655),
    .Y(io_outs_right_1[34]));
 BUFx2_ASAP7_75t_R output1655 (.A(net1654),
    .Y(io_outs_right_1[33]));
 BUFx2_ASAP7_75t_R output1654 (.A(net1653),
    .Y(io_outs_right_1[32]));
 BUFx2_ASAP7_75t_R output1653 (.A(net1652),
    .Y(io_outs_right_1[31]));
 BUFx2_ASAP7_75t_R output1652 (.A(net1651),
    .Y(io_outs_right_1[30]));
 BUFx2_ASAP7_75t_R output1651 (.A(net1650),
    .Y(io_outs_right_1[2]));
 BUFx2_ASAP7_75t_R output1650 (.A(net1649),
    .Y(io_outs_right_1[29]));
 BUFx2_ASAP7_75t_R output1649 (.A(net1648),
    .Y(io_outs_right_1[28]));
 BUFx2_ASAP7_75t_R output1648 (.A(net1647),
    .Y(io_outs_right_1[27]));
 BUFx2_ASAP7_75t_R output1647 (.A(net1646),
    .Y(io_outs_right_1[26]));
 BUFx2_ASAP7_75t_R output1646 (.A(net1645),
    .Y(io_outs_right_1[25]));
 BUFx2_ASAP7_75t_R output1645 (.A(net1644),
    .Y(io_outs_right_1[24]));
 BUFx2_ASAP7_75t_R output1644 (.A(net1643),
    .Y(io_outs_right_1[23]));
 BUFx2_ASAP7_75t_R output1643 (.A(net1642),
    .Y(io_outs_right_1[22]));
 BUFx2_ASAP7_75t_R output1642 (.A(net1641),
    .Y(io_outs_right_1[21]));
 BUFx2_ASAP7_75t_R output1641 (.A(net1640),
    .Y(io_outs_right_1[20]));
 BUFx2_ASAP7_75t_R output1640 (.A(net1639),
    .Y(io_outs_right_1[1]));
 BUFx2_ASAP7_75t_R output1639 (.A(net1638),
    .Y(io_outs_right_1[19]));
 BUFx2_ASAP7_75t_R output1638 (.A(net1637),
    .Y(io_outs_right_1[18]));
 BUFx2_ASAP7_75t_R output1637 (.A(net1636),
    .Y(io_outs_right_1[17]));
 BUFx2_ASAP7_75t_R output1636 (.A(net1635),
    .Y(io_outs_right_1[16]));
 BUFx2_ASAP7_75t_R output1635 (.A(net1634),
    .Y(io_outs_right_1[15]));
 BUFx2_ASAP7_75t_R output1634 (.A(net1633),
    .Y(io_outs_right_1[14]));
 BUFx2_ASAP7_75t_R output1633 (.A(net1632),
    .Y(io_outs_right_1[13]));
 BUFx2_ASAP7_75t_R output1632 (.A(net1631),
    .Y(io_outs_right_1[12]));
 BUFx2_ASAP7_75t_R output1631 (.A(net1630),
    .Y(io_outs_right_1[11]));
 BUFx2_ASAP7_75t_R output1630 (.A(net1629),
    .Y(io_outs_right_1[10]));
 BUFx2_ASAP7_75t_R output1629 (.A(net1628),
    .Y(io_outs_right_1[0]));
 BUFx2_ASAP7_75t_R output1628 (.A(net1627),
    .Y(io_outs_right_0[9]));
 BUFx2_ASAP7_75t_R output1627 (.A(net1626),
    .Y(io_outs_right_0[8]));
 BUFx2_ASAP7_75t_R output1626 (.A(net1625),
    .Y(io_outs_right_0[7]));
 BUFx2_ASAP7_75t_R output1625 (.A(net1624),
    .Y(io_outs_right_0[6]));
 BUFx2_ASAP7_75t_R output1624 (.A(net1623),
    .Y(io_outs_right_0[63]));
 BUFx2_ASAP7_75t_R output1623 (.A(net1622),
    .Y(io_outs_right_0[62]));
 BUFx2_ASAP7_75t_R output1622 (.A(net1621),
    .Y(io_outs_right_0[61]));
 BUFx2_ASAP7_75t_R output1621 (.A(net1620),
    .Y(io_outs_right_0[60]));
 BUFx2_ASAP7_75t_R output1620 (.A(net1619),
    .Y(io_outs_right_0[5]));
 BUFx2_ASAP7_75t_R output1619 (.A(net1618),
    .Y(io_outs_right_0[59]));
 BUFx2_ASAP7_75t_R output1618 (.A(net1617),
    .Y(io_outs_right_0[58]));
 BUFx2_ASAP7_75t_R output1617 (.A(net1616),
    .Y(io_outs_right_0[57]));
 BUFx2_ASAP7_75t_R output1616 (.A(net1615),
    .Y(io_outs_right_0[56]));
 BUFx2_ASAP7_75t_R output1615 (.A(net1614),
    .Y(io_outs_right_0[55]));
 BUFx2_ASAP7_75t_R output1614 (.A(net1613),
    .Y(io_outs_right_0[54]));
 BUFx2_ASAP7_75t_R output1613 (.A(net1612),
    .Y(io_outs_right_0[53]));
 BUFx2_ASAP7_75t_R output1612 (.A(net1611),
    .Y(io_outs_right_0[52]));
 BUFx2_ASAP7_75t_R output1611 (.A(net1610),
    .Y(io_outs_right_0[51]));
 BUFx2_ASAP7_75t_R output1610 (.A(net1609),
    .Y(io_outs_right_0[50]));
 BUFx2_ASAP7_75t_R output1609 (.A(net1608),
    .Y(io_outs_right_0[4]));
 BUFx2_ASAP7_75t_R output1608 (.A(net1607),
    .Y(io_outs_right_0[49]));
 BUFx2_ASAP7_75t_R output1607 (.A(net1606),
    .Y(io_outs_right_0[48]));
 BUFx2_ASAP7_75t_R output1606 (.A(net1605),
    .Y(io_outs_right_0[47]));
 BUFx2_ASAP7_75t_R output1605 (.A(net1604),
    .Y(io_outs_right_0[46]));
 BUFx2_ASAP7_75t_R output1604 (.A(net1603),
    .Y(io_outs_right_0[45]));
 BUFx2_ASAP7_75t_R output1603 (.A(net1602),
    .Y(io_outs_right_0[44]));
 BUFx2_ASAP7_75t_R output1602 (.A(net1601),
    .Y(io_outs_right_0[43]));
 BUFx2_ASAP7_75t_R output1601 (.A(net1600),
    .Y(io_outs_right_0[42]));
 BUFx2_ASAP7_75t_R output1600 (.A(net1599),
    .Y(io_outs_right_0[41]));
 BUFx2_ASAP7_75t_R output1599 (.A(net1598),
    .Y(io_outs_right_0[40]));
 BUFx2_ASAP7_75t_R output1598 (.A(net1597),
    .Y(io_outs_right_0[3]));
 BUFx2_ASAP7_75t_R output1597 (.A(net1596),
    .Y(io_outs_right_0[39]));
 BUFx2_ASAP7_75t_R output1596 (.A(net1595),
    .Y(io_outs_right_0[38]));
 BUFx2_ASAP7_75t_R output1595 (.A(net1594),
    .Y(io_outs_right_0[37]));
 BUFx2_ASAP7_75t_R output1594 (.A(net1593),
    .Y(io_outs_right_0[36]));
 BUFx2_ASAP7_75t_R output1593 (.A(net1592),
    .Y(io_outs_right_0[35]));
 BUFx2_ASAP7_75t_R output1592 (.A(net1591),
    .Y(io_outs_right_0[34]));
 BUFx2_ASAP7_75t_R output1591 (.A(net1590),
    .Y(io_outs_right_0[33]));
 BUFx2_ASAP7_75t_R output1590 (.A(net1589),
    .Y(io_outs_right_0[32]));
 BUFx2_ASAP7_75t_R output1589 (.A(net1588),
    .Y(io_outs_right_0[31]));
 BUFx2_ASAP7_75t_R output1588 (.A(net1587),
    .Y(io_outs_right_0[30]));
 BUFx2_ASAP7_75t_R output1587 (.A(net1586),
    .Y(io_outs_right_0[2]));
 BUFx2_ASAP7_75t_R output1586 (.A(net1585),
    .Y(io_outs_right_0[29]));
 BUFx2_ASAP7_75t_R output1585 (.A(net1584),
    .Y(io_outs_right_0[28]));
 BUFx2_ASAP7_75t_R output1584 (.A(net1583),
    .Y(io_outs_right_0[27]));
 BUFx2_ASAP7_75t_R output1583 (.A(net1582),
    .Y(io_outs_right_0[26]));
 BUFx2_ASAP7_75t_R output1582 (.A(net1581),
    .Y(io_outs_right_0[25]));
 BUFx2_ASAP7_75t_R output1581 (.A(net1580),
    .Y(io_outs_right_0[24]));
 BUFx2_ASAP7_75t_R output1580 (.A(net1579),
    .Y(io_outs_right_0[23]));
 BUFx2_ASAP7_75t_R output1579 (.A(net1578),
    .Y(io_outs_right_0[22]));
 BUFx2_ASAP7_75t_R output1578 (.A(net1577),
    .Y(io_outs_right_0[21]));
 BUFx2_ASAP7_75t_R output1577 (.A(net1576),
    .Y(io_outs_right_0[20]));
 BUFx2_ASAP7_75t_R output1576 (.A(net1575),
    .Y(io_outs_right_0[1]));
 BUFx2_ASAP7_75t_R output1575 (.A(net1574),
    .Y(io_outs_right_0[19]));
 BUFx2_ASAP7_75t_R output1574 (.A(net1573),
    .Y(io_outs_right_0[18]));
 BUFx2_ASAP7_75t_R output1573 (.A(net1572),
    .Y(io_outs_right_0[17]));
 BUFx2_ASAP7_75t_R output1572 (.A(net1571),
    .Y(io_outs_right_0[16]));
 BUFx2_ASAP7_75t_R output1571 (.A(net1570),
    .Y(io_outs_right_0[15]));
 BUFx2_ASAP7_75t_R output1570 (.A(net1569),
    .Y(io_outs_right_0[14]));
 BUFx2_ASAP7_75t_R output1569 (.A(net1568),
    .Y(io_outs_right_0[13]));
 BUFx2_ASAP7_75t_R output1568 (.A(net1567),
    .Y(io_outs_right_0[12]));
 BUFx2_ASAP7_75t_R output1567 (.A(net1566),
    .Y(io_outs_right_0[11]));
 BUFx2_ASAP7_75t_R output1566 (.A(net1565),
    .Y(io_outs_right_0[10]));
 BUFx2_ASAP7_75t_R output1565 (.A(net1564),
    .Y(io_outs_right_0[0]));
 BUFx2_ASAP7_75t_R output1564 (.A(net1563),
    .Y(io_outs_left_3[9]));
 BUFx2_ASAP7_75t_R output1563 (.A(net1562),
    .Y(io_outs_left_3[8]));
 BUFx2_ASAP7_75t_R output1562 (.A(net1561),
    .Y(io_outs_left_3[7]));
 BUFx2_ASAP7_75t_R output1561 (.A(net1560),
    .Y(io_outs_left_3[6]));
 BUFx2_ASAP7_75t_R output1560 (.A(net1559),
    .Y(io_outs_left_3[63]));
 BUFx2_ASAP7_75t_R output1559 (.A(net1558),
    .Y(io_outs_left_3[62]));
 BUFx2_ASAP7_75t_R output1558 (.A(net1557),
    .Y(io_outs_left_3[61]));
 BUFx2_ASAP7_75t_R output1557 (.A(net1556),
    .Y(io_outs_left_3[60]));
 BUFx2_ASAP7_75t_R output1556 (.A(net1555),
    .Y(io_outs_left_3[5]));
 BUFx2_ASAP7_75t_R output1555 (.A(net1554),
    .Y(io_outs_left_3[59]));
 BUFx2_ASAP7_75t_R output1554 (.A(net1553),
    .Y(io_outs_left_3[58]));
 BUFx2_ASAP7_75t_R output1553 (.A(net1552),
    .Y(io_outs_left_3[57]));
 BUFx2_ASAP7_75t_R output1552 (.A(net1551),
    .Y(io_outs_left_3[56]));
 BUFx2_ASAP7_75t_R output1551 (.A(net1550),
    .Y(io_outs_left_3[55]));
 BUFx2_ASAP7_75t_R output1550 (.A(net1549),
    .Y(io_outs_left_3[54]));
 BUFx2_ASAP7_75t_R output1549 (.A(net1548),
    .Y(io_outs_left_3[53]));
 BUFx2_ASAP7_75t_R output1548 (.A(net1547),
    .Y(io_outs_left_3[52]));
 BUFx2_ASAP7_75t_R output1547 (.A(net1546),
    .Y(io_outs_left_3[51]));
 BUFx2_ASAP7_75t_R output1546 (.A(net1545),
    .Y(io_outs_left_3[50]));
 BUFx2_ASAP7_75t_R output1545 (.A(net1544),
    .Y(io_outs_left_3[4]));
 BUFx2_ASAP7_75t_R output1544 (.A(net1543),
    .Y(io_outs_left_3[49]));
 BUFx2_ASAP7_75t_R output1543 (.A(net1542),
    .Y(io_outs_left_3[48]));
 BUFx2_ASAP7_75t_R output1542 (.A(net1541),
    .Y(io_outs_left_3[47]));
 BUFx2_ASAP7_75t_R output1541 (.A(net1540),
    .Y(io_outs_left_3[46]));
 BUFx2_ASAP7_75t_R output1540 (.A(net1539),
    .Y(io_outs_left_3[45]));
 BUFx2_ASAP7_75t_R output1539 (.A(net1538),
    .Y(io_outs_left_3[44]));
 BUFx2_ASAP7_75t_R output1538 (.A(net1537),
    .Y(io_outs_left_3[43]));
 BUFx2_ASAP7_75t_R output1537 (.A(net1536),
    .Y(io_outs_left_3[42]));
 BUFx2_ASAP7_75t_R output1536 (.A(net1535),
    .Y(io_outs_left_3[41]));
 BUFx2_ASAP7_75t_R output1535 (.A(net1534),
    .Y(io_outs_left_3[40]));
 BUFx2_ASAP7_75t_R output1534 (.A(net1533),
    .Y(io_outs_left_3[3]));
 BUFx2_ASAP7_75t_R output1533 (.A(net1532),
    .Y(io_outs_left_3[39]));
 BUFx2_ASAP7_75t_R output1532 (.A(net1531),
    .Y(io_outs_left_3[38]));
 BUFx2_ASAP7_75t_R output1531 (.A(net1530),
    .Y(io_outs_left_3[37]));
 BUFx2_ASAP7_75t_R output1530 (.A(net1529),
    .Y(io_outs_left_3[36]));
 BUFx2_ASAP7_75t_R output1529 (.A(net1528),
    .Y(io_outs_left_3[35]));
 BUFx2_ASAP7_75t_R output1528 (.A(net1527),
    .Y(io_outs_left_3[34]));
 BUFx2_ASAP7_75t_R output1527 (.A(net1526),
    .Y(io_outs_left_3[33]));
 BUFx2_ASAP7_75t_R output1526 (.A(net1525),
    .Y(io_outs_left_3[32]));
 BUFx2_ASAP7_75t_R output1525 (.A(net1524),
    .Y(io_outs_left_3[31]));
 BUFx2_ASAP7_75t_R output1524 (.A(net1523),
    .Y(io_outs_left_3[30]));
 BUFx2_ASAP7_75t_R output1523 (.A(net1522),
    .Y(io_outs_left_3[2]));
 BUFx2_ASAP7_75t_R output1522 (.A(net1521),
    .Y(io_outs_left_3[29]));
 BUFx2_ASAP7_75t_R output1521 (.A(net1520),
    .Y(io_outs_left_3[28]));
 BUFx2_ASAP7_75t_R output1520 (.A(net1519),
    .Y(io_outs_left_3[27]));
 BUFx2_ASAP7_75t_R output1519 (.A(net1518),
    .Y(io_outs_left_3[26]));
 BUFx2_ASAP7_75t_R output1518 (.A(net1517),
    .Y(io_outs_left_3[25]));
 BUFx2_ASAP7_75t_R output1517 (.A(net1516),
    .Y(io_outs_left_3[24]));
 BUFx2_ASAP7_75t_R output1516 (.A(net1515),
    .Y(io_outs_left_3[23]));
 BUFx2_ASAP7_75t_R output1515 (.A(net1514),
    .Y(io_outs_left_3[22]));
 BUFx2_ASAP7_75t_R output1514 (.A(net1513),
    .Y(io_outs_left_3[21]));
 BUFx2_ASAP7_75t_R output1513 (.A(net1512),
    .Y(io_outs_left_3[20]));
 BUFx2_ASAP7_75t_R output1512 (.A(net1511),
    .Y(io_outs_left_3[1]));
 BUFx2_ASAP7_75t_R output1511 (.A(net1510),
    .Y(io_outs_left_3[19]));
 BUFx2_ASAP7_75t_R output1510 (.A(net1509),
    .Y(io_outs_left_3[18]));
 BUFx2_ASAP7_75t_R output1509 (.A(net1508),
    .Y(io_outs_left_3[17]));
 BUFx2_ASAP7_75t_R output1508 (.A(net1507),
    .Y(io_outs_left_3[16]));
 BUFx2_ASAP7_75t_R output1507 (.A(net1506),
    .Y(io_outs_left_3[15]));
 BUFx2_ASAP7_75t_R output1506 (.A(net1505),
    .Y(io_outs_left_3[14]));
 BUFx2_ASAP7_75t_R output1505 (.A(net1504),
    .Y(io_outs_left_3[13]));
 BUFx2_ASAP7_75t_R output1504 (.A(net1503),
    .Y(io_outs_left_3[12]));
 BUFx2_ASAP7_75t_R output1503 (.A(net1502),
    .Y(io_outs_left_3[11]));
 BUFx2_ASAP7_75t_R output1502 (.A(net1501),
    .Y(io_outs_left_3[10]));
 BUFx2_ASAP7_75t_R output1501 (.A(net1500),
    .Y(io_outs_left_3[0]));
 BUFx2_ASAP7_75t_R output1500 (.A(net1499),
    .Y(io_outs_left_2[9]));
 BUFx2_ASAP7_75t_R output1499 (.A(net1498),
    .Y(io_outs_left_2[8]));
 BUFx2_ASAP7_75t_R output1498 (.A(net1497),
    .Y(io_outs_left_2[7]));
 BUFx2_ASAP7_75t_R output1497 (.A(net1496),
    .Y(io_outs_left_2[6]));
 BUFx2_ASAP7_75t_R output1496 (.A(net1495),
    .Y(io_outs_left_2[63]));
 BUFx2_ASAP7_75t_R output1495 (.A(net1494),
    .Y(io_outs_left_2[62]));
 BUFx2_ASAP7_75t_R output1494 (.A(net1493),
    .Y(io_outs_left_2[61]));
 BUFx2_ASAP7_75t_R output1493 (.A(net1492),
    .Y(io_outs_left_2[60]));
 BUFx2_ASAP7_75t_R output1492 (.A(net1491),
    .Y(io_outs_left_2[5]));
 BUFx2_ASAP7_75t_R output1491 (.A(net1490),
    .Y(io_outs_left_2[59]));
 BUFx2_ASAP7_75t_R output1490 (.A(net1489),
    .Y(io_outs_left_2[58]));
 BUFx2_ASAP7_75t_R output1489 (.A(net1488),
    .Y(io_outs_left_2[57]));
 BUFx2_ASAP7_75t_R output1488 (.A(net1487),
    .Y(io_outs_left_2[56]));
 BUFx2_ASAP7_75t_R output1487 (.A(net1486),
    .Y(io_outs_left_2[55]));
 BUFx2_ASAP7_75t_R output1486 (.A(net1485),
    .Y(io_outs_left_2[54]));
 BUFx2_ASAP7_75t_R output1485 (.A(net1484),
    .Y(io_outs_left_2[53]));
 BUFx2_ASAP7_75t_R output1484 (.A(net1483),
    .Y(io_outs_left_2[52]));
 BUFx2_ASAP7_75t_R output1483 (.A(net1482),
    .Y(io_outs_left_2[51]));
 BUFx2_ASAP7_75t_R output1482 (.A(net1481),
    .Y(io_outs_left_2[50]));
 BUFx2_ASAP7_75t_R output1481 (.A(net1480),
    .Y(io_outs_left_2[4]));
 BUFx2_ASAP7_75t_R output1480 (.A(net1479),
    .Y(io_outs_left_2[49]));
 BUFx2_ASAP7_75t_R output1479 (.A(net1478),
    .Y(io_outs_left_2[48]));
 BUFx2_ASAP7_75t_R output1478 (.A(net1477),
    .Y(io_outs_left_2[47]));
 BUFx2_ASAP7_75t_R output1477 (.A(net1476),
    .Y(io_outs_left_2[46]));
 BUFx2_ASAP7_75t_R output1476 (.A(net1475),
    .Y(io_outs_left_2[45]));
 BUFx2_ASAP7_75t_R output1475 (.A(net1474),
    .Y(io_outs_left_2[44]));
 BUFx2_ASAP7_75t_R output1474 (.A(net1473),
    .Y(io_outs_left_2[43]));
 BUFx2_ASAP7_75t_R output1473 (.A(net1472),
    .Y(io_outs_left_2[42]));
 BUFx2_ASAP7_75t_R output1472 (.A(net1471),
    .Y(io_outs_left_2[41]));
 BUFx2_ASAP7_75t_R output1471 (.A(net1470),
    .Y(io_outs_left_2[40]));
 BUFx2_ASAP7_75t_R output1470 (.A(net1469),
    .Y(io_outs_left_2[3]));
 BUFx2_ASAP7_75t_R output1469 (.A(net1468),
    .Y(io_outs_left_2[39]));
 BUFx2_ASAP7_75t_R output1468 (.A(net1467),
    .Y(io_outs_left_2[38]));
 BUFx2_ASAP7_75t_R output1467 (.A(net1466),
    .Y(io_outs_left_2[37]));
 BUFx2_ASAP7_75t_R output1466 (.A(net1465),
    .Y(io_outs_left_2[36]));
 BUFx2_ASAP7_75t_R output1465 (.A(net1464),
    .Y(io_outs_left_2[35]));
 BUFx2_ASAP7_75t_R output1464 (.A(net1463),
    .Y(io_outs_left_2[34]));
 BUFx2_ASAP7_75t_R output1463 (.A(net1462),
    .Y(io_outs_left_2[33]));
 BUFx2_ASAP7_75t_R output1462 (.A(net1461),
    .Y(io_outs_left_2[32]));
 BUFx2_ASAP7_75t_R output1461 (.A(net1460),
    .Y(io_outs_left_2[31]));
 BUFx2_ASAP7_75t_R output1460 (.A(net1459),
    .Y(io_outs_left_2[30]));
 BUFx2_ASAP7_75t_R output1459 (.A(net1458),
    .Y(io_outs_left_2[2]));
 BUFx2_ASAP7_75t_R output1458 (.A(net1457),
    .Y(io_outs_left_2[29]));
 BUFx2_ASAP7_75t_R output1457 (.A(net1456),
    .Y(io_outs_left_2[28]));
 BUFx2_ASAP7_75t_R output1456 (.A(net1455),
    .Y(io_outs_left_2[27]));
 BUFx2_ASAP7_75t_R output1455 (.A(net1454),
    .Y(io_outs_left_2[26]));
 BUFx2_ASAP7_75t_R output1454 (.A(net1453),
    .Y(io_outs_left_2[25]));
 BUFx2_ASAP7_75t_R output1453 (.A(net1452),
    .Y(io_outs_left_2[24]));
 BUFx2_ASAP7_75t_R output1452 (.A(net1451),
    .Y(io_outs_left_2[23]));
 BUFx2_ASAP7_75t_R output1451 (.A(net1450),
    .Y(io_outs_left_2[22]));
 BUFx2_ASAP7_75t_R output1450 (.A(net1449),
    .Y(io_outs_left_2[21]));
 BUFx2_ASAP7_75t_R output1449 (.A(net1448),
    .Y(io_outs_left_2[20]));
 BUFx2_ASAP7_75t_R output1448 (.A(net1447),
    .Y(io_outs_left_2[1]));
 BUFx2_ASAP7_75t_R output1447 (.A(net1446),
    .Y(io_outs_left_2[19]));
 BUFx2_ASAP7_75t_R output1446 (.A(net1445),
    .Y(io_outs_left_2[18]));
 BUFx2_ASAP7_75t_R output1445 (.A(net1444),
    .Y(io_outs_left_2[17]));
 BUFx2_ASAP7_75t_R output1444 (.A(net1443),
    .Y(io_outs_left_2[16]));
 BUFx2_ASAP7_75t_R output1443 (.A(net1442),
    .Y(io_outs_left_2[15]));
 BUFx2_ASAP7_75t_R output1442 (.A(net1441),
    .Y(io_outs_left_2[14]));
 BUFx2_ASAP7_75t_R output1441 (.A(net1440),
    .Y(io_outs_left_2[13]));
 BUFx2_ASAP7_75t_R output1440 (.A(net1439),
    .Y(io_outs_left_2[12]));
 BUFx2_ASAP7_75t_R output1439 (.A(net1438),
    .Y(io_outs_left_2[11]));
 BUFx2_ASAP7_75t_R output1438 (.A(net1437),
    .Y(io_outs_left_2[10]));
 BUFx2_ASAP7_75t_R output1437 (.A(net1436),
    .Y(io_outs_left_2[0]));
 BUFx2_ASAP7_75t_R output1436 (.A(net1435),
    .Y(io_outs_left_1[9]));
 BUFx2_ASAP7_75t_R output1435 (.A(net1434),
    .Y(io_outs_left_1[8]));
 BUFx2_ASAP7_75t_R output1434 (.A(net1433),
    .Y(io_outs_left_1[7]));
 BUFx2_ASAP7_75t_R output1433 (.A(net1432),
    .Y(io_outs_left_1[6]));
 BUFx2_ASAP7_75t_R output1432 (.A(net1431),
    .Y(io_outs_left_1[63]));
 BUFx2_ASAP7_75t_R output1431 (.A(net1430),
    .Y(io_outs_left_1[62]));
 BUFx2_ASAP7_75t_R output1430 (.A(net1429),
    .Y(io_outs_left_1[61]));
 BUFx2_ASAP7_75t_R output1429 (.A(net1428),
    .Y(io_outs_left_1[60]));
 BUFx2_ASAP7_75t_R output1428 (.A(net1427),
    .Y(io_outs_left_1[5]));
 BUFx2_ASAP7_75t_R output1427 (.A(net1426),
    .Y(io_outs_left_1[59]));
 BUFx2_ASAP7_75t_R output1426 (.A(net1425),
    .Y(io_outs_left_1[58]));
 BUFx2_ASAP7_75t_R output1425 (.A(net1424),
    .Y(io_outs_left_1[57]));
 BUFx2_ASAP7_75t_R output1424 (.A(net1423),
    .Y(io_outs_left_1[56]));
 BUFx2_ASAP7_75t_R output1423 (.A(net1422),
    .Y(io_outs_left_1[55]));
 BUFx2_ASAP7_75t_R output1422 (.A(net1421),
    .Y(io_outs_left_1[54]));
 BUFx2_ASAP7_75t_R output1421 (.A(net1420),
    .Y(io_outs_left_1[53]));
 BUFx2_ASAP7_75t_R output1420 (.A(net1419),
    .Y(io_outs_left_1[52]));
 BUFx2_ASAP7_75t_R output1419 (.A(net1418),
    .Y(io_outs_left_1[51]));
 BUFx2_ASAP7_75t_R output1418 (.A(net1417),
    .Y(io_outs_left_1[50]));
 BUFx2_ASAP7_75t_R output1417 (.A(net1416),
    .Y(io_outs_left_1[4]));
 BUFx2_ASAP7_75t_R output1416 (.A(net1415),
    .Y(io_outs_left_1[49]));
 BUFx2_ASAP7_75t_R output1415 (.A(net1414),
    .Y(io_outs_left_1[48]));
 BUFx2_ASAP7_75t_R output1414 (.A(net1413),
    .Y(io_outs_left_1[47]));
 BUFx2_ASAP7_75t_R output1413 (.A(net1412),
    .Y(io_outs_left_1[46]));
 BUFx2_ASAP7_75t_R output1412 (.A(net1411),
    .Y(io_outs_left_1[45]));
 BUFx2_ASAP7_75t_R output1411 (.A(net1410),
    .Y(io_outs_left_1[44]));
 BUFx2_ASAP7_75t_R output1410 (.A(net1409),
    .Y(io_outs_left_1[43]));
 BUFx2_ASAP7_75t_R output1409 (.A(net1408),
    .Y(io_outs_left_1[42]));
 BUFx2_ASAP7_75t_R output1408 (.A(net1407),
    .Y(io_outs_left_1[41]));
 BUFx2_ASAP7_75t_R output1407 (.A(net1406),
    .Y(io_outs_left_1[40]));
 BUFx2_ASAP7_75t_R output1406 (.A(net1405),
    .Y(io_outs_left_1[3]));
 BUFx2_ASAP7_75t_R output1405 (.A(net1404),
    .Y(io_outs_left_1[39]));
 BUFx2_ASAP7_75t_R output1404 (.A(net1403),
    .Y(io_outs_left_1[38]));
 BUFx2_ASAP7_75t_R output1403 (.A(net1402),
    .Y(io_outs_left_1[37]));
 BUFx2_ASAP7_75t_R output1402 (.A(net1401),
    .Y(io_outs_left_1[36]));
 BUFx2_ASAP7_75t_R output1401 (.A(net1400),
    .Y(io_outs_left_1[35]));
 BUFx2_ASAP7_75t_R output1400 (.A(net1399),
    .Y(io_outs_left_1[34]));
 BUFx2_ASAP7_75t_R output1399 (.A(net1398),
    .Y(io_outs_left_1[33]));
 BUFx2_ASAP7_75t_R output1398 (.A(net1397),
    .Y(io_outs_left_1[32]));
 BUFx2_ASAP7_75t_R output1397 (.A(net1396),
    .Y(io_outs_left_1[31]));
 BUFx2_ASAP7_75t_R output1396 (.A(net1395),
    .Y(io_outs_left_1[30]));
 BUFx2_ASAP7_75t_R output1395 (.A(net1394),
    .Y(io_outs_left_1[2]));
 BUFx2_ASAP7_75t_R output1394 (.A(net1393),
    .Y(io_outs_left_1[29]));
 BUFx2_ASAP7_75t_R output1393 (.A(net1392),
    .Y(io_outs_left_1[28]));
 BUFx2_ASAP7_75t_R output1392 (.A(net1391),
    .Y(io_outs_left_1[27]));
 BUFx2_ASAP7_75t_R output1391 (.A(net1390),
    .Y(io_outs_left_1[26]));
 BUFx2_ASAP7_75t_R output1390 (.A(net1389),
    .Y(io_outs_left_1[25]));
 BUFx2_ASAP7_75t_R output1389 (.A(net1388),
    .Y(io_outs_left_1[24]));
 BUFx2_ASAP7_75t_R output1388 (.A(net1387),
    .Y(io_outs_left_1[23]));
 BUFx2_ASAP7_75t_R output1387 (.A(net1386),
    .Y(io_outs_left_1[22]));
 BUFx2_ASAP7_75t_R output1386 (.A(net1385),
    .Y(io_outs_left_1[21]));
 BUFx2_ASAP7_75t_R output1385 (.A(net1384),
    .Y(io_outs_left_1[20]));
 BUFx2_ASAP7_75t_R output1384 (.A(net1383),
    .Y(io_outs_left_1[1]));
 BUFx2_ASAP7_75t_R output1383 (.A(net1382),
    .Y(io_outs_left_1[19]));
 BUFx2_ASAP7_75t_R output1382 (.A(net1381),
    .Y(io_outs_left_1[18]));
 BUFx2_ASAP7_75t_R output1381 (.A(net1380),
    .Y(io_outs_left_1[17]));
 BUFx2_ASAP7_75t_R output1380 (.A(net1379),
    .Y(io_outs_left_1[16]));
 BUFx2_ASAP7_75t_R output1379 (.A(net1378),
    .Y(io_outs_left_1[15]));
 BUFx2_ASAP7_75t_R output1378 (.A(net1377),
    .Y(io_outs_left_1[14]));
 BUFx2_ASAP7_75t_R output1377 (.A(net1376),
    .Y(io_outs_left_1[13]));
 BUFx2_ASAP7_75t_R output1376 (.A(net1375),
    .Y(io_outs_left_1[12]));
 BUFx2_ASAP7_75t_R output1375 (.A(net1374),
    .Y(io_outs_left_1[11]));
 BUFx2_ASAP7_75t_R output1374 (.A(net1373),
    .Y(io_outs_left_1[10]));
 BUFx2_ASAP7_75t_R output1373 (.A(net1372),
    .Y(io_outs_left_1[0]));
 BUFx2_ASAP7_75t_R output1372 (.A(net1371),
    .Y(io_outs_left_0[9]));
 BUFx2_ASAP7_75t_R output1371 (.A(net1370),
    .Y(io_outs_left_0[8]));
 BUFx2_ASAP7_75t_R output1370 (.A(net1369),
    .Y(io_outs_left_0[7]));
 BUFx2_ASAP7_75t_R output1369 (.A(net1368),
    .Y(io_outs_left_0[6]));
 BUFx2_ASAP7_75t_R output1368 (.A(net1367),
    .Y(io_outs_left_0[63]));
 BUFx2_ASAP7_75t_R output1367 (.A(net1366),
    .Y(io_outs_left_0[62]));
 BUFx2_ASAP7_75t_R output1366 (.A(net1365),
    .Y(io_outs_left_0[61]));
 BUFx2_ASAP7_75t_R output1365 (.A(net1364),
    .Y(io_outs_left_0[60]));
 BUFx2_ASAP7_75t_R output1364 (.A(net1363),
    .Y(io_outs_left_0[5]));
 BUFx2_ASAP7_75t_R output1363 (.A(net1362),
    .Y(io_outs_left_0[59]));
 BUFx2_ASAP7_75t_R output1362 (.A(net1361),
    .Y(io_outs_left_0[58]));
 BUFx2_ASAP7_75t_R output1361 (.A(net1360),
    .Y(io_outs_left_0[57]));
 BUFx2_ASAP7_75t_R output1360 (.A(net1359),
    .Y(io_outs_left_0[56]));
 BUFx2_ASAP7_75t_R output1359 (.A(net1358),
    .Y(io_outs_left_0[55]));
 BUFx2_ASAP7_75t_R output1358 (.A(net1357),
    .Y(io_outs_left_0[54]));
 BUFx2_ASAP7_75t_R output1357 (.A(net1356),
    .Y(io_outs_left_0[53]));
 BUFx2_ASAP7_75t_R output1356 (.A(net1355),
    .Y(io_outs_left_0[52]));
 BUFx2_ASAP7_75t_R output1355 (.A(net1354),
    .Y(io_outs_left_0[51]));
 BUFx2_ASAP7_75t_R output1354 (.A(net1353),
    .Y(io_outs_left_0[50]));
 BUFx2_ASAP7_75t_R output1353 (.A(net1352),
    .Y(io_outs_left_0[4]));
 BUFx2_ASAP7_75t_R output1352 (.A(net1351),
    .Y(io_outs_left_0[49]));
 BUFx2_ASAP7_75t_R output1351 (.A(net1350),
    .Y(io_outs_left_0[48]));
 BUFx2_ASAP7_75t_R output1350 (.A(net1349),
    .Y(io_outs_left_0[47]));
 BUFx2_ASAP7_75t_R output1349 (.A(net1348),
    .Y(io_outs_left_0[46]));
 BUFx2_ASAP7_75t_R output1348 (.A(net1347),
    .Y(io_outs_left_0[45]));
 BUFx2_ASAP7_75t_R output1347 (.A(net1346),
    .Y(io_outs_left_0[44]));
 BUFx2_ASAP7_75t_R output1346 (.A(net1345),
    .Y(io_outs_left_0[43]));
 BUFx2_ASAP7_75t_R output1345 (.A(net1344),
    .Y(io_outs_left_0[42]));
 BUFx2_ASAP7_75t_R output1344 (.A(net1343),
    .Y(io_outs_left_0[41]));
 BUFx2_ASAP7_75t_R output1343 (.A(net1342),
    .Y(io_outs_left_0[40]));
 BUFx2_ASAP7_75t_R output1342 (.A(net1341),
    .Y(io_outs_left_0[3]));
 BUFx2_ASAP7_75t_R output1341 (.A(net1340),
    .Y(io_outs_left_0[39]));
 BUFx2_ASAP7_75t_R output1340 (.A(net1339),
    .Y(io_outs_left_0[38]));
 BUFx2_ASAP7_75t_R output1339 (.A(net1338),
    .Y(io_outs_left_0[37]));
 BUFx2_ASAP7_75t_R output1338 (.A(net1337),
    .Y(io_outs_left_0[36]));
 BUFx2_ASAP7_75t_R output1337 (.A(net1336),
    .Y(io_outs_left_0[35]));
 BUFx2_ASAP7_75t_R output1336 (.A(net1335),
    .Y(io_outs_left_0[34]));
 BUFx2_ASAP7_75t_R output1335 (.A(net1334),
    .Y(io_outs_left_0[33]));
 BUFx2_ASAP7_75t_R output1334 (.A(net1333),
    .Y(io_outs_left_0[32]));
 BUFx2_ASAP7_75t_R output1333 (.A(net1332),
    .Y(io_outs_left_0[31]));
 BUFx2_ASAP7_75t_R output1332 (.A(net1331),
    .Y(io_outs_left_0[30]));
 BUFx2_ASAP7_75t_R output1331 (.A(net1330),
    .Y(io_outs_left_0[2]));
 BUFx2_ASAP7_75t_R output1330 (.A(net1329),
    .Y(io_outs_left_0[29]));
 BUFx2_ASAP7_75t_R output1329 (.A(net1328),
    .Y(io_outs_left_0[28]));
 BUFx2_ASAP7_75t_R output1328 (.A(net1327),
    .Y(io_outs_left_0[27]));
 BUFx2_ASAP7_75t_R output1327 (.A(net1326),
    .Y(io_outs_left_0[26]));
 BUFx2_ASAP7_75t_R output1326 (.A(net1325),
    .Y(io_outs_left_0[25]));
 BUFx2_ASAP7_75t_R output1325 (.A(net1324),
    .Y(io_outs_left_0[24]));
 BUFx2_ASAP7_75t_R output1324 (.A(net1323),
    .Y(io_outs_left_0[23]));
 BUFx2_ASAP7_75t_R output1323 (.A(net1322),
    .Y(io_outs_left_0[22]));
 BUFx2_ASAP7_75t_R output1322 (.A(net1321),
    .Y(io_outs_left_0[21]));
 BUFx2_ASAP7_75t_R output1321 (.A(net1320),
    .Y(io_outs_left_0[20]));
 BUFx2_ASAP7_75t_R output1320 (.A(net1319),
    .Y(io_outs_left_0[1]));
 BUFx2_ASAP7_75t_R output1319 (.A(net1318),
    .Y(io_outs_left_0[19]));
 BUFx2_ASAP7_75t_R output1318 (.A(net1317),
    .Y(io_outs_left_0[18]));
 BUFx2_ASAP7_75t_R output1317 (.A(net1316),
    .Y(io_outs_left_0[17]));
 BUFx2_ASAP7_75t_R output1316 (.A(net1315),
    .Y(io_outs_left_0[16]));
 BUFx2_ASAP7_75t_R output1315 (.A(net1314),
    .Y(io_outs_left_0[15]));
 BUFx2_ASAP7_75t_R output1314 (.A(net1313),
    .Y(io_outs_left_0[14]));
 BUFx2_ASAP7_75t_R output1313 (.A(net1312),
    .Y(io_outs_left_0[13]));
 BUFx2_ASAP7_75t_R output1312 (.A(net1311),
    .Y(io_outs_left_0[12]));
 BUFx2_ASAP7_75t_R output1311 (.A(net1310),
    .Y(io_outs_left_0[11]));
 BUFx2_ASAP7_75t_R output1310 (.A(net1309),
    .Y(io_outs_left_0[10]));
 BUFx2_ASAP7_75t_R output1309 (.A(net1308),
    .Y(io_outs_left_0[0]));
 BUFx2_ASAP7_75t_R output1308 (.A(net1307),
    .Y(io_outs_down_3[9]));
 BUFx2_ASAP7_75t_R output1307 (.A(net1306),
    .Y(io_outs_down_3[8]));
 BUFx2_ASAP7_75t_R output1306 (.A(net1305),
    .Y(io_outs_down_3[7]));
 BUFx2_ASAP7_75t_R output1305 (.A(net1304),
    .Y(io_outs_down_3[6]));
 BUFx2_ASAP7_75t_R output1304 (.A(net1303),
    .Y(io_outs_down_3[63]));
 BUFx2_ASAP7_75t_R output1303 (.A(net1302),
    .Y(io_outs_down_3[62]));
 BUFx2_ASAP7_75t_R output1302 (.A(net1301),
    .Y(io_outs_down_3[61]));
 BUFx2_ASAP7_75t_R output1301 (.A(net1300),
    .Y(io_outs_down_3[60]));
 BUFx2_ASAP7_75t_R output1300 (.A(net1299),
    .Y(io_outs_down_3[5]));
 BUFx2_ASAP7_75t_R output1299 (.A(net1298),
    .Y(io_outs_down_3[59]));
 BUFx2_ASAP7_75t_R output1298 (.A(net1297),
    .Y(io_outs_down_3[58]));
 BUFx2_ASAP7_75t_R output1297 (.A(net1296),
    .Y(io_outs_down_3[57]));
 BUFx2_ASAP7_75t_R output1296 (.A(net1295),
    .Y(io_outs_down_3[56]));
 BUFx2_ASAP7_75t_R output1295 (.A(net1294),
    .Y(io_outs_down_3[55]));
 BUFx2_ASAP7_75t_R output1294 (.A(net1293),
    .Y(io_outs_down_3[54]));
 BUFx2_ASAP7_75t_R output1293 (.A(net1292),
    .Y(io_outs_down_3[53]));
 BUFx2_ASAP7_75t_R output1292 (.A(net1291),
    .Y(io_outs_down_3[52]));
 BUFx2_ASAP7_75t_R output1291 (.A(net1290),
    .Y(io_outs_down_3[51]));
 BUFx2_ASAP7_75t_R output1290 (.A(net1289),
    .Y(io_outs_down_3[50]));
 BUFx2_ASAP7_75t_R output1289 (.A(net1288),
    .Y(io_outs_down_3[4]));
 BUFx2_ASAP7_75t_R output1288 (.A(net1287),
    .Y(io_outs_down_3[49]));
 BUFx2_ASAP7_75t_R output1287 (.A(net1286),
    .Y(io_outs_down_3[48]));
 BUFx2_ASAP7_75t_R output1286 (.A(net1285),
    .Y(io_outs_down_3[47]));
 BUFx2_ASAP7_75t_R output1285 (.A(net1284),
    .Y(io_outs_down_3[46]));
 BUFx2_ASAP7_75t_R output1284 (.A(net1283),
    .Y(io_outs_down_3[45]));
 BUFx2_ASAP7_75t_R output1283 (.A(net1282),
    .Y(io_outs_down_3[44]));
 BUFx2_ASAP7_75t_R output1282 (.A(net1281),
    .Y(io_outs_down_3[43]));
 BUFx2_ASAP7_75t_R output1281 (.A(net1280),
    .Y(io_outs_down_3[42]));
 BUFx2_ASAP7_75t_R output1280 (.A(net1279),
    .Y(io_outs_down_3[41]));
 BUFx2_ASAP7_75t_R output1279 (.A(net1278),
    .Y(io_outs_down_3[40]));
 BUFx2_ASAP7_75t_R output1278 (.A(net1277),
    .Y(io_outs_down_3[3]));
 BUFx2_ASAP7_75t_R output1277 (.A(net1276),
    .Y(io_outs_down_3[39]));
 BUFx2_ASAP7_75t_R output1276 (.A(net1275),
    .Y(io_outs_down_3[38]));
 BUFx2_ASAP7_75t_R output1275 (.A(net1274),
    .Y(io_outs_down_3[37]));
 BUFx2_ASAP7_75t_R output1274 (.A(net1273),
    .Y(io_outs_down_3[36]));
 BUFx2_ASAP7_75t_R output1273 (.A(net1272),
    .Y(io_outs_down_3[35]));
 BUFx2_ASAP7_75t_R output1272 (.A(net1271),
    .Y(io_outs_down_3[34]));
 BUFx2_ASAP7_75t_R output1271 (.A(net1270),
    .Y(io_outs_down_3[33]));
 BUFx2_ASAP7_75t_R output1270 (.A(net1269),
    .Y(io_outs_down_3[32]));
 BUFx2_ASAP7_75t_R output1269 (.A(net1268),
    .Y(io_outs_down_3[31]));
 BUFx2_ASAP7_75t_R output1268 (.A(net1267),
    .Y(io_outs_down_3[30]));
 BUFx2_ASAP7_75t_R output1267 (.A(net1266),
    .Y(io_outs_down_3[2]));
 BUFx2_ASAP7_75t_R output1266 (.A(net1265),
    .Y(io_outs_down_3[29]));
 BUFx2_ASAP7_75t_R output1265 (.A(net1264),
    .Y(io_outs_down_3[28]));
 BUFx2_ASAP7_75t_R output1264 (.A(net1263),
    .Y(io_outs_down_3[27]));
 BUFx2_ASAP7_75t_R output1263 (.A(net1262),
    .Y(io_outs_down_3[26]));
 BUFx2_ASAP7_75t_R output1262 (.A(net1261),
    .Y(io_outs_down_3[25]));
 BUFx2_ASAP7_75t_R output1261 (.A(net1260),
    .Y(io_outs_down_3[24]));
 BUFx2_ASAP7_75t_R output1260 (.A(net1259),
    .Y(io_outs_down_3[23]));
 BUFx2_ASAP7_75t_R output1259 (.A(net1258),
    .Y(io_outs_down_3[22]));
 BUFx2_ASAP7_75t_R output1258 (.A(net1257),
    .Y(io_outs_down_3[21]));
 BUFx2_ASAP7_75t_R output1257 (.A(net1256),
    .Y(io_outs_down_3[20]));
 BUFx2_ASAP7_75t_R output1256 (.A(net1255),
    .Y(io_outs_down_3[1]));
 BUFx2_ASAP7_75t_R output1255 (.A(net1254),
    .Y(io_outs_down_3[19]));
 BUFx2_ASAP7_75t_R output1254 (.A(net1253),
    .Y(io_outs_down_3[18]));
 BUFx2_ASAP7_75t_R output1253 (.A(net1252),
    .Y(io_outs_down_3[17]));
 BUFx2_ASAP7_75t_R output1252 (.A(net1251),
    .Y(io_outs_down_3[16]));
 BUFx2_ASAP7_75t_R output1251 (.A(net1250),
    .Y(io_outs_down_3[15]));
 BUFx2_ASAP7_75t_R output1250 (.A(net1249),
    .Y(io_outs_down_3[14]));
 BUFx2_ASAP7_75t_R output1249 (.A(net1248),
    .Y(io_outs_down_3[13]));
 BUFx2_ASAP7_75t_R output1248 (.A(net1247),
    .Y(io_outs_down_3[12]));
 BUFx2_ASAP7_75t_R output1247 (.A(net1246),
    .Y(io_outs_down_3[11]));
 BUFx2_ASAP7_75t_R output1246 (.A(net1245),
    .Y(io_outs_down_3[10]));
 BUFx2_ASAP7_75t_R output1245 (.A(net1244),
    .Y(io_outs_down_3[0]));
 BUFx2_ASAP7_75t_R output1244 (.A(net1243),
    .Y(io_outs_down_2[9]));
 BUFx2_ASAP7_75t_R output1243 (.A(net1242),
    .Y(io_outs_down_2[8]));
 BUFx2_ASAP7_75t_R output1242 (.A(net1241),
    .Y(io_outs_down_2[7]));
 BUFx2_ASAP7_75t_R output1241 (.A(net1240),
    .Y(io_outs_down_2[6]));
 BUFx2_ASAP7_75t_R output1240 (.A(net1239),
    .Y(io_outs_down_2[63]));
 BUFx2_ASAP7_75t_R output1239 (.A(net1238),
    .Y(io_outs_down_2[62]));
 BUFx2_ASAP7_75t_R output1238 (.A(net1237),
    .Y(io_outs_down_2[61]));
 BUFx2_ASAP7_75t_R output1237 (.A(net1236),
    .Y(io_outs_down_2[60]));
 BUFx2_ASAP7_75t_R output1236 (.A(net1235),
    .Y(io_outs_down_2[5]));
 BUFx2_ASAP7_75t_R output1235 (.A(net1234),
    .Y(io_outs_down_2[59]));
 BUFx2_ASAP7_75t_R output1234 (.A(net1233),
    .Y(io_outs_down_2[58]));
 BUFx2_ASAP7_75t_R output1233 (.A(net1232),
    .Y(io_outs_down_2[57]));
 BUFx2_ASAP7_75t_R output1232 (.A(net1231),
    .Y(io_outs_down_2[56]));
 BUFx2_ASAP7_75t_R output1231 (.A(net1230),
    .Y(io_outs_down_2[55]));
 BUFx2_ASAP7_75t_R output1230 (.A(net1229),
    .Y(io_outs_down_2[54]));
 BUFx2_ASAP7_75t_R output1229 (.A(net1228),
    .Y(io_outs_down_2[53]));
 BUFx2_ASAP7_75t_R output1228 (.A(net1227),
    .Y(io_outs_down_2[52]));
 BUFx2_ASAP7_75t_R output1227 (.A(net1226),
    .Y(io_outs_down_2[51]));
 BUFx2_ASAP7_75t_R output1226 (.A(net1225),
    .Y(io_outs_down_2[50]));
 BUFx2_ASAP7_75t_R output1225 (.A(net1224),
    .Y(io_outs_down_2[4]));
 BUFx2_ASAP7_75t_R output1224 (.A(net1223),
    .Y(io_outs_down_2[49]));
 BUFx2_ASAP7_75t_R output1223 (.A(net1222),
    .Y(io_outs_down_2[48]));
 BUFx2_ASAP7_75t_R output1222 (.A(net1221),
    .Y(io_outs_down_2[47]));
 BUFx2_ASAP7_75t_R output1221 (.A(net1220),
    .Y(io_outs_down_2[46]));
 BUFx2_ASAP7_75t_R output1220 (.A(net1219),
    .Y(io_outs_down_2[45]));
 BUFx2_ASAP7_75t_R output1219 (.A(net1218),
    .Y(io_outs_down_2[44]));
 BUFx2_ASAP7_75t_R output1218 (.A(net1217),
    .Y(io_outs_down_2[43]));
 BUFx2_ASAP7_75t_R output1217 (.A(net1216),
    .Y(io_outs_down_2[42]));
 BUFx2_ASAP7_75t_R output1216 (.A(net1215),
    .Y(io_outs_down_2[41]));
 BUFx2_ASAP7_75t_R output1215 (.A(net1214),
    .Y(io_outs_down_2[40]));
 BUFx2_ASAP7_75t_R output1214 (.A(net1213),
    .Y(io_outs_down_2[3]));
 BUFx2_ASAP7_75t_R output1213 (.A(net1212),
    .Y(io_outs_down_2[39]));
 BUFx2_ASAP7_75t_R output1212 (.A(net1211),
    .Y(io_outs_down_2[38]));
 BUFx2_ASAP7_75t_R output1211 (.A(net1210),
    .Y(io_outs_down_2[37]));
 BUFx2_ASAP7_75t_R output1210 (.A(net1209),
    .Y(io_outs_down_2[36]));
 BUFx2_ASAP7_75t_R output1209 (.A(net1208),
    .Y(io_outs_down_2[35]));
 BUFx2_ASAP7_75t_R output1208 (.A(net1207),
    .Y(io_outs_down_2[34]));
 BUFx2_ASAP7_75t_R output1207 (.A(net1206),
    .Y(io_outs_down_2[33]));
 BUFx2_ASAP7_75t_R output1206 (.A(net1205),
    .Y(io_outs_down_2[32]));
 BUFx2_ASAP7_75t_R output1205 (.A(net1204),
    .Y(io_outs_down_2[31]));
 BUFx2_ASAP7_75t_R output1204 (.A(net1203),
    .Y(io_outs_down_2[30]));
 BUFx2_ASAP7_75t_R output1203 (.A(net1202),
    .Y(io_outs_down_2[2]));
 BUFx2_ASAP7_75t_R output1202 (.A(net1201),
    .Y(io_outs_down_2[29]));
 BUFx2_ASAP7_75t_R output1201 (.A(net1200),
    .Y(io_outs_down_2[28]));
 BUFx2_ASAP7_75t_R output1200 (.A(net1199),
    .Y(io_outs_down_2[27]));
 BUFx2_ASAP7_75t_R output1199 (.A(net1198),
    .Y(io_outs_down_2[26]));
 BUFx2_ASAP7_75t_R output1198 (.A(net1197),
    .Y(io_outs_down_2[25]));
 BUFx2_ASAP7_75t_R output1197 (.A(net1196),
    .Y(io_outs_down_2[24]));
 BUFx2_ASAP7_75t_R output1196 (.A(net1195),
    .Y(io_outs_down_2[23]));
 BUFx2_ASAP7_75t_R output1195 (.A(net1194),
    .Y(io_outs_down_2[22]));
 BUFx2_ASAP7_75t_R output1194 (.A(net1193),
    .Y(io_outs_down_2[21]));
 BUFx2_ASAP7_75t_R output1193 (.A(net1192),
    .Y(io_outs_down_2[20]));
 BUFx2_ASAP7_75t_R output1192 (.A(net1191),
    .Y(io_outs_down_2[1]));
 BUFx2_ASAP7_75t_R output1191 (.A(net1190),
    .Y(io_outs_down_2[19]));
 BUFx2_ASAP7_75t_R output1190 (.A(net1189),
    .Y(io_outs_down_2[18]));
 BUFx2_ASAP7_75t_R output1189 (.A(net1188),
    .Y(io_outs_down_2[17]));
 BUFx2_ASAP7_75t_R output1188 (.A(net1187),
    .Y(io_outs_down_2[16]));
 BUFx2_ASAP7_75t_R output1187 (.A(net1186),
    .Y(io_outs_down_2[15]));
 BUFx2_ASAP7_75t_R output1186 (.A(net1185),
    .Y(io_outs_down_2[14]));
 BUFx2_ASAP7_75t_R output1185 (.A(net1184),
    .Y(io_outs_down_2[13]));
 BUFx2_ASAP7_75t_R output1184 (.A(net1183),
    .Y(io_outs_down_2[12]));
 BUFx2_ASAP7_75t_R output1183 (.A(net1182),
    .Y(io_outs_down_2[11]));
 BUFx2_ASAP7_75t_R output1182 (.A(net1181),
    .Y(io_outs_down_2[10]));
 BUFx2_ASAP7_75t_R output1181 (.A(net1180),
    .Y(io_outs_down_2[0]));
 BUFx2_ASAP7_75t_R output1180 (.A(net1179),
    .Y(io_outs_down_1[9]));
 BUFx2_ASAP7_75t_R output1179 (.A(net1178),
    .Y(io_outs_down_1[8]));
 BUFx2_ASAP7_75t_R output1178 (.A(net1177),
    .Y(io_outs_down_1[7]));
 BUFx2_ASAP7_75t_R output1177 (.A(net1176),
    .Y(io_outs_down_1[6]));
 BUFx2_ASAP7_75t_R output1176 (.A(net1175),
    .Y(io_outs_down_1[63]));
 BUFx2_ASAP7_75t_R output1175 (.A(net1174),
    .Y(io_outs_down_1[62]));
 BUFx2_ASAP7_75t_R output1174 (.A(net1173),
    .Y(io_outs_down_1[61]));
 BUFx2_ASAP7_75t_R output1173 (.A(net1172),
    .Y(io_outs_down_1[60]));
 BUFx2_ASAP7_75t_R output1172 (.A(net1171),
    .Y(io_outs_down_1[5]));
 BUFx2_ASAP7_75t_R output1171 (.A(net1170),
    .Y(io_outs_down_1[59]));
 BUFx2_ASAP7_75t_R output1170 (.A(net1169),
    .Y(io_outs_down_1[58]));
 BUFx2_ASAP7_75t_R output1169 (.A(net1168),
    .Y(io_outs_down_1[57]));
 BUFx2_ASAP7_75t_R output1168 (.A(net1167),
    .Y(io_outs_down_1[56]));
 BUFx2_ASAP7_75t_R output1167 (.A(net1166),
    .Y(io_outs_down_1[55]));
 BUFx2_ASAP7_75t_R output1166 (.A(net1165),
    .Y(io_outs_down_1[54]));
 BUFx2_ASAP7_75t_R output1165 (.A(net1164),
    .Y(io_outs_down_1[53]));
 BUFx2_ASAP7_75t_R output1164 (.A(net1163),
    .Y(io_outs_down_1[52]));
 BUFx2_ASAP7_75t_R output1163 (.A(net1162),
    .Y(io_outs_down_1[51]));
 BUFx2_ASAP7_75t_R output1162 (.A(net1161),
    .Y(io_outs_down_1[50]));
 BUFx2_ASAP7_75t_R output1161 (.A(net1160),
    .Y(io_outs_down_1[4]));
 BUFx2_ASAP7_75t_R output1160 (.A(net1159),
    .Y(io_outs_down_1[49]));
 BUFx2_ASAP7_75t_R output1159 (.A(net1158),
    .Y(io_outs_down_1[48]));
 BUFx2_ASAP7_75t_R output1158 (.A(net1157),
    .Y(io_outs_down_1[47]));
 BUFx2_ASAP7_75t_R output1157 (.A(net1156),
    .Y(io_outs_down_1[46]));
 BUFx2_ASAP7_75t_R output1156 (.A(net1155),
    .Y(io_outs_down_1[45]));
 BUFx2_ASAP7_75t_R output1155 (.A(net1154),
    .Y(io_outs_down_1[44]));
 BUFx2_ASAP7_75t_R output1154 (.A(net1153),
    .Y(io_outs_down_1[43]));
 BUFx2_ASAP7_75t_R output1153 (.A(net1152),
    .Y(io_outs_down_1[42]));
 BUFx2_ASAP7_75t_R output1152 (.A(net1151),
    .Y(io_outs_down_1[41]));
 BUFx2_ASAP7_75t_R output1151 (.A(net1150),
    .Y(io_outs_down_1[40]));
 BUFx2_ASAP7_75t_R output1150 (.A(net1149),
    .Y(io_outs_down_1[3]));
 BUFx2_ASAP7_75t_R output1149 (.A(net1148),
    .Y(io_outs_down_1[39]));
 BUFx2_ASAP7_75t_R output1148 (.A(net1147),
    .Y(io_outs_down_1[38]));
 BUFx2_ASAP7_75t_R output1147 (.A(net1146),
    .Y(io_outs_down_1[37]));
 BUFx2_ASAP7_75t_R output1146 (.A(net1145),
    .Y(io_outs_down_1[36]));
 BUFx2_ASAP7_75t_R output1145 (.A(net1144),
    .Y(io_outs_down_1[35]));
 BUFx2_ASAP7_75t_R output1144 (.A(net1143),
    .Y(io_outs_down_1[34]));
 BUFx2_ASAP7_75t_R output1143 (.A(net1142),
    .Y(io_outs_down_1[33]));
 BUFx2_ASAP7_75t_R output1142 (.A(net1141),
    .Y(io_outs_down_1[32]));
 BUFx2_ASAP7_75t_R output1141 (.A(net1140),
    .Y(io_outs_down_1[31]));
 BUFx2_ASAP7_75t_R output1140 (.A(net1139),
    .Y(io_outs_down_1[30]));
 BUFx2_ASAP7_75t_R output1139 (.A(net1138),
    .Y(io_outs_down_1[2]));
 BUFx2_ASAP7_75t_R output1138 (.A(net1137),
    .Y(io_outs_down_1[29]));
 BUFx2_ASAP7_75t_R output1137 (.A(net1136),
    .Y(io_outs_down_1[28]));
 BUFx2_ASAP7_75t_R output1136 (.A(net1135),
    .Y(io_outs_down_1[27]));
 BUFx2_ASAP7_75t_R output1135 (.A(net1134),
    .Y(io_outs_down_1[26]));
 BUFx2_ASAP7_75t_R output1134 (.A(net1133),
    .Y(io_outs_down_1[25]));
 BUFx2_ASAP7_75t_R output1133 (.A(net1132),
    .Y(io_outs_down_1[24]));
 BUFx2_ASAP7_75t_R output1132 (.A(net1131),
    .Y(io_outs_down_1[23]));
 BUFx2_ASAP7_75t_R output1131 (.A(net1130),
    .Y(io_outs_down_1[22]));
 BUFx2_ASAP7_75t_R output1130 (.A(net1129),
    .Y(io_outs_down_1[21]));
 BUFx2_ASAP7_75t_R output1129 (.A(net1128),
    .Y(io_outs_down_1[20]));
 BUFx2_ASAP7_75t_R output1128 (.A(net1127),
    .Y(io_outs_down_1[1]));
 BUFx2_ASAP7_75t_R output1127 (.A(net1126),
    .Y(io_outs_down_1[19]));
 BUFx2_ASAP7_75t_R output1126 (.A(net1125),
    .Y(io_outs_down_1[18]));
 BUFx2_ASAP7_75t_R output1125 (.A(net1124),
    .Y(io_outs_down_1[17]));
 BUFx2_ASAP7_75t_R output1124 (.A(net1123),
    .Y(io_outs_down_1[16]));
 BUFx2_ASAP7_75t_R output1123 (.A(net1122),
    .Y(io_outs_down_1[15]));
 BUFx2_ASAP7_75t_R output1122 (.A(net1121),
    .Y(io_outs_down_1[14]));
 BUFx2_ASAP7_75t_R output1121 (.A(net1120),
    .Y(io_outs_down_1[13]));
 BUFx2_ASAP7_75t_R output1120 (.A(net1119),
    .Y(io_outs_down_1[12]));
 BUFx2_ASAP7_75t_R output1119 (.A(net1118),
    .Y(io_outs_down_1[11]));
 BUFx2_ASAP7_75t_R output1118 (.A(net1117),
    .Y(io_outs_down_1[10]));
 BUFx2_ASAP7_75t_R output1117 (.A(net1116),
    .Y(io_outs_down_1[0]));
 BUFx2_ASAP7_75t_R output1116 (.A(net1115),
    .Y(io_outs_down_0[9]));
 BUFx2_ASAP7_75t_R output1115 (.A(net1114),
    .Y(io_outs_down_0[8]));
 BUFx2_ASAP7_75t_R output1114 (.A(net1113),
    .Y(io_outs_down_0[7]));
 BUFx2_ASAP7_75t_R output1113 (.A(net1112),
    .Y(io_outs_down_0[6]));
 BUFx2_ASAP7_75t_R output1112 (.A(net1111),
    .Y(io_outs_down_0[63]));
 BUFx2_ASAP7_75t_R output1111 (.A(net1110),
    .Y(io_outs_down_0[62]));
 BUFx2_ASAP7_75t_R output1110 (.A(net1109),
    .Y(io_outs_down_0[61]));
 BUFx2_ASAP7_75t_R output1109 (.A(net1108),
    .Y(io_outs_down_0[60]));
 BUFx2_ASAP7_75t_R output1108 (.A(net1107),
    .Y(io_outs_down_0[5]));
 BUFx2_ASAP7_75t_R output1107 (.A(net1106),
    .Y(io_outs_down_0[59]));
 BUFx2_ASAP7_75t_R output1106 (.A(net1105),
    .Y(io_outs_down_0[58]));
 BUFx2_ASAP7_75t_R output1105 (.A(net1104),
    .Y(io_outs_down_0[57]));
 BUFx2_ASAP7_75t_R output1104 (.A(net1103),
    .Y(io_outs_down_0[56]));
 BUFx2_ASAP7_75t_R output1103 (.A(net1102),
    .Y(io_outs_down_0[55]));
 BUFx2_ASAP7_75t_R output1102 (.A(net1101),
    .Y(io_outs_down_0[54]));
 BUFx2_ASAP7_75t_R output1101 (.A(net1100),
    .Y(io_outs_down_0[53]));
 BUFx2_ASAP7_75t_R output1100 (.A(net1099),
    .Y(io_outs_down_0[52]));
 BUFx2_ASAP7_75t_R output1099 (.A(net1098),
    .Y(io_outs_down_0[51]));
 BUFx2_ASAP7_75t_R output1098 (.A(net1097),
    .Y(io_outs_down_0[50]));
 BUFx2_ASAP7_75t_R output1097 (.A(net1096),
    .Y(io_outs_down_0[4]));
 BUFx2_ASAP7_75t_R output1096 (.A(net1095),
    .Y(io_outs_down_0[49]));
 BUFx2_ASAP7_75t_R output1095 (.A(net1094),
    .Y(io_outs_down_0[48]));
 BUFx2_ASAP7_75t_R output1094 (.A(net1093),
    .Y(io_outs_down_0[47]));
 BUFx2_ASAP7_75t_R output1093 (.A(net1092),
    .Y(io_outs_down_0[46]));
 BUFx2_ASAP7_75t_R output1092 (.A(net1091),
    .Y(io_outs_down_0[45]));
 BUFx2_ASAP7_75t_R output1091 (.A(net1090),
    .Y(io_outs_down_0[44]));
 BUFx2_ASAP7_75t_R output1090 (.A(net1089),
    .Y(io_outs_down_0[43]));
 BUFx2_ASAP7_75t_R output1089 (.A(net1088),
    .Y(io_outs_down_0[42]));
 BUFx2_ASAP7_75t_R output1088 (.A(net1087),
    .Y(io_outs_down_0[41]));
 BUFx2_ASAP7_75t_R output1087 (.A(net1086),
    .Y(io_outs_down_0[40]));
 BUFx2_ASAP7_75t_R output1086 (.A(net1085),
    .Y(io_outs_down_0[3]));
 BUFx2_ASAP7_75t_R output1085 (.A(net1084),
    .Y(io_outs_down_0[39]));
 BUFx2_ASAP7_75t_R output1084 (.A(net1083),
    .Y(io_outs_down_0[38]));
 BUFx2_ASAP7_75t_R output1083 (.A(net1082),
    .Y(io_outs_down_0[37]));
 BUFx2_ASAP7_75t_R output1082 (.A(net1081),
    .Y(io_outs_down_0[36]));
 BUFx2_ASAP7_75t_R output1081 (.A(net1080),
    .Y(io_outs_down_0[35]));
 BUFx2_ASAP7_75t_R output1080 (.A(net1079),
    .Y(io_outs_down_0[34]));
 BUFx2_ASAP7_75t_R output1079 (.A(net1078),
    .Y(io_outs_down_0[33]));
 BUFx2_ASAP7_75t_R output1078 (.A(net1077),
    .Y(io_outs_down_0[32]));
 BUFx2_ASAP7_75t_R output1077 (.A(net1076),
    .Y(io_outs_down_0[31]));
 BUFx2_ASAP7_75t_R output1076 (.A(net1075),
    .Y(io_outs_down_0[30]));
 BUFx2_ASAP7_75t_R output1075 (.A(net1074),
    .Y(io_outs_down_0[2]));
 BUFx2_ASAP7_75t_R output1074 (.A(net1073),
    .Y(io_outs_down_0[29]));
 BUFx2_ASAP7_75t_R output1073 (.A(net1072),
    .Y(io_outs_down_0[28]));
 BUFx2_ASAP7_75t_R output1072 (.A(net1071),
    .Y(io_outs_down_0[27]));
 BUFx2_ASAP7_75t_R output1071 (.A(net1070),
    .Y(io_outs_down_0[26]));
 BUFx2_ASAP7_75t_R output1070 (.A(net1069),
    .Y(io_outs_down_0[25]));
 BUFx2_ASAP7_75t_R output1069 (.A(net1068),
    .Y(io_outs_down_0[24]));
 BUFx2_ASAP7_75t_R output1068 (.A(net1067),
    .Y(io_outs_down_0[23]));
 BUFx2_ASAP7_75t_R output1067 (.A(net1066),
    .Y(io_outs_down_0[22]));
 BUFx2_ASAP7_75t_R output1066 (.A(net1065),
    .Y(io_outs_down_0[21]));
 BUFx2_ASAP7_75t_R output1065 (.A(net1064),
    .Y(io_outs_down_0[20]));
 BUFx2_ASAP7_75t_R output1064 (.A(net1063),
    .Y(io_outs_down_0[1]));
 BUFx2_ASAP7_75t_R output1063 (.A(net1062),
    .Y(io_outs_down_0[19]));
 BUFx2_ASAP7_75t_R output1062 (.A(net1061),
    .Y(io_outs_down_0[18]));
 BUFx2_ASAP7_75t_R output1061 (.A(net1060),
    .Y(io_outs_down_0[17]));
 BUFx2_ASAP7_75t_R output1060 (.A(net1059),
    .Y(io_outs_down_0[16]));
 BUFx2_ASAP7_75t_R output1059 (.A(net1058),
    .Y(io_outs_down_0[15]));
 BUFx2_ASAP7_75t_R output1058 (.A(net1057),
    .Y(io_outs_down_0[14]));
 BUFx2_ASAP7_75t_R output1057 (.A(net1056),
    .Y(io_outs_down_0[13]));
 BUFx2_ASAP7_75t_R output1056 (.A(net1055),
    .Y(io_outs_down_0[12]));
 BUFx2_ASAP7_75t_R output1055 (.A(net1054),
    .Y(io_outs_down_0[11]));
 BUFx2_ASAP7_75t_R output1054 (.A(net1053),
    .Y(io_outs_down_0[10]));
 BUFx2_ASAP7_75t_R output1053 (.A(net1052),
    .Y(io_outs_down_0[0]));
 BUFx2_ASAP7_75t_R output1052 (.A(net1051),
    .Y(io_lsbs_9));
 BUFx2_ASAP7_75t_R output1051 (.A(net1050),
    .Y(io_lsbs_8));
 BUFx2_ASAP7_75t_R output1050 (.A(net1049),
    .Y(io_lsbs_7));
 BUFx2_ASAP7_75t_R output1049 (.A(net1048),
    .Y(io_lsbs_6));
 BUFx2_ASAP7_75t_R output1048 (.A(net1047),
    .Y(io_lsbs_5));
 BUFx2_ASAP7_75t_R output1047 (.A(net1046),
    .Y(io_lsbs_4));
 BUFx2_ASAP7_75t_R output1046 (.A(net1045),
    .Y(io_lsbs_3));
 BUFx2_ASAP7_75t_R output1045 (.A(net1044),
    .Y(io_lsbs_2));
 BUFx2_ASAP7_75t_R output1044 (.A(net1043),
    .Y(io_lsbs_15));
 BUFx2_ASAP7_75t_R output1043 (.A(net1042),
    .Y(io_lsbs_14));
 BUFx2_ASAP7_75t_R output1042 (.A(net1041),
    .Y(io_lsbs_13));
 BUFx2_ASAP7_75t_R output1041 (.A(net1040),
    .Y(io_lsbs_12));
 BUFx2_ASAP7_75t_R output1040 (.A(net1039),
    .Y(io_lsbs_11));
 BUFx2_ASAP7_75t_R output1039 (.A(net1038),
    .Y(io_lsbs_10));
 BUFx2_ASAP7_75t_R output1038 (.A(net1037),
    .Y(io_lsbs_1));
 BUFx2_ASAP7_75t_R output1037 (.A(net1036),
    .Y(io_lsbs_0));
 BUFx2_ASAP7_75t_R input1036 (.A(io_ins_up_3[9]),
    .Y(net1035));
 BUFx2_ASAP7_75t_R input1035 (.A(io_ins_up_3[8]),
    .Y(net1034));
 BUFx2_ASAP7_75t_R input1034 (.A(io_ins_up_3[7]),
    .Y(net1033));
 BUFx2_ASAP7_75t_R input1033 (.A(io_ins_up_3[6]),
    .Y(net1032));
 BUFx2_ASAP7_75t_R input1032 (.A(io_ins_up_3[63]),
    .Y(net1031));
 BUFx2_ASAP7_75t_R input1031 (.A(io_ins_up_3[62]),
    .Y(net1030));
 BUFx2_ASAP7_75t_R input1030 (.A(io_ins_up_3[61]),
    .Y(net1029));
 BUFx2_ASAP7_75t_R input1029 (.A(io_ins_up_3[60]),
    .Y(net1028));
 BUFx2_ASAP7_75t_R input1028 (.A(io_ins_up_3[5]),
    .Y(net1027));
 BUFx2_ASAP7_75t_R input1027 (.A(io_ins_up_3[59]),
    .Y(net1026));
 BUFx2_ASAP7_75t_R input1026 (.A(io_ins_up_3[58]),
    .Y(net1025));
 BUFx2_ASAP7_75t_R input1025 (.A(io_ins_up_3[57]),
    .Y(net1024));
 BUFx2_ASAP7_75t_R input1024 (.A(io_ins_up_3[56]),
    .Y(net1023));
 BUFx2_ASAP7_75t_R input1023 (.A(io_ins_up_3[55]),
    .Y(net1022));
 BUFx2_ASAP7_75t_R input1022 (.A(io_ins_up_3[54]),
    .Y(net1021));
 BUFx2_ASAP7_75t_R input1021 (.A(io_ins_up_3[53]),
    .Y(net1020));
 BUFx2_ASAP7_75t_R input1020 (.A(io_ins_up_3[52]),
    .Y(net1019));
 BUFx2_ASAP7_75t_R input1019 (.A(io_ins_up_3[51]),
    .Y(net1018));
 BUFx2_ASAP7_75t_R input1018 (.A(io_ins_up_3[50]),
    .Y(net1017));
 BUFx2_ASAP7_75t_R input1017 (.A(io_ins_up_3[4]),
    .Y(net1016));
 BUFx2_ASAP7_75t_R input1016 (.A(io_ins_up_3[49]),
    .Y(net1015));
 BUFx2_ASAP7_75t_R input1015 (.A(io_ins_up_3[48]),
    .Y(net1014));
 BUFx2_ASAP7_75t_R input1014 (.A(io_ins_up_3[47]),
    .Y(net1013));
 BUFx2_ASAP7_75t_R input1013 (.A(io_ins_up_3[46]),
    .Y(net1012));
 BUFx2_ASAP7_75t_R input1012 (.A(io_ins_up_3[45]),
    .Y(net1011));
 BUFx2_ASAP7_75t_R input1011 (.A(io_ins_up_3[44]),
    .Y(net1010));
 BUFx2_ASAP7_75t_R input1010 (.A(io_ins_up_3[43]),
    .Y(net1009));
 BUFx2_ASAP7_75t_R input1009 (.A(io_ins_up_3[42]),
    .Y(net1008));
 BUFx2_ASAP7_75t_R input1008 (.A(io_ins_up_3[41]),
    .Y(net1007));
 BUFx2_ASAP7_75t_R input1007 (.A(io_ins_up_3[40]),
    .Y(net1006));
 BUFx2_ASAP7_75t_R input1006 (.A(io_ins_up_3[3]),
    .Y(net1005));
 BUFx2_ASAP7_75t_R input1005 (.A(io_ins_up_3[39]),
    .Y(net1004));
 BUFx2_ASAP7_75t_R input1004 (.A(io_ins_up_3[38]),
    .Y(net1003));
 BUFx2_ASAP7_75t_R input1003 (.A(io_ins_up_3[37]),
    .Y(net1002));
 BUFx2_ASAP7_75t_R input1002 (.A(io_ins_up_3[36]),
    .Y(net1001));
 BUFx2_ASAP7_75t_R input1001 (.A(io_ins_up_3[35]),
    .Y(net1000));
 BUFx2_ASAP7_75t_R input1000 (.A(io_ins_up_3[34]),
    .Y(net999));
 BUFx2_ASAP7_75t_R input999 (.A(io_ins_up_3[33]),
    .Y(net998));
 BUFx2_ASAP7_75t_R input998 (.A(io_ins_up_3[32]),
    .Y(net997));
 BUFx2_ASAP7_75t_R input997 (.A(io_ins_up_3[31]),
    .Y(net996));
 BUFx2_ASAP7_75t_R input996 (.A(io_ins_up_3[30]),
    .Y(net995));
 BUFx2_ASAP7_75t_R input995 (.A(io_ins_up_3[2]),
    .Y(net994));
 BUFx2_ASAP7_75t_R input994 (.A(io_ins_up_3[29]),
    .Y(net993));
 BUFx2_ASAP7_75t_R input993 (.A(io_ins_up_3[28]),
    .Y(net992));
 BUFx2_ASAP7_75t_R input992 (.A(io_ins_up_3[27]),
    .Y(net991));
 BUFx2_ASAP7_75t_R input991 (.A(io_ins_up_3[26]),
    .Y(net990));
 BUFx2_ASAP7_75t_R input990 (.A(io_ins_up_3[25]),
    .Y(net989));
 BUFx2_ASAP7_75t_R input989 (.A(io_ins_up_3[24]),
    .Y(net988));
 BUFx2_ASAP7_75t_R input988 (.A(io_ins_up_3[23]),
    .Y(net987));
 BUFx2_ASAP7_75t_R input987 (.A(io_ins_up_3[22]),
    .Y(net986));
 BUFx2_ASAP7_75t_R input986 (.A(io_ins_up_3[21]),
    .Y(net985));
 BUFx2_ASAP7_75t_R input985 (.A(io_ins_up_3[20]),
    .Y(net984));
 BUFx2_ASAP7_75t_R input984 (.A(io_ins_up_3[1]),
    .Y(net983));
 BUFx2_ASAP7_75t_R input983 (.A(io_ins_up_3[19]),
    .Y(net982));
 BUFx2_ASAP7_75t_R input982 (.A(io_ins_up_3[18]),
    .Y(net981));
 BUFx2_ASAP7_75t_R input981 (.A(io_ins_up_3[17]),
    .Y(net980));
 BUFx2_ASAP7_75t_R input980 (.A(io_ins_up_3[16]),
    .Y(net979));
 BUFx2_ASAP7_75t_R input979 (.A(io_ins_up_3[15]),
    .Y(net978));
 BUFx2_ASAP7_75t_R input978 (.A(io_ins_up_3[14]),
    .Y(net977));
 BUFx2_ASAP7_75t_R input977 (.A(io_ins_up_3[13]),
    .Y(net976));
 BUFx2_ASAP7_75t_R input976 (.A(io_ins_up_3[12]),
    .Y(net975));
 BUFx2_ASAP7_75t_R input975 (.A(io_ins_up_3[11]),
    .Y(net974));
 BUFx2_ASAP7_75t_R input974 (.A(io_ins_up_3[10]),
    .Y(net973));
 BUFx2_ASAP7_75t_R input973 (.A(io_ins_up_3[0]),
    .Y(net972));
 BUFx2_ASAP7_75t_R input972 (.A(io_ins_up_2[9]),
    .Y(net971));
 BUFx2_ASAP7_75t_R input971 (.A(io_ins_up_2[8]),
    .Y(net970));
 BUFx2_ASAP7_75t_R input970 (.A(io_ins_up_2[7]),
    .Y(net969));
 BUFx2_ASAP7_75t_R input969 (.A(io_ins_up_2[6]),
    .Y(net968));
 BUFx2_ASAP7_75t_R input968 (.A(io_ins_up_2[63]),
    .Y(net967));
 BUFx2_ASAP7_75t_R input967 (.A(io_ins_up_2[62]),
    .Y(net966));
 BUFx2_ASAP7_75t_R input966 (.A(io_ins_up_2[61]),
    .Y(net965));
 BUFx2_ASAP7_75t_R input965 (.A(io_ins_up_2[60]),
    .Y(net964));
 BUFx2_ASAP7_75t_R input964 (.A(io_ins_up_2[5]),
    .Y(net963));
 BUFx2_ASAP7_75t_R input963 (.A(io_ins_up_2[59]),
    .Y(net962));
 BUFx2_ASAP7_75t_R input962 (.A(io_ins_up_2[58]),
    .Y(net961));
 BUFx2_ASAP7_75t_R input961 (.A(io_ins_up_2[57]),
    .Y(net960));
 BUFx2_ASAP7_75t_R input960 (.A(io_ins_up_2[56]),
    .Y(net959));
 BUFx2_ASAP7_75t_R input959 (.A(io_ins_up_2[55]),
    .Y(net958));
 BUFx2_ASAP7_75t_R input958 (.A(io_ins_up_2[54]),
    .Y(net957));
 BUFx2_ASAP7_75t_R input957 (.A(io_ins_up_2[53]),
    .Y(net956));
 BUFx2_ASAP7_75t_R input956 (.A(io_ins_up_2[52]),
    .Y(net955));
 BUFx2_ASAP7_75t_R input955 (.A(io_ins_up_2[51]),
    .Y(net954));
 BUFx2_ASAP7_75t_R input954 (.A(io_ins_up_2[50]),
    .Y(net953));
 BUFx2_ASAP7_75t_R input953 (.A(io_ins_up_2[4]),
    .Y(net952));
 BUFx2_ASAP7_75t_R input952 (.A(io_ins_up_2[49]),
    .Y(net951));
 BUFx2_ASAP7_75t_R input951 (.A(io_ins_up_2[48]),
    .Y(net950));
 BUFx2_ASAP7_75t_R input950 (.A(io_ins_up_2[47]),
    .Y(net949));
 BUFx2_ASAP7_75t_R input949 (.A(io_ins_up_2[46]),
    .Y(net948));
 BUFx2_ASAP7_75t_R input948 (.A(io_ins_up_2[45]),
    .Y(net947));
 BUFx2_ASAP7_75t_R input947 (.A(io_ins_up_2[44]),
    .Y(net946));
 BUFx2_ASAP7_75t_R input946 (.A(io_ins_up_2[43]),
    .Y(net945));
 BUFx2_ASAP7_75t_R input945 (.A(io_ins_up_2[42]),
    .Y(net944));
 BUFx2_ASAP7_75t_R input944 (.A(io_ins_up_2[41]),
    .Y(net943));
 BUFx2_ASAP7_75t_R input943 (.A(io_ins_up_2[40]),
    .Y(net942));
 BUFx2_ASAP7_75t_R input942 (.A(io_ins_up_2[3]),
    .Y(net941));
 BUFx2_ASAP7_75t_R input941 (.A(io_ins_up_2[39]),
    .Y(net940));
 BUFx2_ASAP7_75t_R input940 (.A(io_ins_up_2[38]),
    .Y(net939));
 BUFx2_ASAP7_75t_R input939 (.A(io_ins_up_2[37]),
    .Y(net938));
 BUFx2_ASAP7_75t_R input938 (.A(io_ins_up_2[36]),
    .Y(net937));
 BUFx2_ASAP7_75t_R input937 (.A(io_ins_up_2[35]),
    .Y(net936));
 BUFx2_ASAP7_75t_R input936 (.A(io_ins_up_2[34]),
    .Y(net935));
 BUFx2_ASAP7_75t_R input935 (.A(io_ins_up_2[33]),
    .Y(net934));
 BUFx2_ASAP7_75t_R input934 (.A(io_ins_up_2[32]),
    .Y(net933));
 BUFx2_ASAP7_75t_R input933 (.A(io_ins_up_2[31]),
    .Y(net932));
 BUFx2_ASAP7_75t_R input932 (.A(io_ins_up_2[30]),
    .Y(net931));
 BUFx2_ASAP7_75t_R input931 (.A(io_ins_up_2[2]),
    .Y(net930));
 BUFx2_ASAP7_75t_R input930 (.A(io_ins_up_2[29]),
    .Y(net929));
 BUFx2_ASAP7_75t_R input929 (.A(io_ins_up_2[28]),
    .Y(net928));
 BUFx2_ASAP7_75t_R input928 (.A(io_ins_up_2[27]),
    .Y(net927));
 BUFx2_ASAP7_75t_R input927 (.A(io_ins_up_2[26]),
    .Y(net926));
 BUFx2_ASAP7_75t_R input926 (.A(io_ins_up_2[25]),
    .Y(net925));
 BUFx2_ASAP7_75t_R input925 (.A(io_ins_up_2[24]),
    .Y(net924));
 BUFx2_ASAP7_75t_R input924 (.A(io_ins_up_2[23]),
    .Y(net923));
 BUFx2_ASAP7_75t_R input923 (.A(io_ins_up_2[22]),
    .Y(net922));
 BUFx2_ASAP7_75t_R input922 (.A(io_ins_up_2[21]),
    .Y(net921));
 BUFx2_ASAP7_75t_R input921 (.A(io_ins_up_2[20]),
    .Y(net920));
 BUFx2_ASAP7_75t_R input920 (.A(io_ins_up_2[1]),
    .Y(net919));
 BUFx2_ASAP7_75t_R input919 (.A(io_ins_up_2[19]),
    .Y(net918));
 BUFx2_ASAP7_75t_R input918 (.A(io_ins_up_2[18]),
    .Y(net917));
 BUFx2_ASAP7_75t_R input917 (.A(io_ins_up_2[17]),
    .Y(net916));
 BUFx2_ASAP7_75t_R input916 (.A(io_ins_up_2[16]),
    .Y(net915));
 BUFx2_ASAP7_75t_R input915 (.A(io_ins_up_2[15]),
    .Y(net914));
 BUFx2_ASAP7_75t_R input914 (.A(io_ins_up_2[14]),
    .Y(net913));
 BUFx2_ASAP7_75t_R input913 (.A(io_ins_up_2[13]),
    .Y(net912));
 BUFx2_ASAP7_75t_R input912 (.A(io_ins_up_2[12]),
    .Y(net911));
 BUFx2_ASAP7_75t_R input911 (.A(io_ins_up_2[11]),
    .Y(net910));
 BUFx2_ASAP7_75t_R input910 (.A(io_ins_up_2[10]),
    .Y(net909));
 BUFx2_ASAP7_75t_R input909 (.A(io_ins_up_2[0]),
    .Y(net908));
 BUFx2_ASAP7_75t_R input908 (.A(io_ins_up_1[9]),
    .Y(net907));
 BUFx2_ASAP7_75t_R input907 (.A(io_ins_up_1[8]),
    .Y(net906));
 BUFx2_ASAP7_75t_R input906 (.A(io_ins_up_1[7]),
    .Y(net905));
 BUFx2_ASAP7_75t_R input905 (.A(io_ins_up_1[6]),
    .Y(net904));
 BUFx2_ASAP7_75t_R input904 (.A(io_ins_up_1[63]),
    .Y(net903));
 BUFx2_ASAP7_75t_R input903 (.A(io_ins_up_1[62]),
    .Y(net902));
 BUFx2_ASAP7_75t_R input902 (.A(io_ins_up_1[61]),
    .Y(net901));
 BUFx2_ASAP7_75t_R input901 (.A(io_ins_up_1[60]),
    .Y(net900));
 BUFx2_ASAP7_75t_R input900 (.A(io_ins_up_1[5]),
    .Y(net899));
 BUFx2_ASAP7_75t_R input899 (.A(io_ins_up_1[59]),
    .Y(net898));
 BUFx2_ASAP7_75t_R input898 (.A(io_ins_up_1[58]),
    .Y(net897));
 BUFx2_ASAP7_75t_R input897 (.A(io_ins_up_1[57]),
    .Y(net896));
 BUFx2_ASAP7_75t_R input896 (.A(io_ins_up_1[56]),
    .Y(net895));
 BUFx2_ASAP7_75t_R input895 (.A(io_ins_up_1[55]),
    .Y(net894));
 BUFx2_ASAP7_75t_R input894 (.A(io_ins_up_1[54]),
    .Y(net893));
 BUFx2_ASAP7_75t_R input893 (.A(io_ins_up_1[53]),
    .Y(net892));
 BUFx2_ASAP7_75t_R input892 (.A(io_ins_up_1[52]),
    .Y(net891));
 BUFx2_ASAP7_75t_R input891 (.A(io_ins_up_1[51]),
    .Y(net890));
 BUFx2_ASAP7_75t_R input890 (.A(io_ins_up_1[50]),
    .Y(net889));
 BUFx2_ASAP7_75t_R input889 (.A(io_ins_up_1[4]),
    .Y(net888));
 BUFx2_ASAP7_75t_R input888 (.A(io_ins_up_1[49]),
    .Y(net887));
 BUFx2_ASAP7_75t_R input887 (.A(io_ins_up_1[48]),
    .Y(net886));
 BUFx2_ASAP7_75t_R input886 (.A(io_ins_up_1[47]),
    .Y(net885));
 BUFx2_ASAP7_75t_R input885 (.A(io_ins_up_1[46]),
    .Y(net884));
 BUFx2_ASAP7_75t_R input884 (.A(io_ins_up_1[45]),
    .Y(net883));
 BUFx2_ASAP7_75t_R input883 (.A(io_ins_up_1[44]),
    .Y(net882));
 BUFx2_ASAP7_75t_R input882 (.A(io_ins_up_1[43]),
    .Y(net881));
 BUFx2_ASAP7_75t_R input881 (.A(io_ins_up_1[42]),
    .Y(net880));
 BUFx2_ASAP7_75t_R input880 (.A(io_ins_up_1[41]),
    .Y(net879));
 BUFx2_ASAP7_75t_R input879 (.A(io_ins_up_1[40]),
    .Y(net878));
 BUFx2_ASAP7_75t_R input878 (.A(io_ins_up_1[3]),
    .Y(net877));
 BUFx2_ASAP7_75t_R input877 (.A(io_ins_up_1[39]),
    .Y(net876));
 BUFx2_ASAP7_75t_R input876 (.A(io_ins_up_1[38]),
    .Y(net875));
 BUFx2_ASAP7_75t_R input875 (.A(io_ins_up_1[37]),
    .Y(net874));
 BUFx2_ASAP7_75t_R input874 (.A(io_ins_up_1[36]),
    .Y(net873));
 BUFx2_ASAP7_75t_R input873 (.A(io_ins_up_1[35]),
    .Y(net872));
 BUFx2_ASAP7_75t_R input872 (.A(io_ins_up_1[34]),
    .Y(net871));
 BUFx2_ASAP7_75t_R input871 (.A(io_ins_up_1[33]),
    .Y(net870));
 BUFx2_ASAP7_75t_R input870 (.A(io_ins_up_1[32]),
    .Y(net869));
 BUFx2_ASAP7_75t_R input869 (.A(io_ins_up_1[31]),
    .Y(net868));
 BUFx2_ASAP7_75t_R input868 (.A(io_ins_up_1[30]),
    .Y(net867));
 BUFx2_ASAP7_75t_R input867 (.A(io_ins_up_1[2]),
    .Y(net866));
 BUFx2_ASAP7_75t_R input866 (.A(io_ins_up_1[29]),
    .Y(net865));
 BUFx2_ASAP7_75t_R input865 (.A(io_ins_up_1[28]),
    .Y(net864));
 BUFx2_ASAP7_75t_R input864 (.A(io_ins_up_1[27]),
    .Y(net863));
 BUFx2_ASAP7_75t_R input863 (.A(io_ins_up_1[26]),
    .Y(net862));
 BUFx2_ASAP7_75t_R input862 (.A(io_ins_up_1[25]),
    .Y(net861));
 BUFx2_ASAP7_75t_R input861 (.A(io_ins_up_1[24]),
    .Y(net860));
 BUFx2_ASAP7_75t_R input860 (.A(io_ins_up_1[23]),
    .Y(net859));
 BUFx2_ASAP7_75t_R input859 (.A(io_ins_up_1[22]),
    .Y(net858));
 BUFx2_ASAP7_75t_R input858 (.A(io_ins_up_1[21]),
    .Y(net857));
 BUFx2_ASAP7_75t_R input857 (.A(io_ins_up_1[20]),
    .Y(net856));
 BUFx2_ASAP7_75t_R input856 (.A(io_ins_up_1[1]),
    .Y(net855));
 BUFx2_ASAP7_75t_R input855 (.A(io_ins_up_1[19]),
    .Y(net854));
 BUFx2_ASAP7_75t_R input854 (.A(io_ins_up_1[18]),
    .Y(net853));
 BUFx2_ASAP7_75t_R input853 (.A(io_ins_up_1[17]),
    .Y(net852));
 BUFx2_ASAP7_75t_R input852 (.A(io_ins_up_1[16]),
    .Y(net851));
 BUFx2_ASAP7_75t_R input851 (.A(io_ins_up_1[15]),
    .Y(net850));
 BUFx2_ASAP7_75t_R input850 (.A(io_ins_up_1[14]),
    .Y(net849));
 BUFx2_ASAP7_75t_R input849 (.A(io_ins_up_1[13]),
    .Y(net848));
 BUFx2_ASAP7_75t_R input848 (.A(io_ins_up_1[12]),
    .Y(net847));
 BUFx2_ASAP7_75t_R input847 (.A(io_ins_up_1[11]),
    .Y(net846));
 BUFx2_ASAP7_75t_R input846 (.A(io_ins_up_1[10]),
    .Y(net845));
 BUFx2_ASAP7_75t_R input845 (.A(io_ins_up_1[0]),
    .Y(net844));
 BUFx2_ASAP7_75t_R input844 (.A(io_ins_up_0[9]),
    .Y(net843));
 BUFx2_ASAP7_75t_R input843 (.A(io_ins_up_0[8]),
    .Y(net842));
 BUFx2_ASAP7_75t_R input842 (.A(io_ins_up_0[7]),
    .Y(net841));
 BUFx2_ASAP7_75t_R input841 (.A(io_ins_up_0[6]),
    .Y(net840));
 BUFx2_ASAP7_75t_R input840 (.A(io_ins_up_0[63]),
    .Y(net839));
 BUFx2_ASAP7_75t_R input839 (.A(io_ins_up_0[62]),
    .Y(net838));
 BUFx2_ASAP7_75t_R input838 (.A(io_ins_up_0[61]),
    .Y(net837));
 BUFx2_ASAP7_75t_R input837 (.A(io_ins_up_0[60]),
    .Y(net836));
 BUFx2_ASAP7_75t_R input836 (.A(io_ins_up_0[5]),
    .Y(net835));
 BUFx2_ASAP7_75t_R input835 (.A(io_ins_up_0[59]),
    .Y(net834));
 BUFx2_ASAP7_75t_R input834 (.A(io_ins_up_0[58]),
    .Y(net833));
 BUFx2_ASAP7_75t_R input833 (.A(io_ins_up_0[57]),
    .Y(net832));
 BUFx2_ASAP7_75t_R input832 (.A(io_ins_up_0[56]),
    .Y(net831));
 BUFx2_ASAP7_75t_R input831 (.A(io_ins_up_0[55]),
    .Y(net830));
 BUFx2_ASAP7_75t_R input830 (.A(io_ins_up_0[54]),
    .Y(net829));
 BUFx2_ASAP7_75t_R input829 (.A(io_ins_up_0[53]),
    .Y(net828));
 BUFx2_ASAP7_75t_R input828 (.A(io_ins_up_0[52]),
    .Y(net827));
 BUFx2_ASAP7_75t_R input827 (.A(io_ins_up_0[51]),
    .Y(net826));
 BUFx2_ASAP7_75t_R input826 (.A(io_ins_up_0[50]),
    .Y(net825));
 BUFx2_ASAP7_75t_R input825 (.A(io_ins_up_0[4]),
    .Y(net824));
 BUFx2_ASAP7_75t_R input824 (.A(io_ins_up_0[49]),
    .Y(net823));
 BUFx2_ASAP7_75t_R input823 (.A(io_ins_up_0[48]),
    .Y(net822));
 BUFx2_ASAP7_75t_R input822 (.A(io_ins_up_0[47]),
    .Y(net821));
 BUFx2_ASAP7_75t_R input821 (.A(io_ins_up_0[46]),
    .Y(net820));
 BUFx2_ASAP7_75t_R input820 (.A(io_ins_up_0[45]),
    .Y(net819));
 BUFx2_ASAP7_75t_R input819 (.A(io_ins_up_0[44]),
    .Y(net818));
 BUFx2_ASAP7_75t_R input818 (.A(io_ins_up_0[43]),
    .Y(net817));
 BUFx2_ASAP7_75t_R input817 (.A(io_ins_up_0[42]),
    .Y(net816));
 BUFx2_ASAP7_75t_R input816 (.A(io_ins_up_0[41]),
    .Y(net815));
 BUFx2_ASAP7_75t_R input815 (.A(io_ins_up_0[40]),
    .Y(net814));
 BUFx2_ASAP7_75t_R input814 (.A(io_ins_up_0[3]),
    .Y(net813));
 BUFx2_ASAP7_75t_R input813 (.A(io_ins_up_0[39]),
    .Y(net812));
 BUFx2_ASAP7_75t_R input812 (.A(io_ins_up_0[38]),
    .Y(net811));
 BUFx2_ASAP7_75t_R input811 (.A(io_ins_up_0[37]),
    .Y(net810));
 BUFx2_ASAP7_75t_R input810 (.A(io_ins_up_0[36]),
    .Y(net809));
 BUFx2_ASAP7_75t_R input809 (.A(io_ins_up_0[35]),
    .Y(net808));
 BUFx2_ASAP7_75t_R input808 (.A(io_ins_up_0[34]),
    .Y(net807));
 BUFx2_ASAP7_75t_R input807 (.A(io_ins_up_0[33]),
    .Y(net806));
 BUFx2_ASAP7_75t_R input806 (.A(io_ins_up_0[32]),
    .Y(net805));
 BUFx2_ASAP7_75t_R input805 (.A(io_ins_up_0[31]),
    .Y(net804));
 BUFx2_ASAP7_75t_R input804 (.A(io_ins_up_0[30]),
    .Y(net803));
 BUFx2_ASAP7_75t_R input803 (.A(io_ins_up_0[2]),
    .Y(net802));
 BUFx2_ASAP7_75t_R input802 (.A(io_ins_up_0[29]),
    .Y(net801));
 BUFx2_ASAP7_75t_R input801 (.A(io_ins_up_0[28]),
    .Y(net800));
 BUFx2_ASAP7_75t_R input800 (.A(io_ins_up_0[27]),
    .Y(net799));
 BUFx2_ASAP7_75t_R input799 (.A(io_ins_up_0[26]),
    .Y(net798));
 BUFx2_ASAP7_75t_R input798 (.A(io_ins_up_0[25]),
    .Y(net797));
 BUFx2_ASAP7_75t_R input797 (.A(io_ins_up_0[24]),
    .Y(net796));
 BUFx2_ASAP7_75t_R input796 (.A(io_ins_up_0[23]),
    .Y(net795));
 BUFx2_ASAP7_75t_R input795 (.A(io_ins_up_0[22]),
    .Y(net794));
 BUFx2_ASAP7_75t_R input794 (.A(io_ins_up_0[21]),
    .Y(net793));
 BUFx2_ASAP7_75t_R input793 (.A(io_ins_up_0[20]),
    .Y(net792));
 BUFx2_ASAP7_75t_R input792 (.A(io_ins_up_0[1]),
    .Y(net791));
 BUFx2_ASAP7_75t_R input791 (.A(io_ins_up_0[19]),
    .Y(net790));
 BUFx2_ASAP7_75t_R input790 (.A(io_ins_up_0[18]),
    .Y(net789));
 BUFx2_ASAP7_75t_R input789 (.A(io_ins_up_0[17]),
    .Y(net788));
 BUFx2_ASAP7_75t_R input788 (.A(io_ins_up_0[16]),
    .Y(net787));
 BUFx2_ASAP7_75t_R input787 (.A(io_ins_up_0[15]),
    .Y(net786));
 BUFx2_ASAP7_75t_R input786 (.A(io_ins_up_0[14]),
    .Y(net785));
 BUFx2_ASAP7_75t_R input785 (.A(io_ins_up_0[13]),
    .Y(net784));
 BUFx2_ASAP7_75t_R input784 (.A(io_ins_up_0[12]),
    .Y(net783));
 BUFx2_ASAP7_75t_R input783 (.A(io_ins_up_0[11]),
    .Y(net782));
 BUFx2_ASAP7_75t_R input782 (.A(io_ins_up_0[10]),
    .Y(net781));
 BUFx2_ASAP7_75t_R input781 (.A(io_ins_up_0[0]),
    .Y(net780));
 BUFx2_ASAP7_75t_R input780 (.A(io_ins_right_3[9]),
    .Y(net779));
 BUFx2_ASAP7_75t_R input779 (.A(io_ins_right_3[8]),
    .Y(net778));
 BUFx2_ASAP7_75t_R input778 (.A(io_ins_right_3[7]),
    .Y(net777));
 BUFx2_ASAP7_75t_R input777 (.A(io_ins_right_3[6]),
    .Y(net776));
 BUFx2_ASAP7_75t_R input776 (.A(io_ins_right_3[63]),
    .Y(net775));
 BUFx2_ASAP7_75t_R input775 (.A(io_ins_right_3[62]),
    .Y(net774));
 BUFx2_ASAP7_75t_R input774 (.A(io_ins_right_3[61]),
    .Y(net773));
 BUFx2_ASAP7_75t_R input773 (.A(io_ins_right_3[60]),
    .Y(net772));
 BUFx2_ASAP7_75t_R input772 (.A(io_ins_right_3[5]),
    .Y(net771));
 BUFx2_ASAP7_75t_R input771 (.A(io_ins_right_3[59]),
    .Y(net770));
 BUFx2_ASAP7_75t_R input770 (.A(io_ins_right_3[58]),
    .Y(net769));
 BUFx2_ASAP7_75t_R input769 (.A(io_ins_right_3[57]),
    .Y(net768));
 BUFx2_ASAP7_75t_R input768 (.A(io_ins_right_3[56]),
    .Y(net767));
 BUFx2_ASAP7_75t_R input767 (.A(io_ins_right_3[55]),
    .Y(net766));
 BUFx2_ASAP7_75t_R input766 (.A(io_ins_right_3[54]),
    .Y(net765));
 BUFx2_ASAP7_75t_R input765 (.A(io_ins_right_3[53]),
    .Y(net764));
 BUFx2_ASAP7_75t_R input764 (.A(io_ins_right_3[52]),
    .Y(net763));
 BUFx2_ASAP7_75t_R input763 (.A(io_ins_right_3[51]),
    .Y(net762));
 BUFx2_ASAP7_75t_R input762 (.A(io_ins_right_3[50]),
    .Y(net761));
 BUFx2_ASAP7_75t_R input761 (.A(io_ins_right_3[4]),
    .Y(net760));
 BUFx2_ASAP7_75t_R input760 (.A(io_ins_right_3[49]),
    .Y(net759));
 BUFx2_ASAP7_75t_R input759 (.A(io_ins_right_3[48]),
    .Y(net758));
 BUFx2_ASAP7_75t_R input758 (.A(io_ins_right_3[47]),
    .Y(net757));
 BUFx2_ASAP7_75t_R input757 (.A(io_ins_right_3[46]),
    .Y(net756));
 BUFx2_ASAP7_75t_R input756 (.A(io_ins_right_3[45]),
    .Y(net755));
 BUFx2_ASAP7_75t_R input755 (.A(io_ins_right_3[44]),
    .Y(net754));
 BUFx2_ASAP7_75t_R input754 (.A(io_ins_right_3[43]),
    .Y(net753));
 BUFx2_ASAP7_75t_R input753 (.A(io_ins_right_3[42]),
    .Y(net752));
 BUFx2_ASAP7_75t_R input752 (.A(io_ins_right_3[41]),
    .Y(net751));
 BUFx2_ASAP7_75t_R input751 (.A(io_ins_right_3[40]),
    .Y(net750));
 BUFx2_ASAP7_75t_R input750 (.A(io_ins_right_3[3]),
    .Y(net749));
 BUFx2_ASAP7_75t_R input749 (.A(io_ins_right_3[39]),
    .Y(net748));
 BUFx2_ASAP7_75t_R input748 (.A(io_ins_right_3[38]),
    .Y(net747));
 BUFx2_ASAP7_75t_R input747 (.A(io_ins_right_3[37]),
    .Y(net746));
 BUFx2_ASAP7_75t_R input746 (.A(io_ins_right_3[36]),
    .Y(net745));
 BUFx2_ASAP7_75t_R input745 (.A(io_ins_right_3[35]),
    .Y(net744));
 BUFx2_ASAP7_75t_R input744 (.A(io_ins_right_3[34]),
    .Y(net743));
 BUFx2_ASAP7_75t_R input743 (.A(io_ins_right_3[33]),
    .Y(net742));
 BUFx2_ASAP7_75t_R input742 (.A(io_ins_right_3[32]),
    .Y(net741));
 BUFx2_ASAP7_75t_R input741 (.A(io_ins_right_3[31]),
    .Y(net740));
 BUFx2_ASAP7_75t_R input740 (.A(io_ins_right_3[30]),
    .Y(net739));
 BUFx2_ASAP7_75t_R input739 (.A(io_ins_right_3[2]),
    .Y(net738));
 BUFx2_ASAP7_75t_R input738 (.A(io_ins_right_3[29]),
    .Y(net737));
 BUFx2_ASAP7_75t_R input737 (.A(io_ins_right_3[28]),
    .Y(net736));
 BUFx2_ASAP7_75t_R input736 (.A(io_ins_right_3[27]),
    .Y(net735));
 BUFx2_ASAP7_75t_R input735 (.A(io_ins_right_3[26]),
    .Y(net734));
 BUFx2_ASAP7_75t_R input734 (.A(io_ins_right_3[25]),
    .Y(net733));
 BUFx2_ASAP7_75t_R input733 (.A(io_ins_right_3[24]),
    .Y(net732));
 BUFx2_ASAP7_75t_R input732 (.A(io_ins_right_3[23]),
    .Y(net731));
 BUFx2_ASAP7_75t_R input731 (.A(io_ins_right_3[22]),
    .Y(net730));
 BUFx2_ASAP7_75t_R input730 (.A(io_ins_right_3[21]),
    .Y(net729));
 BUFx2_ASAP7_75t_R input729 (.A(io_ins_right_3[20]),
    .Y(net728));
 BUFx2_ASAP7_75t_R input728 (.A(io_ins_right_3[1]),
    .Y(net727));
 BUFx2_ASAP7_75t_R input727 (.A(io_ins_right_3[19]),
    .Y(net726));
 BUFx2_ASAP7_75t_R input726 (.A(io_ins_right_3[18]),
    .Y(net725));
 BUFx2_ASAP7_75t_R input725 (.A(io_ins_right_3[17]),
    .Y(net724));
 BUFx2_ASAP7_75t_R input724 (.A(io_ins_right_3[16]),
    .Y(net723));
 BUFx2_ASAP7_75t_R input723 (.A(io_ins_right_3[15]),
    .Y(net722));
 BUFx2_ASAP7_75t_R input722 (.A(io_ins_right_3[14]),
    .Y(net721));
 BUFx2_ASAP7_75t_R input721 (.A(io_ins_right_3[13]),
    .Y(net720));
 BUFx2_ASAP7_75t_R input720 (.A(io_ins_right_3[12]),
    .Y(net719));
 BUFx2_ASAP7_75t_R input719 (.A(io_ins_right_3[11]),
    .Y(net718));
 BUFx2_ASAP7_75t_R input718 (.A(io_ins_right_3[10]),
    .Y(net717));
 BUFx2_ASAP7_75t_R input717 (.A(io_ins_right_3[0]),
    .Y(net716));
 BUFx2_ASAP7_75t_R input716 (.A(io_ins_right_2[9]),
    .Y(net715));
 BUFx2_ASAP7_75t_R input715 (.A(io_ins_right_2[8]),
    .Y(net714));
 BUFx2_ASAP7_75t_R input714 (.A(io_ins_right_2[7]),
    .Y(net713));
 BUFx2_ASAP7_75t_R input713 (.A(io_ins_right_2[6]),
    .Y(net712));
 BUFx2_ASAP7_75t_R input712 (.A(io_ins_right_2[63]),
    .Y(net711));
 BUFx2_ASAP7_75t_R input711 (.A(io_ins_right_2[62]),
    .Y(net710));
 BUFx2_ASAP7_75t_R input710 (.A(io_ins_right_2[61]),
    .Y(net709));
 BUFx2_ASAP7_75t_R input709 (.A(io_ins_right_2[60]),
    .Y(net708));
 BUFx2_ASAP7_75t_R input708 (.A(io_ins_right_2[5]),
    .Y(net707));
 BUFx2_ASAP7_75t_R input707 (.A(io_ins_right_2[59]),
    .Y(net706));
 BUFx2_ASAP7_75t_R input706 (.A(io_ins_right_2[58]),
    .Y(net705));
 BUFx2_ASAP7_75t_R input705 (.A(io_ins_right_2[57]),
    .Y(net704));
 BUFx2_ASAP7_75t_R input704 (.A(io_ins_right_2[56]),
    .Y(net703));
 BUFx2_ASAP7_75t_R input703 (.A(io_ins_right_2[55]),
    .Y(net702));
 BUFx2_ASAP7_75t_R input702 (.A(io_ins_right_2[54]),
    .Y(net701));
 BUFx2_ASAP7_75t_R input701 (.A(io_ins_right_2[53]),
    .Y(net700));
 BUFx2_ASAP7_75t_R input700 (.A(io_ins_right_2[52]),
    .Y(net699));
 BUFx2_ASAP7_75t_R input699 (.A(io_ins_right_2[51]),
    .Y(net698));
 BUFx2_ASAP7_75t_R input698 (.A(io_ins_right_2[50]),
    .Y(net697));
 BUFx2_ASAP7_75t_R input697 (.A(io_ins_right_2[4]),
    .Y(net696));
 BUFx2_ASAP7_75t_R input696 (.A(io_ins_right_2[49]),
    .Y(net695));
 BUFx2_ASAP7_75t_R input695 (.A(io_ins_right_2[48]),
    .Y(net694));
 BUFx2_ASAP7_75t_R input694 (.A(io_ins_right_2[47]),
    .Y(net693));
 BUFx2_ASAP7_75t_R input693 (.A(io_ins_right_2[46]),
    .Y(net692));
 BUFx2_ASAP7_75t_R input692 (.A(io_ins_right_2[45]),
    .Y(net691));
 BUFx2_ASAP7_75t_R input691 (.A(io_ins_right_2[44]),
    .Y(net690));
 BUFx2_ASAP7_75t_R input690 (.A(io_ins_right_2[43]),
    .Y(net689));
 BUFx2_ASAP7_75t_R input689 (.A(io_ins_right_2[42]),
    .Y(net688));
 BUFx2_ASAP7_75t_R input688 (.A(io_ins_right_2[41]),
    .Y(net687));
 BUFx2_ASAP7_75t_R input687 (.A(io_ins_right_2[40]),
    .Y(net686));
 BUFx2_ASAP7_75t_R input686 (.A(io_ins_right_2[3]),
    .Y(net685));
 BUFx2_ASAP7_75t_R input685 (.A(io_ins_right_2[39]),
    .Y(net684));
 BUFx2_ASAP7_75t_R input684 (.A(io_ins_right_2[38]),
    .Y(net683));
 BUFx2_ASAP7_75t_R input683 (.A(io_ins_right_2[37]),
    .Y(net682));
 BUFx2_ASAP7_75t_R input682 (.A(io_ins_right_2[36]),
    .Y(net681));
 BUFx2_ASAP7_75t_R input681 (.A(io_ins_right_2[35]),
    .Y(net680));
 BUFx2_ASAP7_75t_R input680 (.A(io_ins_right_2[34]),
    .Y(net679));
 BUFx2_ASAP7_75t_R input679 (.A(io_ins_right_2[33]),
    .Y(net678));
 BUFx2_ASAP7_75t_R input678 (.A(io_ins_right_2[32]),
    .Y(net677));
 BUFx2_ASAP7_75t_R input677 (.A(io_ins_right_2[31]),
    .Y(net676));
 BUFx2_ASAP7_75t_R input676 (.A(io_ins_right_2[30]),
    .Y(net675));
 BUFx2_ASAP7_75t_R input675 (.A(io_ins_right_2[2]),
    .Y(net674));
 BUFx2_ASAP7_75t_R input674 (.A(io_ins_right_2[29]),
    .Y(net673));
 BUFx2_ASAP7_75t_R input673 (.A(io_ins_right_2[28]),
    .Y(net672));
 BUFx2_ASAP7_75t_R input672 (.A(io_ins_right_2[27]),
    .Y(net671));
 BUFx2_ASAP7_75t_R input671 (.A(io_ins_right_2[26]),
    .Y(net670));
 BUFx2_ASAP7_75t_R input670 (.A(io_ins_right_2[25]),
    .Y(net669));
 BUFx2_ASAP7_75t_R input669 (.A(io_ins_right_2[24]),
    .Y(net668));
 BUFx2_ASAP7_75t_R input668 (.A(io_ins_right_2[23]),
    .Y(net667));
 BUFx2_ASAP7_75t_R input667 (.A(io_ins_right_2[22]),
    .Y(net666));
 BUFx2_ASAP7_75t_R input666 (.A(io_ins_right_2[21]),
    .Y(net665));
 BUFx2_ASAP7_75t_R input665 (.A(io_ins_right_2[20]),
    .Y(net664));
 BUFx2_ASAP7_75t_R input664 (.A(io_ins_right_2[1]),
    .Y(net663));
 BUFx2_ASAP7_75t_R input663 (.A(io_ins_right_2[19]),
    .Y(net662));
 BUFx2_ASAP7_75t_R input662 (.A(io_ins_right_2[18]),
    .Y(net661));
 BUFx2_ASAP7_75t_R input661 (.A(io_ins_right_2[17]),
    .Y(net660));
 BUFx2_ASAP7_75t_R input660 (.A(io_ins_right_2[16]),
    .Y(net659));
 BUFx2_ASAP7_75t_R input659 (.A(io_ins_right_2[15]),
    .Y(net658));
 BUFx2_ASAP7_75t_R input658 (.A(io_ins_right_2[14]),
    .Y(net657));
 BUFx2_ASAP7_75t_R input657 (.A(io_ins_right_2[13]),
    .Y(net656));
 BUFx2_ASAP7_75t_R input656 (.A(io_ins_right_2[12]),
    .Y(net655));
 BUFx2_ASAP7_75t_R input655 (.A(io_ins_right_2[11]),
    .Y(net654));
 BUFx2_ASAP7_75t_R input654 (.A(io_ins_right_2[10]),
    .Y(net653));
 BUFx2_ASAP7_75t_R input653 (.A(io_ins_right_2[0]),
    .Y(net652));
 BUFx2_ASAP7_75t_R input652 (.A(io_ins_right_1[9]),
    .Y(net651));
 BUFx2_ASAP7_75t_R input651 (.A(io_ins_right_1[8]),
    .Y(net650));
 BUFx2_ASAP7_75t_R input650 (.A(io_ins_right_1[7]),
    .Y(net649));
 BUFx2_ASAP7_75t_R input649 (.A(io_ins_right_1[6]),
    .Y(net648));
 BUFx2_ASAP7_75t_R input648 (.A(io_ins_right_1[63]),
    .Y(net647));
 BUFx2_ASAP7_75t_R input647 (.A(io_ins_right_1[62]),
    .Y(net646));
 BUFx2_ASAP7_75t_R input646 (.A(io_ins_right_1[61]),
    .Y(net645));
 BUFx2_ASAP7_75t_R input645 (.A(io_ins_right_1[60]),
    .Y(net644));
 BUFx2_ASAP7_75t_R input644 (.A(io_ins_right_1[5]),
    .Y(net643));
 BUFx2_ASAP7_75t_R input643 (.A(io_ins_right_1[59]),
    .Y(net642));
 BUFx2_ASAP7_75t_R input642 (.A(io_ins_right_1[58]),
    .Y(net641));
 BUFx2_ASAP7_75t_R input641 (.A(io_ins_right_1[57]),
    .Y(net640));
 BUFx2_ASAP7_75t_R input640 (.A(io_ins_right_1[56]),
    .Y(net639));
 BUFx2_ASAP7_75t_R input639 (.A(io_ins_right_1[55]),
    .Y(net638));
 BUFx2_ASAP7_75t_R input638 (.A(io_ins_right_1[54]),
    .Y(net637));
 BUFx2_ASAP7_75t_R input637 (.A(io_ins_right_1[53]),
    .Y(net636));
 BUFx2_ASAP7_75t_R input636 (.A(io_ins_right_1[52]),
    .Y(net635));
 BUFx2_ASAP7_75t_R input635 (.A(io_ins_right_1[51]),
    .Y(net634));
 BUFx2_ASAP7_75t_R input634 (.A(io_ins_right_1[50]),
    .Y(net633));
 BUFx2_ASAP7_75t_R input633 (.A(io_ins_right_1[4]),
    .Y(net632));
 BUFx2_ASAP7_75t_R input632 (.A(io_ins_right_1[49]),
    .Y(net631));
 BUFx2_ASAP7_75t_R input631 (.A(io_ins_right_1[48]),
    .Y(net630));
 BUFx2_ASAP7_75t_R input630 (.A(io_ins_right_1[47]),
    .Y(net629));
 BUFx2_ASAP7_75t_R input629 (.A(io_ins_right_1[46]),
    .Y(net628));
 BUFx2_ASAP7_75t_R input628 (.A(io_ins_right_1[45]),
    .Y(net627));
 BUFx2_ASAP7_75t_R input627 (.A(io_ins_right_1[44]),
    .Y(net626));
 BUFx2_ASAP7_75t_R input626 (.A(io_ins_right_1[43]),
    .Y(net625));
 BUFx2_ASAP7_75t_R input625 (.A(io_ins_right_1[42]),
    .Y(net624));
 BUFx2_ASAP7_75t_R input624 (.A(io_ins_right_1[41]),
    .Y(net623));
 BUFx2_ASAP7_75t_R input623 (.A(io_ins_right_1[40]),
    .Y(net622));
 BUFx2_ASAP7_75t_R input622 (.A(io_ins_right_1[3]),
    .Y(net621));
 BUFx2_ASAP7_75t_R input621 (.A(io_ins_right_1[39]),
    .Y(net620));
 BUFx2_ASAP7_75t_R input620 (.A(io_ins_right_1[38]),
    .Y(net619));
 BUFx2_ASAP7_75t_R input619 (.A(io_ins_right_1[37]),
    .Y(net618));
 BUFx2_ASAP7_75t_R input618 (.A(io_ins_right_1[36]),
    .Y(net617));
 BUFx2_ASAP7_75t_R input617 (.A(io_ins_right_1[35]),
    .Y(net616));
 BUFx2_ASAP7_75t_R input616 (.A(io_ins_right_1[34]),
    .Y(net615));
 BUFx2_ASAP7_75t_R input615 (.A(io_ins_right_1[33]),
    .Y(net614));
 BUFx2_ASAP7_75t_R input614 (.A(io_ins_right_1[32]),
    .Y(net613));
 BUFx2_ASAP7_75t_R input613 (.A(io_ins_right_1[31]),
    .Y(net612));
 BUFx2_ASAP7_75t_R input612 (.A(io_ins_right_1[30]),
    .Y(net611));
 BUFx2_ASAP7_75t_R input611 (.A(io_ins_right_1[2]),
    .Y(net610));
 BUFx2_ASAP7_75t_R input610 (.A(io_ins_right_1[29]),
    .Y(net609));
 BUFx2_ASAP7_75t_R input609 (.A(io_ins_right_1[28]),
    .Y(net608));
 BUFx2_ASAP7_75t_R input608 (.A(io_ins_right_1[27]),
    .Y(net607));
 BUFx2_ASAP7_75t_R input607 (.A(io_ins_right_1[26]),
    .Y(net606));
 BUFx2_ASAP7_75t_R input606 (.A(io_ins_right_1[25]),
    .Y(net605));
 BUFx2_ASAP7_75t_R input605 (.A(io_ins_right_1[24]),
    .Y(net604));
 BUFx2_ASAP7_75t_R input604 (.A(io_ins_right_1[23]),
    .Y(net603));
 BUFx2_ASAP7_75t_R input603 (.A(io_ins_right_1[22]),
    .Y(net602));
 BUFx2_ASAP7_75t_R input602 (.A(io_ins_right_1[21]),
    .Y(net601));
 BUFx2_ASAP7_75t_R input601 (.A(io_ins_right_1[20]),
    .Y(net600));
 BUFx2_ASAP7_75t_R input600 (.A(io_ins_right_1[1]),
    .Y(net599));
 BUFx2_ASAP7_75t_R input599 (.A(io_ins_right_1[19]),
    .Y(net598));
 BUFx2_ASAP7_75t_R input598 (.A(io_ins_right_1[18]),
    .Y(net597));
 BUFx2_ASAP7_75t_R input597 (.A(io_ins_right_1[17]),
    .Y(net596));
 BUFx2_ASAP7_75t_R input596 (.A(io_ins_right_1[16]),
    .Y(net595));
 BUFx2_ASAP7_75t_R input595 (.A(io_ins_right_1[15]),
    .Y(net594));
 BUFx2_ASAP7_75t_R input594 (.A(io_ins_right_1[14]),
    .Y(net593));
 BUFx2_ASAP7_75t_R input593 (.A(io_ins_right_1[13]),
    .Y(net592));
 BUFx2_ASAP7_75t_R input592 (.A(io_ins_right_1[12]),
    .Y(net591));
 BUFx2_ASAP7_75t_R input591 (.A(io_ins_right_1[11]),
    .Y(net590));
 BUFx2_ASAP7_75t_R input590 (.A(io_ins_right_1[10]),
    .Y(net589));
 BUFx2_ASAP7_75t_R input589 (.A(io_ins_right_1[0]),
    .Y(net588));
 BUFx2_ASAP7_75t_R input588 (.A(io_ins_right_0[9]),
    .Y(net587));
 BUFx2_ASAP7_75t_R input587 (.A(io_ins_right_0[8]),
    .Y(net586));
 BUFx2_ASAP7_75t_R input586 (.A(io_ins_right_0[7]),
    .Y(net585));
 BUFx2_ASAP7_75t_R input585 (.A(io_ins_right_0[6]),
    .Y(net584));
 BUFx2_ASAP7_75t_R input584 (.A(io_ins_right_0[63]),
    .Y(net583));
 BUFx2_ASAP7_75t_R input583 (.A(io_ins_right_0[62]),
    .Y(net582));
 BUFx2_ASAP7_75t_R input582 (.A(io_ins_right_0[61]),
    .Y(net581));
 BUFx2_ASAP7_75t_R input581 (.A(io_ins_right_0[60]),
    .Y(net580));
 BUFx2_ASAP7_75t_R input580 (.A(io_ins_right_0[5]),
    .Y(net579));
 BUFx2_ASAP7_75t_R input579 (.A(io_ins_right_0[59]),
    .Y(net578));
 BUFx2_ASAP7_75t_R input578 (.A(io_ins_right_0[58]),
    .Y(net577));
 BUFx2_ASAP7_75t_R input577 (.A(io_ins_right_0[57]),
    .Y(net576));
 BUFx2_ASAP7_75t_R input576 (.A(io_ins_right_0[56]),
    .Y(net575));
 BUFx2_ASAP7_75t_R input575 (.A(io_ins_right_0[55]),
    .Y(net574));
 BUFx2_ASAP7_75t_R input574 (.A(io_ins_right_0[54]),
    .Y(net573));
 BUFx2_ASAP7_75t_R input573 (.A(io_ins_right_0[53]),
    .Y(net572));
 BUFx2_ASAP7_75t_R input572 (.A(io_ins_right_0[52]),
    .Y(net571));
 BUFx2_ASAP7_75t_R input571 (.A(io_ins_right_0[51]),
    .Y(net570));
 BUFx2_ASAP7_75t_R input570 (.A(io_ins_right_0[50]),
    .Y(net569));
 BUFx2_ASAP7_75t_R input569 (.A(io_ins_right_0[4]),
    .Y(net568));
 BUFx2_ASAP7_75t_R input568 (.A(io_ins_right_0[49]),
    .Y(net567));
 BUFx2_ASAP7_75t_R input567 (.A(io_ins_right_0[48]),
    .Y(net566));
 BUFx2_ASAP7_75t_R input566 (.A(io_ins_right_0[47]),
    .Y(net565));
 BUFx2_ASAP7_75t_R input565 (.A(io_ins_right_0[46]),
    .Y(net564));
 BUFx2_ASAP7_75t_R input564 (.A(io_ins_right_0[45]),
    .Y(net563));
 BUFx2_ASAP7_75t_R input563 (.A(io_ins_right_0[44]),
    .Y(net562));
 BUFx2_ASAP7_75t_R input562 (.A(io_ins_right_0[43]),
    .Y(net561));
 BUFx2_ASAP7_75t_R input561 (.A(io_ins_right_0[42]),
    .Y(net560));
 BUFx2_ASAP7_75t_R input560 (.A(io_ins_right_0[41]),
    .Y(net559));
 BUFx2_ASAP7_75t_R input559 (.A(io_ins_right_0[40]),
    .Y(net558));
 BUFx2_ASAP7_75t_R input558 (.A(io_ins_right_0[3]),
    .Y(net557));
 BUFx2_ASAP7_75t_R input557 (.A(io_ins_right_0[39]),
    .Y(net556));
 BUFx2_ASAP7_75t_R input556 (.A(io_ins_right_0[38]),
    .Y(net555));
 BUFx2_ASAP7_75t_R input555 (.A(io_ins_right_0[37]),
    .Y(net554));
 BUFx2_ASAP7_75t_R input554 (.A(io_ins_right_0[36]),
    .Y(net553));
 BUFx2_ASAP7_75t_R input553 (.A(io_ins_right_0[35]),
    .Y(net552));
 BUFx2_ASAP7_75t_R input552 (.A(io_ins_right_0[34]),
    .Y(net551));
 BUFx2_ASAP7_75t_R input551 (.A(io_ins_right_0[33]),
    .Y(net550));
 BUFx2_ASAP7_75t_R input550 (.A(io_ins_right_0[32]),
    .Y(net549));
 BUFx2_ASAP7_75t_R input549 (.A(io_ins_right_0[31]),
    .Y(net548));
 BUFx2_ASAP7_75t_R input548 (.A(io_ins_right_0[30]),
    .Y(net547));
 BUFx2_ASAP7_75t_R input547 (.A(io_ins_right_0[2]),
    .Y(net546));
 BUFx2_ASAP7_75t_R input546 (.A(io_ins_right_0[29]),
    .Y(net545));
 BUFx2_ASAP7_75t_R input545 (.A(io_ins_right_0[28]),
    .Y(net544));
 BUFx2_ASAP7_75t_R input544 (.A(io_ins_right_0[27]),
    .Y(net543));
 BUFx2_ASAP7_75t_R input543 (.A(io_ins_right_0[26]),
    .Y(net542));
 BUFx2_ASAP7_75t_R input542 (.A(io_ins_right_0[25]),
    .Y(net541));
 BUFx2_ASAP7_75t_R input541 (.A(io_ins_right_0[24]),
    .Y(net540));
 BUFx2_ASAP7_75t_R input540 (.A(io_ins_right_0[23]),
    .Y(net539));
 BUFx2_ASAP7_75t_R input539 (.A(io_ins_right_0[22]),
    .Y(net538));
 BUFx2_ASAP7_75t_R input538 (.A(io_ins_right_0[21]),
    .Y(net537));
 BUFx2_ASAP7_75t_R input537 (.A(io_ins_right_0[20]),
    .Y(net536));
 BUFx2_ASAP7_75t_R input536 (.A(io_ins_right_0[1]),
    .Y(net535));
 BUFx2_ASAP7_75t_R input535 (.A(io_ins_right_0[19]),
    .Y(net534));
 BUFx2_ASAP7_75t_R input534 (.A(io_ins_right_0[18]),
    .Y(net533));
 BUFx2_ASAP7_75t_R input533 (.A(io_ins_right_0[17]),
    .Y(net532));
 BUFx2_ASAP7_75t_R input532 (.A(io_ins_right_0[16]),
    .Y(net531));
 BUFx2_ASAP7_75t_R input531 (.A(io_ins_right_0[15]),
    .Y(net530));
 BUFx2_ASAP7_75t_R input530 (.A(io_ins_right_0[14]),
    .Y(net529));
 BUFx2_ASAP7_75t_R input529 (.A(io_ins_right_0[13]),
    .Y(net528));
 BUFx2_ASAP7_75t_R input528 (.A(io_ins_right_0[12]),
    .Y(net527));
 BUFx2_ASAP7_75t_R input527 (.A(io_ins_right_0[11]),
    .Y(net526));
 BUFx2_ASAP7_75t_R input526 (.A(io_ins_right_0[10]),
    .Y(net525));
 BUFx2_ASAP7_75t_R input525 (.A(io_ins_right_0[0]),
    .Y(net524));
 BUFx2_ASAP7_75t_R input524 (.A(io_ins_left_3[9]),
    .Y(net523));
 BUFx2_ASAP7_75t_R input523 (.A(io_ins_left_3[8]),
    .Y(net522));
 BUFx2_ASAP7_75t_R input522 (.A(io_ins_left_3[7]),
    .Y(net521));
 BUFx2_ASAP7_75t_R input521 (.A(io_ins_left_3[6]),
    .Y(net520));
 BUFx2_ASAP7_75t_R input520 (.A(io_ins_left_3[63]),
    .Y(net519));
 BUFx2_ASAP7_75t_R input519 (.A(io_ins_left_3[62]),
    .Y(net518));
 BUFx2_ASAP7_75t_R input518 (.A(io_ins_left_3[61]),
    .Y(net517));
 BUFx2_ASAP7_75t_R input517 (.A(io_ins_left_3[60]),
    .Y(net516));
 BUFx2_ASAP7_75t_R input516 (.A(io_ins_left_3[5]),
    .Y(net515));
 BUFx2_ASAP7_75t_R input515 (.A(io_ins_left_3[59]),
    .Y(net514));
 BUFx2_ASAP7_75t_R input514 (.A(io_ins_left_3[58]),
    .Y(net513));
 BUFx2_ASAP7_75t_R input513 (.A(io_ins_left_3[57]),
    .Y(net512));
 BUFx2_ASAP7_75t_R input512 (.A(io_ins_left_3[56]),
    .Y(net511));
 BUFx2_ASAP7_75t_R input511 (.A(io_ins_left_3[55]),
    .Y(net510));
 BUFx2_ASAP7_75t_R input510 (.A(io_ins_left_3[54]),
    .Y(net509));
 BUFx2_ASAP7_75t_R input509 (.A(io_ins_left_3[53]),
    .Y(net508));
 BUFx2_ASAP7_75t_R input508 (.A(io_ins_left_3[52]),
    .Y(net507));
 BUFx2_ASAP7_75t_R input507 (.A(io_ins_left_3[51]),
    .Y(net506));
 BUFx2_ASAP7_75t_R input506 (.A(io_ins_left_3[50]),
    .Y(net505));
 BUFx2_ASAP7_75t_R input505 (.A(io_ins_left_3[4]),
    .Y(net504));
 BUFx2_ASAP7_75t_R input504 (.A(io_ins_left_3[49]),
    .Y(net503));
 BUFx2_ASAP7_75t_R input503 (.A(io_ins_left_3[48]),
    .Y(net502));
 BUFx2_ASAP7_75t_R input502 (.A(io_ins_left_3[47]),
    .Y(net501));
 BUFx2_ASAP7_75t_R input501 (.A(io_ins_left_3[46]),
    .Y(net500));
 BUFx2_ASAP7_75t_R input500 (.A(io_ins_left_3[45]),
    .Y(net499));
 BUFx2_ASAP7_75t_R input499 (.A(io_ins_left_3[44]),
    .Y(net498));
 BUFx2_ASAP7_75t_R input498 (.A(io_ins_left_3[43]),
    .Y(net497));
 BUFx2_ASAP7_75t_R input497 (.A(io_ins_left_3[42]),
    .Y(net496));
 BUFx2_ASAP7_75t_R input496 (.A(io_ins_left_3[41]),
    .Y(net495));
 BUFx2_ASAP7_75t_R input495 (.A(io_ins_left_3[40]),
    .Y(net494));
 BUFx2_ASAP7_75t_R input494 (.A(io_ins_left_3[3]),
    .Y(net493));
 BUFx2_ASAP7_75t_R input493 (.A(io_ins_left_3[39]),
    .Y(net492));
 BUFx2_ASAP7_75t_R input492 (.A(io_ins_left_3[38]),
    .Y(net491));
 BUFx2_ASAP7_75t_R input491 (.A(io_ins_left_3[37]),
    .Y(net490));
 BUFx2_ASAP7_75t_R input490 (.A(io_ins_left_3[36]),
    .Y(net489));
 BUFx2_ASAP7_75t_R input489 (.A(io_ins_left_3[35]),
    .Y(net488));
 BUFx2_ASAP7_75t_R input488 (.A(io_ins_left_3[34]),
    .Y(net487));
 BUFx2_ASAP7_75t_R input487 (.A(io_ins_left_3[33]),
    .Y(net486));
 BUFx2_ASAP7_75t_R input486 (.A(io_ins_left_3[32]),
    .Y(net485));
 BUFx2_ASAP7_75t_R input485 (.A(io_ins_left_3[31]),
    .Y(net484));
 BUFx2_ASAP7_75t_R input484 (.A(io_ins_left_3[30]),
    .Y(net483));
 BUFx2_ASAP7_75t_R input483 (.A(io_ins_left_3[2]),
    .Y(net482));
 BUFx2_ASAP7_75t_R input482 (.A(io_ins_left_3[29]),
    .Y(net481));
 BUFx2_ASAP7_75t_R input481 (.A(io_ins_left_3[28]),
    .Y(net480));
 BUFx2_ASAP7_75t_R input480 (.A(io_ins_left_3[27]),
    .Y(net479));
 BUFx2_ASAP7_75t_R input479 (.A(io_ins_left_3[26]),
    .Y(net478));
 BUFx2_ASAP7_75t_R input478 (.A(io_ins_left_3[25]),
    .Y(net477));
 BUFx2_ASAP7_75t_R input477 (.A(io_ins_left_3[24]),
    .Y(net476));
 BUFx2_ASAP7_75t_R input476 (.A(io_ins_left_3[23]),
    .Y(net475));
 BUFx2_ASAP7_75t_R input475 (.A(io_ins_left_3[22]),
    .Y(net474));
 BUFx2_ASAP7_75t_R input474 (.A(io_ins_left_3[21]),
    .Y(net473));
 BUFx2_ASAP7_75t_R input473 (.A(io_ins_left_3[20]),
    .Y(net472));
 BUFx2_ASAP7_75t_R input472 (.A(io_ins_left_3[1]),
    .Y(net471));
 BUFx2_ASAP7_75t_R input471 (.A(io_ins_left_3[19]),
    .Y(net470));
 BUFx2_ASAP7_75t_R input470 (.A(io_ins_left_3[18]),
    .Y(net469));
 BUFx2_ASAP7_75t_R input469 (.A(io_ins_left_3[17]),
    .Y(net468));
 BUFx2_ASAP7_75t_R input468 (.A(io_ins_left_3[16]),
    .Y(net467));
 BUFx2_ASAP7_75t_R input467 (.A(io_ins_left_3[15]),
    .Y(net466));
 BUFx2_ASAP7_75t_R input466 (.A(io_ins_left_3[14]),
    .Y(net465));
 BUFx2_ASAP7_75t_R input465 (.A(io_ins_left_3[13]),
    .Y(net464));
 BUFx2_ASAP7_75t_R input464 (.A(io_ins_left_3[12]),
    .Y(net463));
 BUFx2_ASAP7_75t_R input463 (.A(io_ins_left_3[11]),
    .Y(net462));
 BUFx2_ASAP7_75t_R input462 (.A(io_ins_left_3[10]),
    .Y(net461));
 BUFx2_ASAP7_75t_R input461 (.A(io_ins_left_3[0]),
    .Y(net460));
 BUFx2_ASAP7_75t_R input460 (.A(io_ins_left_2[9]),
    .Y(net459));
 BUFx2_ASAP7_75t_R input459 (.A(io_ins_left_2[8]),
    .Y(net458));
 BUFx2_ASAP7_75t_R input458 (.A(io_ins_left_2[7]),
    .Y(net457));
 BUFx2_ASAP7_75t_R input457 (.A(io_ins_left_2[6]),
    .Y(net456));
 BUFx2_ASAP7_75t_R input456 (.A(io_ins_left_2[63]),
    .Y(net455));
 BUFx2_ASAP7_75t_R input455 (.A(io_ins_left_2[62]),
    .Y(net454));
 BUFx2_ASAP7_75t_R input454 (.A(io_ins_left_2[61]),
    .Y(net453));
 BUFx2_ASAP7_75t_R input453 (.A(io_ins_left_2[60]),
    .Y(net452));
 BUFx2_ASAP7_75t_R input452 (.A(io_ins_left_2[5]),
    .Y(net451));
 BUFx2_ASAP7_75t_R input451 (.A(io_ins_left_2[59]),
    .Y(net450));
 BUFx2_ASAP7_75t_R input450 (.A(io_ins_left_2[58]),
    .Y(net449));
 BUFx2_ASAP7_75t_R input449 (.A(io_ins_left_2[57]),
    .Y(net448));
 BUFx2_ASAP7_75t_R input448 (.A(io_ins_left_2[56]),
    .Y(net447));
 BUFx2_ASAP7_75t_R input447 (.A(io_ins_left_2[55]),
    .Y(net446));
 BUFx2_ASAP7_75t_R input446 (.A(io_ins_left_2[54]),
    .Y(net445));
 BUFx2_ASAP7_75t_R input445 (.A(io_ins_left_2[53]),
    .Y(net444));
 BUFx2_ASAP7_75t_R input444 (.A(io_ins_left_2[52]),
    .Y(net443));
 BUFx2_ASAP7_75t_R input443 (.A(io_ins_left_2[51]),
    .Y(net442));
 BUFx2_ASAP7_75t_R input442 (.A(io_ins_left_2[50]),
    .Y(net441));
 BUFx2_ASAP7_75t_R input441 (.A(io_ins_left_2[4]),
    .Y(net440));
 BUFx2_ASAP7_75t_R input440 (.A(io_ins_left_2[49]),
    .Y(net439));
 BUFx2_ASAP7_75t_R input439 (.A(io_ins_left_2[48]),
    .Y(net438));
 BUFx2_ASAP7_75t_R input438 (.A(io_ins_left_2[47]),
    .Y(net437));
 BUFx2_ASAP7_75t_R input437 (.A(io_ins_left_2[46]),
    .Y(net436));
 BUFx2_ASAP7_75t_R input436 (.A(io_ins_left_2[45]),
    .Y(net435));
 BUFx2_ASAP7_75t_R input435 (.A(io_ins_left_2[44]),
    .Y(net434));
 BUFx2_ASAP7_75t_R input434 (.A(io_ins_left_2[43]),
    .Y(net433));
 BUFx2_ASAP7_75t_R input433 (.A(io_ins_left_2[42]),
    .Y(net432));
 BUFx2_ASAP7_75t_R input432 (.A(io_ins_left_2[41]),
    .Y(net431));
 BUFx2_ASAP7_75t_R input431 (.A(io_ins_left_2[40]),
    .Y(net430));
 BUFx2_ASAP7_75t_R input430 (.A(io_ins_left_2[3]),
    .Y(net429));
 BUFx2_ASAP7_75t_R input429 (.A(io_ins_left_2[39]),
    .Y(net428));
 BUFx2_ASAP7_75t_R input428 (.A(io_ins_left_2[38]),
    .Y(net427));
 BUFx2_ASAP7_75t_R input427 (.A(io_ins_left_2[37]),
    .Y(net426));
 BUFx2_ASAP7_75t_R input426 (.A(io_ins_left_2[36]),
    .Y(net425));
 BUFx2_ASAP7_75t_R input425 (.A(io_ins_left_2[35]),
    .Y(net424));
 BUFx2_ASAP7_75t_R input424 (.A(io_ins_left_2[34]),
    .Y(net423));
 BUFx2_ASAP7_75t_R input423 (.A(io_ins_left_2[33]),
    .Y(net422));
 BUFx2_ASAP7_75t_R input422 (.A(io_ins_left_2[32]),
    .Y(net421));
 BUFx2_ASAP7_75t_R input421 (.A(io_ins_left_2[31]),
    .Y(net420));
 BUFx2_ASAP7_75t_R input420 (.A(io_ins_left_2[30]),
    .Y(net419));
 BUFx2_ASAP7_75t_R input419 (.A(io_ins_left_2[2]),
    .Y(net418));
 BUFx2_ASAP7_75t_R input418 (.A(io_ins_left_2[29]),
    .Y(net417));
 BUFx2_ASAP7_75t_R input417 (.A(io_ins_left_2[28]),
    .Y(net416));
 BUFx2_ASAP7_75t_R input416 (.A(io_ins_left_2[27]),
    .Y(net415));
 BUFx2_ASAP7_75t_R input415 (.A(io_ins_left_2[26]),
    .Y(net414));
 BUFx2_ASAP7_75t_R input414 (.A(io_ins_left_2[25]),
    .Y(net413));
 BUFx2_ASAP7_75t_R input413 (.A(io_ins_left_2[24]),
    .Y(net412));
 BUFx2_ASAP7_75t_R input412 (.A(io_ins_left_2[23]),
    .Y(net411));
 BUFx2_ASAP7_75t_R input411 (.A(io_ins_left_2[22]),
    .Y(net410));
 BUFx2_ASAP7_75t_R input410 (.A(io_ins_left_2[21]),
    .Y(net409));
 BUFx2_ASAP7_75t_R input409 (.A(io_ins_left_2[20]),
    .Y(net408));
 BUFx2_ASAP7_75t_R input408 (.A(io_ins_left_2[1]),
    .Y(net407));
 BUFx2_ASAP7_75t_R input407 (.A(io_ins_left_2[19]),
    .Y(net406));
 BUFx2_ASAP7_75t_R input406 (.A(io_ins_left_2[18]),
    .Y(net405));
 BUFx2_ASAP7_75t_R input405 (.A(io_ins_left_2[17]),
    .Y(net404));
 BUFx2_ASAP7_75t_R input404 (.A(io_ins_left_2[16]),
    .Y(net403));
 BUFx2_ASAP7_75t_R input403 (.A(io_ins_left_2[15]),
    .Y(net402));
 BUFx2_ASAP7_75t_R input402 (.A(io_ins_left_2[14]),
    .Y(net401));
 BUFx2_ASAP7_75t_R input401 (.A(io_ins_left_2[13]),
    .Y(net400));
 BUFx2_ASAP7_75t_R input400 (.A(io_ins_left_2[12]),
    .Y(net399));
 BUFx2_ASAP7_75t_R input399 (.A(io_ins_left_2[11]),
    .Y(net398));
 BUFx2_ASAP7_75t_R input398 (.A(io_ins_left_2[10]),
    .Y(net397));
 BUFx2_ASAP7_75t_R input397 (.A(io_ins_left_2[0]),
    .Y(net396));
 BUFx2_ASAP7_75t_R input396 (.A(io_ins_left_1[9]),
    .Y(net395));
 BUFx2_ASAP7_75t_R input395 (.A(io_ins_left_1[8]),
    .Y(net394));
 BUFx2_ASAP7_75t_R input394 (.A(io_ins_left_1[7]),
    .Y(net393));
 BUFx2_ASAP7_75t_R input393 (.A(io_ins_left_1[6]),
    .Y(net392));
 BUFx2_ASAP7_75t_R input392 (.A(io_ins_left_1[63]),
    .Y(net391));
 BUFx2_ASAP7_75t_R input391 (.A(io_ins_left_1[62]),
    .Y(net390));
 BUFx2_ASAP7_75t_R input390 (.A(io_ins_left_1[61]),
    .Y(net389));
 BUFx2_ASAP7_75t_R input389 (.A(io_ins_left_1[60]),
    .Y(net388));
 BUFx2_ASAP7_75t_R input388 (.A(io_ins_left_1[5]),
    .Y(net387));
 BUFx2_ASAP7_75t_R input387 (.A(io_ins_left_1[59]),
    .Y(net386));
 BUFx2_ASAP7_75t_R input386 (.A(io_ins_left_1[58]),
    .Y(net385));
 BUFx2_ASAP7_75t_R input385 (.A(io_ins_left_1[57]),
    .Y(net384));
 BUFx2_ASAP7_75t_R input384 (.A(io_ins_left_1[56]),
    .Y(net383));
 BUFx2_ASAP7_75t_R input383 (.A(io_ins_left_1[55]),
    .Y(net382));
 BUFx2_ASAP7_75t_R input382 (.A(io_ins_left_1[54]),
    .Y(net381));
 BUFx2_ASAP7_75t_R input381 (.A(io_ins_left_1[53]),
    .Y(net380));
 BUFx2_ASAP7_75t_R input380 (.A(io_ins_left_1[52]),
    .Y(net379));
 BUFx2_ASAP7_75t_R input379 (.A(io_ins_left_1[51]),
    .Y(net378));
 BUFx2_ASAP7_75t_R input378 (.A(io_ins_left_1[50]),
    .Y(net377));
 BUFx2_ASAP7_75t_R input377 (.A(io_ins_left_1[4]),
    .Y(net376));
 BUFx2_ASAP7_75t_R input376 (.A(io_ins_left_1[49]),
    .Y(net375));
 BUFx2_ASAP7_75t_R input375 (.A(io_ins_left_1[48]),
    .Y(net374));
 BUFx2_ASAP7_75t_R input374 (.A(io_ins_left_1[47]),
    .Y(net373));
 BUFx2_ASAP7_75t_R input373 (.A(io_ins_left_1[46]),
    .Y(net372));
 BUFx2_ASAP7_75t_R input372 (.A(io_ins_left_1[45]),
    .Y(net371));
 BUFx2_ASAP7_75t_R input371 (.A(io_ins_left_1[44]),
    .Y(net370));
 BUFx2_ASAP7_75t_R input370 (.A(io_ins_left_1[43]),
    .Y(net369));
 BUFx2_ASAP7_75t_R input369 (.A(io_ins_left_1[42]),
    .Y(net368));
 BUFx2_ASAP7_75t_R input368 (.A(io_ins_left_1[41]),
    .Y(net367));
 BUFx2_ASAP7_75t_R input367 (.A(io_ins_left_1[40]),
    .Y(net366));
 BUFx2_ASAP7_75t_R input366 (.A(io_ins_left_1[3]),
    .Y(net365));
 BUFx2_ASAP7_75t_R input365 (.A(io_ins_left_1[39]),
    .Y(net364));
 BUFx2_ASAP7_75t_R input364 (.A(io_ins_left_1[38]),
    .Y(net363));
 BUFx2_ASAP7_75t_R input363 (.A(io_ins_left_1[37]),
    .Y(net362));
 BUFx2_ASAP7_75t_R input362 (.A(io_ins_left_1[36]),
    .Y(net361));
 BUFx2_ASAP7_75t_R input361 (.A(io_ins_left_1[35]),
    .Y(net360));
 BUFx2_ASAP7_75t_R input360 (.A(io_ins_left_1[34]),
    .Y(net359));
 BUFx2_ASAP7_75t_R input359 (.A(io_ins_left_1[33]),
    .Y(net358));
 BUFx2_ASAP7_75t_R input358 (.A(io_ins_left_1[32]),
    .Y(net357));
 BUFx2_ASAP7_75t_R input357 (.A(io_ins_left_1[31]),
    .Y(net356));
 BUFx2_ASAP7_75t_R input356 (.A(io_ins_left_1[30]),
    .Y(net355));
 BUFx2_ASAP7_75t_R input355 (.A(io_ins_left_1[2]),
    .Y(net354));
 BUFx2_ASAP7_75t_R input354 (.A(io_ins_left_1[29]),
    .Y(net353));
 BUFx2_ASAP7_75t_R input353 (.A(io_ins_left_1[28]),
    .Y(net352));
 BUFx2_ASAP7_75t_R input352 (.A(io_ins_left_1[27]),
    .Y(net351));
 BUFx2_ASAP7_75t_R input351 (.A(io_ins_left_1[26]),
    .Y(net350));
 BUFx2_ASAP7_75t_R input350 (.A(io_ins_left_1[25]),
    .Y(net349));
 BUFx2_ASAP7_75t_R input349 (.A(io_ins_left_1[24]),
    .Y(net348));
 BUFx2_ASAP7_75t_R input348 (.A(io_ins_left_1[23]),
    .Y(net347));
 BUFx2_ASAP7_75t_R input347 (.A(io_ins_left_1[22]),
    .Y(net346));
 BUFx2_ASAP7_75t_R input346 (.A(io_ins_left_1[21]),
    .Y(net345));
 BUFx2_ASAP7_75t_R input345 (.A(io_ins_left_1[20]),
    .Y(net344));
 BUFx2_ASAP7_75t_R input344 (.A(io_ins_left_1[1]),
    .Y(net343));
 BUFx2_ASAP7_75t_R input343 (.A(io_ins_left_1[19]),
    .Y(net342));
 BUFx2_ASAP7_75t_R input342 (.A(io_ins_left_1[18]),
    .Y(net341));
 BUFx2_ASAP7_75t_R input341 (.A(io_ins_left_1[17]),
    .Y(net340));
 BUFx2_ASAP7_75t_R input340 (.A(io_ins_left_1[16]),
    .Y(net339));
 BUFx2_ASAP7_75t_R input339 (.A(io_ins_left_1[15]),
    .Y(net338));
 BUFx2_ASAP7_75t_R input338 (.A(io_ins_left_1[14]),
    .Y(net337));
 BUFx2_ASAP7_75t_R input337 (.A(io_ins_left_1[13]),
    .Y(net336));
 BUFx2_ASAP7_75t_R input336 (.A(io_ins_left_1[12]),
    .Y(net335));
 BUFx2_ASAP7_75t_R input335 (.A(io_ins_left_1[11]),
    .Y(net334));
 BUFx2_ASAP7_75t_R input334 (.A(io_ins_left_1[10]),
    .Y(net333));
 BUFx2_ASAP7_75t_R input333 (.A(io_ins_left_1[0]),
    .Y(net332));
 BUFx2_ASAP7_75t_R input332 (.A(io_ins_left_0[9]),
    .Y(net331));
 BUFx2_ASAP7_75t_R input331 (.A(io_ins_left_0[8]),
    .Y(net330));
 BUFx2_ASAP7_75t_R input330 (.A(io_ins_left_0[7]),
    .Y(net329));
 BUFx2_ASAP7_75t_R input329 (.A(io_ins_left_0[6]),
    .Y(net328));
 BUFx2_ASAP7_75t_R input328 (.A(io_ins_left_0[63]),
    .Y(net327));
 BUFx2_ASAP7_75t_R input327 (.A(io_ins_left_0[62]),
    .Y(net326));
 BUFx2_ASAP7_75t_R input326 (.A(io_ins_left_0[61]),
    .Y(net325));
 BUFx2_ASAP7_75t_R input325 (.A(io_ins_left_0[60]),
    .Y(net324));
 BUFx2_ASAP7_75t_R input324 (.A(io_ins_left_0[5]),
    .Y(net323));
 BUFx2_ASAP7_75t_R input323 (.A(io_ins_left_0[59]),
    .Y(net322));
 BUFx2_ASAP7_75t_R input322 (.A(io_ins_left_0[58]),
    .Y(net321));
 BUFx2_ASAP7_75t_R input321 (.A(io_ins_left_0[57]),
    .Y(net320));
 BUFx2_ASAP7_75t_R input320 (.A(io_ins_left_0[56]),
    .Y(net319));
 BUFx2_ASAP7_75t_R input319 (.A(io_ins_left_0[55]),
    .Y(net318));
 BUFx2_ASAP7_75t_R input318 (.A(io_ins_left_0[54]),
    .Y(net317));
 BUFx2_ASAP7_75t_R input317 (.A(io_ins_left_0[53]),
    .Y(net316));
 BUFx2_ASAP7_75t_R input316 (.A(io_ins_left_0[52]),
    .Y(net315));
 BUFx2_ASAP7_75t_R input315 (.A(io_ins_left_0[51]),
    .Y(net314));
 BUFx2_ASAP7_75t_R input314 (.A(io_ins_left_0[50]),
    .Y(net313));
 BUFx2_ASAP7_75t_R input313 (.A(io_ins_left_0[4]),
    .Y(net312));
 BUFx2_ASAP7_75t_R input312 (.A(io_ins_left_0[49]),
    .Y(net311));
 BUFx2_ASAP7_75t_R input311 (.A(io_ins_left_0[48]),
    .Y(net310));
 BUFx2_ASAP7_75t_R input310 (.A(io_ins_left_0[47]),
    .Y(net309));
 BUFx2_ASAP7_75t_R input309 (.A(io_ins_left_0[46]),
    .Y(net308));
 BUFx2_ASAP7_75t_R input308 (.A(io_ins_left_0[45]),
    .Y(net307));
 BUFx2_ASAP7_75t_R input307 (.A(io_ins_left_0[44]),
    .Y(net306));
 BUFx2_ASAP7_75t_R input306 (.A(io_ins_left_0[43]),
    .Y(net305));
 BUFx2_ASAP7_75t_R input305 (.A(io_ins_left_0[42]),
    .Y(net304));
 BUFx2_ASAP7_75t_R input304 (.A(io_ins_left_0[41]),
    .Y(net303));
 BUFx2_ASAP7_75t_R input303 (.A(io_ins_left_0[40]),
    .Y(net302));
 BUFx2_ASAP7_75t_R input302 (.A(io_ins_left_0[3]),
    .Y(net301));
 BUFx2_ASAP7_75t_R input301 (.A(io_ins_left_0[39]),
    .Y(net300));
 BUFx2_ASAP7_75t_R input300 (.A(io_ins_left_0[38]),
    .Y(net299));
 BUFx2_ASAP7_75t_R input299 (.A(io_ins_left_0[37]),
    .Y(net298));
 BUFx2_ASAP7_75t_R input298 (.A(io_ins_left_0[36]),
    .Y(net297));
 BUFx2_ASAP7_75t_R input297 (.A(io_ins_left_0[35]),
    .Y(net296));
 BUFx2_ASAP7_75t_R input296 (.A(io_ins_left_0[34]),
    .Y(net295));
 BUFx2_ASAP7_75t_R input295 (.A(io_ins_left_0[33]),
    .Y(net294));
 BUFx2_ASAP7_75t_R input294 (.A(io_ins_left_0[32]),
    .Y(net293));
 BUFx2_ASAP7_75t_R input293 (.A(io_ins_left_0[31]),
    .Y(net292));
 BUFx2_ASAP7_75t_R input292 (.A(io_ins_left_0[30]),
    .Y(net291));
 BUFx2_ASAP7_75t_R input291 (.A(io_ins_left_0[2]),
    .Y(net290));
 BUFx2_ASAP7_75t_R input290 (.A(io_ins_left_0[29]),
    .Y(net289));
 BUFx2_ASAP7_75t_R input289 (.A(io_ins_left_0[28]),
    .Y(net288));
 BUFx2_ASAP7_75t_R input288 (.A(io_ins_left_0[27]),
    .Y(net287));
 BUFx2_ASAP7_75t_R input287 (.A(io_ins_left_0[26]),
    .Y(net286));
 BUFx2_ASAP7_75t_R input286 (.A(io_ins_left_0[25]),
    .Y(net285));
 BUFx2_ASAP7_75t_R input285 (.A(io_ins_left_0[24]),
    .Y(net284));
 BUFx2_ASAP7_75t_R input284 (.A(io_ins_left_0[23]),
    .Y(net283));
 BUFx2_ASAP7_75t_R input283 (.A(io_ins_left_0[22]),
    .Y(net282));
 BUFx2_ASAP7_75t_R input282 (.A(io_ins_left_0[21]),
    .Y(net281));
 BUFx2_ASAP7_75t_R input281 (.A(io_ins_left_0[20]),
    .Y(net280));
 BUFx2_ASAP7_75t_R input280 (.A(io_ins_left_0[1]),
    .Y(net279));
 BUFx2_ASAP7_75t_R input279 (.A(io_ins_left_0[19]),
    .Y(net278));
 BUFx2_ASAP7_75t_R input278 (.A(io_ins_left_0[18]),
    .Y(net277));
 BUFx2_ASAP7_75t_R input277 (.A(io_ins_left_0[17]),
    .Y(net276));
 BUFx2_ASAP7_75t_R input276 (.A(io_ins_left_0[16]),
    .Y(net275));
 BUFx2_ASAP7_75t_R input275 (.A(io_ins_left_0[15]),
    .Y(net274));
 BUFx2_ASAP7_75t_R input274 (.A(io_ins_left_0[14]),
    .Y(net273));
 BUFx2_ASAP7_75t_R input273 (.A(io_ins_left_0[13]),
    .Y(net272));
 BUFx2_ASAP7_75t_R input272 (.A(io_ins_left_0[12]),
    .Y(net271));
 BUFx2_ASAP7_75t_R input271 (.A(io_ins_left_0[11]),
    .Y(net270));
 BUFx2_ASAP7_75t_R input270 (.A(io_ins_left_0[10]),
    .Y(net269));
 BUFx2_ASAP7_75t_R input269 (.A(io_ins_left_0[0]),
    .Y(net268));
 BUFx2_ASAP7_75t_R input268 (.A(io_ins_down_3[9]),
    .Y(net267));
 BUFx2_ASAP7_75t_R input267 (.A(io_ins_down_3[8]),
    .Y(net266));
 BUFx2_ASAP7_75t_R input266 (.A(io_ins_down_3[7]),
    .Y(net265));
 BUFx2_ASAP7_75t_R input265 (.A(io_ins_down_3[6]),
    .Y(net264));
 BUFx2_ASAP7_75t_R input264 (.A(io_ins_down_3[63]),
    .Y(net263));
 BUFx2_ASAP7_75t_R input263 (.A(io_ins_down_3[62]),
    .Y(net262));
 BUFx2_ASAP7_75t_R input262 (.A(io_ins_down_3[61]),
    .Y(net261));
 BUFx2_ASAP7_75t_R input261 (.A(io_ins_down_3[60]),
    .Y(net260));
 BUFx2_ASAP7_75t_R input260 (.A(io_ins_down_3[5]),
    .Y(net259));
 BUFx2_ASAP7_75t_R input259 (.A(io_ins_down_3[59]),
    .Y(net258));
 BUFx2_ASAP7_75t_R input258 (.A(io_ins_down_3[58]),
    .Y(net257));
 BUFx2_ASAP7_75t_R input257 (.A(io_ins_down_3[57]),
    .Y(net256));
 BUFx2_ASAP7_75t_R input256 (.A(io_ins_down_3[56]),
    .Y(net255));
 BUFx2_ASAP7_75t_R input255 (.A(io_ins_down_3[55]),
    .Y(net254));
 BUFx2_ASAP7_75t_R input254 (.A(io_ins_down_3[54]),
    .Y(net253));
 BUFx2_ASAP7_75t_R input253 (.A(io_ins_down_3[53]),
    .Y(net252));
 BUFx2_ASAP7_75t_R input252 (.A(io_ins_down_3[52]),
    .Y(net251));
 BUFx2_ASAP7_75t_R input251 (.A(io_ins_down_3[51]),
    .Y(net250));
 BUFx2_ASAP7_75t_R input250 (.A(io_ins_down_3[50]),
    .Y(net249));
 BUFx2_ASAP7_75t_R input249 (.A(io_ins_down_3[4]),
    .Y(net248));
 BUFx2_ASAP7_75t_R input248 (.A(io_ins_down_3[49]),
    .Y(net247));
 BUFx2_ASAP7_75t_R input247 (.A(io_ins_down_3[48]),
    .Y(net246));
 BUFx2_ASAP7_75t_R input246 (.A(io_ins_down_3[47]),
    .Y(net245));
 BUFx2_ASAP7_75t_R input245 (.A(io_ins_down_3[46]),
    .Y(net244));
 BUFx2_ASAP7_75t_R input244 (.A(io_ins_down_3[45]),
    .Y(net243));
 BUFx2_ASAP7_75t_R input243 (.A(io_ins_down_3[44]),
    .Y(net242));
 BUFx2_ASAP7_75t_R input242 (.A(io_ins_down_3[43]),
    .Y(net241));
 BUFx2_ASAP7_75t_R input241 (.A(io_ins_down_3[42]),
    .Y(net240));
 BUFx2_ASAP7_75t_R input240 (.A(io_ins_down_3[41]),
    .Y(net239));
 BUFx2_ASAP7_75t_R input239 (.A(io_ins_down_3[40]),
    .Y(net238));
 BUFx2_ASAP7_75t_R input238 (.A(io_ins_down_3[3]),
    .Y(net237));
 BUFx2_ASAP7_75t_R input237 (.A(io_ins_down_3[39]),
    .Y(net236));
 BUFx2_ASAP7_75t_R input236 (.A(io_ins_down_3[38]),
    .Y(net235));
 BUFx2_ASAP7_75t_R input235 (.A(io_ins_down_3[37]),
    .Y(net234));
 BUFx2_ASAP7_75t_R input234 (.A(io_ins_down_3[36]),
    .Y(net233));
 BUFx2_ASAP7_75t_R input233 (.A(io_ins_down_3[35]),
    .Y(net232));
 BUFx2_ASAP7_75t_R input232 (.A(io_ins_down_3[34]),
    .Y(net231));
 BUFx2_ASAP7_75t_R input231 (.A(io_ins_down_3[33]),
    .Y(net230));
 BUFx2_ASAP7_75t_R input230 (.A(io_ins_down_3[32]),
    .Y(net229));
 BUFx2_ASAP7_75t_R input229 (.A(io_ins_down_3[31]),
    .Y(net228));
 BUFx2_ASAP7_75t_R input228 (.A(io_ins_down_3[30]),
    .Y(net227));
 BUFx2_ASAP7_75t_R input227 (.A(io_ins_down_3[2]),
    .Y(net226));
 BUFx2_ASAP7_75t_R input226 (.A(io_ins_down_3[29]),
    .Y(net225));
 BUFx2_ASAP7_75t_R input225 (.A(io_ins_down_3[28]),
    .Y(net224));
 BUFx2_ASAP7_75t_R input224 (.A(io_ins_down_3[27]),
    .Y(net223));
 BUFx2_ASAP7_75t_R input223 (.A(io_ins_down_3[26]),
    .Y(net222));
 BUFx2_ASAP7_75t_R input222 (.A(io_ins_down_3[25]),
    .Y(net221));
 BUFx2_ASAP7_75t_R input221 (.A(io_ins_down_3[24]),
    .Y(net220));
 BUFx2_ASAP7_75t_R input220 (.A(io_ins_down_3[23]),
    .Y(net219));
 BUFx2_ASAP7_75t_R input219 (.A(io_ins_down_3[22]),
    .Y(net218));
 BUFx2_ASAP7_75t_R input218 (.A(io_ins_down_3[21]),
    .Y(net217));
 BUFx2_ASAP7_75t_R input217 (.A(io_ins_down_3[20]),
    .Y(net216));
 BUFx2_ASAP7_75t_R input216 (.A(io_ins_down_3[1]),
    .Y(net215));
 BUFx2_ASAP7_75t_R input215 (.A(io_ins_down_3[19]),
    .Y(net214));
 BUFx2_ASAP7_75t_R input214 (.A(io_ins_down_3[18]),
    .Y(net213));
 BUFx2_ASAP7_75t_R input213 (.A(io_ins_down_3[17]),
    .Y(net212));
 BUFx2_ASAP7_75t_R input212 (.A(io_ins_down_3[16]),
    .Y(net211));
 BUFx2_ASAP7_75t_R input211 (.A(io_ins_down_3[15]),
    .Y(net210));
 BUFx2_ASAP7_75t_R input210 (.A(io_ins_down_3[14]),
    .Y(net209));
 BUFx2_ASAP7_75t_R input209 (.A(io_ins_down_3[13]),
    .Y(net208));
 BUFx2_ASAP7_75t_R input208 (.A(io_ins_down_3[12]),
    .Y(net207));
 BUFx2_ASAP7_75t_R input207 (.A(io_ins_down_3[11]),
    .Y(net206));
 BUFx2_ASAP7_75t_R input206 (.A(io_ins_down_3[10]),
    .Y(net205));
 BUFx2_ASAP7_75t_R input205 (.A(io_ins_down_3[0]),
    .Y(net204));
 BUFx2_ASAP7_75t_R input204 (.A(io_ins_down_2[9]),
    .Y(net203));
 BUFx2_ASAP7_75t_R input203 (.A(io_ins_down_2[8]),
    .Y(net202));
 BUFx2_ASAP7_75t_R input202 (.A(io_ins_down_2[7]),
    .Y(net201));
 BUFx2_ASAP7_75t_R input201 (.A(io_ins_down_2[6]),
    .Y(net200));
 BUFx2_ASAP7_75t_R input200 (.A(io_ins_down_2[63]),
    .Y(net199));
 BUFx2_ASAP7_75t_R input199 (.A(io_ins_down_2[62]),
    .Y(net198));
 BUFx2_ASAP7_75t_R input198 (.A(io_ins_down_2[61]),
    .Y(net197));
 BUFx2_ASAP7_75t_R input197 (.A(io_ins_down_2[60]),
    .Y(net196));
 BUFx2_ASAP7_75t_R input196 (.A(io_ins_down_2[5]),
    .Y(net195));
 BUFx2_ASAP7_75t_R input195 (.A(io_ins_down_2[59]),
    .Y(net194));
 BUFx2_ASAP7_75t_R input194 (.A(io_ins_down_2[58]),
    .Y(net193));
 BUFx2_ASAP7_75t_R input193 (.A(io_ins_down_2[57]),
    .Y(net192));
 BUFx2_ASAP7_75t_R input192 (.A(io_ins_down_2[56]),
    .Y(net191));
 BUFx2_ASAP7_75t_R input191 (.A(io_ins_down_2[55]),
    .Y(net190));
 BUFx2_ASAP7_75t_R input190 (.A(io_ins_down_2[54]),
    .Y(net189));
 BUFx2_ASAP7_75t_R input189 (.A(io_ins_down_2[53]),
    .Y(net188));
 BUFx2_ASAP7_75t_R input188 (.A(io_ins_down_2[52]),
    .Y(net187));
 BUFx2_ASAP7_75t_R input187 (.A(io_ins_down_2[51]),
    .Y(net186));
 BUFx2_ASAP7_75t_R input186 (.A(io_ins_down_2[50]),
    .Y(net185));
 BUFx2_ASAP7_75t_R input185 (.A(io_ins_down_2[4]),
    .Y(net184));
 BUFx2_ASAP7_75t_R input184 (.A(io_ins_down_2[49]),
    .Y(net183));
 BUFx2_ASAP7_75t_R input183 (.A(io_ins_down_2[48]),
    .Y(net182));
 BUFx2_ASAP7_75t_R input182 (.A(io_ins_down_2[47]),
    .Y(net181));
 BUFx2_ASAP7_75t_R input181 (.A(io_ins_down_2[46]),
    .Y(net180));
 BUFx2_ASAP7_75t_R input180 (.A(io_ins_down_2[45]),
    .Y(net179));
 BUFx2_ASAP7_75t_R input179 (.A(io_ins_down_2[44]),
    .Y(net178));
 BUFx2_ASAP7_75t_R input178 (.A(io_ins_down_2[43]),
    .Y(net177));
 BUFx2_ASAP7_75t_R input177 (.A(io_ins_down_2[42]),
    .Y(net176));
 BUFx2_ASAP7_75t_R input176 (.A(io_ins_down_2[41]),
    .Y(net175));
 BUFx2_ASAP7_75t_R input175 (.A(io_ins_down_2[40]),
    .Y(net174));
 BUFx2_ASAP7_75t_R input174 (.A(io_ins_down_2[3]),
    .Y(net173));
 BUFx2_ASAP7_75t_R input173 (.A(io_ins_down_2[39]),
    .Y(net172));
 BUFx2_ASAP7_75t_R input172 (.A(io_ins_down_2[38]),
    .Y(net171));
 BUFx2_ASAP7_75t_R input171 (.A(io_ins_down_2[37]),
    .Y(net170));
 BUFx2_ASAP7_75t_R input170 (.A(io_ins_down_2[36]),
    .Y(net169));
 BUFx2_ASAP7_75t_R input169 (.A(io_ins_down_2[35]),
    .Y(net168));
 BUFx2_ASAP7_75t_R input168 (.A(io_ins_down_2[34]),
    .Y(net167));
 BUFx2_ASAP7_75t_R input167 (.A(io_ins_down_2[33]),
    .Y(net166));
 BUFx2_ASAP7_75t_R input166 (.A(io_ins_down_2[32]),
    .Y(net165));
 BUFx2_ASAP7_75t_R input165 (.A(io_ins_down_2[31]),
    .Y(net164));
 BUFx2_ASAP7_75t_R input164 (.A(io_ins_down_2[30]),
    .Y(net163));
 BUFx2_ASAP7_75t_R input163 (.A(io_ins_down_2[2]),
    .Y(net162));
 BUFx2_ASAP7_75t_R input162 (.A(io_ins_down_2[29]),
    .Y(net161));
 BUFx2_ASAP7_75t_R input161 (.A(io_ins_down_2[28]),
    .Y(net160));
 BUFx2_ASAP7_75t_R input160 (.A(io_ins_down_2[27]),
    .Y(net159));
 BUFx2_ASAP7_75t_R input159 (.A(io_ins_down_2[26]),
    .Y(net158));
 BUFx2_ASAP7_75t_R input158 (.A(io_ins_down_2[25]),
    .Y(net157));
 BUFx2_ASAP7_75t_R input157 (.A(io_ins_down_2[24]),
    .Y(net156));
 BUFx2_ASAP7_75t_R input156 (.A(io_ins_down_2[23]),
    .Y(net155));
 BUFx2_ASAP7_75t_R input155 (.A(io_ins_down_2[22]),
    .Y(net154));
 BUFx2_ASAP7_75t_R input154 (.A(io_ins_down_2[21]),
    .Y(net153));
 BUFx2_ASAP7_75t_R input153 (.A(io_ins_down_2[20]),
    .Y(net152));
 BUFx2_ASAP7_75t_R input152 (.A(io_ins_down_2[1]),
    .Y(net151));
 BUFx2_ASAP7_75t_R input151 (.A(io_ins_down_2[19]),
    .Y(net150));
 BUFx2_ASAP7_75t_R input150 (.A(io_ins_down_2[18]),
    .Y(net149));
 BUFx2_ASAP7_75t_R input149 (.A(io_ins_down_2[17]),
    .Y(net148));
 BUFx2_ASAP7_75t_R input148 (.A(io_ins_down_2[16]),
    .Y(net147));
 BUFx2_ASAP7_75t_R input147 (.A(io_ins_down_2[15]),
    .Y(net146));
 BUFx2_ASAP7_75t_R input146 (.A(io_ins_down_2[14]),
    .Y(net145));
 BUFx2_ASAP7_75t_R input145 (.A(io_ins_down_2[13]),
    .Y(net144));
 BUFx2_ASAP7_75t_R input144 (.A(io_ins_down_2[12]),
    .Y(net143));
 BUFx2_ASAP7_75t_R input143 (.A(io_ins_down_2[11]),
    .Y(net142));
 BUFx2_ASAP7_75t_R input142 (.A(io_ins_down_2[10]),
    .Y(net141));
 BUFx2_ASAP7_75t_R input141 (.A(io_ins_down_2[0]),
    .Y(net140));
 BUFx2_ASAP7_75t_R input140 (.A(io_ins_down_1[9]),
    .Y(net139));
 BUFx2_ASAP7_75t_R input139 (.A(io_ins_down_1[8]),
    .Y(net138));
 BUFx2_ASAP7_75t_R input138 (.A(io_ins_down_1[7]),
    .Y(net137));
 BUFx2_ASAP7_75t_R input137 (.A(io_ins_down_1[6]),
    .Y(net136));
 BUFx2_ASAP7_75t_R input136 (.A(io_ins_down_1[63]),
    .Y(net135));
 BUFx2_ASAP7_75t_R input135 (.A(io_ins_down_1[62]),
    .Y(net134));
 BUFx2_ASAP7_75t_R input134 (.A(io_ins_down_1[61]),
    .Y(net133));
 BUFx2_ASAP7_75t_R input133 (.A(io_ins_down_1[60]),
    .Y(net132));
 BUFx2_ASAP7_75t_R input132 (.A(io_ins_down_1[5]),
    .Y(net131));
 BUFx2_ASAP7_75t_R input131 (.A(io_ins_down_1[59]),
    .Y(net130));
 BUFx2_ASAP7_75t_R input130 (.A(io_ins_down_1[58]),
    .Y(net129));
 BUFx2_ASAP7_75t_R input129 (.A(io_ins_down_1[57]),
    .Y(net128));
 BUFx2_ASAP7_75t_R input128 (.A(io_ins_down_1[56]),
    .Y(net127));
 BUFx2_ASAP7_75t_R input127 (.A(io_ins_down_1[55]),
    .Y(net126));
 BUFx2_ASAP7_75t_R input126 (.A(io_ins_down_1[54]),
    .Y(net125));
 BUFx2_ASAP7_75t_R input125 (.A(io_ins_down_1[53]),
    .Y(net124));
 BUFx2_ASAP7_75t_R input124 (.A(io_ins_down_1[52]),
    .Y(net123));
 BUFx2_ASAP7_75t_R input123 (.A(io_ins_down_1[51]),
    .Y(net122));
 BUFx2_ASAP7_75t_R input122 (.A(io_ins_down_1[50]),
    .Y(net121));
 BUFx2_ASAP7_75t_R input121 (.A(io_ins_down_1[4]),
    .Y(net120));
 BUFx2_ASAP7_75t_R input120 (.A(io_ins_down_1[49]),
    .Y(net119));
 BUFx2_ASAP7_75t_R input119 (.A(io_ins_down_1[48]),
    .Y(net118));
 BUFx2_ASAP7_75t_R input118 (.A(io_ins_down_1[47]),
    .Y(net117));
 BUFx2_ASAP7_75t_R input117 (.A(io_ins_down_1[46]),
    .Y(net116));
 BUFx2_ASAP7_75t_R input116 (.A(io_ins_down_1[45]),
    .Y(net115));
 BUFx2_ASAP7_75t_R input115 (.A(io_ins_down_1[44]),
    .Y(net114));
 BUFx2_ASAP7_75t_R input114 (.A(io_ins_down_1[43]),
    .Y(net113));
 BUFx2_ASAP7_75t_R input113 (.A(io_ins_down_1[42]),
    .Y(net112));
 BUFx2_ASAP7_75t_R input112 (.A(io_ins_down_1[41]),
    .Y(net111));
 BUFx2_ASAP7_75t_R input111 (.A(io_ins_down_1[40]),
    .Y(net110));
 BUFx2_ASAP7_75t_R input110 (.A(io_ins_down_1[3]),
    .Y(net109));
 BUFx2_ASAP7_75t_R input109 (.A(io_ins_down_1[39]),
    .Y(net108));
 BUFx2_ASAP7_75t_R input108 (.A(io_ins_down_1[38]),
    .Y(net107));
 BUFx2_ASAP7_75t_R input107 (.A(io_ins_down_1[37]),
    .Y(net106));
 BUFx2_ASAP7_75t_R input106 (.A(io_ins_down_1[36]),
    .Y(net105));
 BUFx2_ASAP7_75t_R input105 (.A(io_ins_down_1[35]),
    .Y(net104));
 BUFx2_ASAP7_75t_R input104 (.A(io_ins_down_1[34]),
    .Y(net103));
 BUFx2_ASAP7_75t_R input103 (.A(io_ins_down_1[33]),
    .Y(net102));
 BUFx2_ASAP7_75t_R input102 (.A(io_ins_down_1[32]),
    .Y(net101));
 BUFx2_ASAP7_75t_R input101 (.A(io_ins_down_1[31]),
    .Y(net100));
 BUFx2_ASAP7_75t_R input100 (.A(io_ins_down_1[30]),
    .Y(net99));
 BUFx2_ASAP7_75t_R input99 (.A(io_ins_down_1[2]),
    .Y(net98));
 BUFx2_ASAP7_75t_R input98 (.A(io_ins_down_1[29]),
    .Y(net97));
 BUFx2_ASAP7_75t_R input97 (.A(io_ins_down_1[28]),
    .Y(net96));
 BUFx2_ASAP7_75t_R input96 (.A(io_ins_down_1[27]),
    .Y(net95));
 BUFx2_ASAP7_75t_R input95 (.A(io_ins_down_1[26]),
    .Y(net94));
 BUFx2_ASAP7_75t_R input94 (.A(io_ins_down_1[25]),
    .Y(net93));
 BUFx2_ASAP7_75t_R input93 (.A(io_ins_down_1[24]),
    .Y(net92));
 BUFx2_ASAP7_75t_R input92 (.A(io_ins_down_1[23]),
    .Y(net91));
 BUFx2_ASAP7_75t_R input91 (.A(io_ins_down_1[22]),
    .Y(net90));
 BUFx2_ASAP7_75t_R input90 (.A(io_ins_down_1[21]),
    .Y(net89));
 BUFx2_ASAP7_75t_R input89 (.A(io_ins_down_1[20]),
    .Y(net88));
 BUFx2_ASAP7_75t_R input88 (.A(io_ins_down_1[1]),
    .Y(net87));
 BUFx2_ASAP7_75t_R input87 (.A(io_ins_down_1[19]),
    .Y(net86));
 BUFx2_ASAP7_75t_R input86 (.A(io_ins_down_1[18]),
    .Y(net85));
 BUFx2_ASAP7_75t_R input85 (.A(io_ins_down_1[17]),
    .Y(net84));
 BUFx2_ASAP7_75t_R input84 (.A(io_ins_down_1[16]),
    .Y(net83));
 BUFx2_ASAP7_75t_R input83 (.A(io_ins_down_1[15]),
    .Y(net82));
 BUFx2_ASAP7_75t_R input82 (.A(io_ins_down_1[14]),
    .Y(net81));
 BUFx2_ASAP7_75t_R input81 (.A(io_ins_down_1[13]),
    .Y(net80));
 BUFx2_ASAP7_75t_R input80 (.A(io_ins_down_1[12]),
    .Y(net79));
 BUFx2_ASAP7_75t_R input79 (.A(io_ins_down_1[11]),
    .Y(net78));
 BUFx2_ASAP7_75t_R input78 (.A(io_ins_down_1[10]),
    .Y(net77));
 BUFx2_ASAP7_75t_R input77 (.A(io_ins_down_1[0]),
    .Y(net76));
 BUFx2_ASAP7_75t_R input76 (.A(io_ins_down_0[9]),
    .Y(net75));
 BUFx2_ASAP7_75t_R input75 (.A(io_ins_down_0[8]),
    .Y(net74));
 BUFx2_ASAP7_75t_R input74 (.A(io_ins_down_0[7]),
    .Y(net73));
 BUFx2_ASAP7_75t_R input73 (.A(io_ins_down_0[6]),
    .Y(net72));
 BUFx2_ASAP7_75t_R input72 (.A(io_ins_down_0[63]),
    .Y(net71));
 BUFx2_ASAP7_75t_R input71 (.A(io_ins_down_0[62]),
    .Y(net70));
 BUFx2_ASAP7_75t_R input70 (.A(io_ins_down_0[61]),
    .Y(net69));
 BUFx2_ASAP7_75t_R input69 (.A(io_ins_down_0[60]),
    .Y(net68));
 BUFx2_ASAP7_75t_R input68 (.A(io_ins_down_0[5]),
    .Y(net67));
 BUFx2_ASAP7_75t_R input67 (.A(io_ins_down_0[59]),
    .Y(net66));
 BUFx2_ASAP7_75t_R input66 (.A(io_ins_down_0[58]),
    .Y(net65));
 BUFx2_ASAP7_75t_R input65 (.A(io_ins_down_0[57]),
    .Y(net64));
 BUFx2_ASAP7_75t_R input64 (.A(io_ins_down_0[56]),
    .Y(net63));
 BUFx2_ASAP7_75t_R input63 (.A(io_ins_down_0[55]),
    .Y(net62));
 BUFx2_ASAP7_75t_R input62 (.A(io_ins_down_0[54]),
    .Y(net61));
 BUFx2_ASAP7_75t_R input61 (.A(io_ins_down_0[53]),
    .Y(net60));
 BUFx2_ASAP7_75t_R input60 (.A(io_ins_down_0[52]),
    .Y(net59));
 BUFx2_ASAP7_75t_R input59 (.A(io_ins_down_0[51]),
    .Y(net58));
 BUFx2_ASAP7_75t_R input58 (.A(io_ins_down_0[50]),
    .Y(net57));
 BUFx2_ASAP7_75t_R input57 (.A(io_ins_down_0[4]),
    .Y(net56));
 BUFx2_ASAP7_75t_R input56 (.A(io_ins_down_0[49]),
    .Y(net55));
 BUFx2_ASAP7_75t_R input55 (.A(io_ins_down_0[48]),
    .Y(net54));
 BUFx2_ASAP7_75t_R input54 (.A(io_ins_down_0[47]),
    .Y(net53));
 BUFx2_ASAP7_75t_R input53 (.A(io_ins_down_0[46]),
    .Y(net52));
 BUFx2_ASAP7_75t_R input52 (.A(io_ins_down_0[45]),
    .Y(net51));
 BUFx2_ASAP7_75t_R input51 (.A(io_ins_down_0[44]),
    .Y(net50));
 BUFx2_ASAP7_75t_R input50 (.A(io_ins_down_0[43]),
    .Y(net49));
 BUFx2_ASAP7_75t_R input49 (.A(io_ins_down_0[42]),
    .Y(net48));
 BUFx2_ASAP7_75t_R input48 (.A(io_ins_down_0[41]),
    .Y(net47));
 BUFx2_ASAP7_75t_R input47 (.A(io_ins_down_0[40]),
    .Y(net46));
 BUFx2_ASAP7_75t_R input46 (.A(io_ins_down_0[3]),
    .Y(net45));
 BUFx2_ASAP7_75t_R input45 (.A(io_ins_down_0[39]),
    .Y(net44));
 BUFx2_ASAP7_75t_R input44 (.A(io_ins_down_0[38]),
    .Y(net43));
 BUFx2_ASAP7_75t_R input43 (.A(io_ins_down_0[37]),
    .Y(net42));
 BUFx2_ASAP7_75t_R input42 (.A(io_ins_down_0[36]),
    .Y(net41));
 BUFx2_ASAP7_75t_R input41 (.A(io_ins_down_0[35]),
    .Y(net40));
 BUFx2_ASAP7_75t_R input40 (.A(io_ins_down_0[34]),
    .Y(net39));
 BUFx2_ASAP7_75t_R input39 (.A(io_ins_down_0[33]),
    .Y(net38));
 BUFx2_ASAP7_75t_R input38 (.A(io_ins_down_0[32]),
    .Y(net37));
 BUFx2_ASAP7_75t_R input37 (.A(io_ins_down_0[31]),
    .Y(net36));
 BUFx2_ASAP7_75t_R input36 (.A(io_ins_down_0[30]),
    .Y(net35));
 BUFx2_ASAP7_75t_R input35 (.A(io_ins_down_0[2]),
    .Y(net34));
 BUFx2_ASAP7_75t_R input34 (.A(io_ins_down_0[29]),
    .Y(net33));
 BUFx2_ASAP7_75t_R input33 (.A(io_ins_down_0[28]),
    .Y(net32));
 BUFx2_ASAP7_75t_R input32 (.A(io_ins_down_0[27]),
    .Y(net31));
 BUFx2_ASAP7_75t_R input31 (.A(io_ins_down_0[26]),
    .Y(net30));
 BUFx2_ASAP7_75t_R input30 (.A(io_ins_down_0[25]),
    .Y(net29));
 BUFx2_ASAP7_75t_R input29 (.A(io_ins_down_0[24]),
    .Y(net28));
 BUFx2_ASAP7_75t_R input28 (.A(io_ins_down_0[23]),
    .Y(net27));
 BUFx2_ASAP7_75t_R input27 (.A(io_ins_down_0[22]),
    .Y(net26));
 BUFx2_ASAP7_75t_R input26 (.A(io_ins_down_0[21]),
    .Y(net25));
 BUFx2_ASAP7_75t_R input25 (.A(io_ins_down_0[20]),
    .Y(net24));
 BUFx2_ASAP7_75t_R input24 (.A(io_ins_down_0[1]),
    .Y(net23));
 BUFx2_ASAP7_75t_R input23 (.A(io_ins_down_0[19]),
    .Y(net22));
 BUFx2_ASAP7_75t_R input22 (.A(io_ins_down_0[18]),
    .Y(net21));
 BUFx2_ASAP7_75t_R input21 (.A(io_ins_down_0[17]),
    .Y(net20));
 BUFx2_ASAP7_75t_R input20 (.A(io_ins_down_0[16]),
    .Y(net19));
 BUFx2_ASAP7_75t_R input19 (.A(io_ins_down_0[15]),
    .Y(net18));
 BUFx2_ASAP7_75t_R input18 (.A(io_ins_down_0[14]),
    .Y(net17));
 BUFx2_ASAP7_75t_R input17 (.A(io_ins_down_0[13]),
    .Y(net16));
 BUFx2_ASAP7_75t_R input16 (.A(io_ins_down_0[12]),
    .Y(net15));
 BUFx2_ASAP7_75t_R input15 (.A(io_ins_down_0[11]),
    .Y(net14));
 BUFx2_ASAP7_75t_R input14 (.A(io_ins_down_0[10]),
    .Y(net13));
 BUFx2_ASAP7_75t_R input13 (.A(io_ins_down_0[0]),
    .Y(net12));
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_335_1326 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_335_1325 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_335_1324 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_334_1323 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_334_1322 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_333_1321 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_332_1320 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_332_1319 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_331_1318 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_330_1317 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_330_1316 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_329_1315 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_328_1314 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_328_1313 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_327_1312 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_326_1311 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_326_1310 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_325_1309 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_324_1308 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_324_1307 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_323_1306 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_322_1305 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_322_1304 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_322_1303 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_253_1302 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_253_1301 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_253_1300 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_252_1299 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_252_1298 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_251_1297 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_250_1296 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_250_1295 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_249_1294 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_248_1293 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_248_1292 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_247_1291 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_246_1290 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_246_1289 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_245_1288 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_244_1287 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_244_1286 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_243_1285 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_242_1284 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_242_1283 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_242_1282 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_173_1281 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_173_1280 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_173_1279 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_172_1278 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_172_1277 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_171_1276 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_170_1275 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_170_1274 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_169_1273 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_168_1272 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_168_1271 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_167_1270 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_166_1269 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_166_1268 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_165_1267 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_164_1266 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_164_1265 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_163_1264 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_162_1263 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_162_1262 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_162_1261 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_93_1260 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_93_1259 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_93_1258 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_92_1257 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_92_1256 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_91_1255 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_90_1254 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_90_1253 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_89_1252 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_88_1251 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_88_1250 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_87_1249 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_86_1248 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_86_1247 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_85_1246 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_84_1245 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_84_1244 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_83_1243 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_82_1242 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_82_1241 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_82_1240 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_13_1239 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_13_1238 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_13_1237 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_12_1236 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_12_1235 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_11_1234 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_10_1233 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_10_1232 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_9_1231 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_8_1230 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_8_1229 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_7_1228 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_6_1227 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_6_1226 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_5_1225 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_4_1224 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_4_1223 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_3_1222 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_2_1221 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_2_1220 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1_1219 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_0_1218 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_0_1217 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_0_1216 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_321_1_Right_1215 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_320_1_Right_1214 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_319_1_Right_1213 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_318_1_Right_1212 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_317_1_Right_1211 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_316_1_Right_1210 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_315_1_Right_1209 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_314_1_Right_1208 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_313_1_Right_1207 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_312_1_Right_1206 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_311_1_Right_1205 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_310_1_Right_1204 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_309_1_Right_1203 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_308_1_Right_1202 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_307_1_Right_1201 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_306_1_Right_1200 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_305_1_Right_1199 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_304_1_Right_1198 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_303_1_Right_1197 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_302_1_Right_1196 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_301_1_Right_1195 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_300_1_Right_1194 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_299_1_Right_1193 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_298_1_Right_1192 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_297_1_Right_1191 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_296_1_Right_1190 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_295_1_Right_1189 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_294_1_Right_1188 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_293_1_Right_1187 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_292_1_Right_1186 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_291_1_Right_1185 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_290_1_Right_1184 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_289_1_Right_1183 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_288_1_Right_1182 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_287_1_Right_1181 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_286_1_Right_1180 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_285_1_Right_1179 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_284_1_Right_1178 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_283_1_Right_1177 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_282_1_Right_1176 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_281_1_Right_1175 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_280_1_Right_1174 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_279_1_Right_1173 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_278_1_Right_1172 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_277_1_Right_1171 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_276_1_Right_1170 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_275_1_Right_1169 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_274_1_Right_1168 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_273_1_Right_1167 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_272_1_Right_1166 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_271_1_Right_1165 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_270_1_Right_1164 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_269_1_Right_1163 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_268_1_Right_1162 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_267_1_Right_1161 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_266_1_Right_1160 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_265_1_Right_1159 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_264_1_Right_1158 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_263_1_Right_1157 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_262_1_Right_1156 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_261_1_Right_1155 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_260_1_Right_1154 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_259_1_Right_1153 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_258_1_Right_1152 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_257_1_Right_1151 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_256_1_Right_1150 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_255_1_Right_1149 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_254_1_Right_1148 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_321_5_Left_1147 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_320_5_Left_1146 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_319_5_Left_1145 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_318_5_Left_1144 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_317_5_Left_1143 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_316_5_Left_1142 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_315_5_Left_1141 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_314_5_Left_1140 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_313_5_Left_1139 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_312_5_Left_1138 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_311_5_Left_1137 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_310_5_Left_1136 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_309_5_Left_1135 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_308_5_Left_1134 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_307_5_Left_1133 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_306_5_Left_1132 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_305_5_Left_1131 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_304_5_Left_1130 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_303_5_Left_1129 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_302_5_Left_1128 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_301_5_Left_1127 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_300_5_Left_1126 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_299_5_Left_1125 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_298_5_Left_1124 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_297_5_Left_1123 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_296_5_Left_1122 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_295_5_Left_1121 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_294_5_Left_1120 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_293_5_Left_1119 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_292_5_Left_1118 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_291_5_Left_1117 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_290_5_Left_1116 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_289_5_Left_1115 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_288_5_Left_1114 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_287_5_Left_1113 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_286_5_Left_1112 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_285_5_Left_1111 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_284_5_Left_1110 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_283_5_Left_1109 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_282_5_Left_1108 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_281_5_Left_1107 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_280_5_Left_1106 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_279_5_Left_1105 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_278_5_Left_1104 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_277_5_Left_1103 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_276_5_Left_1102 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_275_5_Left_1101 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_274_5_Left_1100 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_273_5_Left_1099 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_272_5_Left_1098 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_271_5_Left_1097 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_270_5_Left_1096 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_269_5_Left_1095 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_268_5_Left_1094 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_267_5_Left_1093 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_266_5_Left_1092 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_265_5_Left_1091 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_264_5_Left_1090 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_263_5_Left_1089 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_262_5_Left_1088 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_261_5_Left_1087 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_260_5_Left_1086 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_259_5_Left_1085 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_258_5_Left_1084 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_257_5_Left_1083 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_256_5_Left_1082 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_255_5_Left_1081 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_254_5_Left_1080 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_241_1_Right_1079 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_240_1_Right_1078 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_239_1_Right_1077 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_238_1_Right_1076 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_237_1_Right_1075 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_236_1_Right_1074 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_235_1_Right_1073 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_234_1_Right_1072 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_233_1_Right_1071 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_232_1_Right_1070 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_231_1_Right_1069 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_230_1_Right_1068 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_229_1_Right_1067 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_228_1_Right_1066 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_227_1_Right_1065 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_226_1_Right_1064 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_225_1_Right_1063 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_224_1_Right_1062 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_223_1_Right_1061 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_222_1_Right_1060 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_221_1_Right_1059 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_220_1_Right_1058 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_219_1_Right_1057 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_218_1_Right_1056 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_217_1_Right_1055 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_216_1_Right_1054 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_215_1_Right_1053 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_214_1_Right_1052 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_213_1_Right_1051 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_212_1_Right_1050 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_211_1_Right_1049 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_210_1_Right_1048 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_209_1_Right_1047 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_208_1_Right_1046 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_207_1_Right_1045 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_206_1_Right_1044 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_205_1_Right_1043 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_204_1_Right_1042 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_203_1_Right_1041 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_202_1_Right_1040 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_201_1_Right_1039 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_200_1_Right_1038 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_199_1_Right_1037 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_198_1_Right_1036 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_197_1_Right_1035 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_196_1_Right_1034 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_195_1_Right_1033 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_194_1_Right_1032 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_193_1_Right_1031 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_192_1_Right_1030 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_191_1_Right_1029 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_190_1_Right_1028 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_189_1_Right_1027 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_188_1_Right_1026 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_187_1_Right_1025 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_186_1_Right_1024 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_185_1_Right_1023 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_184_1_Right_1022 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_183_1_Right_1021 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_182_1_Right_1020 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_181_1_Right_1019 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_180_1_Right_1018 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_179_1_Right_1017 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_178_1_Right_1016 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_177_1_Right_1015 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_176_1_Right_1014 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_175_1_Right_1013 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_174_1_Right_1012 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_241_5_Left_1011 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_240_5_Left_1010 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_239_5_Left_1009 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_238_5_Left_1008 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_237_5_Left_1007 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_236_5_Left_1006 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_235_5_Left_1005 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_234_5_Left_1004 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_233_5_Left_1003 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_232_5_Left_1002 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_231_5_Left_1001 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_230_5_Left_1000 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_229_5_Left_999 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_228_5_Left_998 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_227_5_Left_997 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_226_5_Left_996 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_225_5_Left_995 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_224_5_Left_994 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_223_5_Left_993 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_222_5_Left_992 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_221_5_Left_991 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_220_5_Left_990 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_219_5_Left_989 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_218_5_Left_988 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_217_5_Left_987 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_216_5_Left_986 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_215_5_Left_985 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_214_5_Left_984 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_213_5_Left_983 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_212_5_Left_982 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_211_5_Left_981 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_210_5_Left_980 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_209_5_Left_979 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_208_5_Left_978 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_207_5_Left_977 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_206_5_Left_976 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_205_5_Left_975 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_204_5_Left_974 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_203_5_Left_973 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_202_5_Left_972 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_201_5_Left_971 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_200_5_Left_970 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_199_5_Left_969 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_198_5_Left_968 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_197_5_Left_967 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_196_5_Left_966 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_195_5_Left_965 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_194_5_Left_964 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_193_5_Left_963 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_192_5_Left_962 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_191_5_Left_961 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_190_5_Left_960 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_189_5_Left_959 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_188_5_Left_958 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_187_5_Left_957 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_186_5_Left_956 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_185_5_Left_955 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_184_5_Left_954 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_183_5_Left_953 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_182_5_Left_952 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_181_5_Left_951 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_180_5_Left_950 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_179_5_Left_949 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_178_5_Left_948 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_177_5_Left_947 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_176_5_Left_946 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_175_5_Left_945 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_174_5_Left_944 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_161_1_Right_943 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_160_1_Right_942 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_159_1_Right_941 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_158_1_Right_940 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_157_1_Right_939 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_156_1_Right_938 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_155_1_Right_937 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_154_1_Right_936 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_153_1_Right_935 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_152_1_Right_934 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_151_1_Right_933 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_150_1_Right_932 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_149_1_Right_931 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_148_1_Right_930 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_147_1_Right_929 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_146_1_Right_928 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_145_1_Right_927 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_144_1_Right_926 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_143_1_Right_925 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_142_1_Right_924 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_141_1_Right_923 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_140_1_Right_922 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_139_1_Right_921 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_138_1_Right_920 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_137_1_Right_919 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_136_1_Right_918 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_135_1_Right_917 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_134_1_Right_916 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_133_1_Right_915 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_132_1_Right_914 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_131_1_Right_913 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_130_1_Right_912 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_129_1_Right_911 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_128_1_Right_910 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_127_1_Right_909 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_126_1_Right_908 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_125_1_Right_907 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_124_1_Right_906 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_123_1_Right_905 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_122_1_Right_904 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_121_1_Right_903 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_120_1_Right_902 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_119_1_Right_901 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_118_1_Right_900 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_117_1_Right_899 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_116_1_Right_898 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_115_1_Right_897 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_114_1_Right_896 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_113_1_Right_895 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_112_1_Right_894 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_111_1_Right_893 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_110_1_Right_892 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_109_1_Right_891 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_108_1_Right_890 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_107_1_Right_889 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_106_1_Right_888 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_105_1_Right_887 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_104_1_Right_886 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_103_1_Right_885 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_102_1_Right_884 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_101_1_Right_883 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_100_1_Right_882 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_99_1_Right_881 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_98_1_Right_880 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_97_1_Right_879 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_96_1_Right_878 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_95_1_Right_877 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_94_1_Right_876 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_161_5_Left_875 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_160_5_Left_874 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_159_5_Left_873 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_158_5_Left_872 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_157_5_Left_871 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_156_5_Left_870 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_155_5_Left_869 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_154_5_Left_868 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_153_5_Left_867 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_152_5_Left_866 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_151_5_Left_865 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_150_5_Left_864 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_149_5_Left_863 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_148_5_Left_862 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_147_5_Left_861 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_146_5_Left_860 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_145_5_Left_859 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_144_5_Left_858 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_143_5_Left_857 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_142_5_Left_856 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_141_5_Left_855 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_140_5_Left_854 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_139_5_Left_853 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_138_5_Left_852 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_137_5_Left_851 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_136_5_Left_850 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_135_5_Left_849 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_134_5_Left_848 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_133_5_Left_847 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_132_5_Left_846 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_131_5_Left_845 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_130_5_Left_844 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_129_5_Left_843 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_128_5_Left_842 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_127_5_Left_841 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_126_5_Left_840 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_125_5_Left_839 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_124_5_Left_838 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_123_5_Left_837 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_122_5_Left_836 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_121_5_Left_835 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_120_5_Left_834 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_119_5_Left_833 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_118_5_Left_832 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_117_5_Left_831 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_116_5_Left_830 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_115_5_Left_829 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_114_5_Left_828 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_113_5_Left_827 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_112_5_Left_826 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_111_5_Left_825 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_110_5_Left_824 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_109_5_Left_823 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_108_5_Left_822 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_107_5_Left_821 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_106_5_Left_820 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_105_5_Left_819 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_104_5_Left_818 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_103_5_Left_817 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_102_5_Left_816 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_101_5_Left_815 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_100_5_Left_814 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_99_5_Left_813 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_98_5_Left_812 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_97_5_Left_811 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_96_5_Left_810 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_95_5_Left_809 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_94_5_Left_808 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_1_Right_807 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_81_1_Right_806 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_80_1_Right_805 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_79_1_Right_804 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_78_1_Right_803 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_77_1_Right_802 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_76_1_Right_801 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_75_1_Right_800 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_74_1_Right_799 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_73_1_Right_798 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_72_1_Right_797 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_71_1_Right_796 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_70_1_Right_795 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_69_1_Right_794 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_68_1_Right_793 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_67_1_Right_792 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_66_1_Right_791 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_65_1_Right_790 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_64_1_Right_789 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_63_1_Right_788 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_62_1_Right_787 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_61_1_Right_786 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_60_1_Right_785 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_59_1_Right_784 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_58_1_Right_783 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_57_1_Right_782 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_56_1_Right_781 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_55_1_Right_780 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_1_Right_779 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_1_Right_778 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_1_Right_777 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_1_Right_776 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_1_Right_775 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_1_Right_774 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_1_Right_773 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_1_Right_772 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_1_Right_771 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_1_Right_770 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_1_Right_769 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_1_Right_768 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_1_Right_767 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_1_Right_766 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_1_Right_765 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_1_Right_764 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_1_Right_763 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_1_Right_762 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_1_Right_761 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_1_Right_760 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_1_Right_759 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_1_Right_758 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_1_Right_757 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_1_Right_756 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_1_Right_755 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_1_Right_754 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_1_Right_753 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_1_Right_752 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_1_Right_751 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_1_Right_750 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_1_Right_749 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_1_Right_748 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_1_Right_747 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_1_Right_746 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_1_Right_745 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_1_Right_744 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_1_Right_743 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_1_Right_742 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_1_Right_741 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_1_Right_740 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_81_5_Left_739 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_80_5_Left_738 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_79_5_Left_737 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_78_5_Left_736 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_77_5_Left_735 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_76_5_Left_734 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_75_5_Left_733 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_74_5_Left_732 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_73_5_Left_731 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_72_5_Left_730 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_71_5_Left_729 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_70_5_Left_728 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_69_5_Left_727 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_68_5_Left_726 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_67_5_Left_725 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_66_5_Left_724 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_65_5_Left_723 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_64_5_Left_722 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_63_5_Left_721 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_62_5_Left_720 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_61_5_Left_719 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_60_5_Left_718 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_59_5_Left_717 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_58_5_Left_716 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_57_5_Left_715 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_56_5_Left_714 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_55_5_Left_713 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_5_Left_712 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_5_Left_711 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_5_Left_710 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_5_Left_709 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_5_Left_708 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_5_Left_707 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_5_Left_706 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_5_Left_705 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_5_Left_704 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_5_Left_703 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_5_Left_702 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_5_Left_701 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_5_Left_700 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_5_Left_699 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_5_Left_698 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_5_Left_697 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_5_Left_696 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_5_Left_695 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_5_Left_694 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_5_Left_693 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_5_Left_692 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_5_Left_691 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_5_Left_690 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_5_Left_689 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_5_Left_688 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_5_Left_687 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_5_Left_686 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_5_Left_685 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_5_Left_684 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_5_Left_683 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_5_Left_682 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_5_Left_681 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_5_Left_680 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_5_Left_679 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_5_Left_678 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_5_Left_677 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_5_Left_676 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_5_Left_675 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_5_Left_674 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_5_Left_673 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_5_Left_672 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_1_Left_671 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_335_Left_670 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_334_Left_669 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_333_Left_668 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_332_Left_667 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_331_Left_666 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_330_Left_665 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_329_Left_664 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_328_Left_663 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_327_Left_662 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_326_Left_661 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_325_Left_660 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_324_Left_659 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_323_Left_658 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_322_Left_657 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_321_1_Left_656 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_320_1_Left_655 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_319_1_Left_654 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_318_1_Left_653 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_317_1_Left_652 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_316_1_Left_651 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_315_1_Left_650 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_314_1_Left_649 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_313_1_Left_648 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_312_1_Left_647 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_311_1_Left_646 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_310_1_Left_645 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_309_1_Left_644 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_308_1_Left_643 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_307_1_Left_642 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_306_1_Left_641 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_305_1_Left_640 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_304_1_Left_639 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_303_1_Left_638 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_302_1_Left_637 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_301_1_Left_636 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_300_1_Left_635 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_299_1_Left_634 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_298_1_Left_633 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_297_1_Left_632 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_296_1_Left_631 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_295_1_Left_630 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_294_1_Left_629 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_293_1_Left_628 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_292_1_Left_627 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_291_1_Left_626 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_290_1_Left_625 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_289_1_Left_624 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_288_1_Left_623 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_287_1_Left_622 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_286_1_Left_621 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_285_1_Left_620 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_284_1_Left_619 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_283_1_Left_618 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_282_1_Left_617 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_281_1_Left_616 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_280_1_Left_615 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_279_1_Left_614 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_278_1_Left_613 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_277_1_Left_612 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_276_1_Left_611 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_275_1_Left_610 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_274_1_Left_609 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_273_1_Left_608 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_272_1_Left_607 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_271_1_Left_606 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_270_1_Left_605 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_269_1_Left_604 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_268_1_Left_603 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_267_1_Left_602 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_266_1_Left_601 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_265_1_Left_600 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_264_1_Left_599 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_263_1_Left_598 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_262_1_Left_597 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_261_1_Left_596 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_260_1_Left_595 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_259_1_Left_594 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_258_1_Left_593 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_257_1_Left_592 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_256_1_Left_591 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_255_1_Left_590 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_253_Left_589 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_252_Left_588 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_251_Left_587 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_250_Left_586 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_249_Left_585 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_248_Left_584 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_247_Left_583 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_246_Left_582 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_245_Left_581 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_244_Left_580 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_243_Left_579 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_242_Left_578 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_254_1_Left_577 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_241_1_Left_576 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_240_1_Left_575 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_239_1_Left_574 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_238_1_Left_573 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_237_1_Left_572 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_236_1_Left_571 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_235_1_Left_570 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_234_1_Left_569 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_233_1_Left_568 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_232_1_Left_567 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_231_1_Left_566 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_230_1_Left_565 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_229_1_Left_564 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_228_1_Left_563 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_227_1_Left_562 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_226_1_Left_561 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_225_1_Left_560 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_224_1_Left_559 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_223_1_Left_558 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_222_1_Left_557 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_221_1_Left_556 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_220_1_Left_555 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_219_1_Left_554 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_218_1_Left_553 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_217_1_Left_552 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_216_1_Left_551 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_215_1_Left_550 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_214_1_Left_549 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_213_1_Left_548 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_212_1_Left_547 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_211_1_Left_546 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_210_1_Left_545 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_209_1_Left_544 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_208_1_Left_543 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_207_1_Left_542 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_206_1_Left_541 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_205_1_Left_540 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_204_1_Left_539 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_203_1_Left_538 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_202_1_Left_537 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_201_1_Left_536 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_200_1_Left_535 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_199_1_Left_534 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_198_1_Left_533 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_197_1_Left_532 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_196_1_Left_531 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_195_1_Left_530 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_194_1_Left_529 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_193_1_Left_528 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_192_1_Left_527 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_191_1_Left_526 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_190_1_Left_525 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_189_1_Left_524 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_188_1_Left_523 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_187_1_Left_522 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_186_1_Left_521 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_185_1_Left_520 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_184_1_Left_519 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_183_1_Left_518 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_182_1_Left_517 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_181_1_Left_516 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_180_1_Left_515 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_179_1_Left_514 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_178_1_Left_513 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_177_1_Left_512 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_176_1_Left_511 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_175_1_Left_510 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_173_Left_509 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_172_Left_508 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_171_Left_507 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_170_Left_506 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_169_Left_505 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_168_Left_504 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_167_Left_503 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_166_Left_502 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_165_Left_501 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_164_Left_500 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_163_Left_499 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_162_Left_498 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_174_1_Left_497 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_161_1_Left_496 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_160_1_Left_495 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_159_1_Left_494 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_158_1_Left_493 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_157_1_Left_492 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_156_1_Left_491 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_155_1_Left_490 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_154_1_Left_489 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_153_1_Left_488 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_152_1_Left_487 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_151_1_Left_486 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_150_1_Left_485 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_149_1_Left_484 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_148_1_Left_483 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_147_1_Left_482 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_146_1_Left_481 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_145_1_Left_480 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_144_1_Left_479 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_143_1_Left_478 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_142_1_Left_477 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_141_1_Left_476 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_140_1_Left_475 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_139_1_Left_474 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_138_1_Left_473 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_137_1_Left_472 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_136_1_Left_471 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_135_1_Left_470 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_134_1_Left_469 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_133_1_Left_468 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_132_1_Left_467 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_131_1_Left_466 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_130_1_Left_465 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_129_1_Left_464 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_128_1_Left_463 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_127_1_Left_462 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_126_1_Left_461 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_125_1_Left_460 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_124_1_Left_459 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_123_1_Left_458 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_122_1_Left_457 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_121_1_Left_456 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_120_1_Left_455 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_119_1_Left_454 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_118_1_Left_453 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_117_1_Left_452 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_116_1_Left_451 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_115_1_Left_450 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_114_1_Left_449 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_113_1_Left_448 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_112_1_Left_447 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_111_1_Left_446 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_110_1_Left_445 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_109_1_Left_444 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_108_1_Left_443 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_107_1_Left_442 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_106_1_Left_441 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_105_1_Left_440 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_104_1_Left_439 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_103_1_Left_438 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_102_1_Left_437 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_101_1_Left_436 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_100_1_Left_435 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_99_1_Left_434 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_98_1_Left_433 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_97_1_Left_432 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_96_1_Left_431 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_95_1_Left_430 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_93_Left_429 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_92_Left_428 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_91_Left_427 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_90_Left_426 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_89_Left_425 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_88_Left_424 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_87_Left_423 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_86_Left_422 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_85_Left_421 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_84_Left_420 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_83_Left_419 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_82_Left_418 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_94_1_Left_417 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_81_1_Left_416 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_80_1_Left_415 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_79_1_Left_414 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_78_1_Left_413 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_77_1_Left_412 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_76_1_Left_411 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_75_1_Left_410 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_74_1_Left_409 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_73_1_Left_408 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_72_1_Left_407 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_71_1_Left_406 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_70_1_Left_405 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_69_1_Left_404 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_68_1_Left_403 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_67_1_Left_402 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_66_1_Left_401 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_65_1_Left_400 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_64_1_Left_399 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_63_1_Left_398 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_62_1_Left_397 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_61_1_Left_396 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_60_1_Left_395 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_59_1_Left_394 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_58_1_Left_393 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_57_1_Left_392 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_56_1_Left_391 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_55_1_Left_390 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_1_Left_389 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_1_Left_388 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_1_Left_387 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_1_Left_386 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_1_Left_385 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_1_Left_384 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_1_Left_383 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_1_Left_382 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_1_Left_381 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_1_Left_380 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_1_Left_379 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_1_Left_378 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_1_Left_377 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_1_Left_376 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_1_Left_375 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_1_Left_374 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_1_Left_373 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_1_Left_372 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_1_Left_371 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_1_Left_370 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_1_Left_369 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_1_Left_368 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_1_Left_367 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_1_Left_366 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_1_Left_365 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_1_Left_364 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_1_Left_363 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_1_Left_362 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_1_Left_361 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_1_Left_360 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_1_Left_359 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_1_Left_358 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_1_Left_357 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_1_Left_356 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_1_Left_355 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_1_Left_354 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_1_Left_353 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_1_Left_352 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_1_Left_351 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_1_Left_350 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Left_349 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Left_348 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Left_347 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Left_346 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Left_345 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Left_344 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Left_343 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Left_342 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Left_341 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Left_340 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Left_339 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Left_338 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Left_337 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Left_336 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_321_5_Right_335 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_320_5_Right_334 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_319_5_Right_333 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_318_5_Right_332 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_317_5_Right_331 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_316_5_Right_330 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_315_5_Right_329 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_314_5_Right_328 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_313_5_Right_327 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_312_5_Right_326 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_311_5_Right_325 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_310_5_Right_324 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_309_5_Right_323 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_308_5_Right_322 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_307_5_Right_321 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_306_5_Right_320 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_305_5_Right_319 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_304_5_Right_318 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_303_5_Right_317 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_302_5_Right_316 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_301_5_Right_315 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_300_5_Right_314 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_299_5_Right_313 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_298_5_Right_312 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_297_5_Right_311 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_296_5_Right_310 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_295_5_Right_309 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_294_5_Right_308 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_293_5_Right_307 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_292_5_Right_306 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_291_5_Right_305 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_290_5_Right_304 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_289_5_Right_303 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_288_5_Right_302 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_287_5_Right_301 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_286_5_Right_300 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_285_5_Right_299 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_284_5_Right_298 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_283_5_Right_297 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_282_5_Right_296 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_281_5_Right_295 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_280_5_Right_294 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_279_5_Right_293 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_278_5_Right_292 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_277_5_Right_291 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_276_5_Right_290 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_275_5_Right_289 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_274_5_Right_288 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_273_5_Right_287 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_272_5_Right_286 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_271_5_Right_285 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_270_5_Right_284 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_269_5_Right_283 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_268_5_Right_282 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_267_5_Right_281 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_266_5_Right_280 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_265_5_Right_279 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_264_5_Right_278 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_263_5_Right_277 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_262_5_Right_276 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_261_5_Right_275 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_260_5_Right_274 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_259_5_Right_273 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_258_5_Right_272 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_257_5_Right_271 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_256_5_Right_270 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_255_5_Right_269 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_254_5_Right_268 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_241_5_Right_267 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_240_5_Right_266 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_239_5_Right_265 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_238_5_Right_264 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_237_5_Right_263 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_236_5_Right_262 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_235_5_Right_261 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_234_5_Right_260 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_233_5_Right_259 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_232_5_Right_258 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_231_5_Right_257 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_230_5_Right_256 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_229_5_Right_255 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_228_5_Right_254 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_227_5_Right_253 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_226_5_Right_252 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_225_5_Right_251 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_224_5_Right_250 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_223_5_Right_249 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_222_5_Right_248 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_221_5_Right_247 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_220_5_Right_246 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_219_5_Right_245 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_218_5_Right_244 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_217_5_Right_243 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_216_5_Right_242 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_215_5_Right_241 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_214_5_Right_240 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_213_5_Right_239 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_212_5_Right_238 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_211_5_Right_237 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_210_5_Right_236 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_209_5_Right_235 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_208_5_Right_234 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_207_5_Right_233 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_206_5_Right_232 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_205_5_Right_231 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_204_5_Right_230 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_203_5_Right_229 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_202_5_Right_228 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_201_5_Right_227 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_200_5_Right_226 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_199_5_Right_225 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_198_5_Right_224 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_197_5_Right_223 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_196_5_Right_222 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_195_5_Right_221 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_194_5_Right_220 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_193_5_Right_219 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_192_5_Right_218 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_191_5_Right_217 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_190_5_Right_216 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_189_5_Right_215 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_188_5_Right_214 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_187_5_Right_213 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_186_5_Right_212 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_185_5_Right_211 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_184_5_Right_210 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_183_5_Right_209 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_182_5_Right_208 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_181_5_Right_207 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_180_5_Right_206 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_179_5_Right_205 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_178_5_Right_204 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_177_5_Right_203 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_176_5_Right_202 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_175_5_Right_201 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_174_5_Right_200 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_161_5_Right_199 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_160_5_Right_198 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_159_5_Right_197 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_158_5_Right_196 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_157_5_Right_195 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_156_5_Right_194 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_155_5_Right_193 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_154_5_Right_192 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_153_5_Right_191 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_152_5_Right_190 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_151_5_Right_189 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_150_5_Right_188 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_149_5_Right_187 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_148_5_Right_186 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_147_5_Right_185 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_146_5_Right_184 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_145_5_Right_183 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_144_5_Right_182 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_143_5_Right_181 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_142_5_Right_180 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_141_5_Right_179 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_140_5_Right_178 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_139_5_Right_177 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_138_5_Right_176 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_137_5_Right_175 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_136_5_Right_174 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_135_5_Right_173 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_134_5_Right_172 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_133_5_Right_171 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_132_5_Right_170 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_131_5_Right_169 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_130_5_Right_168 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_129_5_Right_167 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_128_5_Right_166 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_127_5_Right_165 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_126_5_Right_164 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_125_5_Right_163 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_124_5_Right_162 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_123_5_Right_161 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_122_5_Right_160 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_121_5_Right_159 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_120_5_Right_158 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_119_5_Right_157 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_118_5_Right_156 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_117_5_Right_155 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_116_5_Right_154 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_115_5_Right_153 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_114_5_Right_152 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_113_5_Right_151 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_112_5_Right_150 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_111_5_Right_149 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_110_5_Right_148 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_109_5_Right_147 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_108_5_Right_146 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_107_5_Right_145 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_106_5_Right_144 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_105_5_Right_143 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_104_5_Right_142 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_103_5_Right_141 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_102_5_Right_140 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_101_5_Right_139 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_100_5_Right_138 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_99_5_Right_137 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_98_5_Right_136 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_97_5_Right_135 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_96_5_Right_134 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_95_5_Right_133 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_94_5_Right_132 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_81_5_Right_131 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_80_5_Right_130 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_79_5_Right_129 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_78_5_Right_128 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_77_5_Right_127 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_76_5_Right_126 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_75_5_Right_125 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_74_5_Right_124 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_73_5_Right_123 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_72_5_Right_122 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_71_5_Right_121 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_70_5_Right_120 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_69_5_Right_119 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_68_5_Right_118 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_67_5_Right_117 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_66_5_Right_116 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_65_5_Right_115 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_64_5_Right_114 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_63_5_Right_113 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_62_5_Right_112 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_61_5_Right_111 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_60_5_Right_110 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_59_5_Right_109 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_58_5_Right_108 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_57_5_Right_107 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_56_5_Right_106 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_55_5_Right_105 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_5_Right_104 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_5_Right_103 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_5_Right_102 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_5_Right_101 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_5_Right_100 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_5_Right_99 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_5_Right_98 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_5_Right_97 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_5_Right_96 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_5_Right_95 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_5_Right_94 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_5_Right_93 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_5_Right_92 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_5_Right_91 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_5_Right_90 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_5_Right_89 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_5_Right_88 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_5_Right_87 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_5_Right_86 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_5_Right_85 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_5_Right_84 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_5_Right_83 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_5_Right_82 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_5_Right_81 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_5_Right_80 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_5_Right_79 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_5_Right_78 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_5_Right_77 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_5_Right_76 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_5_Right_75 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_5_Right_74 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_5_Right_73 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_5_Right_72 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_5_Right_71 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_5_Right_70 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_5_Right_69 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_5_Right_68 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_5_Right_67 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_5_Right_66 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_5_Right_65 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_5_Right_64 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_335_Right_63 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_334_Right_62 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_333_Right_61 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_332_Right_60 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_331_Right_59 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_330_Right_58 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_329_Right_57 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_328_Right_56 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_327_Right_55 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_326_Right_54 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_325_Right_53 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_324_Right_52 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_323_Right_51 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_322_Right_50 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_253_Right_49 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_252_Right_48 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_251_Right_47 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_250_Right_46 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_249_Right_45 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_248_Right_44 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_247_Right_43 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_246_Right_42 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_245_Right_41 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_244_Right_40 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_243_Right_39 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_242_Right_38 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_173_Right_37 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_172_Right_36 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_171_Right_35 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_170_Right_34 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_169_Right_33 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_168_Right_32 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_167_Right_31 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_166_Right_30 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_165_Right_29 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_164_Right_28 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_163_Right_27 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_162_Right_26 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_93_Right_25 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_92_Right_24 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_91_Right_23 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_90_Right_22 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_89_Right_21 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_88_Right_20 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_87_Right_19 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_86_Right_18 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_85_Right_17 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_84_Right_16 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_83_Right_15 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_82_Right_14 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Right_0 ();
 TIELOx1_ASAP7_75t_R ces_3_0_12 (.L(net11));
 TIELOx1_ASAP7_75t_R ces_3_0_11 (.L(net10));
 TIELOx1_ASAP7_75t_R ces_3_0_10 (.L(net9));
 TIELOx1_ASAP7_75t_R ces_2_0_9 (.L(net8));
 TIELOx1_ASAP7_75t_R ces_2_0_8 (.L(net7));
 TIELOx1_ASAP7_75t_R ces_2_0_7 (.L(net6));
 TIELOx1_ASAP7_75t_R ces_1_0_6 (.L(net5));
 TIELOx1_ASAP7_75t_R ces_1_0_5 (.L(net4));
 TIELOx1_ASAP7_75t_R ces_1_0_4 (.L(net3));
 TIELOx1_ASAP7_75t_R ces_0_0_3 (.L(net2));
 TIELOx1_ASAP7_75t_R ces_0_0_2 (.L(net1));
 TIELOx1_ASAP7_75t_R ces_0_0_1 (.L(net));
 DFFHQNx1_ASAP7_75t_R \REG_0$_DFF_P_  (.CLK(clknet_1_0__leaf_clock_regs),
    .D(_ces_0_3_io_lsbOuts_0),
    .QN(_01_));
 DFFHQNx1_ASAP7_75t_R \REG_1$_DFF_P_  (.CLK(clknet_1_0__leaf_clock_regs),
    .D(_ces_0_3_io_lsbOuts_1),
    .QN(_02_));
 DFFHQNx1_ASAP7_75t_R \REG_10$_DFF_P_  (.CLK(clknet_1_1__leaf_clock_regs),
    .D(_ces_2_3_io_lsbOuts_2),
    .QN(_03_));
 DFFHQNx1_ASAP7_75t_R \REG_11$_DFF_P_  (.CLK(clknet_1_1__leaf_clock_regs),
    .D(_ces_2_3_io_lsbOuts_3),
    .QN(_04_));
 DFFHQNx1_ASAP7_75t_R \REG_12$_DFF_P_  (.CLK(clknet_1_1__leaf_clock_regs),
    .D(_ces_3_3_io_lsbOuts_0),
    .QN(_05_));
 DFFHQNx1_ASAP7_75t_R \REG_13$_DFF_P_  (.CLK(clknet_1_1__leaf_clock_regs),
    .D(_ces_3_3_io_lsbOuts_1),
    .QN(_06_));
 DFFHQNx1_ASAP7_75t_R \REG_14$_DFF_P_  (.CLK(clknet_1_1__leaf_clock_regs),
    .D(_ces_3_3_io_lsbOuts_2),
    .QN(_07_));
 DFFHQNx1_ASAP7_75t_R \REG_15$_DFF_P_  (.CLK(clknet_1_1__leaf_clock_regs),
    .D(_ces_3_3_io_lsbOuts_3),
    .QN(_08_));
 DFFHQNx1_ASAP7_75t_R \REG_2$_DFF_P_  (.CLK(clknet_1_0__leaf_clock_regs),
    .D(_ces_0_3_io_lsbOuts_2),
    .QN(_09_));
 DFFHQNx1_ASAP7_75t_R \REG_3$_DFF_P_  (.CLK(clknet_1_0__leaf_clock_regs),
    .D(_ces_0_3_io_lsbOuts_3),
    .QN(_10_));
 DFFHQNx1_ASAP7_75t_R \REG_4$_DFF_P_  (.CLK(clknet_1_0__leaf_clock_regs),
    .D(_ces_1_3_io_lsbOuts_0),
    .QN(_11_));
 DFFHQNx1_ASAP7_75t_R \REG_5$_DFF_P_  (.CLK(clknet_1_0__leaf_clock_regs),
    .D(_ces_1_3_io_lsbOuts_1),
    .QN(_12_));
 DFFHQNx1_ASAP7_75t_R \REG_6$_DFF_P_  (.CLK(clknet_1_0__leaf_clock_regs),
    .D(_ces_1_3_io_lsbOuts_2),
    .QN(_13_));
 DFFHQNx1_ASAP7_75t_R \REG_7$_DFF_P_  (.CLK(clknet_1_0__leaf_clock_regs),
    .D(_ces_1_3_io_lsbOuts_3),
    .QN(_14_));
 DFFHQNx1_ASAP7_75t_R \REG_8$_DFF_P_  (.CLK(clknet_1_1__leaf_clock_regs),
    .D(_ces_2_3_io_lsbOuts_0),
    .QN(_15_));
 DFFHQNx1_ASAP7_75t_R \REG_9$_DFF_P_  (.CLK(clknet_1_1__leaf_clock_regs),
    .D(_ces_2_3_io_lsbOuts_1),
    .QN(_00_));
 INVx3_ASAP7_75t_R _17_ (.A(_00_),
    .Y(net1051));
 INVx3_ASAP7_75t_R _18_ (.A(_01_),
    .Y(net1036));
 INVx3_ASAP7_75t_R _19_ (.A(_02_),
    .Y(net1037));
 INVx3_ASAP7_75t_R _20_ (.A(_03_),
    .Y(net1038));
 INVx3_ASAP7_75t_R _21_ (.A(_04_),
    .Y(net1039));
 INVx3_ASAP7_75t_R _22_ (.A(_05_),
    .Y(net1040));
 INVx3_ASAP7_75t_R _23_ (.A(_06_),
    .Y(net1041));
 INVx3_ASAP7_75t_R _24_ (.A(_07_),
    .Y(net1042));
 INVx3_ASAP7_75t_R _25_ (.A(_08_),
    .Y(net1043));
 INVx3_ASAP7_75t_R _26_ (.A(_09_),
    .Y(net1044));
 INVx3_ASAP7_75t_R _27_ (.A(_10_),
    .Y(net1045));
 INVx3_ASAP7_75t_R _28_ (.A(_11_),
    .Y(net1046));
 INVx3_ASAP7_75t_R _29_ (.A(_12_),
    .Y(net1047));
 INVx3_ASAP7_75t_R _30_ (.A(_13_),
    .Y(net1048));
 INVx3_ASAP7_75t_R _31_ (.A(_14_),
    .Y(net1049));
 INVx3_ASAP7_75t_R _32_ (.A(_15_),
    .Y(net1050));
 Element ces_0_0 (.clock(clknet_leaf_3_clock),
    .io_lsbIns_1(net),
    .io_lsbIns_2(net1),
    .io_lsbIns_3(net2),
    .io_lsbOuts_1(_ces_0_0_io_lsbOuts_1),
    .io_lsbOuts_2(_ces_0_0_io_lsbOuts_2),
    .io_lsbOuts_3(_ces_0_0_io_lsbOuts_3),
    .io_ins_down({\_ces_1_0_io_outs_down[63] ,
    \_ces_1_0_io_outs_down[62] ,
    \_ces_1_0_io_outs_down[61] ,
    \_ces_1_0_io_outs_down[60] ,
    \_ces_1_0_io_outs_down[59] ,
    \_ces_1_0_io_outs_down[58] ,
    \_ces_1_0_io_outs_down[57] ,
    \_ces_1_0_io_outs_down[56] ,
    \_ces_1_0_io_outs_down[55] ,
    \_ces_1_0_io_outs_down[54] ,
    \_ces_1_0_io_outs_down[53] ,
    \_ces_1_0_io_outs_down[52] ,
    \_ces_1_0_io_outs_down[51] ,
    \_ces_1_0_io_outs_down[50] ,
    \_ces_1_0_io_outs_down[49] ,
    \_ces_1_0_io_outs_down[48] ,
    \_ces_1_0_io_outs_down[47] ,
    \_ces_1_0_io_outs_down[46] ,
    \_ces_1_0_io_outs_down[45] ,
    \_ces_1_0_io_outs_down[44] ,
    \_ces_1_0_io_outs_down[43] ,
    \_ces_1_0_io_outs_down[42] ,
    \_ces_1_0_io_outs_down[41] ,
    \_ces_1_0_io_outs_down[40] ,
    \_ces_1_0_io_outs_down[39] ,
    \_ces_1_0_io_outs_down[38] ,
    \_ces_1_0_io_outs_down[37] ,
    \_ces_1_0_io_outs_down[36] ,
    \_ces_1_0_io_outs_down[35] ,
    \_ces_1_0_io_outs_down[34] ,
    \_ces_1_0_io_outs_down[33] ,
    \_ces_1_0_io_outs_down[32] ,
    \_ces_1_0_io_outs_down[31] ,
    \_ces_1_0_io_outs_down[30] ,
    \_ces_1_0_io_outs_down[29] ,
    \_ces_1_0_io_outs_down[28] ,
    \_ces_1_0_io_outs_down[27] ,
    \_ces_1_0_io_outs_down[26] ,
    \_ces_1_0_io_outs_down[25] ,
    \_ces_1_0_io_outs_down[24] ,
    \_ces_1_0_io_outs_down[23] ,
    \_ces_1_0_io_outs_down[22] ,
    \_ces_1_0_io_outs_down[21] ,
    \_ces_1_0_io_outs_down[20] ,
    \_ces_1_0_io_outs_down[19] ,
    \_ces_1_0_io_outs_down[18] ,
    \_ces_1_0_io_outs_down[17] ,
    \_ces_1_0_io_outs_down[16] ,
    \_ces_1_0_io_outs_down[15] ,
    \_ces_1_0_io_outs_down[14] ,
    \_ces_1_0_io_outs_down[13] ,
    \_ces_1_0_io_outs_down[12] ,
    \_ces_1_0_io_outs_down[11] ,
    \_ces_1_0_io_outs_down[10] ,
    \_ces_1_0_io_outs_down[9] ,
    \_ces_1_0_io_outs_down[8] ,
    \_ces_1_0_io_outs_down[7] ,
    \_ces_1_0_io_outs_down[6] ,
    \_ces_1_0_io_outs_down[5] ,
    \_ces_1_0_io_outs_down[4] ,
    \_ces_1_0_io_outs_down[3] ,
    \_ces_1_0_io_outs_down[2] ,
    \_ces_1_0_io_outs_down[1] ,
    \_ces_1_0_io_outs_down[0] }),
    .io_ins_left({\_ces_0_1_io_outs_left[63] ,
    \_ces_0_1_io_outs_left[62] ,
    \_ces_0_1_io_outs_left[61] ,
    \_ces_0_1_io_outs_left[60] ,
    \_ces_0_1_io_outs_left[59] ,
    \_ces_0_1_io_outs_left[58] ,
    \_ces_0_1_io_outs_left[57] ,
    \_ces_0_1_io_outs_left[56] ,
    \_ces_0_1_io_outs_left[55] ,
    \_ces_0_1_io_outs_left[54] ,
    \_ces_0_1_io_outs_left[53] ,
    \_ces_0_1_io_outs_left[52] ,
    \_ces_0_1_io_outs_left[51] ,
    \_ces_0_1_io_outs_left[50] ,
    \_ces_0_1_io_outs_left[49] ,
    \_ces_0_1_io_outs_left[48] ,
    \_ces_0_1_io_outs_left[47] ,
    \_ces_0_1_io_outs_left[46] ,
    \_ces_0_1_io_outs_left[45] ,
    \_ces_0_1_io_outs_left[44] ,
    \_ces_0_1_io_outs_left[43] ,
    \_ces_0_1_io_outs_left[42] ,
    \_ces_0_1_io_outs_left[41] ,
    \_ces_0_1_io_outs_left[40] ,
    \_ces_0_1_io_outs_left[39] ,
    \_ces_0_1_io_outs_left[38] ,
    \_ces_0_1_io_outs_left[37] ,
    \_ces_0_1_io_outs_left[36] ,
    \_ces_0_1_io_outs_left[35] ,
    \_ces_0_1_io_outs_left[34] ,
    \_ces_0_1_io_outs_left[33] ,
    \_ces_0_1_io_outs_left[32] ,
    \_ces_0_1_io_outs_left[31] ,
    \_ces_0_1_io_outs_left[30] ,
    \_ces_0_1_io_outs_left[29] ,
    \_ces_0_1_io_outs_left[28] ,
    \_ces_0_1_io_outs_left[27] ,
    \_ces_0_1_io_outs_left[26] ,
    \_ces_0_1_io_outs_left[25] ,
    \_ces_0_1_io_outs_left[24] ,
    \_ces_0_1_io_outs_left[23] ,
    \_ces_0_1_io_outs_left[22] ,
    \_ces_0_1_io_outs_left[21] ,
    \_ces_0_1_io_outs_left[20] ,
    \_ces_0_1_io_outs_left[19] ,
    \_ces_0_1_io_outs_left[18] ,
    \_ces_0_1_io_outs_left[17] ,
    \_ces_0_1_io_outs_left[16] ,
    \_ces_0_1_io_outs_left[15] ,
    \_ces_0_1_io_outs_left[14] ,
    \_ces_0_1_io_outs_left[13] ,
    \_ces_0_1_io_outs_left[12] ,
    \_ces_0_1_io_outs_left[11] ,
    \_ces_0_1_io_outs_left[10] ,
    \_ces_0_1_io_outs_left[9] ,
    \_ces_0_1_io_outs_left[8] ,
    \_ces_0_1_io_outs_left[7] ,
    \_ces_0_1_io_outs_left[6] ,
    \_ces_0_1_io_outs_left[5] ,
    \_ces_0_1_io_outs_left[4] ,
    \_ces_0_1_io_outs_left[3] ,
    \_ces_0_1_io_outs_left[2] ,
    \_ces_0_1_io_outs_left[1] ,
    \_ces_0_1_io_outs_left[0] }),
    .io_ins_right({net583,
    net582,
    net581,
    net580,
    net578,
    net577,
    net576,
    net575,
    net574,
    net573,
    net572,
    net571,
    net570,
    net569,
    net567,
    net566,
    net565,
    net564,
    net563,
    net562,
    net561,
    net560,
    net559,
    net558,
    net556,
    net555,
    net554,
    net553,
    net552,
    net551,
    net550,
    net549,
    net548,
    net547,
    net545,
    net544,
    net543,
    net542,
    net541,
    net540,
    net539,
    net538,
    net537,
    net536,
    net534,
    net533,
    net532,
    net531,
    net530,
    net529,
    net528,
    net527,
    net526,
    net525,
    net587,
    net586,
    net585,
    net584,
    net579,
    net568,
    net557,
    net546,
    net535,
    net524}),
    .io_ins_up({net839,
    net838,
    net837,
    net836,
    net834,
    net833,
    net832,
    net831,
    net830,
    net829,
    net828,
    net827,
    net826,
    net825,
    net823,
    net822,
    net821,
    net820,
    net819,
    net818,
    net817,
    net816,
    net815,
    net814,
    net812,
    net811,
    net810,
    net809,
    net808,
    net807,
    net806,
    net805,
    net804,
    net803,
    net801,
    net800,
    net799,
    net798,
    net797,
    net796,
    net795,
    net794,
    net793,
    net792,
    net790,
    net789,
    net788,
    net787,
    net786,
    net785,
    net784,
    net783,
    net782,
    net781,
    net843,
    net842,
    net841,
    net840,
    net835,
    net824,
    net813,
    net802,
    net791,
    net780}),
    .io_outs_down({net1111,
    net1110,
    net1109,
    net1108,
    net1106,
    net1105,
    net1104,
    net1103,
    net1102,
    net1101,
    net1100,
    net1099,
    net1098,
    net1097,
    net1095,
    net1094,
    net1093,
    net1092,
    net1091,
    net1090,
    net1089,
    net1088,
    net1087,
    net1086,
    net1084,
    net1083,
    net1082,
    net1081,
    net1080,
    net1079,
    net1078,
    net1077,
    net1076,
    net1075,
    net1073,
    net1072,
    net1071,
    net1070,
    net1069,
    net1068,
    net1067,
    net1066,
    net1065,
    net1064,
    net1062,
    net1061,
    net1060,
    net1059,
    net1058,
    net1057,
    net1056,
    net1055,
    net1054,
    net1053,
    net1115,
    net1114,
    net1113,
    net1112,
    net1107,
    net1096,
    net1085,
    net1074,
    net1063,
    net1052}),
    .io_outs_left({net1367,
    net1366,
    net1365,
    net1364,
    net1362,
    net1361,
    net1360,
    net1359,
    net1358,
    net1357,
    net1356,
    net1355,
    net1354,
    net1353,
    net1351,
    net1350,
    net1349,
    net1348,
    net1347,
    net1346,
    net1345,
    net1344,
    net1343,
    net1342,
    net1340,
    net1339,
    net1338,
    net1337,
    net1336,
    net1335,
    net1334,
    net1333,
    net1332,
    net1331,
    net1329,
    net1328,
    net1327,
    net1326,
    net1325,
    net1324,
    net1323,
    net1322,
    net1321,
    net1320,
    net1318,
    net1317,
    net1316,
    net1315,
    net1314,
    net1313,
    net1312,
    net1311,
    net1310,
    net1309,
    net1371,
    net1370,
    net1369,
    net1368,
    net1363,
    net1352,
    net1341,
    net1330,
    net1319,
    net1308}),
    .io_outs_right({\_ces_0_0_io_outs_right[63] ,
    \_ces_0_0_io_outs_right[62] ,
    \_ces_0_0_io_outs_right[61] ,
    \_ces_0_0_io_outs_right[60] ,
    \_ces_0_0_io_outs_right[59] ,
    \_ces_0_0_io_outs_right[58] ,
    \_ces_0_0_io_outs_right[57] ,
    \_ces_0_0_io_outs_right[56] ,
    \_ces_0_0_io_outs_right[55] ,
    \_ces_0_0_io_outs_right[54] ,
    \_ces_0_0_io_outs_right[53] ,
    \_ces_0_0_io_outs_right[52] ,
    \_ces_0_0_io_outs_right[51] ,
    \_ces_0_0_io_outs_right[50] ,
    \_ces_0_0_io_outs_right[49] ,
    \_ces_0_0_io_outs_right[48] ,
    \_ces_0_0_io_outs_right[47] ,
    \_ces_0_0_io_outs_right[46] ,
    \_ces_0_0_io_outs_right[45] ,
    \_ces_0_0_io_outs_right[44] ,
    \_ces_0_0_io_outs_right[43] ,
    \_ces_0_0_io_outs_right[42] ,
    \_ces_0_0_io_outs_right[41] ,
    \_ces_0_0_io_outs_right[40] ,
    \_ces_0_0_io_outs_right[39] ,
    \_ces_0_0_io_outs_right[38] ,
    \_ces_0_0_io_outs_right[37] ,
    \_ces_0_0_io_outs_right[36] ,
    \_ces_0_0_io_outs_right[35] ,
    \_ces_0_0_io_outs_right[34] ,
    \_ces_0_0_io_outs_right[33] ,
    \_ces_0_0_io_outs_right[32] ,
    \_ces_0_0_io_outs_right[31] ,
    \_ces_0_0_io_outs_right[30] ,
    \_ces_0_0_io_outs_right[29] ,
    \_ces_0_0_io_outs_right[28] ,
    \_ces_0_0_io_outs_right[27] ,
    \_ces_0_0_io_outs_right[26] ,
    \_ces_0_0_io_outs_right[25] ,
    \_ces_0_0_io_outs_right[24] ,
    \_ces_0_0_io_outs_right[23] ,
    \_ces_0_0_io_outs_right[22] ,
    \_ces_0_0_io_outs_right[21] ,
    \_ces_0_0_io_outs_right[20] ,
    \_ces_0_0_io_outs_right[19] ,
    \_ces_0_0_io_outs_right[18] ,
    \_ces_0_0_io_outs_right[17] ,
    \_ces_0_0_io_outs_right[16] ,
    \_ces_0_0_io_outs_right[15] ,
    \_ces_0_0_io_outs_right[14] ,
    \_ces_0_0_io_outs_right[13] ,
    \_ces_0_0_io_outs_right[12] ,
    \_ces_0_0_io_outs_right[11] ,
    \_ces_0_0_io_outs_right[10] ,
    \_ces_0_0_io_outs_right[9] ,
    \_ces_0_0_io_outs_right[8] ,
    \_ces_0_0_io_outs_right[7] ,
    \_ces_0_0_io_outs_right[6] ,
    \_ces_0_0_io_outs_right[5] ,
    \_ces_0_0_io_outs_right[4] ,
    \_ces_0_0_io_outs_right[3] ,
    \_ces_0_0_io_outs_right[2] ,
    \_ces_0_0_io_outs_right[1] ,
    \_ces_0_0_io_outs_right[0] }),
    .io_outs_up({\_ces_0_0_io_outs_up[63] ,
    \_ces_0_0_io_outs_up[62] ,
    \_ces_0_0_io_outs_up[61] ,
    \_ces_0_0_io_outs_up[60] ,
    \_ces_0_0_io_outs_up[59] ,
    \_ces_0_0_io_outs_up[58] ,
    \_ces_0_0_io_outs_up[57] ,
    \_ces_0_0_io_outs_up[56] ,
    \_ces_0_0_io_outs_up[55] ,
    \_ces_0_0_io_outs_up[54] ,
    \_ces_0_0_io_outs_up[53] ,
    \_ces_0_0_io_outs_up[52] ,
    \_ces_0_0_io_outs_up[51] ,
    \_ces_0_0_io_outs_up[50] ,
    \_ces_0_0_io_outs_up[49] ,
    \_ces_0_0_io_outs_up[48] ,
    \_ces_0_0_io_outs_up[47] ,
    \_ces_0_0_io_outs_up[46] ,
    \_ces_0_0_io_outs_up[45] ,
    \_ces_0_0_io_outs_up[44] ,
    \_ces_0_0_io_outs_up[43] ,
    \_ces_0_0_io_outs_up[42] ,
    \_ces_0_0_io_outs_up[41] ,
    \_ces_0_0_io_outs_up[40] ,
    \_ces_0_0_io_outs_up[39] ,
    \_ces_0_0_io_outs_up[38] ,
    \_ces_0_0_io_outs_up[37] ,
    \_ces_0_0_io_outs_up[36] ,
    \_ces_0_0_io_outs_up[35] ,
    \_ces_0_0_io_outs_up[34] ,
    \_ces_0_0_io_outs_up[33] ,
    \_ces_0_0_io_outs_up[32] ,
    \_ces_0_0_io_outs_up[31] ,
    \_ces_0_0_io_outs_up[30] ,
    \_ces_0_0_io_outs_up[29] ,
    \_ces_0_0_io_outs_up[28] ,
    \_ces_0_0_io_outs_up[27] ,
    \_ces_0_0_io_outs_up[26] ,
    \_ces_0_0_io_outs_up[25] ,
    \_ces_0_0_io_outs_up[24] ,
    \_ces_0_0_io_outs_up[23] ,
    \_ces_0_0_io_outs_up[22] ,
    \_ces_0_0_io_outs_up[21] ,
    \_ces_0_0_io_outs_up[20] ,
    \_ces_0_0_io_outs_up[19] ,
    \_ces_0_0_io_outs_up[18] ,
    \_ces_0_0_io_outs_up[17] ,
    \_ces_0_0_io_outs_up[16] ,
    \_ces_0_0_io_outs_up[15] ,
    \_ces_0_0_io_outs_up[14] ,
    \_ces_0_0_io_outs_up[13] ,
    \_ces_0_0_io_outs_up[12] ,
    \_ces_0_0_io_outs_up[11] ,
    \_ces_0_0_io_outs_up[10] ,
    \_ces_0_0_io_outs_up[9] ,
    \_ces_0_0_io_outs_up[8] ,
    \_ces_0_0_io_outs_up[7] ,
    \_ces_0_0_io_outs_up[6] ,
    \_ces_0_0_io_outs_up[5] ,
    \_ces_0_0_io_outs_up[4] ,
    \_ces_0_0_io_outs_up[3] ,
    \_ces_0_0_io_outs_up[2] ,
    \_ces_0_0_io_outs_up[1] ,
    \_ces_0_0_io_outs_up[0] }));
 Element ces_0_1 (.clock(clknet_leaf_3_clock),
    .io_lsbIns_1(_ces_0_0_io_lsbOuts_1),
    .io_lsbIns_2(_ces_0_0_io_lsbOuts_2),
    .io_lsbIns_3(_ces_0_0_io_lsbOuts_3),
    .io_lsbOuts_1(_ces_0_1_io_lsbOuts_1),
    .io_lsbOuts_2(_ces_0_1_io_lsbOuts_2),
    .io_lsbOuts_3(_ces_0_1_io_lsbOuts_3),
    .io_ins_down({\_ces_1_1_io_outs_down[63] ,
    \_ces_1_1_io_outs_down[62] ,
    \_ces_1_1_io_outs_down[61] ,
    \_ces_1_1_io_outs_down[60] ,
    \_ces_1_1_io_outs_down[59] ,
    \_ces_1_1_io_outs_down[58] ,
    \_ces_1_1_io_outs_down[57] ,
    \_ces_1_1_io_outs_down[56] ,
    \_ces_1_1_io_outs_down[55] ,
    \_ces_1_1_io_outs_down[54] ,
    \_ces_1_1_io_outs_down[53] ,
    \_ces_1_1_io_outs_down[52] ,
    \_ces_1_1_io_outs_down[51] ,
    \_ces_1_1_io_outs_down[50] ,
    \_ces_1_1_io_outs_down[49] ,
    \_ces_1_1_io_outs_down[48] ,
    \_ces_1_1_io_outs_down[47] ,
    \_ces_1_1_io_outs_down[46] ,
    \_ces_1_1_io_outs_down[45] ,
    \_ces_1_1_io_outs_down[44] ,
    \_ces_1_1_io_outs_down[43] ,
    \_ces_1_1_io_outs_down[42] ,
    \_ces_1_1_io_outs_down[41] ,
    \_ces_1_1_io_outs_down[40] ,
    \_ces_1_1_io_outs_down[39] ,
    \_ces_1_1_io_outs_down[38] ,
    \_ces_1_1_io_outs_down[37] ,
    \_ces_1_1_io_outs_down[36] ,
    \_ces_1_1_io_outs_down[35] ,
    \_ces_1_1_io_outs_down[34] ,
    \_ces_1_1_io_outs_down[33] ,
    \_ces_1_1_io_outs_down[32] ,
    \_ces_1_1_io_outs_down[31] ,
    \_ces_1_1_io_outs_down[30] ,
    \_ces_1_1_io_outs_down[29] ,
    \_ces_1_1_io_outs_down[28] ,
    \_ces_1_1_io_outs_down[27] ,
    \_ces_1_1_io_outs_down[26] ,
    \_ces_1_1_io_outs_down[25] ,
    \_ces_1_1_io_outs_down[24] ,
    \_ces_1_1_io_outs_down[23] ,
    \_ces_1_1_io_outs_down[22] ,
    \_ces_1_1_io_outs_down[21] ,
    \_ces_1_1_io_outs_down[20] ,
    \_ces_1_1_io_outs_down[19] ,
    \_ces_1_1_io_outs_down[18] ,
    \_ces_1_1_io_outs_down[17] ,
    \_ces_1_1_io_outs_down[16] ,
    \_ces_1_1_io_outs_down[15] ,
    \_ces_1_1_io_outs_down[14] ,
    \_ces_1_1_io_outs_down[13] ,
    \_ces_1_1_io_outs_down[12] ,
    \_ces_1_1_io_outs_down[11] ,
    \_ces_1_1_io_outs_down[10] ,
    \_ces_1_1_io_outs_down[9] ,
    \_ces_1_1_io_outs_down[8] ,
    \_ces_1_1_io_outs_down[7] ,
    \_ces_1_1_io_outs_down[6] ,
    \_ces_1_1_io_outs_down[5] ,
    \_ces_1_1_io_outs_down[4] ,
    \_ces_1_1_io_outs_down[3] ,
    \_ces_1_1_io_outs_down[2] ,
    \_ces_1_1_io_outs_down[1] ,
    \_ces_1_1_io_outs_down[0] }),
    .io_ins_left({\_ces_0_2_io_outs_left[63] ,
    \_ces_0_2_io_outs_left[62] ,
    \_ces_0_2_io_outs_left[61] ,
    \_ces_0_2_io_outs_left[60] ,
    \_ces_0_2_io_outs_left[59] ,
    \_ces_0_2_io_outs_left[58] ,
    \_ces_0_2_io_outs_left[57] ,
    \_ces_0_2_io_outs_left[56] ,
    \_ces_0_2_io_outs_left[55] ,
    \_ces_0_2_io_outs_left[54] ,
    \_ces_0_2_io_outs_left[53] ,
    \_ces_0_2_io_outs_left[52] ,
    \_ces_0_2_io_outs_left[51] ,
    \_ces_0_2_io_outs_left[50] ,
    \_ces_0_2_io_outs_left[49] ,
    \_ces_0_2_io_outs_left[48] ,
    \_ces_0_2_io_outs_left[47] ,
    \_ces_0_2_io_outs_left[46] ,
    \_ces_0_2_io_outs_left[45] ,
    \_ces_0_2_io_outs_left[44] ,
    \_ces_0_2_io_outs_left[43] ,
    \_ces_0_2_io_outs_left[42] ,
    \_ces_0_2_io_outs_left[41] ,
    \_ces_0_2_io_outs_left[40] ,
    \_ces_0_2_io_outs_left[39] ,
    \_ces_0_2_io_outs_left[38] ,
    \_ces_0_2_io_outs_left[37] ,
    \_ces_0_2_io_outs_left[36] ,
    \_ces_0_2_io_outs_left[35] ,
    \_ces_0_2_io_outs_left[34] ,
    \_ces_0_2_io_outs_left[33] ,
    \_ces_0_2_io_outs_left[32] ,
    \_ces_0_2_io_outs_left[31] ,
    \_ces_0_2_io_outs_left[30] ,
    \_ces_0_2_io_outs_left[29] ,
    \_ces_0_2_io_outs_left[28] ,
    \_ces_0_2_io_outs_left[27] ,
    \_ces_0_2_io_outs_left[26] ,
    \_ces_0_2_io_outs_left[25] ,
    \_ces_0_2_io_outs_left[24] ,
    \_ces_0_2_io_outs_left[23] ,
    \_ces_0_2_io_outs_left[22] ,
    \_ces_0_2_io_outs_left[21] ,
    \_ces_0_2_io_outs_left[20] ,
    \_ces_0_2_io_outs_left[19] ,
    \_ces_0_2_io_outs_left[18] ,
    \_ces_0_2_io_outs_left[17] ,
    \_ces_0_2_io_outs_left[16] ,
    \_ces_0_2_io_outs_left[15] ,
    \_ces_0_2_io_outs_left[14] ,
    \_ces_0_2_io_outs_left[13] ,
    \_ces_0_2_io_outs_left[12] ,
    \_ces_0_2_io_outs_left[11] ,
    \_ces_0_2_io_outs_left[10] ,
    \_ces_0_2_io_outs_left[9] ,
    \_ces_0_2_io_outs_left[8] ,
    \_ces_0_2_io_outs_left[7] ,
    \_ces_0_2_io_outs_left[6] ,
    \_ces_0_2_io_outs_left[5] ,
    \_ces_0_2_io_outs_left[4] ,
    \_ces_0_2_io_outs_left[3] ,
    \_ces_0_2_io_outs_left[2] ,
    \_ces_0_2_io_outs_left[1] ,
    \_ces_0_2_io_outs_left[0] }),
    .io_ins_right({\_ces_0_0_io_outs_right[63] ,
    \_ces_0_0_io_outs_right[62] ,
    \_ces_0_0_io_outs_right[61] ,
    \_ces_0_0_io_outs_right[60] ,
    \_ces_0_0_io_outs_right[59] ,
    \_ces_0_0_io_outs_right[58] ,
    \_ces_0_0_io_outs_right[57] ,
    \_ces_0_0_io_outs_right[56] ,
    \_ces_0_0_io_outs_right[55] ,
    \_ces_0_0_io_outs_right[54] ,
    \_ces_0_0_io_outs_right[53] ,
    \_ces_0_0_io_outs_right[52] ,
    \_ces_0_0_io_outs_right[51] ,
    \_ces_0_0_io_outs_right[50] ,
    \_ces_0_0_io_outs_right[49] ,
    \_ces_0_0_io_outs_right[48] ,
    \_ces_0_0_io_outs_right[47] ,
    \_ces_0_0_io_outs_right[46] ,
    \_ces_0_0_io_outs_right[45] ,
    \_ces_0_0_io_outs_right[44] ,
    \_ces_0_0_io_outs_right[43] ,
    \_ces_0_0_io_outs_right[42] ,
    \_ces_0_0_io_outs_right[41] ,
    \_ces_0_0_io_outs_right[40] ,
    \_ces_0_0_io_outs_right[39] ,
    \_ces_0_0_io_outs_right[38] ,
    \_ces_0_0_io_outs_right[37] ,
    \_ces_0_0_io_outs_right[36] ,
    \_ces_0_0_io_outs_right[35] ,
    \_ces_0_0_io_outs_right[34] ,
    \_ces_0_0_io_outs_right[33] ,
    \_ces_0_0_io_outs_right[32] ,
    \_ces_0_0_io_outs_right[31] ,
    \_ces_0_0_io_outs_right[30] ,
    \_ces_0_0_io_outs_right[29] ,
    \_ces_0_0_io_outs_right[28] ,
    \_ces_0_0_io_outs_right[27] ,
    \_ces_0_0_io_outs_right[26] ,
    \_ces_0_0_io_outs_right[25] ,
    \_ces_0_0_io_outs_right[24] ,
    \_ces_0_0_io_outs_right[23] ,
    \_ces_0_0_io_outs_right[22] ,
    \_ces_0_0_io_outs_right[21] ,
    \_ces_0_0_io_outs_right[20] ,
    \_ces_0_0_io_outs_right[19] ,
    \_ces_0_0_io_outs_right[18] ,
    \_ces_0_0_io_outs_right[17] ,
    \_ces_0_0_io_outs_right[16] ,
    \_ces_0_0_io_outs_right[15] ,
    \_ces_0_0_io_outs_right[14] ,
    \_ces_0_0_io_outs_right[13] ,
    \_ces_0_0_io_outs_right[12] ,
    \_ces_0_0_io_outs_right[11] ,
    \_ces_0_0_io_outs_right[10] ,
    \_ces_0_0_io_outs_right[9] ,
    \_ces_0_0_io_outs_right[8] ,
    \_ces_0_0_io_outs_right[7] ,
    \_ces_0_0_io_outs_right[6] ,
    \_ces_0_0_io_outs_right[5] ,
    \_ces_0_0_io_outs_right[4] ,
    \_ces_0_0_io_outs_right[3] ,
    \_ces_0_0_io_outs_right[2] ,
    \_ces_0_0_io_outs_right[1] ,
    \_ces_0_0_io_outs_right[0] }),
    .io_ins_up({net903,
    net902,
    net901,
    net900,
    net898,
    net897,
    net896,
    net895,
    net894,
    net893,
    net892,
    net891,
    net890,
    net889,
    net887,
    net886,
    net885,
    net884,
    net883,
    net882,
    net881,
    net880,
    net879,
    net878,
    net876,
    net875,
    net874,
    net873,
    net872,
    net871,
    net870,
    net869,
    net868,
    net867,
    net865,
    net864,
    net863,
    net862,
    net861,
    net860,
    net859,
    net858,
    net857,
    net856,
    net854,
    net853,
    net852,
    net851,
    net850,
    net849,
    net848,
    net847,
    net846,
    net845,
    net907,
    net906,
    net905,
    net904,
    net899,
    net888,
    net877,
    net866,
    net855,
    net844}),
    .io_outs_down({net1175,
    net1174,
    net1173,
    net1172,
    net1170,
    net1169,
    net1168,
    net1167,
    net1166,
    net1165,
    net1164,
    net1163,
    net1162,
    net1161,
    net1159,
    net1158,
    net1157,
    net1156,
    net1155,
    net1154,
    net1153,
    net1152,
    net1151,
    net1150,
    net1148,
    net1147,
    net1146,
    net1145,
    net1144,
    net1143,
    net1142,
    net1141,
    net1140,
    net1139,
    net1137,
    net1136,
    net1135,
    net1134,
    net1133,
    net1132,
    net1131,
    net1130,
    net1129,
    net1128,
    net1126,
    net1125,
    net1124,
    net1123,
    net1122,
    net1121,
    net1120,
    net1119,
    net1118,
    net1117,
    net1179,
    net1178,
    net1177,
    net1176,
    net1171,
    net1160,
    net1149,
    net1138,
    net1127,
    net1116}),
    .io_outs_left({\_ces_0_1_io_outs_left[63] ,
    \_ces_0_1_io_outs_left[62] ,
    \_ces_0_1_io_outs_left[61] ,
    \_ces_0_1_io_outs_left[60] ,
    \_ces_0_1_io_outs_left[59] ,
    \_ces_0_1_io_outs_left[58] ,
    \_ces_0_1_io_outs_left[57] ,
    \_ces_0_1_io_outs_left[56] ,
    \_ces_0_1_io_outs_left[55] ,
    \_ces_0_1_io_outs_left[54] ,
    \_ces_0_1_io_outs_left[53] ,
    \_ces_0_1_io_outs_left[52] ,
    \_ces_0_1_io_outs_left[51] ,
    \_ces_0_1_io_outs_left[50] ,
    \_ces_0_1_io_outs_left[49] ,
    \_ces_0_1_io_outs_left[48] ,
    \_ces_0_1_io_outs_left[47] ,
    \_ces_0_1_io_outs_left[46] ,
    \_ces_0_1_io_outs_left[45] ,
    \_ces_0_1_io_outs_left[44] ,
    \_ces_0_1_io_outs_left[43] ,
    \_ces_0_1_io_outs_left[42] ,
    \_ces_0_1_io_outs_left[41] ,
    \_ces_0_1_io_outs_left[40] ,
    \_ces_0_1_io_outs_left[39] ,
    \_ces_0_1_io_outs_left[38] ,
    \_ces_0_1_io_outs_left[37] ,
    \_ces_0_1_io_outs_left[36] ,
    \_ces_0_1_io_outs_left[35] ,
    \_ces_0_1_io_outs_left[34] ,
    \_ces_0_1_io_outs_left[33] ,
    \_ces_0_1_io_outs_left[32] ,
    \_ces_0_1_io_outs_left[31] ,
    \_ces_0_1_io_outs_left[30] ,
    \_ces_0_1_io_outs_left[29] ,
    \_ces_0_1_io_outs_left[28] ,
    \_ces_0_1_io_outs_left[27] ,
    \_ces_0_1_io_outs_left[26] ,
    \_ces_0_1_io_outs_left[25] ,
    \_ces_0_1_io_outs_left[24] ,
    \_ces_0_1_io_outs_left[23] ,
    \_ces_0_1_io_outs_left[22] ,
    \_ces_0_1_io_outs_left[21] ,
    \_ces_0_1_io_outs_left[20] ,
    \_ces_0_1_io_outs_left[19] ,
    \_ces_0_1_io_outs_left[18] ,
    \_ces_0_1_io_outs_left[17] ,
    \_ces_0_1_io_outs_left[16] ,
    \_ces_0_1_io_outs_left[15] ,
    \_ces_0_1_io_outs_left[14] ,
    \_ces_0_1_io_outs_left[13] ,
    \_ces_0_1_io_outs_left[12] ,
    \_ces_0_1_io_outs_left[11] ,
    \_ces_0_1_io_outs_left[10] ,
    \_ces_0_1_io_outs_left[9] ,
    \_ces_0_1_io_outs_left[8] ,
    \_ces_0_1_io_outs_left[7] ,
    \_ces_0_1_io_outs_left[6] ,
    \_ces_0_1_io_outs_left[5] ,
    \_ces_0_1_io_outs_left[4] ,
    \_ces_0_1_io_outs_left[3] ,
    \_ces_0_1_io_outs_left[2] ,
    \_ces_0_1_io_outs_left[1] ,
    \_ces_0_1_io_outs_left[0] }),
    .io_outs_right({\_ces_0_1_io_outs_right[63] ,
    \_ces_0_1_io_outs_right[62] ,
    \_ces_0_1_io_outs_right[61] ,
    \_ces_0_1_io_outs_right[60] ,
    \_ces_0_1_io_outs_right[59] ,
    \_ces_0_1_io_outs_right[58] ,
    \_ces_0_1_io_outs_right[57] ,
    \_ces_0_1_io_outs_right[56] ,
    \_ces_0_1_io_outs_right[55] ,
    \_ces_0_1_io_outs_right[54] ,
    \_ces_0_1_io_outs_right[53] ,
    \_ces_0_1_io_outs_right[52] ,
    \_ces_0_1_io_outs_right[51] ,
    \_ces_0_1_io_outs_right[50] ,
    \_ces_0_1_io_outs_right[49] ,
    \_ces_0_1_io_outs_right[48] ,
    \_ces_0_1_io_outs_right[47] ,
    \_ces_0_1_io_outs_right[46] ,
    \_ces_0_1_io_outs_right[45] ,
    \_ces_0_1_io_outs_right[44] ,
    \_ces_0_1_io_outs_right[43] ,
    \_ces_0_1_io_outs_right[42] ,
    \_ces_0_1_io_outs_right[41] ,
    \_ces_0_1_io_outs_right[40] ,
    \_ces_0_1_io_outs_right[39] ,
    \_ces_0_1_io_outs_right[38] ,
    \_ces_0_1_io_outs_right[37] ,
    \_ces_0_1_io_outs_right[36] ,
    \_ces_0_1_io_outs_right[35] ,
    \_ces_0_1_io_outs_right[34] ,
    \_ces_0_1_io_outs_right[33] ,
    \_ces_0_1_io_outs_right[32] ,
    \_ces_0_1_io_outs_right[31] ,
    \_ces_0_1_io_outs_right[30] ,
    \_ces_0_1_io_outs_right[29] ,
    \_ces_0_1_io_outs_right[28] ,
    \_ces_0_1_io_outs_right[27] ,
    \_ces_0_1_io_outs_right[26] ,
    \_ces_0_1_io_outs_right[25] ,
    \_ces_0_1_io_outs_right[24] ,
    \_ces_0_1_io_outs_right[23] ,
    \_ces_0_1_io_outs_right[22] ,
    \_ces_0_1_io_outs_right[21] ,
    \_ces_0_1_io_outs_right[20] ,
    \_ces_0_1_io_outs_right[19] ,
    \_ces_0_1_io_outs_right[18] ,
    \_ces_0_1_io_outs_right[17] ,
    \_ces_0_1_io_outs_right[16] ,
    \_ces_0_1_io_outs_right[15] ,
    \_ces_0_1_io_outs_right[14] ,
    \_ces_0_1_io_outs_right[13] ,
    \_ces_0_1_io_outs_right[12] ,
    \_ces_0_1_io_outs_right[11] ,
    \_ces_0_1_io_outs_right[10] ,
    \_ces_0_1_io_outs_right[9] ,
    \_ces_0_1_io_outs_right[8] ,
    \_ces_0_1_io_outs_right[7] ,
    \_ces_0_1_io_outs_right[6] ,
    \_ces_0_1_io_outs_right[5] ,
    \_ces_0_1_io_outs_right[4] ,
    \_ces_0_1_io_outs_right[3] ,
    \_ces_0_1_io_outs_right[2] ,
    \_ces_0_1_io_outs_right[1] ,
    \_ces_0_1_io_outs_right[0] }),
    .io_outs_up({\_ces_0_1_io_outs_up[63] ,
    \_ces_0_1_io_outs_up[62] ,
    \_ces_0_1_io_outs_up[61] ,
    \_ces_0_1_io_outs_up[60] ,
    \_ces_0_1_io_outs_up[59] ,
    \_ces_0_1_io_outs_up[58] ,
    \_ces_0_1_io_outs_up[57] ,
    \_ces_0_1_io_outs_up[56] ,
    \_ces_0_1_io_outs_up[55] ,
    \_ces_0_1_io_outs_up[54] ,
    \_ces_0_1_io_outs_up[53] ,
    \_ces_0_1_io_outs_up[52] ,
    \_ces_0_1_io_outs_up[51] ,
    \_ces_0_1_io_outs_up[50] ,
    \_ces_0_1_io_outs_up[49] ,
    \_ces_0_1_io_outs_up[48] ,
    \_ces_0_1_io_outs_up[47] ,
    \_ces_0_1_io_outs_up[46] ,
    \_ces_0_1_io_outs_up[45] ,
    \_ces_0_1_io_outs_up[44] ,
    \_ces_0_1_io_outs_up[43] ,
    \_ces_0_1_io_outs_up[42] ,
    \_ces_0_1_io_outs_up[41] ,
    \_ces_0_1_io_outs_up[40] ,
    \_ces_0_1_io_outs_up[39] ,
    \_ces_0_1_io_outs_up[38] ,
    \_ces_0_1_io_outs_up[37] ,
    \_ces_0_1_io_outs_up[36] ,
    \_ces_0_1_io_outs_up[35] ,
    \_ces_0_1_io_outs_up[34] ,
    \_ces_0_1_io_outs_up[33] ,
    \_ces_0_1_io_outs_up[32] ,
    \_ces_0_1_io_outs_up[31] ,
    \_ces_0_1_io_outs_up[30] ,
    \_ces_0_1_io_outs_up[29] ,
    \_ces_0_1_io_outs_up[28] ,
    \_ces_0_1_io_outs_up[27] ,
    \_ces_0_1_io_outs_up[26] ,
    \_ces_0_1_io_outs_up[25] ,
    \_ces_0_1_io_outs_up[24] ,
    \_ces_0_1_io_outs_up[23] ,
    \_ces_0_1_io_outs_up[22] ,
    \_ces_0_1_io_outs_up[21] ,
    \_ces_0_1_io_outs_up[20] ,
    \_ces_0_1_io_outs_up[19] ,
    \_ces_0_1_io_outs_up[18] ,
    \_ces_0_1_io_outs_up[17] ,
    \_ces_0_1_io_outs_up[16] ,
    \_ces_0_1_io_outs_up[15] ,
    \_ces_0_1_io_outs_up[14] ,
    \_ces_0_1_io_outs_up[13] ,
    \_ces_0_1_io_outs_up[12] ,
    \_ces_0_1_io_outs_up[11] ,
    \_ces_0_1_io_outs_up[10] ,
    \_ces_0_1_io_outs_up[9] ,
    \_ces_0_1_io_outs_up[8] ,
    \_ces_0_1_io_outs_up[7] ,
    \_ces_0_1_io_outs_up[6] ,
    \_ces_0_1_io_outs_up[5] ,
    \_ces_0_1_io_outs_up[4] ,
    \_ces_0_1_io_outs_up[3] ,
    \_ces_0_1_io_outs_up[2] ,
    \_ces_0_1_io_outs_up[1] ,
    \_ces_0_1_io_outs_up[0] }));
 Element ces_0_2 (.clock(clknet_leaf_2_clock),
    .io_lsbIns_1(_ces_0_1_io_lsbOuts_1),
    .io_lsbIns_2(_ces_0_1_io_lsbOuts_2),
    .io_lsbIns_3(_ces_0_1_io_lsbOuts_3),
    .io_lsbOuts_1(_ces_0_2_io_lsbOuts_1),
    .io_lsbOuts_2(_ces_0_2_io_lsbOuts_2),
    .io_lsbOuts_3(_ces_0_2_io_lsbOuts_3),
    .io_ins_down({\_ces_1_2_io_outs_down[63] ,
    \_ces_1_2_io_outs_down[62] ,
    \_ces_1_2_io_outs_down[61] ,
    \_ces_1_2_io_outs_down[60] ,
    \_ces_1_2_io_outs_down[59] ,
    \_ces_1_2_io_outs_down[58] ,
    \_ces_1_2_io_outs_down[57] ,
    \_ces_1_2_io_outs_down[56] ,
    \_ces_1_2_io_outs_down[55] ,
    \_ces_1_2_io_outs_down[54] ,
    \_ces_1_2_io_outs_down[53] ,
    \_ces_1_2_io_outs_down[52] ,
    \_ces_1_2_io_outs_down[51] ,
    \_ces_1_2_io_outs_down[50] ,
    \_ces_1_2_io_outs_down[49] ,
    \_ces_1_2_io_outs_down[48] ,
    \_ces_1_2_io_outs_down[47] ,
    \_ces_1_2_io_outs_down[46] ,
    \_ces_1_2_io_outs_down[45] ,
    \_ces_1_2_io_outs_down[44] ,
    \_ces_1_2_io_outs_down[43] ,
    \_ces_1_2_io_outs_down[42] ,
    \_ces_1_2_io_outs_down[41] ,
    \_ces_1_2_io_outs_down[40] ,
    \_ces_1_2_io_outs_down[39] ,
    \_ces_1_2_io_outs_down[38] ,
    \_ces_1_2_io_outs_down[37] ,
    \_ces_1_2_io_outs_down[36] ,
    \_ces_1_2_io_outs_down[35] ,
    \_ces_1_2_io_outs_down[34] ,
    \_ces_1_2_io_outs_down[33] ,
    \_ces_1_2_io_outs_down[32] ,
    \_ces_1_2_io_outs_down[31] ,
    \_ces_1_2_io_outs_down[30] ,
    \_ces_1_2_io_outs_down[29] ,
    \_ces_1_2_io_outs_down[28] ,
    \_ces_1_2_io_outs_down[27] ,
    \_ces_1_2_io_outs_down[26] ,
    \_ces_1_2_io_outs_down[25] ,
    \_ces_1_2_io_outs_down[24] ,
    \_ces_1_2_io_outs_down[23] ,
    \_ces_1_2_io_outs_down[22] ,
    \_ces_1_2_io_outs_down[21] ,
    \_ces_1_2_io_outs_down[20] ,
    \_ces_1_2_io_outs_down[19] ,
    \_ces_1_2_io_outs_down[18] ,
    \_ces_1_2_io_outs_down[17] ,
    \_ces_1_2_io_outs_down[16] ,
    \_ces_1_2_io_outs_down[15] ,
    \_ces_1_2_io_outs_down[14] ,
    \_ces_1_2_io_outs_down[13] ,
    \_ces_1_2_io_outs_down[12] ,
    \_ces_1_2_io_outs_down[11] ,
    \_ces_1_2_io_outs_down[10] ,
    \_ces_1_2_io_outs_down[9] ,
    \_ces_1_2_io_outs_down[8] ,
    \_ces_1_2_io_outs_down[7] ,
    \_ces_1_2_io_outs_down[6] ,
    \_ces_1_2_io_outs_down[5] ,
    \_ces_1_2_io_outs_down[4] ,
    \_ces_1_2_io_outs_down[3] ,
    \_ces_1_2_io_outs_down[2] ,
    \_ces_1_2_io_outs_down[1] ,
    \_ces_1_2_io_outs_down[0] }),
    .io_ins_left({\_ces_0_3_io_outs_left[63] ,
    \_ces_0_3_io_outs_left[62] ,
    \_ces_0_3_io_outs_left[61] ,
    \_ces_0_3_io_outs_left[60] ,
    \_ces_0_3_io_outs_left[59] ,
    \_ces_0_3_io_outs_left[58] ,
    \_ces_0_3_io_outs_left[57] ,
    \_ces_0_3_io_outs_left[56] ,
    \_ces_0_3_io_outs_left[55] ,
    \_ces_0_3_io_outs_left[54] ,
    \_ces_0_3_io_outs_left[53] ,
    \_ces_0_3_io_outs_left[52] ,
    \_ces_0_3_io_outs_left[51] ,
    \_ces_0_3_io_outs_left[50] ,
    \_ces_0_3_io_outs_left[49] ,
    \_ces_0_3_io_outs_left[48] ,
    \_ces_0_3_io_outs_left[47] ,
    \_ces_0_3_io_outs_left[46] ,
    \_ces_0_3_io_outs_left[45] ,
    \_ces_0_3_io_outs_left[44] ,
    \_ces_0_3_io_outs_left[43] ,
    \_ces_0_3_io_outs_left[42] ,
    \_ces_0_3_io_outs_left[41] ,
    \_ces_0_3_io_outs_left[40] ,
    \_ces_0_3_io_outs_left[39] ,
    \_ces_0_3_io_outs_left[38] ,
    \_ces_0_3_io_outs_left[37] ,
    \_ces_0_3_io_outs_left[36] ,
    \_ces_0_3_io_outs_left[35] ,
    \_ces_0_3_io_outs_left[34] ,
    \_ces_0_3_io_outs_left[33] ,
    \_ces_0_3_io_outs_left[32] ,
    \_ces_0_3_io_outs_left[31] ,
    \_ces_0_3_io_outs_left[30] ,
    \_ces_0_3_io_outs_left[29] ,
    \_ces_0_3_io_outs_left[28] ,
    \_ces_0_3_io_outs_left[27] ,
    \_ces_0_3_io_outs_left[26] ,
    \_ces_0_3_io_outs_left[25] ,
    \_ces_0_3_io_outs_left[24] ,
    \_ces_0_3_io_outs_left[23] ,
    \_ces_0_3_io_outs_left[22] ,
    \_ces_0_3_io_outs_left[21] ,
    \_ces_0_3_io_outs_left[20] ,
    \_ces_0_3_io_outs_left[19] ,
    \_ces_0_3_io_outs_left[18] ,
    \_ces_0_3_io_outs_left[17] ,
    \_ces_0_3_io_outs_left[16] ,
    \_ces_0_3_io_outs_left[15] ,
    \_ces_0_3_io_outs_left[14] ,
    \_ces_0_3_io_outs_left[13] ,
    \_ces_0_3_io_outs_left[12] ,
    \_ces_0_3_io_outs_left[11] ,
    \_ces_0_3_io_outs_left[10] ,
    \_ces_0_3_io_outs_left[9] ,
    \_ces_0_3_io_outs_left[8] ,
    \_ces_0_3_io_outs_left[7] ,
    \_ces_0_3_io_outs_left[6] ,
    \_ces_0_3_io_outs_left[5] ,
    \_ces_0_3_io_outs_left[4] ,
    \_ces_0_3_io_outs_left[3] ,
    \_ces_0_3_io_outs_left[2] ,
    \_ces_0_3_io_outs_left[1] ,
    \_ces_0_3_io_outs_left[0] }),
    .io_ins_right({\_ces_0_1_io_outs_right[63] ,
    \_ces_0_1_io_outs_right[62] ,
    \_ces_0_1_io_outs_right[61] ,
    \_ces_0_1_io_outs_right[60] ,
    \_ces_0_1_io_outs_right[59] ,
    \_ces_0_1_io_outs_right[58] ,
    \_ces_0_1_io_outs_right[57] ,
    \_ces_0_1_io_outs_right[56] ,
    \_ces_0_1_io_outs_right[55] ,
    \_ces_0_1_io_outs_right[54] ,
    \_ces_0_1_io_outs_right[53] ,
    \_ces_0_1_io_outs_right[52] ,
    \_ces_0_1_io_outs_right[51] ,
    \_ces_0_1_io_outs_right[50] ,
    \_ces_0_1_io_outs_right[49] ,
    \_ces_0_1_io_outs_right[48] ,
    \_ces_0_1_io_outs_right[47] ,
    \_ces_0_1_io_outs_right[46] ,
    \_ces_0_1_io_outs_right[45] ,
    \_ces_0_1_io_outs_right[44] ,
    \_ces_0_1_io_outs_right[43] ,
    \_ces_0_1_io_outs_right[42] ,
    \_ces_0_1_io_outs_right[41] ,
    \_ces_0_1_io_outs_right[40] ,
    \_ces_0_1_io_outs_right[39] ,
    \_ces_0_1_io_outs_right[38] ,
    \_ces_0_1_io_outs_right[37] ,
    \_ces_0_1_io_outs_right[36] ,
    \_ces_0_1_io_outs_right[35] ,
    \_ces_0_1_io_outs_right[34] ,
    \_ces_0_1_io_outs_right[33] ,
    \_ces_0_1_io_outs_right[32] ,
    \_ces_0_1_io_outs_right[31] ,
    \_ces_0_1_io_outs_right[30] ,
    \_ces_0_1_io_outs_right[29] ,
    \_ces_0_1_io_outs_right[28] ,
    \_ces_0_1_io_outs_right[27] ,
    \_ces_0_1_io_outs_right[26] ,
    \_ces_0_1_io_outs_right[25] ,
    \_ces_0_1_io_outs_right[24] ,
    \_ces_0_1_io_outs_right[23] ,
    \_ces_0_1_io_outs_right[22] ,
    \_ces_0_1_io_outs_right[21] ,
    \_ces_0_1_io_outs_right[20] ,
    \_ces_0_1_io_outs_right[19] ,
    \_ces_0_1_io_outs_right[18] ,
    \_ces_0_1_io_outs_right[17] ,
    \_ces_0_1_io_outs_right[16] ,
    \_ces_0_1_io_outs_right[15] ,
    \_ces_0_1_io_outs_right[14] ,
    \_ces_0_1_io_outs_right[13] ,
    \_ces_0_1_io_outs_right[12] ,
    \_ces_0_1_io_outs_right[11] ,
    \_ces_0_1_io_outs_right[10] ,
    \_ces_0_1_io_outs_right[9] ,
    \_ces_0_1_io_outs_right[8] ,
    \_ces_0_1_io_outs_right[7] ,
    \_ces_0_1_io_outs_right[6] ,
    \_ces_0_1_io_outs_right[5] ,
    \_ces_0_1_io_outs_right[4] ,
    \_ces_0_1_io_outs_right[3] ,
    \_ces_0_1_io_outs_right[2] ,
    \_ces_0_1_io_outs_right[1] ,
    \_ces_0_1_io_outs_right[0] }),
    .io_ins_up({net967,
    net966,
    net965,
    net964,
    net962,
    net961,
    net960,
    net959,
    net958,
    net957,
    net956,
    net955,
    net954,
    net953,
    net951,
    net950,
    net949,
    net948,
    net947,
    net946,
    net945,
    net944,
    net943,
    net942,
    net940,
    net939,
    net938,
    net937,
    net936,
    net935,
    net934,
    net933,
    net932,
    net931,
    net929,
    net928,
    net927,
    net926,
    net925,
    net924,
    net923,
    net922,
    net921,
    net920,
    net918,
    net917,
    net916,
    net915,
    net914,
    net913,
    net912,
    net911,
    net910,
    net909,
    net971,
    net970,
    net969,
    net968,
    net963,
    net952,
    net941,
    net930,
    net919,
    net908}),
    .io_outs_down({net1239,
    net1238,
    net1237,
    net1236,
    net1234,
    net1233,
    net1232,
    net1231,
    net1230,
    net1229,
    net1228,
    net1227,
    net1226,
    net1225,
    net1223,
    net1222,
    net1221,
    net1220,
    net1219,
    net1218,
    net1217,
    net1216,
    net1215,
    net1214,
    net1212,
    net1211,
    net1210,
    net1209,
    net1208,
    net1207,
    net1206,
    net1205,
    net1204,
    net1203,
    net1201,
    net1200,
    net1199,
    net1198,
    net1197,
    net1196,
    net1195,
    net1194,
    net1193,
    net1192,
    net1190,
    net1189,
    net1188,
    net1187,
    net1186,
    net1185,
    net1184,
    net1183,
    net1182,
    net1181,
    net1243,
    net1242,
    net1241,
    net1240,
    net1235,
    net1224,
    net1213,
    net1202,
    net1191,
    net1180}),
    .io_outs_left({\_ces_0_2_io_outs_left[63] ,
    \_ces_0_2_io_outs_left[62] ,
    \_ces_0_2_io_outs_left[61] ,
    \_ces_0_2_io_outs_left[60] ,
    \_ces_0_2_io_outs_left[59] ,
    \_ces_0_2_io_outs_left[58] ,
    \_ces_0_2_io_outs_left[57] ,
    \_ces_0_2_io_outs_left[56] ,
    \_ces_0_2_io_outs_left[55] ,
    \_ces_0_2_io_outs_left[54] ,
    \_ces_0_2_io_outs_left[53] ,
    \_ces_0_2_io_outs_left[52] ,
    \_ces_0_2_io_outs_left[51] ,
    \_ces_0_2_io_outs_left[50] ,
    \_ces_0_2_io_outs_left[49] ,
    \_ces_0_2_io_outs_left[48] ,
    \_ces_0_2_io_outs_left[47] ,
    \_ces_0_2_io_outs_left[46] ,
    \_ces_0_2_io_outs_left[45] ,
    \_ces_0_2_io_outs_left[44] ,
    \_ces_0_2_io_outs_left[43] ,
    \_ces_0_2_io_outs_left[42] ,
    \_ces_0_2_io_outs_left[41] ,
    \_ces_0_2_io_outs_left[40] ,
    \_ces_0_2_io_outs_left[39] ,
    \_ces_0_2_io_outs_left[38] ,
    \_ces_0_2_io_outs_left[37] ,
    \_ces_0_2_io_outs_left[36] ,
    \_ces_0_2_io_outs_left[35] ,
    \_ces_0_2_io_outs_left[34] ,
    \_ces_0_2_io_outs_left[33] ,
    \_ces_0_2_io_outs_left[32] ,
    \_ces_0_2_io_outs_left[31] ,
    \_ces_0_2_io_outs_left[30] ,
    \_ces_0_2_io_outs_left[29] ,
    \_ces_0_2_io_outs_left[28] ,
    \_ces_0_2_io_outs_left[27] ,
    \_ces_0_2_io_outs_left[26] ,
    \_ces_0_2_io_outs_left[25] ,
    \_ces_0_2_io_outs_left[24] ,
    \_ces_0_2_io_outs_left[23] ,
    \_ces_0_2_io_outs_left[22] ,
    \_ces_0_2_io_outs_left[21] ,
    \_ces_0_2_io_outs_left[20] ,
    \_ces_0_2_io_outs_left[19] ,
    \_ces_0_2_io_outs_left[18] ,
    \_ces_0_2_io_outs_left[17] ,
    \_ces_0_2_io_outs_left[16] ,
    \_ces_0_2_io_outs_left[15] ,
    \_ces_0_2_io_outs_left[14] ,
    \_ces_0_2_io_outs_left[13] ,
    \_ces_0_2_io_outs_left[12] ,
    \_ces_0_2_io_outs_left[11] ,
    \_ces_0_2_io_outs_left[10] ,
    \_ces_0_2_io_outs_left[9] ,
    \_ces_0_2_io_outs_left[8] ,
    \_ces_0_2_io_outs_left[7] ,
    \_ces_0_2_io_outs_left[6] ,
    \_ces_0_2_io_outs_left[5] ,
    \_ces_0_2_io_outs_left[4] ,
    \_ces_0_2_io_outs_left[3] ,
    \_ces_0_2_io_outs_left[2] ,
    \_ces_0_2_io_outs_left[1] ,
    \_ces_0_2_io_outs_left[0] }),
    .io_outs_right({\_ces_0_2_io_outs_right[63] ,
    \_ces_0_2_io_outs_right[62] ,
    \_ces_0_2_io_outs_right[61] ,
    \_ces_0_2_io_outs_right[60] ,
    \_ces_0_2_io_outs_right[59] ,
    \_ces_0_2_io_outs_right[58] ,
    \_ces_0_2_io_outs_right[57] ,
    \_ces_0_2_io_outs_right[56] ,
    \_ces_0_2_io_outs_right[55] ,
    \_ces_0_2_io_outs_right[54] ,
    \_ces_0_2_io_outs_right[53] ,
    \_ces_0_2_io_outs_right[52] ,
    \_ces_0_2_io_outs_right[51] ,
    \_ces_0_2_io_outs_right[50] ,
    \_ces_0_2_io_outs_right[49] ,
    \_ces_0_2_io_outs_right[48] ,
    \_ces_0_2_io_outs_right[47] ,
    \_ces_0_2_io_outs_right[46] ,
    \_ces_0_2_io_outs_right[45] ,
    \_ces_0_2_io_outs_right[44] ,
    \_ces_0_2_io_outs_right[43] ,
    \_ces_0_2_io_outs_right[42] ,
    \_ces_0_2_io_outs_right[41] ,
    \_ces_0_2_io_outs_right[40] ,
    \_ces_0_2_io_outs_right[39] ,
    \_ces_0_2_io_outs_right[38] ,
    \_ces_0_2_io_outs_right[37] ,
    \_ces_0_2_io_outs_right[36] ,
    \_ces_0_2_io_outs_right[35] ,
    \_ces_0_2_io_outs_right[34] ,
    \_ces_0_2_io_outs_right[33] ,
    \_ces_0_2_io_outs_right[32] ,
    \_ces_0_2_io_outs_right[31] ,
    \_ces_0_2_io_outs_right[30] ,
    \_ces_0_2_io_outs_right[29] ,
    \_ces_0_2_io_outs_right[28] ,
    \_ces_0_2_io_outs_right[27] ,
    \_ces_0_2_io_outs_right[26] ,
    \_ces_0_2_io_outs_right[25] ,
    \_ces_0_2_io_outs_right[24] ,
    \_ces_0_2_io_outs_right[23] ,
    \_ces_0_2_io_outs_right[22] ,
    \_ces_0_2_io_outs_right[21] ,
    \_ces_0_2_io_outs_right[20] ,
    \_ces_0_2_io_outs_right[19] ,
    \_ces_0_2_io_outs_right[18] ,
    \_ces_0_2_io_outs_right[17] ,
    \_ces_0_2_io_outs_right[16] ,
    \_ces_0_2_io_outs_right[15] ,
    \_ces_0_2_io_outs_right[14] ,
    \_ces_0_2_io_outs_right[13] ,
    \_ces_0_2_io_outs_right[12] ,
    \_ces_0_2_io_outs_right[11] ,
    \_ces_0_2_io_outs_right[10] ,
    \_ces_0_2_io_outs_right[9] ,
    \_ces_0_2_io_outs_right[8] ,
    \_ces_0_2_io_outs_right[7] ,
    \_ces_0_2_io_outs_right[6] ,
    \_ces_0_2_io_outs_right[5] ,
    \_ces_0_2_io_outs_right[4] ,
    \_ces_0_2_io_outs_right[3] ,
    \_ces_0_2_io_outs_right[2] ,
    \_ces_0_2_io_outs_right[1] ,
    \_ces_0_2_io_outs_right[0] }),
    .io_outs_up({\_ces_0_2_io_outs_up[63] ,
    \_ces_0_2_io_outs_up[62] ,
    \_ces_0_2_io_outs_up[61] ,
    \_ces_0_2_io_outs_up[60] ,
    \_ces_0_2_io_outs_up[59] ,
    \_ces_0_2_io_outs_up[58] ,
    \_ces_0_2_io_outs_up[57] ,
    \_ces_0_2_io_outs_up[56] ,
    \_ces_0_2_io_outs_up[55] ,
    \_ces_0_2_io_outs_up[54] ,
    \_ces_0_2_io_outs_up[53] ,
    \_ces_0_2_io_outs_up[52] ,
    \_ces_0_2_io_outs_up[51] ,
    \_ces_0_2_io_outs_up[50] ,
    \_ces_0_2_io_outs_up[49] ,
    \_ces_0_2_io_outs_up[48] ,
    \_ces_0_2_io_outs_up[47] ,
    \_ces_0_2_io_outs_up[46] ,
    \_ces_0_2_io_outs_up[45] ,
    \_ces_0_2_io_outs_up[44] ,
    \_ces_0_2_io_outs_up[43] ,
    \_ces_0_2_io_outs_up[42] ,
    \_ces_0_2_io_outs_up[41] ,
    \_ces_0_2_io_outs_up[40] ,
    \_ces_0_2_io_outs_up[39] ,
    \_ces_0_2_io_outs_up[38] ,
    \_ces_0_2_io_outs_up[37] ,
    \_ces_0_2_io_outs_up[36] ,
    \_ces_0_2_io_outs_up[35] ,
    \_ces_0_2_io_outs_up[34] ,
    \_ces_0_2_io_outs_up[33] ,
    \_ces_0_2_io_outs_up[32] ,
    \_ces_0_2_io_outs_up[31] ,
    \_ces_0_2_io_outs_up[30] ,
    \_ces_0_2_io_outs_up[29] ,
    \_ces_0_2_io_outs_up[28] ,
    \_ces_0_2_io_outs_up[27] ,
    \_ces_0_2_io_outs_up[26] ,
    \_ces_0_2_io_outs_up[25] ,
    \_ces_0_2_io_outs_up[24] ,
    \_ces_0_2_io_outs_up[23] ,
    \_ces_0_2_io_outs_up[22] ,
    \_ces_0_2_io_outs_up[21] ,
    \_ces_0_2_io_outs_up[20] ,
    \_ces_0_2_io_outs_up[19] ,
    \_ces_0_2_io_outs_up[18] ,
    \_ces_0_2_io_outs_up[17] ,
    \_ces_0_2_io_outs_up[16] ,
    \_ces_0_2_io_outs_up[15] ,
    \_ces_0_2_io_outs_up[14] ,
    \_ces_0_2_io_outs_up[13] ,
    \_ces_0_2_io_outs_up[12] ,
    \_ces_0_2_io_outs_up[11] ,
    \_ces_0_2_io_outs_up[10] ,
    \_ces_0_2_io_outs_up[9] ,
    \_ces_0_2_io_outs_up[8] ,
    \_ces_0_2_io_outs_up[7] ,
    \_ces_0_2_io_outs_up[6] ,
    \_ces_0_2_io_outs_up[5] ,
    \_ces_0_2_io_outs_up[4] ,
    \_ces_0_2_io_outs_up[3] ,
    \_ces_0_2_io_outs_up[2] ,
    \_ces_0_2_io_outs_up[1] ,
    \_ces_0_2_io_outs_up[0] }));
 Element ces_0_3 (.clock(clknet_leaf_2_clock),
    .io_lsbIns_1(_ces_0_2_io_lsbOuts_1),
    .io_lsbIns_2(_ces_0_2_io_lsbOuts_2),
    .io_lsbIns_3(_ces_0_2_io_lsbOuts_3),
    .io_lsbOuts_0(_ces_0_3_io_lsbOuts_0),
    .io_lsbOuts_1(_ces_0_3_io_lsbOuts_1),
    .io_lsbOuts_2(_ces_0_3_io_lsbOuts_2),
    .io_lsbOuts_3(_ces_0_3_io_lsbOuts_3),
    .io_ins_down({\_ces_1_3_io_outs_down[63] ,
    \_ces_1_3_io_outs_down[62] ,
    \_ces_1_3_io_outs_down[61] ,
    \_ces_1_3_io_outs_down[60] ,
    \_ces_1_3_io_outs_down[59] ,
    \_ces_1_3_io_outs_down[58] ,
    \_ces_1_3_io_outs_down[57] ,
    \_ces_1_3_io_outs_down[56] ,
    \_ces_1_3_io_outs_down[55] ,
    \_ces_1_3_io_outs_down[54] ,
    \_ces_1_3_io_outs_down[53] ,
    \_ces_1_3_io_outs_down[52] ,
    \_ces_1_3_io_outs_down[51] ,
    \_ces_1_3_io_outs_down[50] ,
    \_ces_1_3_io_outs_down[49] ,
    \_ces_1_3_io_outs_down[48] ,
    \_ces_1_3_io_outs_down[47] ,
    \_ces_1_3_io_outs_down[46] ,
    \_ces_1_3_io_outs_down[45] ,
    \_ces_1_3_io_outs_down[44] ,
    \_ces_1_3_io_outs_down[43] ,
    \_ces_1_3_io_outs_down[42] ,
    \_ces_1_3_io_outs_down[41] ,
    \_ces_1_3_io_outs_down[40] ,
    \_ces_1_3_io_outs_down[39] ,
    \_ces_1_3_io_outs_down[38] ,
    \_ces_1_3_io_outs_down[37] ,
    \_ces_1_3_io_outs_down[36] ,
    \_ces_1_3_io_outs_down[35] ,
    \_ces_1_3_io_outs_down[34] ,
    \_ces_1_3_io_outs_down[33] ,
    \_ces_1_3_io_outs_down[32] ,
    \_ces_1_3_io_outs_down[31] ,
    \_ces_1_3_io_outs_down[30] ,
    \_ces_1_3_io_outs_down[29] ,
    \_ces_1_3_io_outs_down[28] ,
    \_ces_1_3_io_outs_down[27] ,
    \_ces_1_3_io_outs_down[26] ,
    \_ces_1_3_io_outs_down[25] ,
    \_ces_1_3_io_outs_down[24] ,
    \_ces_1_3_io_outs_down[23] ,
    \_ces_1_3_io_outs_down[22] ,
    \_ces_1_3_io_outs_down[21] ,
    \_ces_1_3_io_outs_down[20] ,
    \_ces_1_3_io_outs_down[19] ,
    \_ces_1_3_io_outs_down[18] ,
    \_ces_1_3_io_outs_down[17] ,
    \_ces_1_3_io_outs_down[16] ,
    \_ces_1_3_io_outs_down[15] ,
    \_ces_1_3_io_outs_down[14] ,
    \_ces_1_3_io_outs_down[13] ,
    \_ces_1_3_io_outs_down[12] ,
    \_ces_1_3_io_outs_down[11] ,
    \_ces_1_3_io_outs_down[10] ,
    \_ces_1_3_io_outs_down[9] ,
    \_ces_1_3_io_outs_down[8] ,
    \_ces_1_3_io_outs_down[7] ,
    \_ces_1_3_io_outs_down[6] ,
    \_ces_1_3_io_outs_down[5] ,
    \_ces_1_3_io_outs_down[4] ,
    \_ces_1_3_io_outs_down[3] ,
    \_ces_1_3_io_outs_down[2] ,
    \_ces_1_3_io_outs_down[1] ,
    \_ces_1_3_io_outs_down[0] }),
    .io_ins_left({net327,
    net326,
    net325,
    net324,
    net322,
    net321,
    net320,
    net319,
    net318,
    net317,
    net316,
    net315,
    net314,
    net313,
    net311,
    net310,
    net309,
    net308,
    net307,
    net306,
    net305,
    net304,
    net303,
    net302,
    net300,
    net299,
    net298,
    net297,
    net296,
    net295,
    net294,
    net293,
    net292,
    net291,
    net289,
    net288,
    net287,
    net286,
    net285,
    net284,
    net283,
    net282,
    net281,
    net280,
    net278,
    net277,
    net276,
    net275,
    net274,
    net273,
    net272,
    net271,
    net270,
    net269,
    net331,
    net330,
    net329,
    net328,
    net323,
    net312,
    net301,
    net290,
    net279,
    net268}),
    .io_ins_right({\_ces_0_2_io_outs_right[63] ,
    \_ces_0_2_io_outs_right[62] ,
    \_ces_0_2_io_outs_right[61] ,
    \_ces_0_2_io_outs_right[60] ,
    \_ces_0_2_io_outs_right[59] ,
    \_ces_0_2_io_outs_right[58] ,
    \_ces_0_2_io_outs_right[57] ,
    \_ces_0_2_io_outs_right[56] ,
    \_ces_0_2_io_outs_right[55] ,
    \_ces_0_2_io_outs_right[54] ,
    \_ces_0_2_io_outs_right[53] ,
    \_ces_0_2_io_outs_right[52] ,
    \_ces_0_2_io_outs_right[51] ,
    \_ces_0_2_io_outs_right[50] ,
    \_ces_0_2_io_outs_right[49] ,
    \_ces_0_2_io_outs_right[48] ,
    \_ces_0_2_io_outs_right[47] ,
    \_ces_0_2_io_outs_right[46] ,
    \_ces_0_2_io_outs_right[45] ,
    \_ces_0_2_io_outs_right[44] ,
    \_ces_0_2_io_outs_right[43] ,
    \_ces_0_2_io_outs_right[42] ,
    \_ces_0_2_io_outs_right[41] ,
    \_ces_0_2_io_outs_right[40] ,
    \_ces_0_2_io_outs_right[39] ,
    \_ces_0_2_io_outs_right[38] ,
    \_ces_0_2_io_outs_right[37] ,
    \_ces_0_2_io_outs_right[36] ,
    \_ces_0_2_io_outs_right[35] ,
    \_ces_0_2_io_outs_right[34] ,
    \_ces_0_2_io_outs_right[33] ,
    \_ces_0_2_io_outs_right[32] ,
    \_ces_0_2_io_outs_right[31] ,
    \_ces_0_2_io_outs_right[30] ,
    \_ces_0_2_io_outs_right[29] ,
    \_ces_0_2_io_outs_right[28] ,
    \_ces_0_2_io_outs_right[27] ,
    \_ces_0_2_io_outs_right[26] ,
    \_ces_0_2_io_outs_right[25] ,
    \_ces_0_2_io_outs_right[24] ,
    \_ces_0_2_io_outs_right[23] ,
    \_ces_0_2_io_outs_right[22] ,
    \_ces_0_2_io_outs_right[21] ,
    \_ces_0_2_io_outs_right[20] ,
    \_ces_0_2_io_outs_right[19] ,
    \_ces_0_2_io_outs_right[18] ,
    \_ces_0_2_io_outs_right[17] ,
    \_ces_0_2_io_outs_right[16] ,
    \_ces_0_2_io_outs_right[15] ,
    \_ces_0_2_io_outs_right[14] ,
    \_ces_0_2_io_outs_right[13] ,
    \_ces_0_2_io_outs_right[12] ,
    \_ces_0_2_io_outs_right[11] ,
    \_ces_0_2_io_outs_right[10] ,
    \_ces_0_2_io_outs_right[9] ,
    \_ces_0_2_io_outs_right[8] ,
    \_ces_0_2_io_outs_right[7] ,
    \_ces_0_2_io_outs_right[6] ,
    \_ces_0_2_io_outs_right[5] ,
    \_ces_0_2_io_outs_right[4] ,
    \_ces_0_2_io_outs_right[3] ,
    \_ces_0_2_io_outs_right[2] ,
    \_ces_0_2_io_outs_right[1] ,
    \_ces_0_2_io_outs_right[0] }),
    .io_ins_up({net1031,
    net1030,
    net1029,
    net1028,
    net1026,
    net1025,
    net1024,
    net1023,
    net1022,
    net1021,
    net1020,
    net1019,
    net1018,
    net1017,
    net1015,
    net1014,
    net1013,
    net1012,
    net1011,
    net1010,
    net1009,
    net1008,
    net1007,
    net1006,
    net1004,
    net1003,
    net1002,
    net1001,
    net1000,
    net999,
    net998,
    net997,
    net996,
    net995,
    net993,
    net992,
    net991,
    net990,
    net989,
    net988,
    net987,
    net986,
    net985,
    net984,
    net982,
    net981,
    net980,
    net979,
    net978,
    net977,
    net976,
    net975,
    net974,
    net973,
    net1035,
    net1034,
    net1033,
    net1032,
    net1027,
    net1016,
    net1005,
    net994,
    net983,
    net972}),
    .io_outs_down({net1303,
    net1302,
    net1301,
    net1300,
    net1298,
    net1297,
    net1296,
    net1295,
    net1294,
    net1293,
    net1292,
    net1291,
    net1290,
    net1289,
    net1287,
    net1286,
    net1285,
    net1284,
    net1283,
    net1282,
    net1281,
    net1280,
    net1279,
    net1278,
    net1276,
    net1275,
    net1274,
    net1273,
    net1272,
    net1271,
    net1270,
    net1269,
    net1268,
    net1267,
    net1265,
    net1264,
    net1263,
    net1262,
    net1261,
    net1260,
    net1259,
    net1258,
    net1257,
    net1256,
    net1254,
    net1253,
    net1252,
    net1251,
    net1250,
    net1249,
    net1248,
    net1247,
    net1246,
    net1245,
    net1307,
    net1306,
    net1305,
    net1304,
    net1299,
    net1288,
    net1277,
    net1266,
    net1255,
    net1244}),
    .io_outs_left({\_ces_0_3_io_outs_left[63] ,
    \_ces_0_3_io_outs_left[62] ,
    \_ces_0_3_io_outs_left[61] ,
    \_ces_0_3_io_outs_left[60] ,
    \_ces_0_3_io_outs_left[59] ,
    \_ces_0_3_io_outs_left[58] ,
    \_ces_0_3_io_outs_left[57] ,
    \_ces_0_3_io_outs_left[56] ,
    \_ces_0_3_io_outs_left[55] ,
    \_ces_0_3_io_outs_left[54] ,
    \_ces_0_3_io_outs_left[53] ,
    \_ces_0_3_io_outs_left[52] ,
    \_ces_0_3_io_outs_left[51] ,
    \_ces_0_3_io_outs_left[50] ,
    \_ces_0_3_io_outs_left[49] ,
    \_ces_0_3_io_outs_left[48] ,
    \_ces_0_3_io_outs_left[47] ,
    \_ces_0_3_io_outs_left[46] ,
    \_ces_0_3_io_outs_left[45] ,
    \_ces_0_3_io_outs_left[44] ,
    \_ces_0_3_io_outs_left[43] ,
    \_ces_0_3_io_outs_left[42] ,
    \_ces_0_3_io_outs_left[41] ,
    \_ces_0_3_io_outs_left[40] ,
    \_ces_0_3_io_outs_left[39] ,
    \_ces_0_3_io_outs_left[38] ,
    \_ces_0_3_io_outs_left[37] ,
    \_ces_0_3_io_outs_left[36] ,
    \_ces_0_3_io_outs_left[35] ,
    \_ces_0_3_io_outs_left[34] ,
    \_ces_0_3_io_outs_left[33] ,
    \_ces_0_3_io_outs_left[32] ,
    \_ces_0_3_io_outs_left[31] ,
    \_ces_0_3_io_outs_left[30] ,
    \_ces_0_3_io_outs_left[29] ,
    \_ces_0_3_io_outs_left[28] ,
    \_ces_0_3_io_outs_left[27] ,
    \_ces_0_3_io_outs_left[26] ,
    \_ces_0_3_io_outs_left[25] ,
    \_ces_0_3_io_outs_left[24] ,
    \_ces_0_3_io_outs_left[23] ,
    \_ces_0_3_io_outs_left[22] ,
    \_ces_0_3_io_outs_left[21] ,
    \_ces_0_3_io_outs_left[20] ,
    \_ces_0_3_io_outs_left[19] ,
    \_ces_0_3_io_outs_left[18] ,
    \_ces_0_3_io_outs_left[17] ,
    \_ces_0_3_io_outs_left[16] ,
    \_ces_0_3_io_outs_left[15] ,
    \_ces_0_3_io_outs_left[14] ,
    \_ces_0_3_io_outs_left[13] ,
    \_ces_0_3_io_outs_left[12] ,
    \_ces_0_3_io_outs_left[11] ,
    \_ces_0_3_io_outs_left[10] ,
    \_ces_0_3_io_outs_left[9] ,
    \_ces_0_3_io_outs_left[8] ,
    \_ces_0_3_io_outs_left[7] ,
    \_ces_0_3_io_outs_left[6] ,
    \_ces_0_3_io_outs_left[5] ,
    \_ces_0_3_io_outs_left[4] ,
    \_ces_0_3_io_outs_left[3] ,
    \_ces_0_3_io_outs_left[2] ,
    \_ces_0_3_io_outs_left[1] ,
    \_ces_0_3_io_outs_left[0] }),
    .io_outs_right({net1623,
    net1622,
    net1621,
    net1620,
    net1618,
    net1617,
    net1616,
    net1615,
    net1614,
    net1613,
    net1612,
    net1611,
    net1610,
    net1609,
    net1607,
    net1606,
    net1605,
    net1604,
    net1603,
    net1602,
    net1601,
    net1600,
    net1599,
    net1598,
    net1596,
    net1595,
    net1594,
    net1593,
    net1592,
    net1591,
    net1590,
    net1589,
    net1588,
    net1587,
    net1585,
    net1584,
    net1583,
    net1582,
    net1581,
    net1580,
    net1579,
    net1578,
    net1577,
    net1576,
    net1574,
    net1573,
    net1572,
    net1571,
    net1570,
    net1569,
    net1568,
    net1567,
    net1566,
    net1565,
    net1627,
    net1626,
    net1625,
    net1624,
    net1619,
    net1608,
    net1597,
    net1586,
    net1575,
    net1564}),
    .io_outs_up({\_ces_0_3_io_outs_up[63] ,
    \_ces_0_3_io_outs_up[62] ,
    \_ces_0_3_io_outs_up[61] ,
    \_ces_0_3_io_outs_up[60] ,
    \_ces_0_3_io_outs_up[59] ,
    \_ces_0_3_io_outs_up[58] ,
    \_ces_0_3_io_outs_up[57] ,
    \_ces_0_3_io_outs_up[56] ,
    \_ces_0_3_io_outs_up[55] ,
    \_ces_0_3_io_outs_up[54] ,
    \_ces_0_3_io_outs_up[53] ,
    \_ces_0_3_io_outs_up[52] ,
    \_ces_0_3_io_outs_up[51] ,
    \_ces_0_3_io_outs_up[50] ,
    \_ces_0_3_io_outs_up[49] ,
    \_ces_0_3_io_outs_up[48] ,
    \_ces_0_3_io_outs_up[47] ,
    \_ces_0_3_io_outs_up[46] ,
    \_ces_0_3_io_outs_up[45] ,
    \_ces_0_3_io_outs_up[44] ,
    \_ces_0_3_io_outs_up[43] ,
    \_ces_0_3_io_outs_up[42] ,
    \_ces_0_3_io_outs_up[41] ,
    \_ces_0_3_io_outs_up[40] ,
    \_ces_0_3_io_outs_up[39] ,
    \_ces_0_3_io_outs_up[38] ,
    \_ces_0_3_io_outs_up[37] ,
    \_ces_0_3_io_outs_up[36] ,
    \_ces_0_3_io_outs_up[35] ,
    \_ces_0_3_io_outs_up[34] ,
    \_ces_0_3_io_outs_up[33] ,
    \_ces_0_3_io_outs_up[32] ,
    \_ces_0_3_io_outs_up[31] ,
    \_ces_0_3_io_outs_up[30] ,
    \_ces_0_3_io_outs_up[29] ,
    \_ces_0_3_io_outs_up[28] ,
    \_ces_0_3_io_outs_up[27] ,
    \_ces_0_3_io_outs_up[26] ,
    \_ces_0_3_io_outs_up[25] ,
    \_ces_0_3_io_outs_up[24] ,
    \_ces_0_3_io_outs_up[23] ,
    \_ces_0_3_io_outs_up[22] ,
    \_ces_0_3_io_outs_up[21] ,
    \_ces_0_3_io_outs_up[20] ,
    \_ces_0_3_io_outs_up[19] ,
    \_ces_0_3_io_outs_up[18] ,
    \_ces_0_3_io_outs_up[17] ,
    \_ces_0_3_io_outs_up[16] ,
    \_ces_0_3_io_outs_up[15] ,
    \_ces_0_3_io_outs_up[14] ,
    \_ces_0_3_io_outs_up[13] ,
    \_ces_0_3_io_outs_up[12] ,
    \_ces_0_3_io_outs_up[11] ,
    \_ces_0_3_io_outs_up[10] ,
    \_ces_0_3_io_outs_up[9] ,
    \_ces_0_3_io_outs_up[8] ,
    \_ces_0_3_io_outs_up[7] ,
    \_ces_0_3_io_outs_up[6] ,
    \_ces_0_3_io_outs_up[5] ,
    \_ces_0_3_io_outs_up[4] ,
    \_ces_0_3_io_outs_up[3] ,
    \_ces_0_3_io_outs_up[2] ,
    \_ces_0_3_io_outs_up[1] ,
    \_ces_0_3_io_outs_up[0] }));
 Element ces_1_0 (.clock(clknet_leaf_3_clock),
    .io_lsbIns_1(net3),
    .io_lsbIns_2(net4),
    .io_lsbIns_3(net5),
    .io_lsbOuts_1(_ces_1_0_io_lsbOuts_1),
    .io_lsbOuts_2(_ces_1_0_io_lsbOuts_2),
    .io_lsbOuts_3(_ces_1_0_io_lsbOuts_3),
    .io_ins_down({\_ces_2_0_io_outs_down[63] ,
    \_ces_2_0_io_outs_down[62] ,
    \_ces_2_0_io_outs_down[61] ,
    \_ces_2_0_io_outs_down[60] ,
    \_ces_2_0_io_outs_down[59] ,
    \_ces_2_0_io_outs_down[58] ,
    \_ces_2_0_io_outs_down[57] ,
    \_ces_2_0_io_outs_down[56] ,
    \_ces_2_0_io_outs_down[55] ,
    \_ces_2_0_io_outs_down[54] ,
    \_ces_2_0_io_outs_down[53] ,
    \_ces_2_0_io_outs_down[52] ,
    \_ces_2_0_io_outs_down[51] ,
    \_ces_2_0_io_outs_down[50] ,
    \_ces_2_0_io_outs_down[49] ,
    \_ces_2_0_io_outs_down[48] ,
    \_ces_2_0_io_outs_down[47] ,
    \_ces_2_0_io_outs_down[46] ,
    \_ces_2_0_io_outs_down[45] ,
    \_ces_2_0_io_outs_down[44] ,
    \_ces_2_0_io_outs_down[43] ,
    \_ces_2_0_io_outs_down[42] ,
    \_ces_2_0_io_outs_down[41] ,
    \_ces_2_0_io_outs_down[40] ,
    \_ces_2_0_io_outs_down[39] ,
    \_ces_2_0_io_outs_down[38] ,
    \_ces_2_0_io_outs_down[37] ,
    \_ces_2_0_io_outs_down[36] ,
    \_ces_2_0_io_outs_down[35] ,
    \_ces_2_0_io_outs_down[34] ,
    \_ces_2_0_io_outs_down[33] ,
    \_ces_2_0_io_outs_down[32] ,
    \_ces_2_0_io_outs_down[31] ,
    \_ces_2_0_io_outs_down[30] ,
    \_ces_2_0_io_outs_down[29] ,
    \_ces_2_0_io_outs_down[28] ,
    \_ces_2_0_io_outs_down[27] ,
    \_ces_2_0_io_outs_down[26] ,
    \_ces_2_0_io_outs_down[25] ,
    \_ces_2_0_io_outs_down[24] ,
    \_ces_2_0_io_outs_down[23] ,
    \_ces_2_0_io_outs_down[22] ,
    \_ces_2_0_io_outs_down[21] ,
    \_ces_2_0_io_outs_down[20] ,
    \_ces_2_0_io_outs_down[19] ,
    \_ces_2_0_io_outs_down[18] ,
    \_ces_2_0_io_outs_down[17] ,
    \_ces_2_0_io_outs_down[16] ,
    \_ces_2_0_io_outs_down[15] ,
    \_ces_2_0_io_outs_down[14] ,
    \_ces_2_0_io_outs_down[13] ,
    \_ces_2_0_io_outs_down[12] ,
    \_ces_2_0_io_outs_down[11] ,
    \_ces_2_0_io_outs_down[10] ,
    \_ces_2_0_io_outs_down[9] ,
    \_ces_2_0_io_outs_down[8] ,
    \_ces_2_0_io_outs_down[7] ,
    \_ces_2_0_io_outs_down[6] ,
    \_ces_2_0_io_outs_down[5] ,
    \_ces_2_0_io_outs_down[4] ,
    \_ces_2_0_io_outs_down[3] ,
    \_ces_2_0_io_outs_down[2] ,
    \_ces_2_0_io_outs_down[1] ,
    \_ces_2_0_io_outs_down[0] }),
    .io_ins_left({\_ces_1_1_io_outs_left[63] ,
    \_ces_1_1_io_outs_left[62] ,
    \_ces_1_1_io_outs_left[61] ,
    \_ces_1_1_io_outs_left[60] ,
    \_ces_1_1_io_outs_left[59] ,
    \_ces_1_1_io_outs_left[58] ,
    \_ces_1_1_io_outs_left[57] ,
    \_ces_1_1_io_outs_left[56] ,
    \_ces_1_1_io_outs_left[55] ,
    \_ces_1_1_io_outs_left[54] ,
    \_ces_1_1_io_outs_left[53] ,
    \_ces_1_1_io_outs_left[52] ,
    \_ces_1_1_io_outs_left[51] ,
    \_ces_1_1_io_outs_left[50] ,
    \_ces_1_1_io_outs_left[49] ,
    \_ces_1_1_io_outs_left[48] ,
    \_ces_1_1_io_outs_left[47] ,
    \_ces_1_1_io_outs_left[46] ,
    \_ces_1_1_io_outs_left[45] ,
    \_ces_1_1_io_outs_left[44] ,
    \_ces_1_1_io_outs_left[43] ,
    \_ces_1_1_io_outs_left[42] ,
    \_ces_1_1_io_outs_left[41] ,
    \_ces_1_1_io_outs_left[40] ,
    \_ces_1_1_io_outs_left[39] ,
    \_ces_1_1_io_outs_left[38] ,
    \_ces_1_1_io_outs_left[37] ,
    \_ces_1_1_io_outs_left[36] ,
    \_ces_1_1_io_outs_left[35] ,
    \_ces_1_1_io_outs_left[34] ,
    \_ces_1_1_io_outs_left[33] ,
    \_ces_1_1_io_outs_left[32] ,
    \_ces_1_1_io_outs_left[31] ,
    \_ces_1_1_io_outs_left[30] ,
    \_ces_1_1_io_outs_left[29] ,
    \_ces_1_1_io_outs_left[28] ,
    \_ces_1_1_io_outs_left[27] ,
    \_ces_1_1_io_outs_left[26] ,
    \_ces_1_1_io_outs_left[25] ,
    \_ces_1_1_io_outs_left[24] ,
    \_ces_1_1_io_outs_left[23] ,
    \_ces_1_1_io_outs_left[22] ,
    \_ces_1_1_io_outs_left[21] ,
    \_ces_1_1_io_outs_left[20] ,
    \_ces_1_1_io_outs_left[19] ,
    \_ces_1_1_io_outs_left[18] ,
    \_ces_1_1_io_outs_left[17] ,
    \_ces_1_1_io_outs_left[16] ,
    \_ces_1_1_io_outs_left[15] ,
    \_ces_1_1_io_outs_left[14] ,
    \_ces_1_1_io_outs_left[13] ,
    \_ces_1_1_io_outs_left[12] ,
    \_ces_1_1_io_outs_left[11] ,
    \_ces_1_1_io_outs_left[10] ,
    \_ces_1_1_io_outs_left[9] ,
    \_ces_1_1_io_outs_left[8] ,
    \_ces_1_1_io_outs_left[7] ,
    \_ces_1_1_io_outs_left[6] ,
    \_ces_1_1_io_outs_left[5] ,
    \_ces_1_1_io_outs_left[4] ,
    \_ces_1_1_io_outs_left[3] ,
    \_ces_1_1_io_outs_left[2] ,
    \_ces_1_1_io_outs_left[1] ,
    \_ces_1_1_io_outs_left[0] }),
    .io_ins_right({net647,
    net646,
    net645,
    net644,
    net642,
    net641,
    net640,
    net639,
    net638,
    net637,
    net636,
    net635,
    net634,
    net633,
    net631,
    net630,
    net629,
    net628,
    net627,
    net626,
    net625,
    net624,
    net623,
    net622,
    net620,
    net619,
    net618,
    net617,
    net616,
    net615,
    net614,
    net613,
    net612,
    net611,
    net609,
    net608,
    net607,
    net606,
    net605,
    net604,
    net603,
    net602,
    net601,
    net600,
    net598,
    net597,
    net596,
    net595,
    net594,
    net593,
    net592,
    net591,
    net590,
    net589,
    net651,
    net650,
    net649,
    net648,
    net643,
    net632,
    net621,
    net610,
    net599,
    net588}),
    .io_ins_up({\_ces_0_0_io_outs_up[63] ,
    \_ces_0_0_io_outs_up[62] ,
    \_ces_0_0_io_outs_up[61] ,
    \_ces_0_0_io_outs_up[60] ,
    \_ces_0_0_io_outs_up[59] ,
    \_ces_0_0_io_outs_up[58] ,
    \_ces_0_0_io_outs_up[57] ,
    \_ces_0_0_io_outs_up[56] ,
    \_ces_0_0_io_outs_up[55] ,
    \_ces_0_0_io_outs_up[54] ,
    \_ces_0_0_io_outs_up[53] ,
    \_ces_0_0_io_outs_up[52] ,
    \_ces_0_0_io_outs_up[51] ,
    \_ces_0_0_io_outs_up[50] ,
    \_ces_0_0_io_outs_up[49] ,
    \_ces_0_0_io_outs_up[48] ,
    \_ces_0_0_io_outs_up[47] ,
    \_ces_0_0_io_outs_up[46] ,
    \_ces_0_0_io_outs_up[45] ,
    \_ces_0_0_io_outs_up[44] ,
    \_ces_0_0_io_outs_up[43] ,
    \_ces_0_0_io_outs_up[42] ,
    \_ces_0_0_io_outs_up[41] ,
    \_ces_0_0_io_outs_up[40] ,
    \_ces_0_0_io_outs_up[39] ,
    \_ces_0_0_io_outs_up[38] ,
    \_ces_0_0_io_outs_up[37] ,
    \_ces_0_0_io_outs_up[36] ,
    \_ces_0_0_io_outs_up[35] ,
    \_ces_0_0_io_outs_up[34] ,
    \_ces_0_0_io_outs_up[33] ,
    \_ces_0_0_io_outs_up[32] ,
    \_ces_0_0_io_outs_up[31] ,
    \_ces_0_0_io_outs_up[30] ,
    \_ces_0_0_io_outs_up[29] ,
    \_ces_0_0_io_outs_up[28] ,
    \_ces_0_0_io_outs_up[27] ,
    \_ces_0_0_io_outs_up[26] ,
    \_ces_0_0_io_outs_up[25] ,
    \_ces_0_0_io_outs_up[24] ,
    \_ces_0_0_io_outs_up[23] ,
    \_ces_0_0_io_outs_up[22] ,
    \_ces_0_0_io_outs_up[21] ,
    \_ces_0_0_io_outs_up[20] ,
    \_ces_0_0_io_outs_up[19] ,
    \_ces_0_0_io_outs_up[18] ,
    \_ces_0_0_io_outs_up[17] ,
    \_ces_0_0_io_outs_up[16] ,
    \_ces_0_0_io_outs_up[15] ,
    \_ces_0_0_io_outs_up[14] ,
    \_ces_0_0_io_outs_up[13] ,
    \_ces_0_0_io_outs_up[12] ,
    \_ces_0_0_io_outs_up[11] ,
    \_ces_0_0_io_outs_up[10] ,
    \_ces_0_0_io_outs_up[9] ,
    \_ces_0_0_io_outs_up[8] ,
    \_ces_0_0_io_outs_up[7] ,
    \_ces_0_0_io_outs_up[6] ,
    \_ces_0_0_io_outs_up[5] ,
    \_ces_0_0_io_outs_up[4] ,
    \_ces_0_0_io_outs_up[3] ,
    \_ces_0_0_io_outs_up[2] ,
    \_ces_0_0_io_outs_up[1] ,
    \_ces_0_0_io_outs_up[0] }),
    .io_outs_down({\_ces_1_0_io_outs_down[63] ,
    \_ces_1_0_io_outs_down[62] ,
    \_ces_1_0_io_outs_down[61] ,
    \_ces_1_0_io_outs_down[60] ,
    \_ces_1_0_io_outs_down[59] ,
    \_ces_1_0_io_outs_down[58] ,
    \_ces_1_0_io_outs_down[57] ,
    \_ces_1_0_io_outs_down[56] ,
    \_ces_1_0_io_outs_down[55] ,
    \_ces_1_0_io_outs_down[54] ,
    \_ces_1_0_io_outs_down[53] ,
    \_ces_1_0_io_outs_down[52] ,
    \_ces_1_0_io_outs_down[51] ,
    \_ces_1_0_io_outs_down[50] ,
    \_ces_1_0_io_outs_down[49] ,
    \_ces_1_0_io_outs_down[48] ,
    \_ces_1_0_io_outs_down[47] ,
    \_ces_1_0_io_outs_down[46] ,
    \_ces_1_0_io_outs_down[45] ,
    \_ces_1_0_io_outs_down[44] ,
    \_ces_1_0_io_outs_down[43] ,
    \_ces_1_0_io_outs_down[42] ,
    \_ces_1_0_io_outs_down[41] ,
    \_ces_1_0_io_outs_down[40] ,
    \_ces_1_0_io_outs_down[39] ,
    \_ces_1_0_io_outs_down[38] ,
    \_ces_1_0_io_outs_down[37] ,
    \_ces_1_0_io_outs_down[36] ,
    \_ces_1_0_io_outs_down[35] ,
    \_ces_1_0_io_outs_down[34] ,
    \_ces_1_0_io_outs_down[33] ,
    \_ces_1_0_io_outs_down[32] ,
    \_ces_1_0_io_outs_down[31] ,
    \_ces_1_0_io_outs_down[30] ,
    \_ces_1_0_io_outs_down[29] ,
    \_ces_1_0_io_outs_down[28] ,
    \_ces_1_0_io_outs_down[27] ,
    \_ces_1_0_io_outs_down[26] ,
    \_ces_1_0_io_outs_down[25] ,
    \_ces_1_0_io_outs_down[24] ,
    \_ces_1_0_io_outs_down[23] ,
    \_ces_1_0_io_outs_down[22] ,
    \_ces_1_0_io_outs_down[21] ,
    \_ces_1_0_io_outs_down[20] ,
    \_ces_1_0_io_outs_down[19] ,
    \_ces_1_0_io_outs_down[18] ,
    \_ces_1_0_io_outs_down[17] ,
    \_ces_1_0_io_outs_down[16] ,
    \_ces_1_0_io_outs_down[15] ,
    \_ces_1_0_io_outs_down[14] ,
    \_ces_1_0_io_outs_down[13] ,
    \_ces_1_0_io_outs_down[12] ,
    \_ces_1_0_io_outs_down[11] ,
    \_ces_1_0_io_outs_down[10] ,
    \_ces_1_0_io_outs_down[9] ,
    \_ces_1_0_io_outs_down[8] ,
    \_ces_1_0_io_outs_down[7] ,
    \_ces_1_0_io_outs_down[6] ,
    \_ces_1_0_io_outs_down[5] ,
    \_ces_1_0_io_outs_down[4] ,
    \_ces_1_0_io_outs_down[3] ,
    \_ces_1_0_io_outs_down[2] ,
    \_ces_1_0_io_outs_down[1] ,
    \_ces_1_0_io_outs_down[0] }),
    .io_outs_left({net1431,
    net1430,
    net1429,
    net1428,
    net1426,
    net1425,
    net1424,
    net1423,
    net1422,
    net1421,
    net1420,
    net1419,
    net1418,
    net1417,
    net1415,
    net1414,
    net1413,
    net1412,
    net1411,
    net1410,
    net1409,
    net1408,
    net1407,
    net1406,
    net1404,
    net1403,
    net1402,
    net1401,
    net1400,
    net1399,
    net1398,
    net1397,
    net1396,
    net1395,
    net1393,
    net1392,
    net1391,
    net1390,
    net1389,
    net1388,
    net1387,
    net1386,
    net1385,
    net1384,
    net1382,
    net1381,
    net1380,
    net1379,
    net1378,
    net1377,
    net1376,
    net1375,
    net1374,
    net1373,
    net1435,
    net1434,
    net1433,
    net1432,
    net1427,
    net1416,
    net1405,
    net1394,
    net1383,
    net1372}),
    .io_outs_right({\_ces_1_0_io_outs_right[63] ,
    \_ces_1_0_io_outs_right[62] ,
    \_ces_1_0_io_outs_right[61] ,
    \_ces_1_0_io_outs_right[60] ,
    \_ces_1_0_io_outs_right[59] ,
    \_ces_1_0_io_outs_right[58] ,
    \_ces_1_0_io_outs_right[57] ,
    \_ces_1_0_io_outs_right[56] ,
    \_ces_1_0_io_outs_right[55] ,
    \_ces_1_0_io_outs_right[54] ,
    \_ces_1_0_io_outs_right[53] ,
    \_ces_1_0_io_outs_right[52] ,
    \_ces_1_0_io_outs_right[51] ,
    \_ces_1_0_io_outs_right[50] ,
    \_ces_1_0_io_outs_right[49] ,
    \_ces_1_0_io_outs_right[48] ,
    \_ces_1_0_io_outs_right[47] ,
    \_ces_1_0_io_outs_right[46] ,
    \_ces_1_0_io_outs_right[45] ,
    \_ces_1_0_io_outs_right[44] ,
    \_ces_1_0_io_outs_right[43] ,
    \_ces_1_0_io_outs_right[42] ,
    \_ces_1_0_io_outs_right[41] ,
    \_ces_1_0_io_outs_right[40] ,
    \_ces_1_0_io_outs_right[39] ,
    \_ces_1_0_io_outs_right[38] ,
    \_ces_1_0_io_outs_right[37] ,
    \_ces_1_0_io_outs_right[36] ,
    \_ces_1_0_io_outs_right[35] ,
    \_ces_1_0_io_outs_right[34] ,
    \_ces_1_0_io_outs_right[33] ,
    \_ces_1_0_io_outs_right[32] ,
    \_ces_1_0_io_outs_right[31] ,
    \_ces_1_0_io_outs_right[30] ,
    \_ces_1_0_io_outs_right[29] ,
    \_ces_1_0_io_outs_right[28] ,
    \_ces_1_0_io_outs_right[27] ,
    \_ces_1_0_io_outs_right[26] ,
    \_ces_1_0_io_outs_right[25] ,
    \_ces_1_0_io_outs_right[24] ,
    \_ces_1_0_io_outs_right[23] ,
    \_ces_1_0_io_outs_right[22] ,
    \_ces_1_0_io_outs_right[21] ,
    \_ces_1_0_io_outs_right[20] ,
    \_ces_1_0_io_outs_right[19] ,
    \_ces_1_0_io_outs_right[18] ,
    \_ces_1_0_io_outs_right[17] ,
    \_ces_1_0_io_outs_right[16] ,
    \_ces_1_0_io_outs_right[15] ,
    \_ces_1_0_io_outs_right[14] ,
    \_ces_1_0_io_outs_right[13] ,
    \_ces_1_0_io_outs_right[12] ,
    \_ces_1_0_io_outs_right[11] ,
    \_ces_1_0_io_outs_right[10] ,
    \_ces_1_0_io_outs_right[9] ,
    \_ces_1_0_io_outs_right[8] ,
    \_ces_1_0_io_outs_right[7] ,
    \_ces_1_0_io_outs_right[6] ,
    \_ces_1_0_io_outs_right[5] ,
    \_ces_1_0_io_outs_right[4] ,
    \_ces_1_0_io_outs_right[3] ,
    \_ces_1_0_io_outs_right[2] ,
    \_ces_1_0_io_outs_right[1] ,
    \_ces_1_0_io_outs_right[0] }),
    .io_outs_up({\_ces_1_0_io_outs_up[63] ,
    \_ces_1_0_io_outs_up[62] ,
    \_ces_1_0_io_outs_up[61] ,
    \_ces_1_0_io_outs_up[60] ,
    \_ces_1_0_io_outs_up[59] ,
    \_ces_1_0_io_outs_up[58] ,
    \_ces_1_0_io_outs_up[57] ,
    \_ces_1_0_io_outs_up[56] ,
    \_ces_1_0_io_outs_up[55] ,
    \_ces_1_0_io_outs_up[54] ,
    \_ces_1_0_io_outs_up[53] ,
    \_ces_1_0_io_outs_up[52] ,
    \_ces_1_0_io_outs_up[51] ,
    \_ces_1_0_io_outs_up[50] ,
    \_ces_1_0_io_outs_up[49] ,
    \_ces_1_0_io_outs_up[48] ,
    \_ces_1_0_io_outs_up[47] ,
    \_ces_1_0_io_outs_up[46] ,
    \_ces_1_0_io_outs_up[45] ,
    \_ces_1_0_io_outs_up[44] ,
    \_ces_1_0_io_outs_up[43] ,
    \_ces_1_0_io_outs_up[42] ,
    \_ces_1_0_io_outs_up[41] ,
    \_ces_1_0_io_outs_up[40] ,
    \_ces_1_0_io_outs_up[39] ,
    \_ces_1_0_io_outs_up[38] ,
    \_ces_1_0_io_outs_up[37] ,
    \_ces_1_0_io_outs_up[36] ,
    \_ces_1_0_io_outs_up[35] ,
    \_ces_1_0_io_outs_up[34] ,
    \_ces_1_0_io_outs_up[33] ,
    \_ces_1_0_io_outs_up[32] ,
    \_ces_1_0_io_outs_up[31] ,
    \_ces_1_0_io_outs_up[30] ,
    \_ces_1_0_io_outs_up[29] ,
    \_ces_1_0_io_outs_up[28] ,
    \_ces_1_0_io_outs_up[27] ,
    \_ces_1_0_io_outs_up[26] ,
    \_ces_1_0_io_outs_up[25] ,
    \_ces_1_0_io_outs_up[24] ,
    \_ces_1_0_io_outs_up[23] ,
    \_ces_1_0_io_outs_up[22] ,
    \_ces_1_0_io_outs_up[21] ,
    \_ces_1_0_io_outs_up[20] ,
    \_ces_1_0_io_outs_up[19] ,
    \_ces_1_0_io_outs_up[18] ,
    \_ces_1_0_io_outs_up[17] ,
    \_ces_1_0_io_outs_up[16] ,
    \_ces_1_0_io_outs_up[15] ,
    \_ces_1_0_io_outs_up[14] ,
    \_ces_1_0_io_outs_up[13] ,
    \_ces_1_0_io_outs_up[12] ,
    \_ces_1_0_io_outs_up[11] ,
    \_ces_1_0_io_outs_up[10] ,
    \_ces_1_0_io_outs_up[9] ,
    \_ces_1_0_io_outs_up[8] ,
    \_ces_1_0_io_outs_up[7] ,
    \_ces_1_0_io_outs_up[6] ,
    \_ces_1_0_io_outs_up[5] ,
    \_ces_1_0_io_outs_up[4] ,
    \_ces_1_0_io_outs_up[3] ,
    \_ces_1_0_io_outs_up[2] ,
    \_ces_1_0_io_outs_up[1] ,
    \_ces_1_0_io_outs_up[0] }));
 Element ces_1_1 (.clock(clknet_leaf_3_clock),
    .io_lsbIns_1(_ces_1_0_io_lsbOuts_1),
    .io_lsbIns_2(_ces_1_0_io_lsbOuts_2),
    .io_lsbIns_3(_ces_1_0_io_lsbOuts_3),
    .io_lsbOuts_1(_ces_1_1_io_lsbOuts_1),
    .io_lsbOuts_2(_ces_1_1_io_lsbOuts_2),
    .io_lsbOuts_3(_ces_1_1_io_lsbOuts_3),
    .io_ins_down({\_ces_2_1_io_outs_down[63] ,
    \_ces_2_1_io_outs_down[62] ,
    \_ces_2_1_io_outs_down[61] ,
    \_ces_2_1_io_outs_down[60] ,
    \_ces_2_1_io_outs_down[59] ,
    \_ces_2_1_io_outs_down[58] ,
    \_ces_2_1_io_outs_down[57] ,
    \_ces_2_1_io_outs_down[56] ,
    \_ces_2_1_io_outs_down[55] ,
    \_ces_2_1_io_outs_down[54] ,
    \_ces_2_1_io_outs_down[53] ,
    \_ces_2_1_io_outs_down[52] ,
    \_ces_2_1_io_outs_down[51] ,
    \_ces_2_1_io_outs_down[50] ,
    \_ces_2_1_io_outs_down[49] ,
    \_ces_2_1_io_outs_down[48] ,
    \_ces_2_1_io_outs_down[47] ,
    \_ces_2_1_io_outs_down[46] ,
    \_ces_2_1_io_outs_down[45] ,
    \_ces_2_1_io_outs_down[44] ,
    \_ces_2_1_io_outs_down[43] ,
    \_ces_2_1_io_outs_down[42] ,
    \_ces_2_1_io_outs_down[41] ,
    \_ces_2_1_io_outs_down[40] ,
    \_ces_2_1_io_outs_down[39] ,
    \_ces_2_1_io_outs_down[38] ,
    \_ces_2_1_io_outs_down[37] ,
    \_ces_2_1_io_outs_down[36] ,
    \_ces_2_1_io_outs_down[35] ,
    \_ces_2_1_io_outs_down[34] ,
    \_ces_2_1_io_outs_down[33] ,
    \_ces_2_1_io_outs_down[32] ,
    \_ces_2_1_io_outs_down[31] ,
    \_ces_2_1_io_outs_down[30] ,
    \_ces_2_1_io_outs_down[29] ,
    \_ces_2_1_io_outs_down[28] ,
    \_ces_2_1_io_outs_down[27] ,
    \_ces_2_1_io_outs_down[26] ,
    \_ces_2_1_io_outs_down[25] ,
    \_ces_2_1_io_outs_down[24] ,
    \_ces_2_1_io_outs_down[23] ,
    \_ces_2_1_io_outs_down[22] ,
    \_ces_2_1_io_outs_down[21] ,
    \_ces_2_1_io_outs_down[20] ,
    \_ces_2_1_io_outs_down[19] ,
    \_ces_2_1_io_outs_down[18] ,
    \_ces_2_1_io_outs_down[17] ,
    \_ces_2_1_io_outs_down[16] ,
    \_ces_2_1_io_outs_down[15] ,
    \_ces_2_1_io_outs_down[14] ,
    \_ces_2_1_io_outs_down[13] ,
    \_ces_2_1_io_outs_down[12] ,
    \_ces_2_1_io_outs_down[11] ,
    \_ces_2_1_io_outs_down[10] ,
    \_ces_2_1_io_outs_down[9] ,
    \_ces_2_1_io_outs_down[8] ,
    \_ces_2_1_io_outs_down[7] ,
    \_ces_2_1_io_outs_down[6] ,
    \_ces_2_1_io_outs_down[5] ,
    \_ces_2_1_io_outs_down[4] ,
    \_ces_2_1_io_outs_down[3] ,
    \_ces_2_1_io_outs_down[2] ,
    \_ces_2_1_io_outs_down[1] ,
    \_ces_2_1_io_outs_down[0] }),
    .io_ins_left({\_ces_1_2_io_outs_left[63] ,
    \_ces_1_2_io_outs_left[62] ,
    \_ces_1_2_io_outs_left[61] ,
    \_ces_1_2_io_outs_left[60] ,
    \_ces_1_2_io_outs_left[59] ,
    \_ces_1_2_io_outs_left[58] ,
    \_ces_1_2_io_outs_left[57] ,
    \_ces_1_2_io_outs_left[56] ,
    \_ces_1_2_io_outs_left[55] ,
    \_ces_1_2_io_outs_left[54] ,
    \_ces_1_2_io_outs_left[53] ,
    \_ces_1_2_io_outs_left[52] ,
    \_ces_1_2_io_outs_left[51] ,
    \_ces_1_2_io_outs_left[50] ,
    \_ces_1_2_io_outs_left[49] ,
    \_ces_1_2_io_outs_left[48] ,
    \_ces_1_2_io_outs_left[47] ,
    \_ces_1_2_io_outs_left[46] ,
    \_ces_1_2_io_outs_left[45] ,
    \_ces_1_2_io_outs_left[44] ,
    \_ces_1_2_io_outs_left[43] ,
    \_ces_1_2_io_outs_left[42] ,
    \_ces_1_2_io_outs_left[41] ,
    \_ces_1_2_io_outs_left[40] ,
    \_ces_1_2_io_outs_left[39] ,
    \_ces_1_2_io_outs_left[38] ,
    \_ces_1_2_io_outs_left[37] ,
    \_ces_1_2_io_outs_left[36] ,
    \_ces_1_2_io_outs_left[35] ,
    \_ces_1_2_io_outs_left[34] ,
    \_ces_1_2_io_outs_left[33] ,
    \_ces_1_2_io_outs_left[32] ,
    \_ces_1_2_io_outs_left[31] ,
    \_ces_1_2_io_outs_left[30] ,
    \_ces_1_2_io_outs_left[29] ,
    \_ces_1_2_io_outs_left[28] ,
    \_ces_1_2_io_outs_left[27] ,
    \_ces_1_2_io_outs_left[26] ,
    \_ces_1_2_io_outs_left[25] ,
    \_ces_1_2_io_outs_left[24] ,
    \_ces_1_2_io_outs_left[23] ,
    \_ces_1_2_io_outs_left[22] ,
    \_ces_1_2_io_outs_left[21] ,
    \_ces_1_2_io_outs_left[20] ,
    \_ces_1_2_io_outs_left[19] ,
    \_ces_1_2_io_outs_left[18] ,
    \_ces_1_2_io_outs_left[17] ,
    \_ces_1_2_io_outs_left[16] ,
    \_ces_1_2_io_outs_left[15] ,
    \_ces_1_2_io_outs_left[14] ,
    \_ces_1_2_io_outs_left[13] ,
    \_ces_1_2_io_outs_left[12] ,
    \_ces_1_2_io_outs_left[11] ,
    \_ces_1_2_io_outs_left[10] ,
    \_ces_1_2_io_outs_left[9] ,
    \_ces_1_2_io_outs_left[8] ,
    \_ces_1_2_io_outs_left[7] ,
    \_ces_1_2_io_outs_left[6] ,
    \_ces_1_2_io_outs_left[5] ,
    \_ces_1_2_io_outs_left[4] ,
    \_ces_1_2_io_outs_left[3] ,
    \_ces_1_2_io_outs_left[2] ,
    \_ces_1_2_io_outs_left[1] ,
    \_ces_1_2_io_outs_left[0] }),
    .io_ins_right({\_ces_1_0_io_outs_right[63] ,
    \_ces_1_0_io_outs_right[62] ,
    \_ces_1_0_io_outs_right[61] ,
    \_ces_1_0_io_outs_right[60] ,
    \_ces_1_0_io_outs_right[59] ,
    \_ces_1_0_io_outs_right[58] ,
    \_ces_1_0_io_outs_right[57] ,
    \_ces_1_0_io_outs_right[56] ,
    \_ces_1_0_io_outs_right[55] ,
    \_ces_1_0_io_outs_right[54] ,
    \_ces_1_0_io_outs_right[53] ,
    \_ces_1_0_io_outs_right[52] ,
    \_ces_1_0_io_outs_right[51] ,
    \_ces_1_0_io_outs_right[50] ,
    \_ces_1_0_io_outs_right[49] ,
    \_ces_1_0_io_outs_right[48] ,
    \_ces_1_0_io_outs_right[47] ,
    \_ces_1_0_io_outs_right[46] ,
    \_ces_1_0_io_outs_right[45] ,
    \_ces_1_0_io_outs_right[44] ,
    \_ces_1_0_io_outs_right[43] ,
    \_ces_1_0_io_outs_right[42] ,
    \_ces_1_0_io_outs_right[41] ,
    \_ces_1_0_io_outs_right[40] ,
    \_ces_1_0_io_outs_right[39] ,
    \_ces_1_0_io_outs_right[38] ,
    \_ces_1_0_io_outs_right[37] ,
    \_ces_1_0_io_outs_right[36] ,
    \_ces_1_0_io_outs_right[35] ,
    \_ces_1_0_io_outs_right[34] ,
    \_ces_1_0_io_outs_right[33] ,
    \_ces_1_0_io_outs_right[32] ,
    \_ces_1_0_io_outs_right[31] ,
    \_ces_1_0_io_outs_right[30] ,
    \_ces_1_0_io_outs_right[29] ,
    \_ces_1_0_io_outs_right[28] ,
    \_ces_1_0_io_outs_right[27] ,
    \_ces_1_0_io_outs_right[26] ,
    \_ces_1_0_io_outs_right[25] ,
    \_ces_1_0_io_outs_right[24] ,
    \_ces_1_0_io_outs_right[23] ,
    \_ces_1_0_io_outs_right[22] ,
    \_ces_1_0_io_outs_right[21] ,
    \_ces_1_0_io_outs_right[20] ,
    \_ces_1_0_io_outs_right[19] ,
    \_ces_1_0_io_outs_right[18] ,
    \_ces_1_0_io_outs_right[17] ,
    \_ces_1_0_io_outs_right[16] ,
    \_ces_1_0_io_outs_right[15] ,
    \_ces_1_0_io_outs_right[14] ,
    \_ces_1_0_io_outs_right[13] ,
    \_ces_1_0_io_outs_right[12] ,
    \_ces_1_0_io_outs_right[11] ,
    \_ces_1_0_io_outs_right[10] ,
    \_ces_1_0_io_outs_right[9] ,
    \_ces_1_0_io_outs_right[8] ,
    \_ces_1_0_io_outs_right[7] ,
    \_ces_1_0_io_outs_right[6] ,
    \_ces_1_0_io_outs_right[5] ,
    \_ces_1_0_io_outs_right[4] ,
    \_ces_1_0_io_outs_right[3] ,
    \_ces_1_0_io_outs_right[2] ,
    \_ces_1_0_io_outs_right[1] ,
    \_ces_1_0_io_outs_right[0] }),
    .io_ins_up({\_ces_0_1_io_outs_up[63] ,
    \_ces_0_1_io_outs_up[62] ,
    \_ces_0_1_io_outs_up[61] ,
    \_ces_0_1_io_outs_up[60] ,
    \_ces_0_1_io_outs_up[59] ,
    \_ces_0_1_io_outs_up[58] ,
    \_ces_0_1_io_outs_up[57] ,
    \_ces_0_1_io_outs_up[56] ,
    \_ces_0_1_io_outs_up[55] ,
    \_ces_0_1_io_outs_up[54] ,
    \_ces_0_1_io_outs_up[53] ,
    \_ces_0_1_io_outs_up[52] ,
    \_ces_0_1_io_outs_up[51] ,
    \_ces_0_1_io_outs_up[50] ,
    \_ces_0_1_io_outs_up[49] ,
    \_ces_0_1_io_outs_up[48] ,
    \_ces_0_1_io_outs_up[47] ,
    \_ces_0_1_io_outs_up[46] ,
    \_ces_0_1_io_outs_up[45] ,
    \_ces_0_1_io_outs_up[44] ,
    \_ces_0_1_io_outs_up[43] ,
    \_ces_0_1_io_outs_up[42] ,
    \_ces_0_1_io_outs_up[41] ,
    \_ces_0_1_io_outs_up[40] ,
    \_ces_0_1_io_outs_up[39] ,
    \_ces_0_1_io_outs_up[38] ,
    \_ces_0_1_io_outs_up[37] ,
    \_ces_0_1_io_outs_up[36] ,
    \_ces_0_1_io_outs_up[35] ,
    \_ces_0_1_io_outs_up[34] ,
    \_ces_0_1_io_outs_up[33] ,
    \_ces_0_1_io_outs_up[32] ,
    \_ces_0_1_io_outs_up[31] ,
    \_ces_0_1_io_outs_up[30] ,
    \_ces_0_1_io_outs_up[29] ,
    \_ces_0_1_io_outs_up[28] ,
    \_ces_0_1_io_outs_up[27] ,
    \_ces_0_1_io_outs_up[26] ,
    \_ces_0_1_io_outs_up[25] ,
    \_ces_0_1_io_outs_up[24] ,
    \_ces_0_1_io_outs_up[23] ,
    \_ces_0_1_io_outs_up[22] ,
    \_ces_0_1_io_outs_up[21] ,
    \_ces_0_1_io_outs_up[20] ,
    \_ces_0_1_io_outs_up[19] ,
    \_ces_0_1_io_outs_up[18] ,
    \_ces_0_1_io_outs_up[17] ,
    \_ces_0_1_io_outs_up[16] ,
    \_ces_0_1_io_outs_up[15] ,
    \_ces_0_1_io_outs_up[14] ,
    \_ces_0_1_io_outs_up[13] ,
    \_ces_0_1_io_outs_up[12] ,
    \_ces_0_1_io_outs_up[11] ,
    \_ces_0_1_io_outs_up[10] ,
    \_ces_0_1_io_outs_up[9] ,
    \_ces_0_1_io_outs_up[8] ,
    \_ces_0_1_io_outs_up[7] ,
    \_ces_0_1_io_outs_up[6] ,
    \_ces_0_1_io_outs_up[5] ,
    \_ces_0_1_io_outs_up[4] ,
    \_ces_0_1_io_outs_up[3] ,
    \_ces_0_1_io_outs_up[2] ,
    \_ces_0_1_io_outs_up[1] ,
    \_ces_0_1_io_outs_up[0] }),
    .io_outs_down({\_ces_1_1_io_outs_down[63] ,
    \_ces_1_1_io_outs_down[62] ,
    \_ces_1_1_io_outs_down[61] ,
    \_ces_1_1_io_outs_down[60] ,
    \_ces_1_1_io_outs_down[59] ,
    \_ces_1_1_io_outs_down[58] ,
    \_ces_1_1_io_outs_down[57] ,
    \_ces_1_1_io_outs_down[56] ,
    \_ces_1_1_io_outs_down[55] ,
    \_ces_1_1_io_outs_down[54] ,
    \_ces_1_1_io_outs_down[53] ,
    \_ces_1_1_io_outs_down[52] ,
    \_ces_1_1_io_outs_down[51] ,
    \_ces_1_1_io_outs_down[50] ,
    \_ces_1_1_io_outs_down[49] ,
    \_ces_1_1_io_outs_down[48] ,
    \_ces_1_1_io_outs_down[47] ,
    \_ces_1_1_io_outs_down[46] ,
    \_ces_1_1_io_outs_down[45] ,
    \_ces_1_1_io_outs_down[44] ,
    \_ces_1_1_io_outs_down[43] ,
    \_ces_1_1_io_outs_down[42] ,
    \_ces_1_1_io_outs_down[41] ,
    \_ces_1_1_io_outs_down[40] ,
    \_ces_1_1_io_outs_down[39] ,
    \_ces_1_1_io_outs_down[38] ,
    \_ces_1_1_io_outs_down[37] ,
    \_ces_1_1_io_outs_down[36] ,
    \_ces_1_1_io_outs_down[35] ,
    \_ces_1_1_io_outs_down[34] ,
    \_ces_1_1_io_outs_down[33] ,
    \_ces_1_1_io_outs_down[32] ,
    \_ces_1_1_io_outs_down[31] ,
    \_ces_1_1_io_outs_down[30] ,
    \_ces_1_1_io_outs_down[29] ,
    \_ces_1_1_io_outs_down[28] ,
    \_ces_1_1_io_outs_down[27] ,
    \_ces_1_1_io_outs_down[26] ,
    \_ces_1_1_io_outs_down[25] ,
    \_ces_1_1_io_outs_down[24] ,
    \_ces_1_1_io_outs_down[23] ,
    \_ces_1_1_io_outs_down[22] ,
    \_ces_1_1_io_outs_down[21] ,
    \_ces_1_1_io_outs_down[20] ,
    \_ces_1_1_io_outs_down[19] ,
    \_ces_1_1_io_outs_down[18] ,
    \_ces_1_1_io_outs_down[17] ,
    \_ces_1_1_io_outs_down[16] ,
    \_ces_1_1_io_outs_down[15] ,
    \_ces_1_1_io_outs_down[14] ,
    \_ces_1_1_io_outs_down[13] ,
    \_ces_1_1_io_outs_down[12] ,
    \_ces_1_1_io_outs_down[11] ,
    \_ces_1_1_io_outs_down[10] ,
    \_ces_1_1_io_outs_down[9] ,
    \_ces_1_1_io_outs_down[8] ,
    \_ces_1_1_io_outs_down[7] ,
    \_ces_1_1_io_outs_down[6] ,
    \_ces_1_1_io_outs_down[5] ,
    \_ces_1_1_io_outs_down[4] ,
    \_ces_1_1_io_outs_down[3] ,
    \_ces_1_1_io_outs_down[2] ,
    \_ces_1_1_io_outs_down[1] ,
    \_ces_1_1_io_outs_down[0] }),
    .io_outs_left({\_ces_1_1_io_outs_left[63] ,
    \_ces_1_1_io_outs_left[62] ,
    \_ces_1_1_io_outs_left[61] ,
    \_ces_1_1_io_outs_left[60] ,
    \_ces_1_1_io_outs_left[59] ,
    \_ces_1_1_io_outs_left[58] ,
    \_ces_1_1_io_outs_left[57] ,
    \_ces_1_1_io_outs_left[56] ,
    \_ces_1_1_io_outs_left[55] ,
    \_ces_1_1_io_outs_left[54] ,
    \_ces_1_1_io_outs_left[53] ,
    \_ces_1_1_io_outs_left[52] ,
    \_ces_1_1_io_outs_left[51] ,
    \_ces_1_1_io_outs_left[50] ,
    \_ces_1_1_io_outs_left[49] ,
    \_ces_1_1_io_outs_left[48] ,
    \_ces_1_1_io_outs_left[47] ,
    \_ces_1_1_io_outs_left[46] ,
    \_ces_1_1_io_outs_left[45] ,
    \_ces_1_1_io_outs_left[44] ,
    \_ces_1_1_io_outs_left[43] ,
    \_ces_1_1_io_outs_left[42] ,
    \_ces_1_1_io_outs_left[41] ,
    \_ces_1_1_io_outs_left[40] ,
    \_ces_1_1_io_outs_left[39] ,
    \_ces_1_1_io_outs_left[38] ,
    \_ces_1_1_io_outs_left[37] ,
    \_ces_1_1_io_outs_left[36] ,
    \_ces_1_1_io_outs_left[35] ,
    \_ces_1_1_io_outs_left[34] ,
    \_ces_1_1_io_outs_left[33] ,
    \_ces_1_1_io_outs_left[32] ,
    \_ces_1_1_io_outs_left[31] ,
    \_ces_1_1_io_outs_left[30] ,
    \_ces_1_1_io_outs_left[29] ,
    \_ces_1_1_io_outs_left[28] ,
    \_ces_1_1_io_outs_left[27] ,
    \_ces_1_1_io_outs_left[26] ,
    \_ces_1_1_io_outs_left[25] ,
    \_ces_1_1_io_outs_left[24] ,
    \_ces_1_1_io_outs_left[23] ,
    \_ces_1_1_io_outs_left[22] ,
    \_ces_1_1_io_outs_left[21] ,
    \_ces_1_1_io_outs_left[20] ,
    \_ces_1_1_io_outs_left[19] ,
    \_ces_1_1_io_outs_left[18] ,
    \_ces_1_1_io_outs_left[17] ,
    \_ces_1_1_io_outs_left[16] ,
    \_ces_1_1_io_outs_left[15] ,
    \_ces_1_1_io_outs_left[14] ,
    \_ces_1_1_io_outs_left[13] ,
    \_ces_1_1_io_outs_left[12] ,
    \_ces_1_1_io_outs_left[11] ,
    \_ces_1_1_io_outs_left[10] ,
    \_ces_1_1_io_outs_left[9] ,
    \_ces_1_1_io_outs_left[8] ,
    \_ces_1_1_io_outs_left[7] ,
    \_ces_1_1_io_outs_left[6] ,
    \_ces_1_1_io_outs_left[5] ,
    \_ces_1_1_io_outs_left[4] ,
    \_ces_1_1_io_outs_left[3] ,
    \_ces_1_1_io_outs_left[2] ,
    \_ces_1_1_io_outs_left[1] ,
    \_ces_1_1_io_outs_left[0] }),
    .io_outs_right({\_ces_1_1_io_outs_right[63] ,
    \_ces_1_1_io_outs_right[62] ,
    \_ces_1_1_io_outs_right[61] ,
    \_ces_1_1_io_outs_right[60] ,
    \_ces_1_1_io_outs_right[59] ,
    \_ces_1_1_io_outs_right[58] ,
    \_ces_1_1_io_outs_right[57] ,
    \_ces_1_1_io_outs_right[56] ,
    \_ces_1_1_io_outs_right[55] ,
    \_ces_1_1_io_outs_right[54] ,
    \_ces_1_1_io_outs_right[53] ,
    \_ces_1_1_io_outs_right[52] ,
    \_ces_1_1_io_outs_right[51] ,
    \_ces_1_1_io_outs_right[50] ,
    \_ces_1_1_io_outs_right[49] ,
    \_ces_1_1_io_outs_right[48] ,
    \_ces_1_1_io_outs_right[47] ,
    \_ces_1_1_io_outs_right[46] ,
    \_ces_1_1_io_outs_right[45] ,
    \_ces_1_1_io_outs_right[44] ,
    \_ces_1_1_io_outs_right[43] ,
    \_ces_1_1_io_outs_right[42] ,
    \_ces_1_1_io_outs_right[41] ,
    \_ces_1_1_io_outs_right[40] ,
    \_ces_1_1_io_outs_right[39] ,
    \_ces_1_1_io_outs_right[38] ,
    \_ces_1_1_io_outs_right[37] ,
    \_ces_1_1_io_outs_right[36] ,
    \_ces_1_1_io_outs_right[35] ,
    \_ces_1_1_io_outs_right[34] ,
    \_ces_1_1_io_outs_right[33] ,
    \_ces_1_1_io_outs_right[32] ,
    \_ces_1_1_io_outs_right[31] ,
    \_ces_1_1_io_outs_right[30] ,
    \_ces_1_1_io_outs_right[29] ,
    \_ces_1_1_io_outs_right[28] ,
    \_ces_1_1_io_outs_right[27] ,
    \_ces_1_1_io_outs_right[26] ,
    \_ces_1_1_io_outs_right[25] ,
    \_ces_1_1_io_outs_right[24] ,
    \_ces_1_1_io_outs_right[23] ,
    \_ces_1_1_io_outs_right[22] ,
    \_ces_1_1_io_outs_right[21] ,
    \_ces_1_1_io_outs_right[20] ,
    \_ces_1_1_io_outs_right[19] ,
    \_ces_1_1_io_outs_right[18] ,
    \_ces_1_1_io_outs_right[17] ,
    \_ces_1_1_io_outs_right[16] ,
    \_ces_1_1_io_outs_right[15] ,
    \_ces_1_1_io_outs_right[14] ,
    \_ces_1_1_io_outs_right[13] ,
    \_ces_1_1_io_outs_right[12] ,
    \_ces_1_1_io_outs_right[11] ,
    \_ces_1_1_io_outs_right[10] ,
    \_ces_1_1_io_outs_right[9] ,
    \_ces_1_1_io_outs_right[8] ,
    \_ces_1_1_io_outs_right[7] ,
    \_ces_1_1_io_outs_right[6] ,
    \_ces_1_1_io_outs_right[5] ,
    \_ces_1_1_io_outs_right[4] ,
    \_ces_1_1_io_outs_right[3] ,
    \_ces_1_1_io_outs_right[2] ,
    \_ces_1_1_io_outs_right[1] ,
    \_ces_1_1_io_outs_right[0] }),
    .io_outs_up({\_ces_1_1_io_outs_up[63] ,
    \_ces_1_1_io_outs_up[62] ,
    \_ces_1_1_io_outs_up[61] ,
    \_ces_1_1_io_outs_up[60] ,
    \_ces_1_1_io_outs_up[59] ,
    \_ces_1_1_io_outs_up[58] ,
    \_ces_1_1_io_outs_up[57] ,
    \_ces_1_1_io_outs_up[56] ,
    \_ces_1_1_io_outs_up[55] ,
    \_ces_1_1_io_outs_up[54] ,
    \_ces_1_1_io_outs_up[53] ,
    \_ces_1_1_io_outs_up[52] ,
    \_ces_1_1_io_outs_up[51] ,
    \_ces_1_1_io_outs_up[50] ,
    \_ces_1_1_io_outs_up[49] ,
    \_ces_1_1_io_outs_up[48] ,
    \_ces_1_1_io_outs_up[47] ,
    \_ces_1_1_io_outs_up[46] ,
    \_ces_1_1_io_outs_up[45] ,
    \_ces_1_1_io_outs_up[44] ,
    \_ces_1_1_io_outs_up[43] ,
    \_ces_1_1_io_outs_up[42] ,
    \_ces_1_1_io_outs_up[41] ,
    \_ces_1_1_io_outs_up[40] ,
    \_ces_1_1_io_outs_up[39] ,
    \_ces_1_1_io_outs_up[38] ,
    \_ces_1_1_io_outs_up[37] ,
    \_ces_1_1_io_outs_up[36] ,
    \_ces_1_1_io_outs_up[35] ,
    \_ces_1_1_io_outs_up[34] ,
    \_ces_1_1_io_outs_up[33] ,
    \_ces_1_1_io_outs_up[32] ,
    \_ces_1_1_io_outs_up[31] ,
    \_ces_1_1_io_outs_up[30] ,
    \_ces_1_1_io_outs_up[29] ,
    \_ces_1_1_io_outs_up[28] ,
    \_ces_1_1_io_outs_up[27] ,
    \_ces_1_1_io_outs_up[26] ,
    \_ces_1_1_io_outs_up[25] ,
    \_ces_1_1_io_outs_up[24] ,
    \_ces_1_1_io_outs_up[23] ,
    \_ces_1_1_io_outs_up[22] ,
    \_ces_1_1_io_outs_up[21] ,
    \_ces_1_1_io_outs_up[20] ,
    \_ces_1_1_io_outs_up[19] ,
    \_ces_1_1_io_outs_up[18] ,
    \_ces_1_1_io_outs_up[17] ,
    \_ces_1_1_io_outs_up[16] ,
    \_ces_1_1_io_outs_up[15] ,
    \_ces_1_1_io_outs_up[14] ,
    \_ces_1_1_io_outs_up[13] ,
    \_ces_1_1_io_outs_up[12] ,
    \_ces_1_1_io_outs_up[11] ,
    \_ces_1_1_io_outs_up[10] ,
    \_ces_1_1_io_outs_up[9] ,
    \_ces_1_1_io_outs_up[8] ,
    \_ces_1_1_io_outs_up[7] ,
    \_ces_1_1_io_outs_up[6] ,
    \_ces_1_1_io_outs_up[5] ,
    \_ces_1_1_io_outs_up[4] ,
    \_ces_1_1_io_outs_up[3] ,
    \_ces_1_1_io_outs_up[2] ,
    \_ces_1_1_io_outs_up[1] ,
    \_ces_1_1_io_outs_up[0] }));
 Element ces_1_2 (.clock(clknet_leaf_2_clock),
    .io_lsbIns_1(_ces_1_1_io_lsbOuts_1),
    .io_lsbIns_2(_ces_1_1_io_lsbOuts_2),
    .io_lsbIns_3(_ces_1_1_io_lsbOuts_3),
    .io_lsbOuts_1(_ces_1_2_io_lsbOuts_1),
    .io_lsbOuts_2(_ces_1_2_io_lsbOuts_2),
    .io_lsbOuts_3(_ces_1_2_io_lsbOuts_3),
    .io_ins_down({\_ces_2_2_io_outs_down[63] ,
    \_ces_2_2_io_outs_down[62] ,
    \_ces_2_2_io_outs_down[61] ,
    \_ces_2_2_io_outs_down[60] ,
    \_ces_2_2_io_outs_down[59] ,
    \_ces_2_2_io_outs_down[58] ,
    \_ces_2_2_io_outs_down[57] ,
    \_ces_2_2_io_outs_down[56] ,
    \_ces_2_2_io_outs_down[55] ,
    \_ces_2_2_io_outs_down[54] ,
    \_ces_2_2_io_outs_down[53] ,
    \_ces_2_2_io_outs_down[52] ,
    \_ces_2_2_io_outs_down[51] ,
    \_ces_2_2_io_outs_down[50] ,
    \_ces_2_2_io_outs_down[49] ,
    \_ces_2_2_io_outs_down[48] ,
    \_ces_2_2_io_outs_down[47] ,
    \_ces_2_2_io_outs_down[46] ,
    \_ces_2_2_io_outs_down[45] ,
    \_ces_2_2_io_outs_down[44] ,
    \_ces_2_2_io_outs_down[43] ,
    \_ces_2_2_io_outs_down[42] ,
    \_ces_2_2_io_outs_down[41] ,
    \_ces_2_2_io_outs_down[40] ,
    \_ces_2_2_io_outs_down[39] ,
    \_ces_2_2_io_outs_down[38] ,
    \_ces_2_2_io_outs_down[37] ,
    \_ces_2_2_io_outs_down[36] ,
    \_ces_2_2_io_outs_down[35] ,
    \_ces_2_2_io_outs_down[34] ,
    \_ces_2_2_io_outs_down[33] ,
    \_ces_2_2_io_outs_down[32] ,
    \_ces_2_2_io_outs_down[31] ,
    \_ces_2_2_io_outs_down[30] ,
    \_ces_2_2_io_outs_down[29] ,
    \_ces_2_2_io_outs_down[28] ,
    \_ces_2_2_io_outs_down[27] ,
    \_ces_2_2_io_outs_down[26] ,
    \_ces_2_2_io_outs_down[25] ,
    \_ces_2_2_io_outs_down[24] ,
    \_ces_2_2_io_outs_down[23] ,
    \_ces_2_2_io_outs_down[22] ,
    \_ces_2_2_io_outs_down[21] ,
    \_ces_2_2_io_outs_down[20] ,
    \_ces_2_2_io_outs_down[19] ,
    \_ces_2_2_io_outs_down[18] ,
    \_ces_2_2_io_outs_down[17] ,
    \_ces_2_2_io_outs_down[16] ,
    \_ces_2_2_io_outs_down[15] ,
    \_ces_2_2_io_outs_down[14] ,
    \_ces_2_2_io_outs_down[13] ,
    \_ces_2_2_io_outs_down[12] ,
    \_ces_2_2_io_outs_down[11] ,
    \_ces_2_2_io_outs_down[10] ,
    \_ces_2_2_io_outs_down[9] ,
    \_ces_2_2_io_outs_down[8] ,
    \_ces_2_2_io_outs_down[7] ,
    \_ces_2_2_io_outs_down[6] ,
    \_ces_2_2_io_outs_down[5] ,
    \_ces_2_2_io_outs_down[4] ,
    \_ces_2_2_io_outs_down[3] ,
    \_ces_2_2_io_outs_down[2] ,
    \_ces_2_2_io_outs_down[1] ,
    \_ces_2_2_io_outs_down[0] }),
    .io_ins_left({\_ces_1_3_io_outs_left[63] ,
    \_ces_1_3_io_outs_left[62] ,
    \_ces_1_3_io_outs_left[61] ,
    \_ces_1_3_io_outs_left[60] ,
    \_ces_1_3_io_outs_left[59] ,
    \_ces_1_3_io_outs_left[58] ,
    \_ces_1_3_io_outs_left[57] ,
    \_ces_1_3_io_outs_left[56] ,
    \_ces_1_3_io_outs_left[55] ,
    \_ces_1_3_io_outs_left[54] ,
    \_ces_1_3_io_outs_left[53] ,
    \_ces_1_3_io_outs_left[52] ,
    \_ces_1_3_io_outs_left[51] ,
    \_ces_1_3_io_outs_left[50] ,
    \_ces_1_3_io_outs_left[49] ,
    \_ces_1_3_io_outs_left[48] ,
    \_ces_1_3_io_outs_left[47] ,
    \_ces_1_3_io_outs_left[46] ,
    \_ces_1_3_io_outs_left[45] ,
    \_ces_1_3_io_outs_left[44] ,
    \_ces_1_3_io_outs_left[43] ,
    \_ces_1_3_io_outs_left[42] ,
    \_ces_1_3_io_outs_left[41] ,
    \_ces_1_3_io_outs_left[40] ,
    \_ces_1_3_io_outs_left[39] ,
    \_ces_1_3_io_outs_left[38] ,
    \_ces_1_3_io_outs_left[37] ,
    \_ces_1_3_io_outs_left[36] ,
    \_ces_1_3_io_outs_left[35] ,
    \_ces_1_3_io_outs_left[34] ,
    \_ces_1_3_io_outs_left[33] ,
    \_ces_1_3_io_outs_left[32] ,
    \_ces_1_3_io_outs_left[31] ,
    \_ces_1_3_io_outs_left[30] ,
    \_ces_1_3_io_outs_left[29] ,
    \_ces_1_3_io_outs_left[28] ,
    \_ces_1_3_io_outs_left[27] ,
    \_ces_1_3_io_outs_left[26] ,
    \_ces_1_3_io_outs_left[25] ,
    \_ces_1_3_io_outs_left[24] ,
    \_ces_1_3_io_outs_left[23] ,
    \_ces_1_3_io_outs_left[22] ,
    \_ces_1_3_io_outs_left[21] ,
    \_ces_1_3_io_outs_left[20] ,
    \_ces_1_3_io_outs_left[19] ,
    \_ces_1_3_io_outs_left[18] ,
    \_ces_1_3_io_outs_left[17] ,
    \_ces_1_3_io_outs_left[16] ,
    \_ces_1_3_io_outs_left[15] ,
    \_ces_1_3_io_outs_left[14] ,
    \_ces_1_3_io_outs_left[13] ,
    \_ces_1_3_io_outs_left[12] ,
    \_ces_1_3_io_outs_left[11] ,
    \_ces_1_3_io_outs_left[10] ,
    \_ces_1_3_io_outs_left[9] ,
    \_ces_1_3_io_outs_left[8] ,
    \_ces_1_3_io_outs_left[7] ,
    \_ces_1_3_io_outs_left[6] ,
    \_ces_1_3_io_outs_left[5] ,
    \_ces_1_3_io_outs_left[4] ,
    \_ces_1_3_io_outs_left[3] ,
    \_ces_1_3_io_outs_left[2] ,
    \_ces_1_3_io_outs_left[1] ,
    \_ces_1_3_io_outs_left[0] }),
    .io_ins_right({\_ces_1_1_io_outs_right[63] ,
    \_ces_1_1_io_outs_right[62] ,
    \_ces_1_1_io_outs_right[61] ,
    \_ces_1_1_io_outs_right[60] ,
    \_ces_1_1_io_outs_right[59] ,
    \_ces_1_1_io_outs_right[58] ,
    \_ces_1_1_io_outs_right[57] ,
    \_ces_1_1_io_outs_right[56] ,
    \_ces_1_1_io_outs_right[55] ,
    \_ces_1_1_io_outs_right[54] ,
    \_ces_1_1_io_outs_right[53] ,
    \_ces_1_1_io_outs_right[52] ,
    \_ces_1_1_io_outs_right[51] ,
    \_ces_1_1_io_outs_right[50] ,
    \_ces_1_1_io_outs_right[49] ,
    \_ces_1_1_io_outs_right[48] ,
    \_ces_1_1_io_outs_right[47] ,
    \_ces_1_1_io_outs_right[46] ,
    \_ces_1_1_io_outs_right[45] ,
    \_ces_1_1_io_outs_right[44] ,
    \_ces_1_1_io_outs_right[43] ,
    \_ces_1_1_io_outs_right[42] ,
    \_ces_1_1_io_outs_right[41] ,
    \_ces_1_1_io_outs_right[40] ,
    \_ces_1_1_io_outs_right[39] ,
    \_ces_1_1_io_outs_right[38] ,
    \_ces_1_1_io_outs_right[37] ,
    \_ces_1_1_io_outs_right[36] ,
    \_ces_1_1_io_outs_right[35] ,
    \_ces_1_1_io_outs_right[34] ,
    \_ces_1_1_io_outs_right[33] ,
    \_ces_1_1_io_outs_right[32] ,
    \_ces_1_1_io_outs_right[31] ,
    \_ces_1_1_io_outs_right[30] ,
    \_ces_1_1_io_outs_right[29] ,
    \_ces_1_1_io_outs_right[28] ,
    \_ces_1_1_io_outs_right[27] ,
    \_ces_1_1_io_outs_right[26] ,
    \_ces_1_1_io_outs_right[25] ,
    \_ces_1_1_io_outs_right[24] ,
    \_ces_1_1_io_outs_right[23] ,
    \_ces_1_1_io_outs_right[22] ,
    \_ces_1_1_io_outs_right[21] ,
    \_ces_1_1_io_outs_right[20] ,
    \_ces_1_1_io_outs_right[19] ,
    \_ces_1_1_io_outs_right[18] ,
    \_ces_1_1_io_outs_right[17] ,
    \_ces_1_1_io_outs_right[16] ,
    \_ces_1_1_io_outs_right[15] ,
    \_ces_1_1_io_outs_right[14] ,
    \_ces_1_1_io_outs_right[13] ,
    \_ces_1_1_io_outs_right[12] ,
    \_ces_1_1_io_outs_right[11] ,
    \_ces_1_1_io_outs_right[10] ,
    \_ces_1_1_io_outs_right[9] ,
    \_ces_1_1_io_outs_right[8] ,
    \_ces_1_1_io_outs_right[7] ,
    \_ces_1_1_io_outs_right[6] ,
    \_ces_1_1_io_outs_right[5] ,
    \_ces_1_1_io_outs_right[4] ,
    \_ces_1_1_io_outs_right[3] ,
    \_ces_1_1_io_outs_right[2] ,
    \_ces_1_1_io_outs_right[1] ,
    \_ces_1_1_io_outs_right[0] }),
    .io_ins_up({\_ces_0_2_io_outs_up[63] ,
    \_ces_0_2_io_outs_up[62] ,
    \_ces_0_2_io_outs_up[61] ,
    \_ces_0_2_io_outs_up[60] ,
    \_ces_0_2_io_outs_up[59] ,
    \_ces_0_2_io_outs_up[58] ,
    \_ces_0_2_io_outs_up[57] ,
    \_ces_0_2_io_outs_up[56] ,
    \_ces_0_2_io_outs_up[55] ,
    \_ces_0_2_io_outs_up[54] ,
    \_ces_0_2_io_outs_up[53] ,
    \_ces_0_2_io_outs_up[52] ,
    \_ces_0_2_io_outs_up[51] ,
    \_ces_0_2_io_outs_up[50] ,
    \_ces_0_2_io_outs_up[49] ,
    \_ces_0_2_io_outs_up[48] ,
    \_ces_0_2_io_outs_up[47] ,
    \_ces_0_2_io_outs_up[46] ,
    \_ces_0_2_io_outs_up[45] ,
    \_ces_0_2_io_outs_up[44] ,
    \_ces_0_2_io_outs_up[43] ,
    \_ces_0_2_io_outs_up[42] ,
    \_ces_0_2_io_outs_up[41] ,
    \_ces_0_2_io_outs_up[40] ,
    \_ces_0_2_io_outs_up[39] ,
    \_ces_0_2_io_outs_up[38] ,
    \_ces_0_2_io_outs_up[37] ,
    \_ces_0_2_io_outs_up[36] ,
    \_ces_0_2_io_outs_up[35] ,
    \_ces_0_2_io_outs_up[34] ,
    \_ces_0_2_io_outs_up[33] ,
    \_ces_0_2_io_outs_up[32] ,
    \_ces_0_2_io_outs_up[31] ,
    \_ces_0_2_io_outs_up[30] ,
    \_ces_0_2_io_outs_up[29] ,
    \_ces_0_2_io_outs_up[28] ,
    \_ces_0_2_io_outs_up[27] ,
    \_ces_0_2_io_outs_up[26] ,
    \_ces_0_2_io_outs_up[25] ,
    \_ces_0_2_io_outs_up[24] ,
    \_ces_0_2_io_outs_up[23] ,
    \_ces_0_2_io_outs_up[22] ,
    \_ces_0_2_io_outs_up[21] ,
    \_ces_0_2_io_outs_up[20] ,
    \_ces_0_2_io_outs_up[19] ,
    \_ces_0_2_io_outs_up[18] ,
    \_ces_0_2_io_outs_up[17] ,
    \_ces_0_2_io_outs_up[16] ,
    \_ces_0_2_io_outs_up[15] ,
    \_ces_0_2_io_outs_up[14] ,
    \_ces_0_2_io_outs_up[13] ,
    \_ces_0_2_io_outs_up[12] ,
    \_ces_0_2_io_outs_up[11] ,
    \_ces_0_2_io_outs_up[10] ,
    \_ces_0_2_io_outs_up[9] ,
    \_ces_0_2_io_outs_up[8] ,
    \_ces_0_2_io_outs_up[7] ,
    \_ces_0_2_io_outs_up[6] ,
    \_ces_0_2_io_outs_up[5] ,
    \_ces_0_2_io_outs_up[4] ,
    \_ces_0_2_io_outs_up[3] ,
    \_ces_0_2_io_outs_up[2] ,
    \_ces_0_2_io_outs_up[1] ,
    \_ces_0_2_io_outs_up[0] }),
    .io_outs_down({\_ces_1_2_io_outs_down[63] ,
    \_ces_1_2_io_outs_down[62] ,
    \_ces_1_2_io_outs_down[61] ,
    \_ces_1_2_io_outs_down[60] ,
    \_ces_1_2_io_outs_down[59] ,
    \_ces_1_2_io_outs_down[58] ,
    \_ces_1_2_io_outs_down[57] ,
    \_ces_1_2_io_outs_down[56] ,
    \_ces_1_2_io_outs_down[55] ,
    \_ces_1_2_io_outs_down[54] ,
    \_ces_1_2_io_outs_down[53] ,
    \_ces_1_2_io_outs_down[52] ,
    \_ces_1_2_io_outs_down[51] ,
    \_ces_1_2_io_outs_down[50] ,
    \_ces_1_2_io_outs_down[49] ,
    \_ces_1_2_io_outs_down[48] ,
    \_ces_1_2_io_outs_down[47] ,
    \_ces_1_2_io_outs_down[46] ,
    \_ces_1_2_io_outs_down[45] ,
    \_ces_1_2_io_outs_down[44] ,
    \_ces_1_2_io_outs_down[43] ,
    \_ces_1_2_io_outs_down[42] ,
    \_ces_1_2_io_outs_down[41] ,
    \_ces_1_2_io_outs_down[40] ,
    \_ces_1_2_io_outs_down[39] ,
    \_ces_1_2_io_outs_down[38] ,
    \_ces_1_2_io_outs_down[37] ,
    \_ces_1_2_io_outs_down[36] ,
    \_ces_1_2_io_outs_down[35] ,
    \_ces_1_2_io_outs_down[34] ,
    \_ces_1_2_io_outs_down[33] ,
    \_ces_1_2_io_outs_down[32] ,
    \_ces_1_2_io_outs_down[31] ,
    \_ces_1_2_io_outs_down[30] ,
    \_ces_1_2_io_outs_down[29] ,
    \_ces_1_2_io_outs_down[28] ,
    \_ces_1_2_io_outs_down[27] ,
    \_ces_1_2_io_outs_down[26] ,
    \_ces_1_2_io_outs_down[25] ,
    \_ces_1_2_io_outs_down[24] ,
    \_ces_1_2_io_outs_down[23] ,
    \_ces_1_2_io_outs_down[22] ,
    \_ces_1_2_io_outs_down[21] ,
    \_ces_1_2_io_outs_down[20] ,
    \_ces_1_2_io_outs_down[19] ,
    \_ces_1_2_io_outs_down[18] ,
    \_ces_1_2_io_outs_down[17] ,
    \_ces_1_2_io_outs_down[16] ,
    \_ces_1_2_io_outs_down[15] ,
    \_ces_1_2_io_outs_down[14] ,
    \_ces_1_2_io_outs_down[13] ,
    \_ces_1_2_io_outs_down[12] ,
    \_ces_1_2_io_outs_down[11] ,
    \_ces_1_2_io_outs_down[10] ,
    \_ces_1_2_io_outs_down[9] ,
    \_ces_1_2_io_outs_down[8] ,
    \_ces_1_2_io_outs_down[7] ,
    \_ces_1_2_io_outs_down[6] ,
    \_ces_1_2_io_outs_down[5] ,
    \_ces_1_2_io_outs_down[4] ,
    \_ces_1_2_io_outs_down[3] ,
    \_ces_1_2_io_outs_down[2] ,
    \_ces_1_2_io_outs_down[1] ,
    \_ces_1_2_io_outs_down[0] }),
    .io_outs_left({\_ces_1_2_io_outs_left[63] ,
    \_ces_1_2_io_outs_left[62] ,
    \_ces_1_2_io_outs_left[61] ,
    \_ces_1_2_io_outs_left[60] ,
    \_ces_1_2_io_outs_left[59] ,
    \_ces_1_2_io_outs_left[58] ,
    \_ces_1_2_io_outs_left[57] ,
    \_ces_1_2_io_outs_left[56] ,
    \_ces_1_2_io_outs_left[55] ,
    \_ces_1_2_io_outs_left[54] ,
    \_ces_1_2_io_outs_left[53] ,
    \_ces_1_2_io_outs_left[52] ,
    \_ces_1_2_io_outs_left[51] ,
    \_ces_1_2_io_outs_left[50] ,
    \_ces_1_2_io_outs_left[49] ,
    \_ces_1_2_io_outs_left[48] ,
    \_ces_1_2_io_outs_left[47] ,
    \_ces_1_2_io_outs_left[46] ,
    \_ces_1_2_io_outs_left[45] ,
    \_ces_1_2_io_outs_left[44] ,
    \_ces_1_2_io_outs_left[43] ,
    \_ces_1_2_io_outs_left[42] ,
    \_ces_1_2_io_outs_left[41] ,
    \_ces_1_2_io_outs_left[40] ,
    \_ces_1_2_io_outs_left[39] ,
    \_ces_1_2_io_outs_left[38] ,
    \_ces_1_2_io_outs_left[37] ,
    \_ces_1_2_io_outs_left[36] ,
    \_ces_1_2_io_outs_left[35] ,
    \_ces_1_2_io_outs_left[34] ,
    \_ces_1_2_io_outs_left[33] ,
    \_ces_1_2_io_outs_left[32] ,
    \_ces_1_2_io_outs_left[31] ,
    \_ces_1_2_io_outs_left[30] ,
    \_ces_1_2_io_outs_left[29] ,
    \_ces_1_2_io_outs_left[28] ,
    \_ces_1_2_io_outs_left[27] ,
    \_ces_1_2_io_outs_left[26] ,
    \_ces_1_2_io_outs_left[25] ,
    \_ces_1_2_io_outs_left[24] ,
    \_ces_1_2_io_outs_left[23] ,
    \_ces_1_2_io_outs_left[22] ,
    \_ces_1_2_io_outs_left[21] ,
    \_ces_1_2_io_outs_left[20] ,
    \_ces_1_2_io_outs_left[19] ,
    \_ces_1_2_io_outs_left[18] ,
    \_ces_1_2_io_outs_left[17] ,
    \_ces_1_2_io_outs_left[16] ,
    \_ces_1_2_io_outs_left[15] ,
    \_ces_1_2_io_outs_left[14] ,
    \_ces_1_2_io_outs_left[13] ,
    \_ces_1_2_io_outs_left[12] ,
    \_ces_1_2_io_outs_left[11] ,
    \_ces_1_2_io_outs_left[10] ,
    \_ces_1_2_io_outs_left[9] ,
    \_ces_1_2_io_outs_left[8] ,
    \_ces_1_2_io_outs_left[7] ,
    \_ces_1_2_io_outs_left[6] ,
    \_ces_1_2_io_outs_left[5] ,
    \_ces_1_2_io_outs_left[4] ,
    \_ces_1_2_io_outs_left[3] ,
    \_ces_1_2_io_outs_left[2] ,
    \_ces_1_2_io_outs_left[1] ,
    \_ces_1_2_io_outs_left[0] }),
    .io_outs_right({\_ces_1_2_io_outs_right[63] ,
    \_ces_1_2_io_outs_right[62] ,
    \_ces_1_2_io_outs_right[61] ,
    \_ces_1_2_io_outs_right[60] ,
    \_ces_1_2_io_outs_right[59] ,
    \_ces_1_2_io_outs_right[58] ,
    \_ces_1_2_io_outs_right[57] ,
    \_ces_1_2_io_outs_right[56] ,
    \_ces_1_2_io_outs_right[55] ,
    \_ces_1_2_io_outs_right[54] ,
    \_ces_1_2_io_outs_right[53] ,
    \_ces_1_2_io_outs_right[52] ,
    \_ces_1_2_io_outs_right[51] ,
    \_ces_1_2_io_outs_right[50] ,
    \_ces_1_2_io_outs_right[49] ,
    \_ces_1_2_io_outs_right[48] ,
    \_ces_1_2_io_outs_right[47] ,
    \_ces_1_2_io_outs_right[46] ,
    \_ces_1_2_io_outs_right[45] ,
    \_ces_1_2_io_outs_right[44] ,
    \_ces_1_2_io_outs_right[43] ,
    \_ces_1_2_io_outs_right[42] ,
    \_ces_1_2_io_outs_right[41] ,
    \_ces_1_2_io_outs_right[40] ,
    \_ces_1_2_io_outs_right[39] ,
    \_ces_1_2_io_outs_right[38] ,
    \_ces_1_2_io_outs_right[37] ,
    \_ces_1_2_io_outs_right[36] ,
    \_ces_1_2_io_outs_right[35] ,
    \_ces_1_2_io_outs_right[34] ,
    \_ces_1_2_io_outs_right[33] ,
    \_ces_1_2_io_outs_right[32] ,
    \_ces_1_2_io_outs_right[31] ,
    \_ces_1_2_io_outs_right[30] ,
    \_ces_1_2_io_outs_right[29] ,
    \_ces_1_2_io_outs_right[28] ,
    \_ces_1_2_io_outs_right[27] ,
    \_ces_1_2_io_outs_right[26] ,
    \_ces_1_2_io_outs_right[25] ,
    \_ces_1_2_io_outs_right[24] ,
    \_ces_1_2_io_outs_right[23] ,
    \_ces_1_2_io_outs_right[22] ,
    \_ces_1_2_io_outs_right[21] ,
    \_ces_1_2_io_outs_right[20] ,
    \_ces_1_2_io_outs_right[19] ,
    \_ces_1_2_io_outs_right[18] ,
    \_ces_1_2_io_outs_right[17] ,
    \_ces_1_2_io_outs_right[16] ,
    \_ces_1_2_io_outs_right[15] ,
    \_ces_1_2_io_outs_right[14] ,
    \_ces_1_2_io_outs_right[13] ,
    \_ces_1_2_io_outs_right[12] ,
    \_ces_1_2_io_outs_right[11] ,
    \_ces_1_2_io_outs_right[10] ,
    \_ces_1_2_io_outs_right[9] ,
    \_ces_1_2_io_outs_right[8] ,
    \_ces_1_2_io_outs_right[7] ,
    \_ces_1_2_io_outs_right[6] ,
    \_ces_1_2_io_outs_right[5] ,
    \_ces_1_2_io_outs_right[4] ,
    \_ces_1_2_io_outs_right[3] ,
    \_ces_1_2_io_outs_right[2] ,
    \_ces_1_2_io_outs_right[1] ,
    \_ces_1_2_io_outs_right[0] }),
    .io_outs_up({\_ces_1_2_io_outs_up[63] ,
    \_ces_1_2_io_outs_up[62] ,
    \_ces_1_2_io_outs_up[61] ,
    \_ces_1_2_io_outs_up[60] ,
    \_ces_1_2_io_outs_up[59] ,
    \_ces_1_2_io_outs_up[58] ,
    \_ces_1_2_io_outs_up[57] ,
    \_ces_1_2_io_outs_up[56] ,
    \_ces_1_2_io_outs_up[55] ,
    \_ces_1_2_io_outs_up[54] ,
    \_ces_1_2_io_outs_up[53] ,
    \_ces_1_2_io_outs_up[52] ,
    \_ces_1_2_io_outs_up[51] ,
    \_ces_1_2_io_outs_up[50] ,
    \_ces_1_2_io_outs_up[49] ,
    \_ces_1_2_io_outs_up[48] ,
    \_ces_1_2_io_outs_up[47] ,
    \_ces_1_2_io_outs_up[46] ,
    \_ces_1_2_io_outs_up[45] ,
    \_ces_1_2_io_outs_up[44] ,
    \_ces_1_2_io_outs_up[43] ,
    \_ces_1_2_io_outs_up[42] ,
    \_ces_1_2_io_outs_up[41] ,
    \_ces_1_2_io_outs_up[40] ,
    \_ces_1_2_io_outs_up[39] ,
    \_ces_1_2_io_outs_up[38] ,
    \_ces_1_2_io_outs_up[37] ,
    \_ces_1_2_io_outs_up[36] ,
    \_ces_1_2_io_outs_up[35] ,
    \_ces_1_2_io_outs_up[34] ,
    \_ces_1_2_io_outs_up[33] ,
    \_ces_1_2_io_outs_up[32] ,
    \_ces_1_2_io_outs_up[31] ,
    \_ces_1_2_io_outs_up[30] ,
    \_ces_1_2_io_outs_up[29] ,
    \_ces_1_2_io_outs_up[28] ,
    \_ces_1_2_io_outs_up[27] ,
    \_ces_1_2_io_outs_up[26] ,
    \_ces_1_2_io_outs_up[25] ,
    \_ces_1_2_io_outs_up[24] ,
    \_ces_1_2_io_outs_up[23] ,
    \_ces_1_2_io_outs_up[22] ,
    \_ces_1_2_io_outs_up[21] ,
    \_ces_1_2_io_outs_up[20] ,
    \_ces_1_2_io_outs_up[19] ,
    \_ces_1_2_io_outs_up[18] ,
    \_ces_1_2_io_outs_up[17] ,
    \_ces_1_2_io_outs_up[16] ,
    \_ces_1_2_io_outs_up[15] ,
    \_ces_1_2_io_outs_up[14] ,
    \_ces_1_2_io_outs_up[13] ,
    \_ces_1_2_io_outs_up[12] ,
    \_ces_1_2_io_outs_up[11] ,
    \_ces_1_2_io_outs_up[10] ,
    \_ces_1_2_io_outs_up[9] ,
    \_ces_1_2_io_outs_up[8] ,
    \_ces_1_2_io_outs_up[7] ,
    \_ces_1_2_io_outs_up[6] ,
    \_ces_1_2_io_outs_up[5] ,
    \_ces_1_2_io_outs_up[4] ,
    \_ces_1_2_io_outs_up[3] ,
    \_ces_1_2_io_outs_up[2] ,
    \_ces_1_2_io_outs_up[1] ,
    \_ces_1_2_io_outs_up[0] }));
 Element ces_1_3 (.clock(clknet_leaf_2_clock),
    .io_lsbIns_1(_ces_1_2_io_lsbOuts_1),
    .io_lsbIns_2(_ces_1_2_io_lsbOuts_2),
    .io_lsbIns_3(_ces_1_2_io_lsbOuts_3),
    .io_lsbOuts_0(_ces_1_3_io_lsbOuts_0),
    .io_lsbOuts_1(_ces_1_3_io_lsbOuts_1),
    .io_lsbOuts_2(_ces_1_3_io_lsbOuts_2),
    .io_lsbOuts_3(_ces_1_3_io_lsbOuts_3),
    .io_ins_down({\_ces_2_3_io_outs_down[63] ,
    \_ces_2_3_io_outs_down[62] ,
    \_ces_2_3_io_outs_down[61] ,
    \_ces_2_3_io_outs_down[60] ,
    \_ces_2_3_io_outs_down[59] ,
    \_ces_2_3_io_outs_down[58] ,
    \_ces_2_3_io_outs_down[57] ,
    \_ces_2_3_io_outs_down[56] ,
    \_ces_2_3_io_outs_down[55] ,
    \_ces_2_3_io_outs_down[54] ,
    \_ces_2_3_io_outs_down[53] ,
    \_ces_2_3_io_outs_down[52] ,
    \_ces_2_3_io_outs_down[51] ,
    \_ces_2_3_io_outs_down[50] ,
    \_ces_2_3_io_outs_down[49] ,
    \_ces_2_3_io_outs_down[48] ,
    \_ces_2_3_io_outs_down[47] ,
    \_ces_2_3_io_outs_down[46] ,
    \_ces_2_3_io_outs_down[45] ,
    \_ces_2_3_io_outs_down[44] ,
    \_ces_2_3_io_outs_down[43] ,
    \_ces_2_3_io_outs_down[42] ,
    \_ces_2_3_io_outs_down[41] ,
    \_ces_2_3_io_outs_down[40] ,
    \_ces_2_3_io_outs_down[39] ,
    \_ces_2_3_io_outs_down[38] ,
    \_ces_2_3_io_outs_down[37] ,
    \_ces_2_3_io_outs_down[36] ,
    \_ces_2_3_io_outs_down[35] ,
    \_ces_2_3_io_outs_down[34] ,
    \_ces_2_3_io_outs_down[33] ,
    \_ces_2_3_io_outs_down[32] ,
    \_ces_2_3_io_outs_down[31] ,
    \_ces_2_3_io_outs_down[30] ,
    \_ces_2_3_io_outs_down[29] ,
    \_ces_2_3_io_outs_down[28] ,
    \_ces_2_3_io_outs_down[27] ,
    \_ces_2_3_io_outs_down[26] ,
    \_ces_2_3_io_outs_down[25] ,
    \_ces_2_3_io_outs_down[24] ,
    \_ces_2_3_io_outs_down[23] ,
    \_ces_2_3_io_outs_down[22] ,
    \_ces_2_3_io_outs_down[21] ,
    \_ces_2_3_io_outs_down[20] ,
    \_ces_2_3_io_outs_down[19] ,
    \_ces_2_3_io_outs_down[18] ,
    \_ces_2_3_io_outs_down[17] ,
    \_ces_2_3_io_outs_down[16] ,
    \_ces_2_3_io_outs_down[15] ,
    \_ces_2_3_io_outs_down[14] ,
    \_ces_2_3_io_outs_down[13] ,
    \_ces_2_3_io_outs_down[12] ,
    \_ces_2_3_io_outs_down[11] ,
    \_ces_2_3_io_outs_down[10] ,
    \_ces_2_3_io_outs_down[9] ,
    \_ces_2_3_io_outs_down[8] ,
    \_ces_2_3_io_outs_down[7] ,
    \_ces_2_3_io_outs_down[6] ,
    \_ces_2_3_io_outs_down[5] ,
    \_ces_2_3_io_outs_down[4] ,
    \_ces_2_3_io_outs_down[3] ,
    \_ces_2_3_io_outs_down[2] ,
    \_ces_2_3_io_outs_down[1] ,
    \_ces_2_3_io_outs_down[0] }),
    .io_ins_left({net391,
    net390,
    net389,
    net388,
    net386,
    net385,
    net384,
    net383,
    net382,
    net381,
    net380,
    net379,
    net378,
    net377,
    net375,
    net374,
    net373,
    net372,
    net371,
    net370,
    net369,
    net368,
    net367,
    net366,
    net364,
    net363,
    net362,
    net361,
    net360,
    net359,
    net358,
    net357,
    net356,
    net355,
    net353,
    net352,
    net351,
    net350,
    net349,
    net348,
    net347,
    net346,
    net345,
    net344,
    net342,
    net341,
    net340,
    net339,
    net338,
    net337,
    net336,
    net335,
    net334,
    net333,
    net395,
    net394,
    net393,
    net392,
    net387,
    net376,
    net365,
    net354,
    net343,
    net332}),
    .io_ins_right({\_ces_1_2_io_outs_right[63] ,
    \_ces_1_2_io_outs_right[62] ,
    \_ces_1_2_io_outs_right[61] ,
    \_ces_1_2_io_outs_right[60] ,
    \_ces_1_2_io_outs_right[59] ,
    \_ces_1_2_io_outs_right[58] ,
    \_ces_1_2_io_outs_right[57] ,
    \_ces_1_2_io_outs_right[56] ,
    \_ces_1_2_io_outs_right[55] ,
    \_ces_1_2_io_outs_right[54] ,
    \_ces_1_2_io_outs_right[53] ,
    \_ces_1_2_io_outs_right[52] ,
    \_ces_1_2_io_outs_right[51] ,
    \_ces_1_2_io_outs_right[50] ,
    \_ces_1_2_io_outs_right[49] ,
    \_ces_1_2_io_outs_right[48] ,
    \_ces_1_2_io_outs_right[47] ,
    \_ces_1_2_io_outs_right[46] ,
    \_ces_1_2_io_outs_right[45] ,
    \_ces_1_2_io_outs_right[44] ,
    \_ces_1_2_io_outs_right[43] ,
    \_ces_1_2_io_outs_right[42] ,
    \_ces_1_2_io_outs_right[41] ,
    \_ces_1_2_io_outs_right[40] ,
    \_ces_1_2_io_outs_right[39] ,
    \_ces_1_2_io_outs_right[38] ,
    \_ces_1_2_io_outs_right[37] ,
    \_ces_1_2_io_outs_right[36] ,
    \_ces_1_2_io_outs_right[35] ,
    \_ces_1_2_io_outs_right[34] ,
    \_ces_1_2_io_outs_right[33] ,
    \_ces_1_2_io_outs_right[32] ,
    \_ces_1_2_io_outs_right[31] ,
    \_ces_1_2_io_outs_right[30] ,
    \_ces_1_2_io_outs_right[29] ,
    \_ces_1_2_io_outs_right[28] ,
    \_ces_1_2_io_outs_right[27] ,
    \_ces_1_2_io_outs_right[26] ,
    \_ces_1_2_io_outs_right[25] ,
    \_ces_1_2_io_outs_right[24] ,
    \_ces_1_2_io_outs_right[23] ,
    \_ces_1_2_io_outs_right[22] ,
    \_ces_1_2_io_outs_right[21] ,
    \_ces_1_2_io_outs_right[20] ,
    \_ces_1_2_io_outs_right[19] ,
    \_ces_1_2_io_outs_right[18] ,
    \_ces_1_2_io_outs_right[17] ,
    \_ces_1_2_io_outs_right[16] ,
    \_ces_1_2_io_outs_right[15] ,
    \_ces_1_2_io_outs_right[14] ,
    \_ces_1_2_io_outs_right[13] ,
    \_ces_1_2_io_outs_right[12] ,
    \_ces_1_2_io_outs_right[11] ,
    \_ces_1_2_io_outs_right[10] ,
    \_ces_1_2_io_outs_right[9] ,
    \_ces_1_2_io_outs_right[8] ,
    \_ces_1_2_io_outs_right[7] ,
    \_ces_1_2_io_outs_right[6] ,
    \_ces_1_2_io_outs_right[5] ,
    \_ces_1_2_io_outs_right[4] ,
    \_ces_1_2_io_outs_right[3] ,
    \_ces_1_2_io_outs_right[2] ,
    \_ces_1_2_io_outs_right[1] ,
    \_ces_1_2_io_outs_right[0] }),
    .io_ins_up({\_ces_0_3_io_outs_up[63] ,
    \_ces_0_3_io_outs_up[62] ,
    \_ces_0_3_io_outs_up[61] ,
    \_ces_0_3_io_outs_up[60] ,
    \_ces_0_3_io_outs_up[59] ,
    \_ces_0_3_io_outs_up[58] ,
    \_ces_0_3_io_outs_up[57] ,
    \_ces_0_3_io_outs_up[56] ,
    \_ces_0_3_io_outs_up[55] ,
    \_ces_0_3_io_outs_up[54] ,
    \_ces_0_3_io_outs_up[53] ,
    \_ces_0_3_io_outs_up[52] ,
    \_ces_0_3_io_outs_up[51] ,
    \_ces_0_3_io_outs_up[50] ,
    \_ces_0_3_io_outs_up[49] ,
    \_ces_0_3_io_outs_up[48] ,
    \_ces_0_3_io_outs_up[47] ,
    \_ces_0_3_io_outs_up[46] ,
    \_ces_0_3_io_outs_up[45] ,
    \_ces_0_3_io_outs_up[44] ,
    \_ces_0_3_io_outs_up[43] ,
    \_ces_0_3_io_outs_up[42] ,
    \_ces_0_3_io_outs_up[41] ,
    \_ces_0_3_io_outs_up[40] ,
    \_ces_0_3_io_outs_up[39] ,
    \_ces_0_3_io_outs_up[38] ,
    \_ces_0_3_io_outs_up[37] ,
    \_ces_0_3_io_outs_up[36] ,
    \_ces_0_3_io_outs_up[35] ,
    \_ces_0_3_io_outs_up[34] ,
    \_ces_0_3_io_outs_up[33] ,
    \_ces_0_3_io_outs_up[32] ,
    \_ces_0_3_io_outs_up[31] ,
    \_ces_0_3_io_outs_up[30] ,
    \_ces_0_3_io_outs_up[29] ,
    \_ces_0_3_io_outs_up[28] ,
    \_ces_0_3_io_outs_up[27] ,
    \_ces_0_3_io_outs_up[26] ,
    \_ces_0_3_io_outs_up[25] ,
    \_ces_0_3_io_outs_up[24] ,
    \_ces_0_3_io_outs_up[23] ,
    \_ces_0_3_io_outs_up[22] ,
    \_ces_0_3_io_outs_up[21] ,
    \_ces_0_3_io_outs_up[20] ,
    \_ces_0_3_io_outs_up[19] ,
    \_ces_0_3_io_outs_up[18] ,
    \_ces_0_3_io_outs_up[17] ,
    \_ces_0_3_io_outs_up[16] ,
    \_ces_0_3_io_outs_up[15] ,
    \_ces_0_3_io_outs_up[14] ,
    \_ces_0_3_io_outs_up[13] ,
    \_ces_0_3_io_outs_up[12] ,
    \_ces_0_3_io_outs_up[11] ,
    \_ces_0_3_io_outs_up[10] ,
    \_ces_0_3_io_outs_up[9] ,
    \_ces_0_3_io_outs_up[8] ,
    \_ces_0_3_io_outs_up[7] ,
    \_ces_0_3_io_outs_up[6] ,
    \_ces_0_3_io_outs_up[5] ,
    \_ces_0_3_io_outs_up[4] ,
    \_ces_0_3_io_outs_up[3] ,
    \_ces_0_3_io_outs_up[2] ,
    \_ces_0_3_io_outs_up[1] ,
    \_ces_0_3_io_outs_up[0] }),
    .io_outs_down({\_ces_1_3_io_outs_down[63] ,
    \_ces_1_3_io_outs_down[62] ,
    \_ces_1_3_io_outs_down[61] ,
    \_ces_1_3_io_outs_down[60] ,
    \_ces_1_3_io_outs_down[59] ,
    \_ces_1_3_io_outs_down[58] ,
    \_ces_1_3_io_outs_down[57] ,
    \_ces_1_3_io_outs_down[56] ,
    \_ces_1_3_io_outs_down[55] ,
    \_ces_1_3_io_outs_down[54] ,
    \_ces_1_3_io_outs_down[53] ,
    \_ces_1_3_io_outs_down[52] ,
    \_ces_1_3_io_outs_down[51] ,
    \_ces_1_3_io_outs_down[50] ,
    \_ces_1_3_io_outs_down[49] ,
    \_ces_1_3_io_outs_down[48] ,
    \_ces_1_3_io_outs_down[47] ,
    \_ces_1_3_io_outs_down[46] ,
    \_ces_1_3_io_outs_down[45] ,
    \_ces_1_3_io_outs_down[44] ,
    \_ces_1_3_io_outs_down[43] ,
    \_ces_1_3_io_outs_down[42] ,
    \_ces_1_3_io_outs_down[41] ,
    \_ces_1_3_io_outs_down[40] ,
    \_ces_1_3_io_outs_down[39] ,
    \_ces_1_3_io_outs_down[38] ,
    \_ces_1_3_io_outs_down[37] ,
    \_ces_1_3_io_outs_down[36] ,
    \_ces_1_3_io_outs_down[35] ,
    \_ces_1_3_io_outs_down[34] ,
    \_ces_1_3_io_outs_down[33] ,
    \_ces_1_3_io_outs_down[32] ,
    \_ces_1_3_io_outs_down[31] ,
    \_ces_1_3_io_outs_down[30] ,
    \_ces_1_3_io_outs_down[29] ,
    \_ces_1_3_io_outs_down[28] ,
    \_ces_1_3_io_outs_down[27] ,
    \_ces_1_3_io_outs_down[26] ,
    \_ces_1_3_io_outs_down[25] ,
    \_ces_1_3_io_outs_down[24] ,
    \_ces_1_3_io_outs_down[23] ,
    \_ces_1_3_io_outs_down[22] ,
    \_ces_1_3_io_outs_down[21] ,
    \_ces_1_3_io_outs_down[20] ,
    \_ces_1_3_io_outs_down[19] ,
    \_ces_1_3_io_outs_down[18] ,
    \_ces_1_3_io_outs_down[17] ,
    \_ces_1_3_io_outs_down[16] ,
    \_ces_1_3_io_outs_down[15] ,
    \_ces_1_3_io_outs_down[14] ,
    \_ces_1_3_io_outs_down[13] ,
    \_ces_1_3_io_outs_down[12] ,
    \_ces_1_3_io_outs_down[11] ,
    \_ces_1_3_io_outs_down[10] ,
    \_ces_1_3_io_outs_down[9] ,
    \_ces_1_3_io_outs_down[8] ,
    \_ces_1_3_io_outs_down[7] ,
    \_ces_1_3_io_outs_down[6] ,
    \_ces_1_3_io_outs_down[5] ,
    \_ces_1_3_io_outs_down[4] ,
    \_ces_1_3_io_outs_down[3] ,
    \_ces_1_3_io_outs_down[2] ,
    \_ces_1_3_io_outs_down[1] ,
    \_ces_1_3_io_outs_down[0] }),
    .io_outs_left({\_ces_1_3_io_outs_left[63] ,
    \_ces_1_3_io_outs_left[62] ,
    \_ces_1_3_io_outs_left[61] ,
    \_ces_1_3_io_outs_left[60] ,
    \_ces_1_3_io_outs_left[59] ,
    \_ces_1_3_io_outs_left[58] ,
    \_ces_1_3_io_outs_left[57] ,
    \_ces_1_3_io_outs_left[56] ,
    \_ces_1_3_io_outs_left[55] ,
    \_ces_1_3_io_outs_left[54] ,
    \_ces_1_3_io_outs_left[53] ,
    \_ces_1_3_io_outs_left[52] ,
    \_ces_1_3_io_outs_left[51] ,
    \_ces_1_3_io_outs_left[50] ,
    \_ces_1_3_io_outs_left[49] ,
    \_ces_1_3_io_outs_left[48] ,
    \_ces_1_3_io_outs_left[47] ,
    \_ces_1_3_io_outs_left[46] ,
    \_ces_1_3_io_outs_left[45] ,
    \_ces_1_3_io_outs_left[44] ,
    \_ces_1_3_io_outs_left[43] ,
    \_ces_1_3_io_outs_left[42] ,
    \_ces_1_3_io_outs_left[41] ,
    \_ces_1_3_io_outs_left[40] ,
    \_ces_1_3_io_outs_left[39] ,
    \_ces_1_3_io_outs_left[38] ,
    \_ces_1_3_io_outs_left[37] ,
    \_ces_1_3_io_outs_left[36] ,
    \_ces_1_3_io_outs_left[35] ,
    \_ces_1_3_io_outs_left[34] ,
    \_ces_1_3_io_outs_left[33] ,
    \_ces_1_3_io_outs_left[32] ,
    \_ces_1_3_io_outs_left[31] ,
    \_ces_1_3_io_outs_left[30] ,
    \_ces_1_3_io_outs_left[29] ,
    \_ces_1_3_io_outs_left[28] ,
    \_ces_1_3_io_outs_left[27] ,
    \_ces_1_3_io_outs_left[26] ,
    \_ces_1_3_io_outs_left[25] ,
    \_ces_1_3_io_outs_left[24] ,
    \_ces_1_3_io_outs_left[23] ,
    \_ces_1_3_io_outs_left[22] ,
    \_ces_1_3_io_outs_left[21] ,
    \_ces_1_3_io_outs_left[20] ,
    \_ces_1_3_io_outs_left[19] ,
    \_ces_1_3_io_outs_left[18] ,
    \_ces_1_3_io_outs_left[17] ,
    \_ces_1_3_io_outs_left[16] ,
    \_ces_1_3_io_outs_left[15] ,
    \_ces_1_3_io_outs_left[14] ,
    \_ces_1_3_io_outs_left[13] ,
    \_ces_1_3_io_outs_left[12] ,
    \_ces_1_3_io_outs_left[11] ,
    \_ces_1_3_io_outs_left[10] ,
    \_ces_1_3_io_outs_left[9] ,
    \_ces_1_3_io_outs_left[8] ,
    \_ces_1_3_io_outs_left[7] ,
    \_ces_1_3_io_outs_left[6] ,
    \_ces_1_3_io_outs_left[5] ,
    \_ces_1_3_io_outs_left[4] ,
    \_ces_1_3_io_outs_left[3] ,
    \_ces_1_3_io_outs_left[2] ,
    \_ces_1_3_io_outs_left[1] ,
    \_ces_1_3_io_outs_left[0] }),
    .io_outs_right({net1687,
    net1686,
    net1685,
    net1684,
    net1682,
    net1681,
    net1680,
    net1679,
    net1678,
    net1677,
    net1676,
    net1675,
    net1674,
    net1673,
    net1671,
    net1670,
    net1669,
    net1668,
    net1667,
    net1666,
    net1665,
    net1664,
    net1663,
    net1662,
    net1660,
    net1659,
    net1658,
    net1657,
    net1656,
    net1655,
    net1654,
    net1653,
    net1652,
    net1651,
    net1649,
    net1648,
    net1647,
    net1646,
    net1645,
    net1644,
    net1643,
    net1642,
    net1641,
    net1640,
    net1638,
    net1637,
    net1636,
    net1635,
    net1634,
    net1633,
    net1632,
    net1631,
    net1630,
    net1629,
    net1691,
    net1690,
    net1689,
    net1688,
    net1683,
    net1672,
    net1661,
    net1650,
    net1639,
    net1628}),
    .io_outs_up({\_ces_1_3_io_outs_up[63] ,
    \_ces_1_3_io_outs_up[62] ,
    \_ces_1_3_io_outs_up[61] ,
    \_ces_1_3_io_outs_up[60] ,
    \_ces_1_3_io_outs_up[59] ,
    \_ces_1_3_io_outs_up[58] ,
    \_ces_1_3_io_outs_up[57] ,
    \_ces_1_3_io_outs_up[56] ,
    \_ces_1_3_io_outs_up[55] ,
    \_ces_1_3_io_outs_up[54] ,
    \_ces_1_3_io_outs_up[53] ,
    \_ces_1_3_io_outs_up[52] ,
    \_ces_1_3_io_outs_up[51] ,
    \_ces_1_3_io_outs_up[50] ,
    \_ces_1_3_io_outs_up[49] ,
    \_ces_1_3_io_outs_up[48] ,
    \_ces_1_3_io_outs_up[47] ,
    \_ces_1_3_io_outs_up[46] ,
    \_ces_1_3_io_outs_up[45] ,
    \_ces_1_3_io_outs_up[44] ,
    \_ces_1_3_io_outs_up[43] ,
    \_ces_1_3_io_outs_up[42] ,
    \_ces_1_3_io_outs_up[41] ,
    \_ces_1_3_io_outs_up[40] ,
    \_ces_1_3_io_outs_up[39] ,
    \_ces_1_3_io_outs_up[38] ,
    \_ces_1_3_io_outs_up[37] ,
    \_ces_1_3_io_outs_up[36] ,
    \_ces_1_3_io_outs_up[35] ,
    \_ces_1_3_io_outs_up[34] ,
    \_ces_1_3_io_outs_up[33] ,
    \_ces_1_3_io_outs_up[32] ,
    \_ces_1_3_io_outs_up[31] ,
    \_ces_1_3_io_outs_up[30] ,
    \_ces_1_3_io_outs_up[29] ,
    \_ces_1_3_io_outs_up[28] ,
    \_ces_1_3_io_outs_up[27] ,
    \_ces_1_3_io_outs_up[26] ,
    \_ces_1_3_io_outs_up[25] ,
    \_ces_1_3_io_outs_up[24] ,
    \_ces_1_3_io_outs_up[23] ,
    \_ces_1_3_io_outs_up[22] ,
    \_ces_1_3_io_outs_up[21] ,
    \_ces_1_3_io_outs_up[20] ,
    \_ces_1_3_io_outs_up[19] ,
    \_ces_1_3_io_outs_up[18] ,
    \_ces_1_3_io_outs_up[17] ,
    \_ces_1_3_io_outs_up[16] ,
    \_ces_1_3_io_outs_up[15] ,
    \_ces_1_3_io_outs_up[14] ,
    \_ces_1_3_io_outs_up[13] ,
    \_ces_1_3_io_outs_up[12] ,
    \_ces_1_3_io_outs_up[11] ,
    \_ces_1_3_io_outs_up[10] ,
    \_ces_1_3_io_outs_up[9] ,
    \_ces_1_3_io_outs_up[8] ,
    \_ces_1_3_io_outs_up[7] ,
    \_ces_1_3_io_outs_up[6] ,
    \_ces_1_3_io_outs_up[5] ,
    \_ces_1_3_io_outs_up[4] ,
    \_ces_1_3_io_outs_up[3] ,
    \_ces_1_3_io_outs_up[2] ,
    \_ces_1_3_io_outs_up[1] ,
    \_ces_1_3_io_outs_up[0] }));
 Element ces_2_0 (.clock(clknet_leaf_0_clock),
    .io_lsbIns_1(net6),
    .io_lsbIns_2(net7),
    .io_lsbIns_3(net8),
    .io_lsbOuts_1(_ces_2_0_io_lsbOuts_1),
    .io_lsbOuts_2(_ces_2_0_io_lsbOuts_2),
    .io_lsbOuts_3(_ces_2_0_io_lsbOuts_3),
    .io_ins_down({\_ces_3_0_io_outs_down[63] ,
    \_ces_3_0_io_outs_down[62] ,
    \_ces_3_0_io_outs_down[61] ,
    \_ces_3_0_io_outs_down[60] ,
    \_ces_3_0_io_outs_down[59] ,
    \_ces_3_0_io_outs_down[58] ,
    \_ces_3_0_io_outs_down[57] ,
    \_ces_3_0_io_outs_down[56] ,
    \_ces_3_0_io_outs_down[55] ,
    \_ces_3_0_io_outs_down[54] ,
    \_ces_3_0_io_outs_down[53] ,
    \_ces_3_0_io_outs_down[52] ,
    \_ces_3_0_io_outs_down[51] ,
    \_ces_3_0_io_outs_down[50] ,
    \_ces_3_0_io_outs_down[49] ,
    \_ces_3_0_io_outs_down[48] ,
    \_ces_3_0_io_outs_down[47] ,
    \_ces_3_0_io_outs_down[46] ,
    \_ces_3_0_io_outs_down[45] ,
    \_ces_3_0_io_outs_down[44] ,
    \_ces_3_0_io_outs_down[43] ,
    \_ces_3_0_io_outs_down[42] ,
    \_ces_3_0_io_outs_down[41] ,
    \_ces_3_0_io_outs_down[40] ,
    \_ces_3_0_io_outs_down[39] ,
    \_ces_3_0_io_outs_down[38] ,
    \_ces_3_0_io_outs_down[37] ,
    \_ces_3_0_io_outs_down[36] ,
    \_ces_3_0_io_outs_down[35] ,
    \_ces_3_0_io_outs_down[34] ,
    \_ces_3_0_io_outs_down[33] ,
    \_ces_3_0_io_outs_down[32] ,
    \_ces_3_0_io_outs_down[31] ,
    \_ces_3_0_io_outs_down[30] ,
    \_ces_3_0_io_outs_down[29] ,
    \_ces_3_0_io_outs_down[28] ,
    \_ces_3_0_io_outs_down[27] ,
    \_ces_3_0_io_outs_down[26] ,
    \_ces_3_0_io_outs_down[25] ,
    \_ces_3_0_io_outs_down[24] ,
    \_ces_3_0_io_outs_down[23] ,
    \_ces_3_0_io_outs_down[22] ,
    \_ces_3_0_io_outs_down[21] ,
    \_ces_3_0_io_outs_down[20] ,
    \_ces_3_0_io_outs_down[19] ,
    \_ces_3_0_io_outs_down[18] ,
    \_ces_3_0_io_outs_down[17] ,
    \_ces_3_0_io_outs_down[16] ,
    \_ces_3_0_io_outs_down[15] ,
    \_ces_3_0_io_outs_down[14] ,
    \_ces_3_0_io_outs_down[13] ,
    \_ces_3_0_io_outs_down[12] ,
    \_ces_3_0_io_outs_down[11] ,
    \_ces_3_0_io_outs_down[10] ,
    \_ces_3_0_io_outs_down[9] ,
    \_ces_3_0_io_outs_down[8] ,
    \_ces_3_0_io_outs_down[7] ,
    \_ces_3_0_io_outs_down[6] ,
    \_ces_3_0_io_outs_down[5] ,
    \_ces_3_0_io_outs_down[4] ,
    \_ces_3_0_io_outs_down[3] ,
    \_ces_3_0_io_outs_down[2] ,
    \_ces_3_0_io_outs_down[1] ,
    \_ces_3_0_io_outs_down[0] }),
    .io_ins_left({\_ces_2_1_io_outs_left[63] ,
    \_ces_2_1_io_outs_left[62] ,
    \_ces_2_1_io_outs_left[61] ,
    \_ces_2_1_io_outs_left[60] ,
    \_ces_2_1_io_outs_left[59] ,
    \_ces_2_1_io_outs_left[58] ,
    \_ces_2_1_io_outs_left[57] ,
    \_ces_2_1_io_outs_left[56] ,
    \_ces_2_1_io_outs_left[55] ,
    \_ces_2_1_io_outs_left[54] ,
    \_ces_2_1_io_outs_left[53] ,
    \_ces_2_1_io_outs_left[52] ,
    \_ces_2_1_io_outs_left[51] ,
    \_ces_2_1_io_outs_left[50] ,
    \_ces_2_1_io_outs_left[49] ,
    \_ces_2_1_io_outs_left[48] ,
    \_ces_2_1_io_outs_left[47] ,
    \_ces_2_1_io_outs_left[46] ,
    \_ces_2_1_io_outs_left[45] ,
    \_ces_2_1_io_outs_left[44] ,
    \_ces_2_1_io_outs_left[43] ,
    \_ces_2_1_io_outs_left[42] ,
    \_ces_2_1_io_outs_left[41] ,
    \_ces_2_1_io_outs_left[40] ,
    \_ces_2_1_io_outs_left[39] ,
    \_ces_2_1_io_outs_left[38] ,
    \_ces_2_1_io_outs_left[37] ,
    \_ces_2_1_io_outs_left[36] ,
    \_ces_2_1_io_outs_left[35] ,
    \_ces_2_1_io_outs_left[34] ,
    \_ces_2_1_io_outs_left[33] ,
    \_ces_2_1_io_outs_left[32] ,
    \_ces_2_1_io_outs_left[31] ,
    \_ces_2_1_io_outs_left[30] ,
    \_ces_2_1_io_outs_left[29] ,
    \_ces_2_1_io_outs_left[28] ,
    \_ces_2_1_io_outs_left[27] ,
    \_ces_2_1_io_outs_left[26] ,
    \_ces_2_1_io_outs_left[25] ,
    \_ces_2_1_io_outs_left[24] ,
    \_ces_2_1_io_outs_left[23] ,
    \_ces_2_1_io_outs_left[22] ,
    \_ces_2_1_io_outs_left[21] ,
    \_ces_2_1_io_outs_left[20] ,
    \_ces_2_1_io_outs_left[19] ,
    \_ces_2_1_io_outs_left[18] ,
    \_ces_2_1_io_outs_left[17] ,
    \_ces_2_1_io_outs_left[16] ,
    \_ces_2_1_io_outs_left[15] ,
    \_ces_2_1_io_outs_left[14] ,
    \_ces_2_1_io_outs_left[13] ,
    \_ces_2_1_io_outs_left[12] ,
    \_ces_2_1_io_outs_left[11] ,
    \_ces_2_1_io_outs_left[10] ,
    \_ces_2_1_io_outs_left[9] ,
    \_ces_2_1_io_outs_left[8] ,
    \_ces_2_1_io_outs_left[7] ,
    \_ces_2_1_io_outs_left[6] ,
    \_ces_2_1_io_outs_left[5] ,
    \_ces_2_1_io_outs_left[4] ,
    \_ces_2_1_io_outs_left[3] ,
    \_ces_2_1_io_outs_left[2] ,
    \_ces_2_1_io_outs_left[1] ,
    \_ces_2_1_io_outs_left[0] }),
    .io_ins_right({net711,
    net710,
    net709,
    net708,
    net706,
    net705,
    net704,
    net703,
    net702,
    net701,
    net700,
    net699,
    net698,
    net697,
    net695,
    net694,
    net693,
    net692,
    net691,
    net690,
    net689,
    net688,
    net687,
    net686,
    net684,
    net683,
    net682,
    net681,
    net680,
    net679,
    net678,
    net677,
    net676,
    net675,
    net673,
    net672,
    net671,
    net670,
    net669,
    net668,
    net667,
    net666,
    net665,
    net664,
    net662,
    net661,
    net660,
    net659,
    net658,
    net657,
    net656,
    net655,
    net654,
    net653,
    net715,
    net714,
    net713,
    net712,
    net707,
    net696,
    net685,
    net674,
    net663,
    net652}),
    .io_ins_up({\_ces_1_0_io_outs_up[63] ,
    \_ces_1_0_io_outs_up[62] ,
    \_ces_1_0_io_outs_up[61] ,
    \_ces_1_0_io_outs_up[60] ,
    \_ces_1_0_io_outs_up[59] ,
    \_ces_1_0_io_outs_up[58] ,
    \_ces_1_0_io_outs_up[57] ,
    \_ces_1_0_io_outs_up[56] ,
    \_ces_1_0_io_outs_up[55] ,
    \_ces_1_0_io_outs_up[54] ,
    \_ces_1_0_io_outs_up[53] ,
    \_ces_1_0_io_outs_up[52] ,
    \_ces_1_0_io_outs_up[51] ,
    \_ces_1_0_io_outs_up[50] ,
    \_ces_1_0_io_outs_up[49] ,
    \_ces_1_0_io_outs_up[48] ,
    \_ces_1_0_io_outs_up[47] ,
    \_ces_1_0_io_outs_up[46] ,
    \_ces_1_0_io_outs_up[45] ,
    \_ces_1_0_io_outs_up[44] ,
    \_ces_1_0_io_outs_up[43] ,
    \_ces_1_0_io_outs_up[42] ,
    \_ces_1_0_io_outs_up[41] ,
    \_ces_1_0_io_outs_up[40] ,
    \_ces_1_0_io_outs_up[39] ,
    \_ces_1_0_io_outs_up[38] ,
    \_ces_1_0_io_outs_up[37] ,
    \_ces_1_0_io_outs_up[36] ,
    \_ces_1_0_io_outs_up[35] ,
    \_ces_1_0_io_outs_up[34] ,
    \_ces_1_0_io_outs_up[33] ,
    \_ces_1_0_io_outs_up[32] ,
    \_ces_1_0_io_outs_up[31] ,
    \_ces_1_0_io_outs_up[30] ,
    \_ces_1_0_io_outs_up[29] ,
    \_ces_1_0_io_outs_up[28] ,
    \_ces_1_0_io_outs_up[27] ,
    \_ces_1_0_io_outs_up[26] ,
    \_ces_1_0_io_outs_up[25] ,
    \_ces_1_0_io_outs_up[24] ,
    \_ces_1_0_io_outs_up[23] ,
    \_ces_1_0_io_outs_up[22] ,
    \_ces_1_0_io_outs_up[21] ,
    \_ces_1_0_io_outs_up[20] ,
    \_ces_1_0_io_outs_up[19] ,
    \_ces_1_0_io_outs_up[18] ,
    \_ces_1_0_io_outs_up[17] ,
    \_ces_1_0_io_outs_up[16] ,
    \_ces_1_0_io_outs_up[15] ,
    \_ces_1_0_io_outs_up[14] ,
    \_ces_1_0_io_outs_up[13] ,
    \_ces_1_0_io_outs_up[12] ,
    \_ces_1_0_io_outs_up[11] ,
    \_ces_1_0_io_outs_up[10] ,
    \_ces_1_0_io_outs_up[9] ,
    \_ces_1_0_io_outs_up[8] ,
    \_ces_1_0_io_outs_up[7] ,
    \_ces_1_0_io_outs_up[6] ,
    \_ces_1_0_io_outs_up[5] ,
    \_ces_1_0_io_outs_up[4] ,
    \_ces_1_0_io_outs_up[3] ,
    \_ces_1_0_io_outs_up[2] ,
    \_ces_1_0_io_outs_up[1] ,
    \_ces_1_0_io_outs_up[0] }),
    .io_outs_down({\_ces_2_0_io_outs_down[63] ,
    \_ces_2_0_io_outs_down[62] ,
    \_ces_2_0_io_outs_down[61] ,
    \_ces_2_0_io_outs_down[60] ,
    \_ces_2_0_io_outs_down[59] ,
    \_ces_2_0_io_outs_down[58] ,
    \_ces_2_0_io_outs_down[57] ,
    \_ces_2_0_io_outs_down[56] ,
    \_ces_2_0_io_outs_down[55] ,
    \_ces_2_0_io_outs_down[54] ,
    \_ces_2_0_io_outs_down[53] ,
    \_ces_2_0_io_outs_down[52] ,
    \_ces_2_0_io_outs_down[51] ,
    \_ces_2_0_io_outs_down[50] ,
    \_ces_2_0_io_outs_down[49] ,
    \_ces_2_0_io_outs_down[48] ,
    \_ces_2_0_io_outs_down[47] ,
    \_ces_2_0_io_outs_down[46] ,
    \_ces_2_0_io_outs_down[45] ,
    \_ces_2_0_io_outs_down[44] ,
    \_ces_2_0_io_outs_down[43] ,
    \_ces_2_0_io_outs_down[42] ,
    \_ces_2_0_io_outs_down[41] ,
    \_ces_2_0_io_outs_down[40] ,
    \_ces_2_0_io_outs_down[39] ,
    \_ces_2_0_io_outs_down[38] ,
    \_ces_2_0_io_outs_down[37] ,
    \_ces_2_0_io_outs_down[36] ,
    \_ces_2_0_io_outs_down[35] ,
    \_ces_2_0_io_outs_down[34] ,
    \_ces_2_0_io_outs_down[33] ,
    \_ces_2_0_io_outs_down[32] ,
    \_ces_2_0_io_outs_down[31] ,
    \_ces_2_0_io_outs_down[30] ,
    \_ces_2_0_io_outs_down[29] ,
    \_ces_2_0_io_outs_down[28] ,
    \_ces_2_0_io_outs_down[27] ,
    \_ces_2_0_io_outs_down[26] ,
    \_ces_2_0_io_outs_down[25] ,
    \_ces_2_0_io_outs_down[24] ,
    \_ces_2_0_io_outs_down[23] ,
    \_ces_2_0_io_outs_down[22] ,
    \_ces_2_0_io_outs_down[21] ,
    \_ces_2_0_io_outs_down[20] ,
    \_ces_2_0_io_outs_down[19] ,
    \_ces_2_0_io_outs_down[18] ,
    \_ces_2_0_io_outs_down[17] ,
    \_ces_2_0_io_outs_down[16] ,
    \_ces_2_0_io_outs_down[15] ,
    \_ces_2_0_io_outs_down[14] ,
    \_ces_2_0_io_outs_down[13] ,
    \_ces_2_0_io_outs_down[12] ,
    \_ces_2_0_io_outs_down[11] ,
    \_ces_2_0_io_outs_down[10] ,
    \_ces_2_0_io_outs_down[9] ,
    \_ces_2_0_io_outs_down[8] ,
    \_ces_2_0_io_outs_down[7] ,
    \_ces_2_0_io_outs_down[6] ,
    \_ces_2_0_io_outs_down[5] ,
    \_ces_2_0_io_outs_down[4] ,
    \_ces_2_0_io_outs_down[3] ,
    \_ces_2_0_io_outs_down[2] ,
    \_ces_2_0_io_outs_down[1] ,
    \_ces_2_0_io_outs_down[0] }),
    .io_outs_left({net1495,
    net1494,
    net1493,
    net1492,
    net1490,
    net1489,
    net1488,
    net1487,
    net1486,
    net1485,
    net1484,
    net1483,
    net1482,
    net1481,
    net1479,
    net1478,
    net1477,
    net1476,
    net1475,
    net1474,
    net1473,
    net1472,
    net1471,
    net1470,
    net1468,
    net1467,
    net1466,
    net1465,
    net1464,
    net1463,
    net1462,
    net1461,
    net1460,
    net1459,
    net1457,
    net1456,
    net1455,
    net1454,
    net1453,
    net1452,
    net1451,
    net1450,
    net1449,
    net1448,
    net1446,
    net1445,
    net1444,
    net1443,
    net1442,
    net1441,
    net1440,
    net1439,
    net1438,
    net1437,
    net1499,
    net1498,
    net1497,
    net1496,
    net1491,
    net1480,
    net1469,
    net1458,
    net1447,
    net1436}),
    .io_outs_right({\_ces_2_0_io_outs_right[63] ,
    \_ces_2_0_io_outs_right[62] ,
    \_ces_2_0_io_outs_right[61] ,
    \_ces_2_0_io_outs_right[60] ,
    \_ces_2_0_io_outs_right[59] ,
    \_ces_2_0_io_outs_right[58] ,
    \_ces_2_0_io_outs_right[57] ,
    \_ces_2_0_io_outs_right[56] ,
    \_ces_2_0_io_outs_right[55] ,
    \_ces_2_0_io_outs_right[54] ,
    \_ces_2_0_io_outs_right[53] ,
    \_ces_2_0_io_outs_right[52] ,
    \_ces_2_0_io_outs_right[51] ,
    \_ces_2_0_io_outs_right[50] ,
    \_ces_2_0_io_outs_right[49] ,
    \_ces_2_0_io_outs_right[48] ,
    \_ces_2_0_io_outs_right[47] ,
    \_ces_2_0_io_outs_right[46] ,
    \_ces_2_0_io_outs_right[45] ,
    \_ces_2_0_io_outs_right[44] ,
    \_ces_2_0_io_outs_right[43] ,
    \_ces_2_0_io_outs_right[42] ,
    \_ces_2_0_io_outs_right[41] ,
    \_ces_2_0_io_outs_right[40] ,
    \_ces_2_0_io_outs_right[39] ,
    \_ces_2_0_io_outs_right[38] ,
    \_ces_2_0_io_outs_right[37] ,
    \_ces_2_0_io_outs_right[36] ,
    \_ces_2_0_io_outs_right[35] ,
    \_ces_2_0_io_outs_right[34] ,
    \_ces_2_0_io_outs_right[33] ,
    \_ces_2_0_io_outs_right[32] ,
    \_ces_2_0_io_outs_right[31] ,
    \_ces_2_0_io_outs_right[30] ,
    \_ces_2_0_io_outs_right[29] ,
    \_ces_2_0_io_outs_right[28] ,
    \_ces_2_0_io_outs_right[27] ,
    \_ces_2_0_io_outs_right[26] ,
    \_ces_2_0_io_outs_right[25] ,
    \_ces_2_0_io_outs_right[24] ,
    \_ces_2_0_io_outs_right[23] ,
    \_ces_2_0_io_outs_right[22] ,
    \_ces_2_0_io_outs_right[21] ,
    \_ces_2_0_io_outs_right[20] ,
    \_ces_2_0_io_outs_right[19] ,
    \_ces_2_0_io_outs_right[18] ,
    \_ces_2_0_io_outs_right[17] ,
    \_ces_2_0_io_outs_right[16] ,
    \_ces_2_0_io_outs_right[15] ,
    \_ces_2_0_io_outs_right[14] ,
    \_ces_2_0_io_outs_right[13] ,
    \_ces_2_0_io_outs_right[12] ,
    \_ces_2_0_io_outs_right[11] ,
    \_ces_2_0_io_outs_right[10] ,
    \_ces_2_0_io_outs_right[9] ,
    \_ces_2_0_io_outs_right[8] ,
    \_ces_2_0_io_outs_right[7] ,
    \_ces_2_0_io_outs_right[6] ,
    \_ces_2_0_io_outs_right[5] ,
    \_ces_2_0_io_outs_right[4] ,
    \_ces_2_0_io_outs_right[3] ,
    \_ces_2_0_io_outs_right[2] ,
    \_ces_2_0_io_outs_right[1] ,
    \_ces_2_0_io_outs_right[0] }),
    .io_outs_up({\_ces_2_0_io_outs_up[63] ,
    \_ces_2_0_io_outs_up[62] ,
    \_ces_2_0_io_outs_up[61] ,
    \_ces_2_0_io_outs_up[60] ,
    \_ces_2_0_io_outs_up[59] ,
    \_ces_2_0_io_outs_up[58] ,
    \_ces_2_0_io_outs_up[57] ,
    \_ces_2_0_io_outs_up[56] ,
    \_ces_2_0_io_outs_up[55] ,
    \_ces_2_0_io_outs_up[54] ,
    \_ces_2_0_io_outs_up[53] ,
    \_ces_2_0_io_outs_up[52] ,
    \_ces_2_0_io_outs_up[51] ,
    \_ces_2_0_io_outs_up[50] ,
    \_ces_2_0_io_outs_up[49] ,
    \_ces_2_0_io_outs_up[48] ,
    \_ces_2_0_io_outs_up[47] ,
    \_ces_2_0_io_outs_up[46] ,
    \_ces_2_0_io_outs_up[45] ,
    \_ces_2_0_io_outs_up[44] ,
    \_ces_2_0_io_outs_up[43] ,
    \_ces_2_0_io_outs_up[42] ,
    \_ces_2_0_io_outs_up[41] ,
    \_ces_2_0_io_outs_up[40] ,
    \_ces_2_0_io_outs_up[39] ,
    \_ces_2_0_io_outs_up[38] ,
    \_ces_2_0_io_outs_up[37] ,
    \_ces_2_0_io_outs_up[36] ,
    \_ces_2_0_io_outs_up[35] ,
    \_ces_2_0_io_outs_up[34] ,
    \_ces_2_0_io_outs_up[33] ,
    \_ces_2_0_io_outs_up[32] ,
    \_ces_2_0_io_outs_up[31] ,
    \_ces_2_0_io_outs_up[30] ,
    \_ces_2_0_io_outs_up[29] ,
    \_ces_2_0_io_outs_up[28] ,
    \_ces_2_0_io_outs_up[27] ,
    \_ces_2_0_io_outs_up[26] ,
    \_ces_2_0_io_outs_up[25] ,
    \_ces_2_0_io_outs_up[24] ,
    \_ces_2_0_io_outs_up[23] ,
    \_ces_2_0_io_outs_up[22] ,
    \_ces_2_0_io_outs_up[21] ,
    \_ces_2_0_io_outs_up[20] ,
    \_ces_2_0_io_outs_up[19] ,
    \_ces_2_0_io_outs_up[18] ,
    \_ces_2_0_io_outs_up[17] ,
    \_ces_2_0_io_outs_up[16] ,
    \_ces_2_0_io_outs_up[15] ,
    \_ces_2_0_io_outs_up[14] ,
    \_ces_2_0_io_outs_up[13] ,
    \_ces_2_0_io_outs_up[12] ,
    \_ces_2_0_io_outs_up[11] ,
    \_ces_2_0_io_outs_up[10] ,
    \_ces_2_0_io_outs_up[9] ,
    \_ces_2_0_io_outs_up[8] ,
    \_ces_2_0_io_outs_up[7] ,
    \_ces_2_0_io_outs_up[6] ,
    \_ces_2_0_io_outs_up[5] ,
    \_ces_2_0_io_outs_up[4] ,
    \_ces_2_0_io_outs_up[3] ,
    \_ces_2_0_io_outs_up[2] ,
    \_ces_2_0_io_outs_up[1] ,
    \_ces_2_0_io_outs_up[0] }));
 Element ces_2_1 (.clock(clknet_leaf_0_clock),
    .io_lsbIns_1(_ces_2_0_io_lsbOuts_1),
    .io_lsbIns_2(_ces_2_0_io_lsbOuts_2),
    .io_lsbIns_3(_ces_2_0_io_lsbOuts_3),
    .io_lsbOuts_1(_ces_2_1_io_lsbOuts_1),
    .io_lsbOuts_2(_ces_2_1_io_lsbOuts_2),
    .io_lsbOuts_3(_ces_2_1_io_lsbOuts_3),
    .io_ins_down({\_ces_3_1_io_outs_down[63] ,
    \_ces_3_1_io_outs_down[62] ,
    \_ces_3_1_io_outs_down[61] ,
    \_ces_3_1_io_outs_down[60] ,
    \_ces_3_1_io_outs_down[59] ,
    \_ces_3_1_io_outs_down[58] ,
    \_ces_3_1_io_outs_down[57] ,
    \_ces_3_1_io_outs_down[56] ,
    \_ces_3_1_io_outs_down[55] ,
    \_ces_3_1_io_outs_down[54] ,
    \_ces_3_1_io_outs_down[53] ,
    \_ces_3_1_io_outs_down[52] ,
    \_ces_3_1_io_outs_down[51] ,
    \_ces_3_1_io_outs_down[50] ,
    \_ces_3_1_io_outs_down[49] ,
    \_ces_3_1_io_outs_down[48] ,
    \_ces_3_1_io_outs_down[47] ,
    \_ces_3_1_io_outs_down[46] ,
    \_ces_3_1_io_outs_down[45] ,
    \_ces_3_1_io_outs_down[44] ,
    \_ces_3_1_io_outs_down[43] ,
    \_ces_3_1_io_outs_down[42] ,
    \_ces_3_1_io_outs_down[41] ,
    \_ces_3_1_io_outs_down[40] ,
    \_ces_3_1_io_outs_down[39] ,
    \_ces_3_1_io_outs_down[38] ,
    \_ces_3_1_io_outs_down[37] ,
    \_ces_3_1_io_outs_down[36] ,
    \_ces_3_1_io_outs_down[35] ,
    \_ces_3_1_io_outs_down[34] ,
    \_ces_3_1_io_outs_down[33] ,
    \_ces_3_1_io_outs_down[32] ,
    \_ces_3_1_io_outs_down[31] ,
    \_ces_3_1_io_outs_down[30] ,
    \_ces_3_1_io_outs_down[29] ,
    \_ces_3_1_io_outs_down[28] ,
    \_ces_3_1_io_outs_down[27] ,
    \_ces_3_1_io_outs_down[26] ,
    \_ces_3_1_io_outs_down[25] ,
    \_ces_3_1_io_outs_down[24] ,
    \_ces_3_1_io_outs_down[23] ,
    \_ces_3_1_io_outs_down[22] ,
    \_ces_3_1_io_outs_down[21] ,
    \_ces_3_1_io_outs_down[20] ,
    \_ces_3_1_io_outs_down[19] ,
    \_ces_3_1_io_outs_down[18] ,
    \_ces_3_1_io_outs_down[17] ,
    \_ces_3_1_io_outs_down[16] ,
    \_ces_3_1_io_outs_down[15] ,
    \_ces_3_1_io_outs_down[14] ,
    \_ces_3_1_io_outs_down[13] ,
    \_ces_3_1_io_outs_down[12] ,
    \_ces_3_1_io_outs_down[11] ,
    \_ces_3_1_io_outs_down[10] ,
    \_ces_3_1_io_outs_down[9] ,
    \_ces_3_1_io_outs_down[8] ,
    \_ces_3_1_io_outs_down[7] ,
    \_ces_3_1_io_outs_down[6] ,
    \_ces_3_1_io_outs_down[5] ,
    \_ces_3_1_io_outs_down[4] ,
    \_ces_3_1_io_outs_down[3] ,
    \_ces_3_1_io_outs_down[2] ,
    \_ces_3_1_io_outs_down[1] ,
    \_ces_3_1_io_outs_down[0] }),
    .io_ins_left({\_ces_2_2_io_outs_left[63] ,
    \_ces_2_2_io_outs_left[62] ,
    \_ces_2_2_io_outs_left[61] ,
    \_ces_2_2_io_outs_left[60] ,
    \_ces_2_2_io_outs_left[59] ,
    \_ces_2_2_io_outs_left[58] ,
    \_ces_2_2_io_outs_left[57] ,
    \_ces_2_2_io_outs_left[56] ,
    \_ces_2_2_io_outs_left[55] ,
    \_ces_2_2_io_outs_left[54] ,
    \_ces_2_2_io_outs_left[53] ,
    \_ces_2_2_io_outs_left[52] ,
    \_ces_2_2_io_outs_left[51] ,
    \_ces_2_2_io_outs_left[50] ,
    \_ces_2_2_io_outs_left[49] ,
    \_ces_2_2_io_outs_left[48] ,
    \_ces_2_2_io_outs_left[47] ,
    \_ces_2_2_io_outs_left[46] ,
    \_ces_2_2_io_outs_left[45] ,
    \_ces_2_2_io_outs_left[44] ,
    \_ces_2_2_io_outs_left[43] ,
    \_ces_2_2_io_outs_left[42] ,
    \_ces_2_2_io_outs_left[41] ,
    \_ces_2_2_io_outs_left[40] ,
    \_ces_2_2_io_outs_left[39] ,
    \_ces_2_2_io_outs_left[38] ,
    \_ces_2_2_io_outs_left[37] ,
    \_ces_2_2_io_outs_left[36] ,
    \_ces_2_2_io_outs_left[35] ,
    \_ces_2_2_io_outs_left[34] ,
    \_ces_2_2_io_outs_left[33] ,
    \_ces_2_2_io_outs_left[32] ,
    \_ces_2_2_io_outs_left[31] ,
    \_ces_2_2_io_outs_left[30] ,
    \_ces_2_2_io_outs_left[29] ,
    \_ces_2_2_io_outs_left[28] ,
    \_ces_2_2_io_outs_left[27] ,
    \_ces_2_2_io_outs_left[26] ,
    \_ces_2_2_io_outs_left[25] ,
    \_ces_2_2_io_outs_left[24] ,
    \_ces_2_2_io_outs_left[23] ,
    \_ces_2_2_io_outs_left[22] ,
    \_ces_2_2_io_outs_left[21] ,
    \_ces_2_2_io_outs_left[20] ,
    \_ces_2_2_io_outs_left[19] ,
    \_ces_2_2_io_outs_left[18] ,
    \_ces_2_2_io_outs_left[17] ,
    \_ces_2_2_io_outs_left[16] ,
    \_ces_2_2_io_outs_left[15] ,
    \_ces_2_2_io_outs_left[14] ,
    \_ces_2_2_io_outs_left[13] ,
    \_ces_2_2_io_outs_left[12] ,
    \_ces_2_2_io_outs_left[11] ,
    \_ces_2_2_io_outs_left[10] ,
    \_ces_2_2_io_outs_left[9] ,
    \_ces_2_2_io_outs_left[8] ,
    \_ces_2_2_io_outs_left[7] ,
    \_ces_2_2_io_outs_left[6] ,
    \_ces_2_2_io_outs_left[5] ,
    \_ces_2_2_io_outs_left[4] ,
    \_ces_2_2_io_outs_left[3] ,
    \_ces_2_2_io_outs_left[2] ,
    \_ces_2_2_io_outs_left[1] ,
    \_ces_2_2_io_outs_left[0] }),
    .io_ins_right({\_ces_2_0_io_outs_right[63] ,
    \_ces_2_0_io_outs_right[62] ,
    \_ces_2_0_io_outs_right[61] ,
    \_ces_2_0_io_outs_right[60] ,
    \_ces_2_0_io_outs_right[59] ,
    \_ces_2_0_io_outs_right[58] ,
    \_ces_2_0_io_outs_right[57] ,
    \_ces_2_0_io_outs_right[56] ,
    \_ces_2_0_io_outs_right[55] ,
    \_ces_2_0_io_outs_right[54] ,
    \_ces_2_0_io_outs_right[53] ,
    \_ces_2_0_io_outs_right[52] ,
    \_ces_2_0_io_outs_right[51] ,
    \_ces_2_0_io_outs_right[50] ,
    \_ces_2_0_io_outs_right[49] ,
    \_ces_2_0_io_outs_right[48] ,
    \_ces_2_0_io_outs_right[47] ,
    \_ces_2_0_io_outs_right[46] ,
    \_ces_2_0_io_outs_right[45] ,
    \_ces_2_0_io_outs_right[44] ,
    \_ces_2_0_io_outs_right[43] ,
    \_ces_2_0_io_outs_right[42] ,
    \_ces_2_0_io_outs_right[41] ,
    \_ces_2_0_io_outs_right[40] ,
    \_ces_2_0_io_outs_right[39] ,
    \_ces_2_0_io_outs_right[38] ,
    \_ces_2_0_io_outs_right[37] ,
    \_ces_2_0_io_outs_right[36] ,
    \_ces_2_0_io_outs_right[35] ,
    \_ces_2_0_io_outs_right[34] ,
    \_ces_2_0_io_outs_right[33] ,
    \_ces_2_0_io_outs_right[32] ,
    \_ces_2_0_io_outs_right[31] ,
    \_ces_2_0_io_outs_right[30] ,
    \_ces_2_0_io_outs_right[29] ,
    \_ces_2_0_io_outs_right[28] ,
    \_ces_2_0_io_outs_right[27] ,
    \_ces_2_0_io_outs_right[26] ,
    \_ces_2_0_io_outs_right[25] ,
    \_ces_2_0_io_outs_right[24] ,
    \_ces_2_0_io_outs_right[23] ,
    \_ces_2_0_io_outs_right[22] ,
    \_ces_2_0_io_outs_right[21] ,
    \_ces_2_0_io_outs_right[20] ,
    \_ces_2_0_io_outs_right[19] ,
    \_ces_2_0_io_outs_right[18] ,
    \_ces_2_0_io_outs_right[17] ,
    \_ces_2_0_io_outs_right[16] ,
    \_ces_2_0_io_outs_right[15] ,
    \_ces_2_0_io_outs_right[14] ,
    \_ces_2_0_io_outs_right[13] ,
    \_ces_2_0_io_outs_right[12] ,
    \_ces_2_0_io_outs_right[11] ,
    \_ces_2_0_io_outs_right[10] ,
    \_ces_2_0_io_outs_right[9] ,
    \_ces_2_0_io_outs_right[8] ,
    \_ces_2_0_io_outs_right[7] ,
    \_ces_2_0_io_outs_right[6] ,
    \_ces_2_0_io_outs_right[5] ,
    \_ces_2_0_io_outs_right[4] ,
    \_ces_2_0_io_outs_right[3] ,
    \_ces_2_0_io_outs_right[2] ,
    \_ces_2_0_io_outs_right[1] ,
    \_ces_2_0_io_outs_right[0] }),
    .io_ins_up({\_ces_1_1_io_outs_up[63] ,
    \_ces_1_1_io_outs_up[62] ,
    \_ces_1_1_io_outs_up[61] ,
    \_ces_1_1_io_outs_up[60] ,
    \_ces_1_1_io_outs_up[59] ,
    \_ces_1_1_io_outs_up[58] ,
    \_ces_1_1_io_outs_up[57] ,
    \_ces_1_1_io_outs_up[56] ,
    \_ces_1_1_io_outs_up[55] ,
    \_ces_1_1_io_outs_up[54] ,
    \_ces_1_1_io_outs_up[53] ,
    \_ces_1_1_io_outs_up[52] ,
    \_ces_1_1_io_outs_up[51] ,
    \_ces_1_1_io_outs_up[50] ,
    \_ces_1_1_io_outs_up[49] ,
    \_ces_1_1_io_outs_up[48] ,
    \_ces_1_1_io_outs_up[47] ,
    \_ces_1_1_io_outs_up[46] ,
    \_ces_1_1_io_outs_up[45] ,
    \_ces_1_1_io_outs_up[44] ,
    \_ces_1_1_io_outs_up[43] ,
    \_ces_1_1_io_outs_up[42] ,
    \_ces_1_1_io_outs_up[41] ,
    \_ces_1_1_io_outs_up[40] ,
    \_ces_1_1_io_outs_up[39] ,
    \_ces_1_1_io_outs_up[38] ,
    \_ces_1_1_io_outs_up[37] ,
    \_ces_1_1_io_outs_up[36] ,
    \_ces_1_1_io_outs_up[35] ,
    \_ces_1_1_io_outs_up[34] ,
    \_ces_1_1_io_outs_up[33] ,
    \_ces_1_1_io_outs_up[32] ,
    \_ces_1_1_io_outs_up[31] ,
    \_ces_1_1_io_outs_up[30] ,
    \_ces_1_1_io_outs_up[29] ,
    \_ces_1_1_io_outs_up[28] ,
    \_ces_1_1_io_outs_up[27] ,
    \_ces_1_1_io_outs_up[26] ,
    \_ces_1_1_io_outs_up[25] ,
    \_ces_1_1_io_outs_up[24] ,
    \_ces_1_1_io_outs_up[23] ,
    \_ces_1_1_io_outs_up[22] ,
    \_ces_1_1_io_outs_up[21] ,
    \_ces_1_1_io_outs_up[20] ,
    \_ces_1_1_io_outs_up[19] ,
    \_ces_1_1_io_outs_up[18] ,
    \_ces_1_1_io_outs_up[17] ,
    \_ces_1_1_io_outs_up[16] ,
    \_ces_1_1_io_outs_up[15] ,
    \_ces_1_1_io_outs_up[14] ,
    \_ces_1_1_io_outs_up[13] ,
    \_ces_1_1_io_outs_up[12] ,
    \_ces_1_1_io_outs_up[11] ,
    \_ces_1_1_io_outs_up[10] ,
    \_ces_1_1_io_outs_up[9] ,
    \_ces_1_1_io_outs_up[8] ,
    \_ces_1_1_io_outs_up[7] ,
    \_ces_1_1_io_outs_up[6] ,
    \_ces_1_1_io_outs_up[5] ,
    \_ces_1_1_io_outs_up[4] ,
    \_ces_1_1_io_outs_up[3] ,
    \_ces_1_1_io_outs_up[2] ,
    \_ces_1_1_io_outs_up[1] ,
    \_ces_1_1_io_outs_up[0] }),
    .io_outs_down({\_ces_2_1_io_outs_down[63] ,
    \_ces_2_1_io_outs_down[62] ,
    \_ces_2_1_io_outs_down[61] ,
    \_ces_2_1_io_outs_down[60] ,
    \_ces_2_1_io_outs_down[59] ,
    \_ces_2_1_io_outs_down[58] ,
    \_ces_2_1_io_outs_down[57] ,
    \_ces_2_1_io_outs_down[56] ,
    \_ces_2_1_io_outs_down[55] ,
    \_ces_2_1_io_outs_down[54] ,
    \_ces_2_1_io_outs_down[53] ,
    \_ces_2_1_io_outs_down[52] ,
    \_ces_2_1_io_outs_down[51] ,
    \_ces_2_1_io_outs_down[50] ,
    \_ces_2_1_io_outs_down[49] ,
    \_ces_2_1_io_outs_down[48] ,
    \_ces_2_1_io_outs_down[47] ,
    \_ces_2_1_io_outs_down[46] ,
    \_ces_2_1_io_outs_down[45] ,
    \_ces_2_1_io_outs_down[44] ,
    \_ces_2_1_io_outs_down[43] ,
    \_ces_2_1_io_outs_down[42] ,
    \_ces_2_1_io_outs_down[41] ,
    \_ces_2_1_io_outs_down[40] ,
    \_ces_2_1_io_outs_down[39] ,
    \_ces_2_1_io_outs_down[38] ,
    \_ces_2_1_io_outs_down[37] ,
    \_ces_2_1_io_outs_down[36] ,
    \_ces_2_1_io_outs_down[35] ,
    \_ces_2_1_io_outs_down[34] ,
    \_ces_2_1_io_outs_down[33] ,
    \_ces_2_1_io_outs_down[32] ,
    \_ces_2_1_io_outs_down[31] ,
    \_ces_2_1_io_outs_down[30] ,
    \_ces_2_1_io_outs_down[29] ,
    \_ces_2_1_io_outs_down[28] ,
    \_ces_2_1_io_outs_down[27] ,
    \_ces_2_1_io_outs_down[26] ,
    \_ces_2_1_io_outs_down[25] ,
    \_ces_2_1_io_outs_down[24] ,
    \_ces_2_1_io_outs_down[23] ,
    \_ces_2_1_io_outs_down[22] ,
    \_ces_2_1_io_outs_down[21] ,
    \_ces_2_1_io_outs_down[20] ,
    \_ces_2_1_io_outs_down[19] ,
    \_ces_2_1_io_outs_down[18] ,
    \_ces_2_1_io_outs_down[17] ,
    \_ces_2_1_io_outs_down[16] ,
    \_ces_2_1_io_outs_down[15] ,
    \_ces_2_1_io_outs_down[14] ,
    \_ces_2_1_io_outs_down[13] ,
    \_ces_2_1_io_outs_down[12] ,
    \_ces_2_1_io_outs_down[11] ,
    \_ces_2_1_io_outs_down[10] ,
    \_ces_2_1_io_outs_down[9] ,
    \_ces_2_1_io_outs_down[8] ,
    \_ces_2_1_io_outs_down[7] ,
    \_ces_2_1_io_outs_down[6] ,
    \_ces_2_1_io_outs_down[5] ,
    \_ces_2_1_io_outs_down[4] ,
    \_ces_2_1_io_outs_down[3] ,
    \_ces_2_1_io_outs_down[2] ,
    \_ces_2_1_io_outs_down[1] ,
    \_ces_2_1_io_outs_down[0] }),
    .io_outs_left({\_ces_2_1_io_outs_left[63] ,
    \_ces_2_1_io_outs_left[62] ,
    \_ces_2_1_io_outs_left[61] ,
    \_ces_2_1_io_outs_left[60] ,
    \_ces_2_1_io_outs_left[59] ,
    \_ces_2_1_io_outs_left[58] ,
    \_ces_2_1_io_outs_left[57] ,
    \_ces_2_1_io_outs_left[56] ,
    \_ces_2_1_io_outs_left[55] ,
    \_ces_2_1_io_outs_left[54] ,
    \_ces_2_1_io_outs_left[53] ,
    \_ces_2_1_io_outs_left[52] ,
    \_ces_2_1_io_outs_left[51] ,
    \_ces_2_1_io_outs_left[50] ,
    \_ces_2_1_io_outs_left[49] ,
    \_ces_2_1_io_outs_left[48] ,
    \_ces_2_1_io_outs_left[47] ,
    \_ces_2_1_io_outs_left[46] ,
    \_ces_2_1_io_outs_left[45] ,
    \_ces_2_1_io_outs_left[44] ,
    \_ces_2_1_io_outs_left[43] ,
    \_ces_2_1_io_outs_left[42] ,
    \_ces_2_1_io_outs_left[41] ,
    \_ces_2_1_io_outs_left[40] ,
    \_ces_2_1_io_outs_left[39] ,
    \_ces_2_1_io_outs_left[38] ,
    \_ces_2_1_io_outs_left[37] ,
    \_ces_2_1_io_outs_left[36] ,
    \_ces_2_1_io_outs_left[35] ,
    \_ces_2_1_io_outs_left[34] ,
    \_ces_2_1_io_outs_left[33] ,
    \_ces_2_1_io_outs_left[32] ,
    \_ces_2_1_io_outs_left[31] ,
    \_ces_2_1_io_outs_left[30] ,
    \_ces_2_1_io_outs_left[29] ,
    \_ces_2_1_io_outs_left[28] ,
    \_ces_2_1_io_outs_left[27] ,
    \_ces_2_1_io_outs_left[26] ,
    \_ces_2_1_io_outs_left[25] ,
    \_ces_2_1_io_outs_left[24] ,
    \_ces_2_1_io_outs_left[23] ,
    \_ces_2_1_io_outs_left[22] ,
    \_ces_2_1_io_outs_left[21] ,
    \_ces_2_1_io_outs_left[20] ,
    \_ces_2_1_io_outs_left[19] ,
    \_ces_2_1_io_outs_left[18] ,
    \_ces_2_1_io_outs_left[17] ,
    \_ces_2_1_io_outs_left[16] ,
    \_ces_2_1_io_outs_left[15] ,
    \_ces_2_1_io_outs_left[14] ,
    \_ces_2_1_io_outs_left[13] ,
    \_ces_2_1_io_outs_left[12] ,
    \_ces_2_1_io_outs_left[11] ,
    \_ces_2_1_io_outs_left[10] ,
    \_ces_2_1_io_outs_left[9] ,
    \_ces_2_1_io_outs_left[8] ,
    \_ces_2_1_io_outs_left[7] ,
    \_ces_2_1_io_outs_left[6] ,
    \_ces_2_1_io_outs_left[5] ,
    \_ces_2_1_io_outs_left[4] ,
    \_ces_2_1_io_outs_left[3] ,
    \_ces_2_1_io_outs_left[2] ,
    \_ces_2_1_io_outs_left[1] ,
    \_ces_2_1_io_outs_left[0] }),
    .io_outs_right({\_ces_2_1_io_outs_right[63] ,
    \_ces_2_1_io_outs_right[62] ,
    \_ces_2_1_io_outs_right[61] ,
    \_ces_2_1_io_outs_right[60] ,
    \_ces_2_1_io_outs_right[59] ,
    \_ces_2_1_io_outs_right[58] ,
    \_ces_2_1_io_outs_right[57] ,
    \_ces_2_1_io_outs_right[56] ,
    \_ces_2_1_io_outs_right[55] ,
    \_ces_2_1_io_outs_right[54] ,
    \_ces_2_1_io_outs_right[53] ,
    \_ces_2_1_io_outs_right[52] ,
    \_ces_2_1_io_outs_right[51] ,
    \_ces_2_1_io_outs_right[50] ,
    \_ces_2_1_io_outs_right[49] ,
    \_ces_2_1_io_outs_right[48] ,
    \_ces_2_1_io_outs_right[47] ,
    \_ces_2_1_io_outs_right[46] ,
    \_ces_2_1_io_outs_right[45] ,
    \_ces_2_1_io_outs_right[44] ,
    \_ces_2_1_io_outs_right[43] ,
    \_ces_2_1_io_outs_right[42] ,
    \_ces_2_1_io_outs_right[41] ,
    \_ces_2_1_io_outs_right[40] ,
    \_ces_2_1_io_outs_right[39] ,
    \_ces_2_1_io_outs_right[38] ,
    \_ces_2_1_io_outs_right[37] ,
    \_ces_2_1_io_outs_right[36] ,
    \_ces_2_1_io_outs_right[35] ,
    \_ces_2_1_io_outs_right[34] ,
    \_ces_2_1_io_outs_right[33] ,
    \_ces_2_1_io_outs_right[32] ,
    \_ces_2_1_io_outs_right[31] ,
    \_ces_2_1_io_outs_right[30] ,
    \_ces_2_1_io_outs_right[29] ,
    \_ces_2_1_io_outs_right[28] ,
    \_ces_2_1_io_outs_right[27] ,
    \_ces_2_1_io_outs_right[26] ,
    \_ces_2_1_io_outs_right[25] ,
    \_ces_2_1_io_outs_right[24] ,
    \_ces_2_1_io_outs_right[23] ,
    \_ces_2_1_io_outs_right[22] ,
    \_ces_2_1_io_outs_right[21] ,
    \_ces_2_1_io_outs_right[20] ,
    \_ces_2_1_io_outs_right[19] ,
    \_ces_2_1_io_outs_right[18] ,
    \_ces_2_1_io_outs_right[17] ,
    \_ces_2_1_io_outs_right[16] ,
    \_ces_2_1_io_outs_right[15] ,
    \_ces_2_1_io_outs_right[14] ,
    \_ces_2_1_io_outs_right[13] ,
    \_ces_2_1_io_outs_right[12] ,
    \_ces_2_1_io_outs_right[11] ,
    \_ces_2_1_io_outs_right[10] ,
    \_ces_2_1_io_outs_right[9] ,
    \_ces_2_1_io_outs_right[8] ,
    \_ces_2_1_io_outs_right[7] ,
    \_ces_2_1_io_outs_right[6] ,
    \_ces_2_1_io_outs_right[5] ,
    \_ces_2_1_io_outs_right[4] ,
    \_ces_2_1_io_outs_right[3] ,
    \_ces_2_1_io_outs_right[2] ,
    \_ces_2_1_io_outs_right[1] ,
    \_ces_2_1_io_outs_right[0] }),
    .io_outs_up({\_ces_2_1_io_outs_up[63] ,
    \_ces_2_1_io_outs_up[62] ,
    \_ces_2_1_io_outs_up[61] ,
    \_ces_2_1_io_outs_up[60] ,
    \_ces_2_1_io_outs_up[59] ,
    \_ces_2_1_io_outs_up[58] ,
    \_ces_2_1_io_outs_up[57] ,
    \_ces_2_1_io_outs_up[56] ,
    \_ces_2_1_io_outs_up[55] ,
    \_ces_2_1_io_outs_up[54] ,
    \_ces_2_1_io_outs_up[53] ,
    \_ces_2_1_io_outs_up[52] ,
    \_ces_2_1_io_outs_up[51] ,
    \_ces_2_1_io_outs_up[50] ,
    \_ces_2_1_io_outs_up[49] ,
    \_ces_2_1_io_outs_up[48] ,
    \_ces_2_1_io_outs_up[47] ,
    \_ces_2_1_io_outs_up[46] ,
    \_ces_2_1_io_outs_up[45] ,
    \_ces_2_1_io_outs_up[44] ,
    \_ces_2_1_io_outs_up[43] ,
    \_ces_2_1_io_outs_up[42] ,
    \_ces_2_1_io_outs_up[41] ,
    \_ces_2_1_io_outs_up[40] ,
    \_ces_2_1_io_outs_up[39] ,
    \_ces_2_1_io_outs_up[38] ,
    \_ces_2_1_io_outs_up[37] ,
    \_ces_2_1_io_outs_up[36] ,
    \_ces_2_1_io_outs_up[35] ,
    \_ces_2_1_io_outs_up[34] ,
    \_ces_2_1_io_outs_up[33] ,
    \_ces_2_1_io_outs_up[32] ,
    \_ces_2_1_io_outs_up[31] ,
    \_ces_2_1_io_outs_up[30] ,
    \_ces_2_1_io_outs_up[29] ,
    \_ces_2_1_io_outs_up[28] ,
    \_ces_2_1_io_outs_up[27] ,
    \_ces_2_1_io_outs_up[26] ,
    \_ces_2_1_io_outs_up[25] ,
    \_ces_2_1_io_outs_up[24] ,
    \_ces_2_1_io_outs_up[23] ,
    \_ces_2_1_io_outs_up[22] ,
    \_ces_2_1_io_outs_up[21] ,
    \_ces_2_1_io_outs_up[20] ,
    \_ces_2_1_io_outs_up[19] ,
    \_ces_2_1_io_outs_up[18] ,
    \_ces_2_1_io_outs_up[17] ,
    \_ces_2_1_io_outs_up[16] ,
    \_ces_2_1_io_outs_up[15] ,
    \_ces_2_1_io_outs_up[14] ,
    \_ces_2_1_io_outs_up[13] ,
    \_ces_2_1_io_outs_up[12] ,
    \_ces_2_1_io_outs_up[11] ,
    \_ces_2_1_io_outs_up[10] ,
    \_ces_2_1_io_outs_up[9] ,
    \_ces_2_1_io_outs_up[8] ,
    \_ces_2_1_io_outs_up[7] ,
    \_ces_2_1_io_outs_up[6] ,
    \_ces_2_1_io_outs_up[5] ,
    \_ces_2_1_io_outs_up[4] ,
    \_ces_2_1_io_outs_up[3] ,
    \_ces_2_1_io_outs_up[2] ,
    \_ces_2_1_io_outs_up[1] ,
    \_ces_2_1_io_outs_up[0] }));
 Element ces_2_2 (.clock(clknet_leaf_1_clock),
    .io_lsbIns_1(_ces_2_1_io_lsbOuts_1),
    .io_lsbIns_2(_ces_2_1_io_lsbOuts_2),
    .io_lsbIns_3(_ces_2_1_io_lsbOuts_3),
    .io_lsbOuts_1(_ces_2_2_io_lsbOuts_1),
    .io_lsbOuts_2(_ces_2_2_io_lsbOuts_2),
    .io_lsbOuts_3(_ces_2_2_io_lsbOuts_3),
    .io_ins_down({\_ces_3_2_io_outs_down[63] ,
    \_ces_3_2_io_outs_down[62] ,
    \_ces_3_2_io_outs_down[61] ,
    \_ces_3_2_io_outs_down[60] ,
    \_ces_3_2_io_outs_down[59] ,
    \_ces_3_2_io_outs_down[58] ,
    \_ces_3_2_io_outs_down[57] ,
    \_ces_3_2_io_outs_down[56] ,
    \_ces_3_2_io_outs_down[55] ,
    \_ces_3_2_io_outs_down[54] ,
    \_ces_3_2_io_outs_down[53] ,
    \_ces_3_2_io_outs_down[52] ,
    \_ces_3_2_io_outs_down[51] ,
    \_ces_3_2_io_outs_down[50] ,
    \_ces_3_2_io_outs_down[49] ,
    \_ces_3_2_io_outs_down[48] ,
    \_ces_3_2_io_outs_down[47] ,
    \_ces_3_2_io_outs_down[46] ,
    \_ces_3_2_io_outs_down[45] ,
    \_ces_3_2_io_outs_down[44] ,
    \_ces_3_2_io_outs_down[43] ,
    \_ces_3_2_io_outs_down[42] ,
    \_ces_3_2_io_outs_down[41] ,
    \_ces_3_2_io_outs_down[40] ,
    \_ces_3_2_io_outs_down[39] ,
    \_ces_3_2_io_outs_down[38] ,
    \_ces_3_2_io_outs_down[37] ,
    \_ces_3_2_io_outs_down[36] ,
    \_ces_3_2_io_outs_down[35] ,
    \_ces_3_2_io_outs_down[34] ,
    \_ces_3_2_io_outs_down[33] ,
    \_ces_3_2_io_outs_down[32] ,
    \_ces_3_2_io_outs_down[31] ,
    \_ces_3_2_io_outs_down[30] ,
    \_ces_3_2_io_outs_down[29] ,
    \_ces_3_2_io_outs_down[28] ,
    \_ces_3_2_io_outs_down[27] ,
    \_ces_3_2_io_outs_down[26] ,
    \_ces_3_2_io_outs_down[25] ,
    \_ces_3_2_io_outs_down[24] ,
    \_ces_3_2_io_outs_down[23] ,
    \_ces_3_2_io_outs_down[22] ,
    \_ces_3_2_io_outs_down[21] ,
    \_ces_3_2_io_outs_down[20] ,
    \_ces_3_2_io_outs_down[19] ,
    \_ces_3_2_io_outs_down[18] ,
    \_ces_3_2_io_outs_down[17] ,
    \_ces_3_2_io_outs_down[16] ,
    \_ces_3_2_io_outs_down[15] ,
    \_ces_3_2_io_outs_down[14] ,
    \_ces_3_2_io_outs_down[13] ,
    \_ces_3_2_io_outs_down[12] ,
    \_ces_3_2_io_outs_down[11] ,
    \_ces_3_2_io_outs_down[10] ,
    \_ces_3_2_io_outs_down[9] ,
    \_ces_3_2_io_outs_down[8] ,
    \_ces_3_2_io_outs_down[7] ,
    \_ces_3_2_io_outs_down[6] ,
    \_ces_3_2_io_outs_down[5] ,
    \_ces_3_2_io_outs_down[4] ,
    \_ces_3_2_io_outs_down[3] ,
    \_ces_3_2_io_outs_down[2] ,
    \_ces_3_2_io_outs_down[1] ,
    \_ces_3_2_io_outs_down[0] }),
    .io_ins_left({\_ces_2_3_io_outs_left[63] ,
    \_ces_2_3_io_outs_left[62] ,
    \_ces_2_3_io_outs_left[61] ,
    \_ces_2_3_io_outs_left[60] ,
    \_ces_2_3_io_outs_left[59] ,
    \_ces_2_3_io_outs_left[58] ,
    \_ces_2_3_io_outs_left[57] ,
    \_ces_2_3_io_outs_left[56] ,
    \_ces_2_3_io_outs_left[55] ,
    \_ces_2_3_io_outs_left[54] ,
    \_ces_2_3_io_outs_left[53] ,
    \_ces_2_3_io_outs_left[52] ,
    \_ces_2_3_io_outs_left[51] ,
    \_ces_2_3_io_outs_left[50] ,
    \_ces_2_3_io_outs_left[49] ,
    \_ces_2_3_io_outs_left[48] ,
    \_ces_2_3_io_outs_left[47] ,
    \_ces_2_3_io_outs_left[46] ,
    \_ces_2_3_io_outs_left[45] ,
    \_ces_2_3_io_outs_left[44] ,
    \_ces_2_3_io_outs_left[43] ,
    \_ces_2_3_io_outs_left[42] ,
    \_ces_2_3_io_outs_left[41] ,
    \_ces_2_3_io_outs_left[40] ,
    \_ces_2_3_io_outs_left[39] ,
    \_ces_2_3_io_outs_left[38] ,
    \_ces_2_3_io_outs_left[37] ,
    \_ces_2_3_io_outs_left[36] ,
    \_ces_2_3_io_outs_left[35] ,
    \_ces_2_3_io_outs_left[34] ,
    \_ces_2_3_io_outs_left[33] ,
    \_ces_2_3_io_outs_left[32] ,
    \_ces_2_3_io_outs_left[31] ,
    \_ces_2_3_io_outs_left[30] ,
    \_ces_2_3_io_outs_left[29] ,
    \_ces_2_3_io_outs_left[28] ,
    \_ces_2_3_io_outs_left[27] ,
    \_ces_2_3_io_outs_left[26] ,
    \_ces_2_3_io_outs_left[25] ,
    \_ces_2_3_io_outs_left[24] ,
    \_ces_2_3_io_outs_left[23] ,
    \_ces_2_3_io_outs_left[22] ,
    \_ces_2_3_io_outs_left[21] ,
    \_ces_2_3_io_outs_left[20] ,
    \_ces_2_3_io_outs_left[19] ,
    \_ces_2_3_io_outs_left[18] ,
    \_ces_2_3_io_outs_left[17] ,
    \_ces_2_3_io_outs_left[16] ,
    \_ces_2_3_io_outs_left[15] ,
    \_ces_2_3_io_outs_left[14] ,
    \_ces_2_3_io_outs_left[13] ,
    \_ces_2_3_io_outs_left[12] ,
    \_ces_2_3_io_outs_left[11] ,
    \_ces_2_3_io_outs_left[10] ,
    \_ces_2_3_io_outs_left[9] ,
    \_ces_2_3_io_outs_left[8] ,
    \_ces_2_3_io_outs_left[7] ,
    \_ces_2_3_io_outs_left[6] ,
    \_ces_2_3_io_outs_left[5] ,
    \_ces_2_3_io_outs_left[4] ,
    \_ces_2_3_io_outs_left[3] ,
    \_ces_2_3_io_outs_left[2] ,
    \_ces_2_3_io_outs_left[1] ,
    \_ces_2_3_io_outs_left[0] }),
    .io_ins_right({\_ces_2_1_io_outs_right[63] ,
    \_ces_2_1_io_outs_right[62] ,
    \_ces_2_1_io_outs_right[61] ,
    \_ces_2_1_io_outs_right[60] ,
    \_ces_2_1_io_outs_right[59] ,
    \_ces_2_1_io_outs_right[58] ,
    \_ces_2_1_io_outs_right[57] ,
    \_ces_2_1_io_outs_right[56] ,
    \_ces_2_1_io_outs_right[55] ,
    \_ces_2_1_io_outs_right[54] ,
    \_ces_2_1_io_outs_right[53] ,
    \_ces_2_1_io_outs_right[52] ,
    \_ces_2_1_io_outs_right[51] ,
    \_ces_2_1_io_outs_right[50] ,
    \_ces_2_1_io_outs_right[49] ,
    \_ces_2_1_io_outs_right[48] ,
    \_ces_2_1_io_outs_right[47] ,
    \_ces_2_1_io_outs_right[46] ,
    \_ces_2_1_io_outs_right[45] ,
    \_ces_2_1_io_outs_right[44] ,
    \_ces_2_1_io_outs_right[43] ,
    \_ces_2_1_io_outs_right[42] ,
    \_ces_2_1_io_outs_right[41] ,
    \_ces_2_1_io_outs_right[40] ,
    \_ces_2_1_io_outs_right[39] ,
    \_ces_2_1_io_outs_right[38] ,
    \_ces_2_1_io_outs_right[37] ,
    \_ces_2_1_io_outs_right[36] ,
    \_ces_2_1_io_outs_right[35] ,
    \_ces_2_1_io_outs_right[34] ,
    \_ces_2_1_io_outs_right[33] ,
    \_ces_2_1_io_outs_right[32] ,
    \_ces_2_1_io_outs_right[31] ,
    \_ces_2_1_io_outs_right[30] ,
    \_ces_2_1_io_outs_right[29] ,
    \_ces_2_1_io_outs_right[28] ,
    \_ces_2_1_io_outs_right[27] ,
    \_ces_2_1_io_outs_right[26] ,
    \_ces_2_1_io_outs_right[25] ,
    \_ces_2_1_io_outs_right[24] ,
    \_ces_2_1_io_outs_right[23] ,
    \_ces_2_1_io_outs_right[22] ,
    \_ces_2_1_io_outs_right[21] ,
    \_ces_2_1_io_outs_right[20] ,
    \_ces_2_1_io_outs_right[19] ,
    \_ces_2_1_io_outs_right[18] ,
    \_ces_2_1_io_outs_right[17] ,
    \_ces_2_1_io_outs_right[16] ,
    \_ces_2_1_io_outs_right[15] ,
    \_ces_2_1_io_outs_right[14] ,
    \_ces_2_1_io_outs_right[13] ,
    \_ces_2_1_io_outs_right[12] ,
    \_ces_2_1_io_outs_right[11] ,
    \_ces_2_1_io_outs_right[10] ,
    \_ces_2_1_io_outs_right[9] ,
    \_ces_2_1_io_outs_right[8] ,
    \_ces_2_1_io_outs_right[7] ,
    \_ces_2_1_io_outs_right[6] ,
    \_ces_2_1_io_outs_right[5] ,
    \_ces_2_1_io_outs_right[4] ,
    \_ces_2_1_io_outs_right[3] ,
    \_ces_2_1_io_outs_right[2] ,
    \_ces_2_1_io_outs_right[1] ,
    \_ces_2_1_io_outs_right[0] }),
    .io_ins_up({\_ces_1_2_io_outs_up[63] ,
    \_ces_1_2_io_outs_up[62] ,
    \_ces_1_2_io_outs_up[61] ,
    \_ces_1_2_io_outs_up[60] ,
    \_ces_1_2_io_outs_up[59] ,
    \_ces_1_2_io_outs_up[58] ,
    \_ces_1_2_io_outs_up[57] ,
    \_ces_1_2_io_outs_up[56] ,
    \_ces_1_2_io_outs_up[55] ,
    \_ces_1_2_io_outs_up[54] ,
    \_ces_1_2_io_outs_up[53] ,
    \_ces_1_2_io_outs_up[52] ,
    \_ces_1_2_io_outs_up[51] ,
    \_ces_1_2_io_outs_up[50] ,
    \_ces_1_2_io_outs_up[49] ,
    \_ces_1_2_io_outs_up[48] ,
    \_ces_1_2_io_outs_up[47] ,
    \_ces_1_2_io_outs_up[46] ,
    \_ces_1_2_io_outs_up[45] ,
    \_ces_1_2_io_outs_up[44] ,
    \_ces_1_2_io_outs_up[43] ,
    \_ces_1_2_io_outs_up[42] ,
    \_ces_1_2_io_outs_up[41] ,
    \_ces_1_2_io_outs_up[40] ,
    \_ces_1_2_io_outs_up[39] ,
    \_ces_1_2_io_outs_up[38] ,
    \_ces_1_2_io_outs_up[37] ,
    \_ces_1_2_io_outs_up[36] ,
    \_ces_1_2_io_outs_up[35] ,
    \_ces_1_2_io_outs_up[34] ,
    \_ces_1_2_io_outs_up[33] ,
    \_ces_1_2_io_outs_up[32] ,
    \_ces_1_2_io_outs_up[31] ,
    \_ces_1_2_io_outs_up[30] ,
    \_ces_1_2_io_outs_up[29] ,
    \_ces_1_2_io_outs_up[28] ,
    \_ces_1_2_io_outs_up[27] ,
    \_ces_1_2_io_outs_up[26] ,
    \_ces_1_2_io_outs_up[25] ,
    \_ces_1_2_io_outs_up[24] ,
    \_ces_1_2_io_outs_up[23] ,
    \_ces_1_2_io_outs_up[22] ,
    \_ces_1_2_io_outs_up[21] ,
    \_ces_1_2_io_outs_up[20] ,
    \_ces_1_2_io_outs_up[19] ,
    \_ces_1_2_io_outs_up[18] ,
    \_ces_1_2_io_outs_up[17] ,
    \_ces_1_2_io_outs_up[16] ,
    \_ces_1_2_io_outs_up[15] ,
    \_ces_1_2_io_outs_up[14] ,
    \_ces_1_2_io_outs_up[13] ,
    \_ces_1_2_io_outs_up[12] ,
    \_ces_1_2_io_outs_up[11] ,
    \_ces_1_2_io_outs_up[10] ,
    \_ces_1_2_io_outs_up[9] ,
    \_ces_1_2_io_outs_up[8] ,
    \_ces_1_2_io_outs_up[7] ,
    \_ces_1_2_io_outs_up[6] ,
    \_ces_1_2_io_outs_up[5] ,
    \_ces_1_2_io_outs_up[4] ,
    \_ces_1_2_io_outs_up[3] ,
    \_ces_1_2_io_outs_up[2] ,
    \_ces_1_2_io_outs_up[1] ,
    \_ces_1_2_io_outs_up[0] }),
    .io_outs_down({\_ces_2_2_io_outs_down[63] ,
    \_ces_2_2_io_outs_down[62] ,
    \_ces_2_2_io_outs_down[61] ,
    \_ces_2_2_io_outs_down[60] ,
    \_ces_2_2_io_outs_down[59] ,
    \_ces_2_2_io_outs_down[58] ,
    \_ces_2_2_io_outs_down[57] ,
    \_ces_2_2_io_outs_down[56] ,
    \_ces_2_2_io_outs_down[55] ,
    \_ces_2_2_io_outs_down[54] ,
    \_ces_2_2_io_outs_down[53] ,
    \_ces_2_2_io_outs_down[52] ,
    \_ces_2_2_io_outs_down[51] ,
    \_ces_2_2_io_outs_down[50] ,
    \_ces_2_2_io_outs_down[49] ,
    \_ces_2_2_io_outs_down[48] ,
    \_ces_2_2_io_outs_down[47] ,
    \_ces_2_2_io_outs_down[46] ,
    \_ces_2_2_io_outs_down[45] ,
    \_ces_2_2_io_outs_down[44] ,
    \_ces_2_2_io_outs_down[43] ,
    \_ces_2_2_io_outs_down[42] ,
    \_ces_2_2_io_outs_down[41] ,
    \_ces_2_2_io_outs_down[40] ,
    \_ces_2_2_io_outs_down[39] ,
    \_ces_2_2_io_outs_down[38] ,
    \_ces_2_2_io_outs_down[37] ,
    \_ces_2_2_io_outs_down[36] ,
    \_ces_2_2_io_outs_down[35] ,
    \_ces_2_2_io_outs_down[34] ,
    \_ces_2_2_io_outs_down[33] ,
    \_ces_2_2_io_outs_down[32] ,
    \_ces_2_2_io_outs_down[31] ,
    \_ces_2_2_io_outs_down[30] ,
    \_ces_2_2_io_outs_down[29] ,
    \_ces_2_2_io_outs_down[28] ,
    \_ces_2_2_io_outs_down[27] ,
    \_ces_2_2_io_outs_down[26] ,
    \_ces_2_2_io_outs_down[25] ,
    \_ces_2_2_io_outs_down[24] ,
    \_ces_2_2_io_outs_down[23] ,
    \_ces_2_2_io_outs_down[22] ,
    \_ces_2_2_io_outs_down[21] ,
    \_ces_2_2_io_outs_down[20] ,
    \_ces_2_2_io_outs_down[19] ,
    \_ces_2_2_io_outs_down[18] ,
    \_ces_2_2_io_outs_down[17] ,
    \_ces_2_2_io_outs_down[16] ,
    \_ces_2_2_io_outs_down[15] ,
    \_ces_2_2_io_outs_down[14] ,
    \_ces_2_2_io_outs_down[13] ,
    \_ces_2_2_io_outs_down[12] ,
    \_ces_2_2_io_outs_down[11] ,
    \_ces_2_2_io_outs_down[10] ,
    \_ces_2_2_io_outs_down[9] ,
    \_ces_2_2_io_outs_down[8] ,
    \_ces_2_2_io_outs_down[7] ,
    \_ces_2_2_io_outs_down[6] ,
    \_ces_2_2_io_outs_down[5] ,
    \_ces_2_2_io_outs_down[4] ,
    \_ces_2_2_io_outs_down[3] ,
    \_ces_2_2_io_outs_down[2] ,
    \_ces_2_2_io_outs_down[1] ,
    \_ces_2_2_io_outs_down[0] }),
    .io_outs_left({\_ces_2_2_io_outs_left[63] ,
    \_ces_2_2_io_outs_left[62] ,
    \_ces_2_2_io_outs_left[61] ,
    \_ces_2_2_io_outs_left[60] ,
    \_ces_2_2_io_outs_left[59] ,
    \_ces_2_2_io_outs_left[58] ,
    \_ces_2_2_io_outs_left[57] ,
    \_ces_2_2_io_outs_left[56] ,
    \_ces_2_2_io_outs_left[55] ,
    \_ces_2_2_io_outs_left[54] ,
    \_ces_2_2_io_outs_left[53] ,
    \_ces_2_2_io_outs_left[52] ,
    \_ces_2_2_io_outs_left[51] ,
    \_ces_2_2_io_outs_left[50] ,
    \_ces_2_2_io_outs_left[49] ,
    \_ces_2_2_io_outs_left[48] ,
    \_ces_2_2_io_outs_left[47] ,
    \_ces_2_2_io_outs_left[46] ,
    \_ces_2_2_io_outs_left[45] ,
    \_ces_2_2_io_outs_left[44] ,
    \_ces_2_2_io_outs_left[43] ,
    \_ces_2_2_io_outs_left[42] ,
    \_ces_2_2_io_outs_left[41] ,
    \_ces_2_2_io_outs_left[40] ,
    \_ces_2_2_io_outs_left[39] ,
    \_ces_2_2_io_outs_left[38] ,
    \_ces_2_2_io_outs_left[37] ,
    \_ces_2_2_io_outs_left[36] ,
    \_ces_2_2_io_outs_left[35] ,
    \_ces_2_2_io_outs_left[34] ,
    \_ces_2_2_io_outs_left[33] ,
    \_ces_2_2_io_outs_left[32] ,
    \_ces_2_2_io_outs_left[31] ,
    \_ces_2_2_io_outs_left[30] ,
    \_ces_2_2_io_outs_left[29] ,
    \_ces_2_2_io_outs_left[28] ,
    \_ces_2_2_io_outs_left[27] ,
    \_ces_2_2_io_outs_left[26] ,
    \_ces_2_2_io_outs_left[25] ,
    \_ces_2_2_io_outs_left[24] ,
    \_ces_2_2_io_outs_left[23] ,
    \_ces_2_2_io_outs_left[22] ,
    \_ces_2_2_io_outs_left[21] ,
    \_ces_2_2_io_outs_left[20] ,
    \_ces_2_2_io_outs_left[19] ,
    \_ces_2_2_io_outs_left[18] ,
    \_ces_2_2_io_outs_left[17] ,
    \_ces_2_2_io_outs_left[16] ,
    \_ces_2_2_io_outs_left[15] ,
    \_ces_2_2_io_outs_left[14] ,
    \_ces_2_2_io_outs_left[13] ,
    \_ces_2_2_io_outs_left[12] ,
    \_ces_2_2_io_outs_left[11] ,
    \_ces_2_2_io_outs_left[10] ,
    \_ces_2_2_io_outs_left[9] ,
    \_ces_2_2_io_outs_left[8] ,
    \_ces_2_2_io_outs_left[7] ,
    \_ces_2_2_io_outs_left[6] ,
    \_ces_2_2_io_outs_left[5] ,
    \_ces_2_2_io_outs_left[4] ,
    \_ces_2_2_io_outs_left[3] ,
    \_ces_2_2_io_outs_left[2] ,
    \_ces_2_2_io_outs_left[1] ,
    \_ces_2_2_io_outs_left[0] }),
    .io_outs_right({\_ces_2_2_io_outs_right[63] ,
    \_ces_2_2_io_outs_right[62] ,
    \_ces_2_2_io_outs_right[61] ,
    \_ces_2_2_io_outs_right[60] ,
    \_ces_2_2_io_outs_right[59] ,
    \_ces_2_2_io_outs_right[58] ,
    \_ces_2_2_io_outs_right[57] ,
    \_ces_2_2_io_outs_right[56] ,
    \_ces_2_2_io_outs_right[55] ,
    \_ces_2_2_io_outs_right[54] ,
    \_ces_2_2_io_outs_right[53] ,
    \_ces_2_2_io_outs_right[52] ,
    \_ces_2_2_io_outs_right[51] ,
    \_ces_2_2_io_outs_right[50] ,
    \_ces_2_2_io_outs_right[49] ,
    \_ces_2_2_io_outs_right[48] ,
    \_ces_2_2_io_outs_right[47] ,
    \_ces_2_2_io_outs_right[46] ,
    \_ces_2_2_io_outs_right[45] ,
    \_ces_2_2_io_outs_right[44] ,
    \_ces_2_2_io_outs_right[43] ,
    \_ces_2_2_io_outs_right[42] ,
    \_ces_2_2_io_outs_right[41] ,
    \_ces_2_2_io_outs_right[40] ,
    \_ces_2_2_io_outs_right[39] ,
    \_ces_2_2_io_outs_right[38] ,
    \_ces_2_2_io_outs_right[37] ,
    \_ces_2_2_io_outs_right[36] ,
    \_ces_2_2_io_outs_right[35] ,
    \_ces_2_2_io_outs_right[34] ,
    \_ces_2_2_io_outs_right[33] ,
    \_ces_2_2_io_outs_right[32] ,
    \_ces_2_2_io_outs_right[31] ,
    \_ces_2_2_io_outs_right[30] ,
    \_ces_2_2_io_outs_right[29] ,
    \_ces_2_2_io_outs_right[28] ,
    \_ces_2_2_io_outs_right[27] ,
    \_ces_2_2_io_outs_right[26] ,
    \_ces_2_2_io_outs_right[25] ,
    \_ces_2_2_io_outs_right[24] ,
    \_ces_2_2_io_outs_right[23] ,
    \_ces_2_2_io_outs_right[22] ,
    \_ces_2_2_io_outs_right[21] ,
    \_ces_2_2_io_outs_right[20] ,
    \_ces_2_2_io_outs_right[19] ,
    \_ces_2_2_io_outs_right[18] ,
    \_ces_2_2_io_outs_right[17] ,
    \_ces_2_2_io_outs_right[16] ,
    \_ces_2_2_io_outs_right[15] ,
    \_ces_2_2_io_outs_right[14] ,
    \_ces_2_2_io_outs_right[13] ,
    \_ces_2_2_io_outs_right[12] ,
    \_ces_2_2_io_outs_right[11] ,
    \_ces_2_2_io_outs_right[10] ,
    \_ces_2_2_io_outs_right[9] ,
    \_ces_2_2_io_outs_right[8] ,
    \_ces_2_2_io_outs_right[7] ,
    \_ces_2_2_io_outs_right[6] ,
    \_ces_2_2_io_outs_right[5] ,
    \_ces_2_2_io_outs_right[4] ,
    \_ces_2_2_io_outs_right[3] ,
    \_ces_2_2_io_outs_right[2] ,
    \_ces_2_2_io_outs_right[1] ,
    \_ces_2_2_io_outs_right[0] }),
    .io_outs_up({\_ces_2_2_io_outs_up[63] ,
    \_ces_2_2_io_outs_up[62] ,
    \_ces_2_2_io_outs_up[61] ,
    \_ces_2_2_io_outs_up[60] ,
    \_ces_2_2_io_outs_up[59] ,
    \_ces_2_2_io_outs_up[58] ,
    \_ces_2_2_io_outs_up[57] ,
    \_ces_2_2_io_outs_up[56] ,
    \_ces_2_2_io_outs_up[55] ,
    \_ces_2_2_io_outs_up[54] ,
    \_ces_2_2_io_outs_up[53] ,
    \_ces_2_2_io_outs_up[52] ,
    \_ces_2_2_io_outs_up[51] ,
    \_ces_2_2_io_outs_up[50] ,
    \_ces_2_2_io_outs_up[49] ,
    \_ces_2_2_io_outs_up[48] ,
    \_ces_2_2_io_outs_up[47] ,
    \_ces_2_2_io_outs_up[46] ,
    \_ces_2_2_io_outs_up[45] ,
    \_ces_2_2_io_outs_up[44] ,
    \_ces_2_2_io_outs_up[43] ,
    \_ces_2_2_io_outs_up[42] ,
    \_ces_2_2_io_outs_up[41] ,
    \_ces_2_2_io_outs_up[40] ,
    \_ces_2_2_io_outs_up[39] ,
    \_ces_2_2_io_outs_up[38] ,
    \_ces_2_2_io_outs_up[37] ,
    \_ces_2_2_io_outs_up[36] ,
    \_ces_2_2_io_outs_up[35] ,
    \_ces_2_2_io_outs_up[34] ,
    \_ces_2_2_io_outs_up[33] ,
    \_ces_2_2_io_outs_up[32] ,
    \_ces_2_2_io_outs_up[31] ,
    \_ces_2_2_io_outs_up[30] ,
    \_ces_2_2_io_outs_up[29] ,
    \_ces_2_2_io_outs_up[28] ,
    \_ces_2_2_io_outs_up[27] ,
    \_ces_2_2_io_outs_up[26] ,
    \_ces_2_2_io_outs_up[25] ,
    \_ces_2_2_io_outs_up[24] ,
    \_ces_2_2_io_outs_up[23] ,
    \_ces_2_2_io_outs_up[22] ,
    \_ces_2_2_io_outs_up[21] ,
    \_ces_2_2_io_outs_up[20] ,
    \_ces_2_2_io_outs_up[19] ,
    \_ces_2_2_io_outs_up[18] ,
    \_ces_2_2_io_outs_up[17] ,
    \_ces_2_2_io_outs_up[16] ,
    \_ces_2_2_io_outs_up[15] ,
    \_ces_2_2_io_outs_up[14] ,
    \_ces_2_2_io_outs_up[13] ,
    \_ces_2_2_io_outs_up[12] ,
    \_ces_2_2_io_outs_up[11] ,
    \_ces_2_2_io_outs_up[10] ,
    \_ces_2_2_io_outs_up[9] ,
    \_ces_2_2_io_outs_up[8] ,
    \_ces_2_2_io_outs_up[7] ,
    \_ces_2_2_io_outs_up[6] ,
    \_ces_2_2_io_outs_up[5] ,
    \_ces_2_2_io_outs_up[4] ,
    \_ces_2_2_io_outs_up[3] ,
    \_ces_2_2_io_outs_up[2] ,
    \_ces_2_2_io_outs_up[1] ,
    \_ces_2_2_io_outs_up[0] }));
 Element ces_2_3 (.clock(clknet_leaf_1_clock),
    .io_lsbIns_1(_ces_2_2_io_lsbOuts_1),
    .io_lsbIns_2(_ces_2_2_io_lsbOuts_2),
    .io_lsbIns_3(_ces_2_2_io_lsbOuts_3),
    .io_lsbOuts_0(_ces_2_3_io_lsbOuts_0),
    .io_lsbOuts_1(_ces_2_3_io_lsbOuts_1),
    .io_lsbOuts_2(_ces_2_3_io_lsbOuts_2),
    .io_lsbOuts_3(_ces_2_3_io_lsbOuts_3),
    .io_ins_down({\_ces_3_3_io_outs_down[63] ,
    \_ces_3_3_io_outs_down[62] ,
    \_ces_3_3_io_outs_down[61] ,
    \_ces_3_3_io_outs_down[60] ,
    \_ces_3_3_io_outs_down[59] ,
    \_ces_3_3_io_outs_down[58] ,
    \_ces_3_3_io_outs_down[57] ,
    \_ces_3_3_io_outs_down[56] ,
    \_ces_3_3_io_outs_down[55] ,
    \_ces_3_3_io_outs_down[54] ,
    \_ces_3_3_io_outs_down[53] ,
    \_ces_3_3_io_outs_down[52] ,
    \_ces_3_3_io_outs_down[51] ,
    \_ces_3_3_io_outs_down[50] ,
    \_ces_3_3_io_outs_down[49] ,
    \_ces_3_3_io_outs_down[48] ,
    \_ces_3_3_io_outs_down[47] ,
    \_ces_3_3_io_outs_down[46] ,
    \_ces_3_3_io_outs_down[45] ,
    \_ces_3_3_io_outs_down[44] ,
    \_ces_3_3_io_outs_down[43] ,
    \_ces_3_3_io_outs_down[42] ,
    \_ces_3_3_io_outs_down[41] ,
    \_ces_3_3_io_outs_down[40] ,
    \_ces_3_3_io_outs_down[39] ,
    \_ces_3_3_io_outs_down[38] ,
    \_ces_3_3_io_outs_down[37] ,
    \_ces_3_3_io_outs_down[36] ,
    \_ces_3_3_io_outs_down[35] ,
    \_ces_3_3_io_outs_down[34] ,
    \_ces_3_3_io_outs_down[33] ,
    \_ces_3_3_io_outs_down[32] ,
    \_ces_3_3_io_outs_down[31] ,
    \_ces_3_3_io_outs_down[30] ,
    \_ces_3_3_io_outs_down[29] ,
    \_ces_3_3_io_outs_down[28] ,
    \_ces_3_3_io_outs_down[27] ,
    \_ces_3_3_io_outs_down[26] ,
    \_ces_3_3_io_outs_down[25] ,
    \_ces_3_3_io_outs_down[24] ,
    \_ces_3_3_io_outs_down[23] ,
    \_ces_3_3_io_outs_down[22] ,
    \_ces_3_3_io_outs_down[21] ,
    \_ces_3_3_io_outs_down[20] ,
    \_ces_3_3_io_outs_down[19] ,
    \_ces_3_3_io_outs_down[18] ,
    \_ces_3_3_io_outs_down[17] ,
    \_ces_3_3_io_outs_down[16] ,
    \_ces_3_3_io_outs_down[15] ,
    \_ces_3_3_io_outs_down[14] ,
    \_ces_3_3_io_outs_down[13] ,
    \_ces_3_3_io_outs_down[12] ,
    \_ces_3_3_io_outs_down[11] ,
    \_ces_3_3_io_outs_down[10] ,
    \_ces_3_3_io_outs_down[9] ,
    \_ces_3_3_io_outs_down[8] ,
    \_ces_3_3_io_outs_down[7] ,
    \_ces_3_3_io_outs_down[6] ,
    \_ces_3_3_io_outs_down[5] ,
    \_ces_3_3_io_outs_down[4] ,
    \_ces_3_3_io_outs_down[3] ,
    \_ces_3_3_io_outs_down[2] ,
    \_ces_3_3_io_outs_down[1] ,
    \_ces_3_3_io_outs_down[0] }),
    .io_ins_left({net455,
    net454,
    net453,
    net452,
    net450,
    net449,
    net448,
    net447,
    net446,
    net445,
    net444,
    net443,
    net442,
    net441,
    net439,
    net438,
    net437,
    net436,
    net435,
    net434,
    net433,
    net432,
    net431,
    net430,
    net428,
    net427,
    net426,
    net425,
    net424,
    net423,
    net422,
    net421,
    net420,
    net419,
    net417,
    net416,
    net415,
    net414,
    net413,
    net412,
    net411,
    net410,
    net409,
    net408,
    net406,
    net405,
    net404,
    net403,
    net402,
    net401,
    net400,
    net399,
    net398,
    net397,
    net459,
    net458,
    net457,
    net456,
    net451,
    net440,
    net429,
    net418,
    net407,
    net396}),
    .io_ins_right({\_ces_2_2_io_outs_right[63] ,
    \_ces_2_2_io_outs_right[62] ,
    \_ces_2_2_io_outs_right[61] ,
    \_ces_2_2_io_outs_right[60] ,
    \_ces_2_2_io_outs_right[59] ,
    \_ces_2_2_io_outs_right[58] ,
    \_ces_2_2_io_outs_right[57] ,
    \_ces_2_2_io_outs_right[56] ,
    \_ces_2_2_io_outs_right[55] ,
    \_ces_2_2_io_outs_right[54] ,
    \_ces_2_2_io_outs_right[53] ,
    \_ces_2_2_io_outs_right[52] ,
    \_ces_2_2_io_outs_right[51] ,
    \_ces_2_2_io_outs_right[50] ,
    \_ces_2_2_io_outs_right[49] ,
    \_ces_2_2_io_outs_right[48] ,
    \_ces_2_2_io_outs_right[47] ,
    \_ces_2_2_io_outs_right[46] ,
    \_ces_2_2_io_outs_right[45] ,
    \_ces_2_2_io_outs_right[44] ,
    \_ces_2_2_io_outs_right[43] ,
    \_ces_2_2_io_outs_right[42] ,
    \_ces_2_2_io_outs_right[41] ,
    \_ces_2_2_io_outs_right[40] ,
    \_ces_2_2_io_outs_right[39] ,
    \_ces_2_2_io_outs_right[38] ,
    \_ces_2_2_io_outs_right[37] ,
    \_ces_2_2_io_outs_right[36] ,
    \_ces_2_2_io_outs_right[35] ,
    \_ces_2_2_io_outs_right[34] ,
    \_ces_2_2_io_outs_right[33] ,
    \_ces_2_2_io_outs_right[32] ,
    \_ces_2_2_io_outs_right[31] ,
    \_ces_2_2_io_outs_right[30] ,
    \_ces_2_2_io_outs_right[29] ,
    \_ces_2_2_io_outs_right[28] ,
    \_ces_2_2_io_outs_right[27] ,
    \_ces_2_2_io_outs_right[26] ,
    \_ces_2_2_io_outs_right[25] ,
    \_ces_2_2_io_outs_right[24] ,
    \_ces_2_2_io_outs_right[23] ,
    \_ces_2_2_io_outs_right[22] ,
    \_ces_2_2_io_outs_right[21] ,
    \_ces_2_2_io_outs_right[20] ,
    \_ces_2_2_io_outs_right[19] ,
    \_ces_2_2_io_outs_right[18] ,
    \_ces_2_2_io_outs_right[17] ,
    \_ces_2_2_io_outs_right[16] ,
    \_ces_2_2_io_outs_right[15] ,
    \_ces_2_2_io_outs_right[14] ,
    \_ces_2_2_io_outs_right[13] ,
    \_ces_2_2_io_outs_right[12] ,
    \_ces_2_2_io_outs_right[11] ,
    \_ces_2_2_io_outs_right[10] ,
    \_ces_2_2_io_outs_right[9] ,
    \_ces_2_2_io_outs_right[8] ,
    \_ces_2_2_io_outs_right[7] ,
    \_ces_2_2_io_outs_right[6] ,
    \_ces_2_2_io_outs_right[5] ,
    \_ces_2_2_io_outs_right[4] ,
    \_ces_2_2_io_outs_right[3] ,
    \_ces_2_2_io_outs_right[2] ,
    \_ces_2_2_io_outs_right[1] ,
    \_ces_2_2_io_outs_right[0] }),
    .io_ins_up({\_ces_1_3_io_outs_up[63] ,
    \_ces_1_3_io_outs_up[62] ,
    \_ces_1_3_io_outs_up[61] ,
    \_ces_1_3_io_outs_up[60] ,
    \_ces_1_3_io_outs_up[59] ,
    \_ces_1_3_io_outs_up[58] ,
    \_ces_1_3_io_outs_up[57] ,
    \_ces_1_3_io_outs_up[56] ,
    \_ces_1_3_io_outs_up[55] ,
    \_ces_1_3_io_outs_up[54] ,
    \_ces_1_3_io_outs_up[53] ,
    \_ces_1_3_io_outs_up[52] ,
    \_ces_1_3_io_outs_up[51] ,
    \_ces_1_3_io_outs_up[50] ,
    \_ces_1_3_io_outs_up[49] ,
    \_ces_1_3_io_outs_up[48] ,
    \_ces_1_3_io_outs_up[47] ,
    \_ces_1_3_io_outs_up[46] ,
    \_ces_1_3_io_outs_up[45] ,
    \_ces_1_3_io_outs_up[44] ,
    \_ces_1_3_io_outs_up[43] ,
    \_ces_1_3_io_outs_up[42] ,
    \_ces_1_3_io_outs_up[41] ,
    \_ces_1_3_io_outs_up[40] ,
    \_ces_1_3_io_outs_up[39] ,
    \_ces_1_3_io_outs_up[38] ,
    \_ces_1_3_io_outs_up[37] ,
    \_ces_1_3_io_outs_up[36] ,
    \_ces_1_3_io_outs_up[35] ,
    \_ces_1_3_io_outs_up[34] ,
    \_ces_1_3_io_outs_up[33] ,
    \_ces_1_3_io_outs_up[32] ,
    \_ces_1_3_io_outs_up[31] ,
    \_ces_1_3_io_outs_up[30] ,
    \_ces_1_3_io_outs_up[29] ,
    \_ces_1_3_io_outs_up[28] ,
    \_ces_1_3_io_outs_up[27] ,
    \_ces_1_3_io_outs_up[26] ,
    \_ces_1_3_io_outs_up[25] ,
    \_ces_1_3_io_outs_up[24] ,
    \_ces_1_3_io_outs_up[23] ,
    \_ces_1_3_io_outs_up[22] ,
    \_ces_1_3_io_outs_up[21] ,
    \_ces_1_3_io_outs_up[20] ,
    \_ces_1_3_io_outs_up[19] ,
    \_ces_1_3_io_outs_up[18] ,
    \_ces_1_3_io_outs_up[17] ,
    \_ces_1_3_io_outs_up[16] ,
    \_ces_1_3_io_outs_up[15] ,
    \_ces_1_3_io_outs_up[14] ,
    \_ces_1_3_io_outs_up[13] ,
    \_ces_1_3_io_outs_up[12] ,
    \_ces_1_3_io_outs_up[11] ,
    \_ces_1_3_io_outs_up[10] ,
    \_ces_1_3_io_outs_up[9] ,
    \_ces_1_3_io_outs_up[8] ,
    \_ces_1_3_io_outs_up[7] ,
    \_ces_1_3_io_outs_up[6] ,
    \_ces_1_3_io_outs_up[5] ,
    \_ces_1_3_io_outs_up[4] ,
    \_ces_1_3_io_outs_up[3] ,
    \_ces_1_3_io_outs_up[2] ,
    \_ces_1_3_io_outs_up[1] ,
    \_ces_1_3_io_outs_up[0] }),
    .io_outs_down({\_ces_2_3_io_outs_down[63] ,
    \_ces_2_3_io_outs_down[62] ,
    \_ces_2_3_io_outs_down[61] ,
    \_ces_2_3_io_outs_down[60] ,
    \_ces_2_3_io_outs_down[59] ,
    \_ces_2_3_io_outs_down[58] ,
    \_ces_2_3_io_outs_down[57] ,
    \_ces_2_3_io_outs_down[56] ,
    \_ces_2_3_io_outs_down[55] ,
    \_ces_2_3_io_outs_down[54] ,
    \_ces_2_3_io_outs_down[53] ,
    \_ces_2_3_io_outs_down[52] ,
    \_ces_2_3_io_outs_down[51] ,
    \_ces_2_3_io_outs_down[50] ,
    \_ces_2_3_io_outs_down[49] ,
    \_ces_2_3_io_outs_down[48] ,
    \_ces_2_3_io_outs_down[47] ,
    \_ces_2_3_io_outs_down[46] ,
    \_ces_2_3_io_outs_down[45] ,
    \_ces_2_3_io_outs_down[44] ,
    \_ces_2_3_io_outs_down[43] ,
    \_ces_2_3_io_outs_down[42] ,
    \_ces_2_3_io_outs_down[41] ,
    \_ces_2_3_io_outs_down[40] ,
    \_ces_2_3_io_outs_down[39] ,
    \_ces_2_3_io_outs_down[38] ,
    \_ces_2_3_io_outs_down[37] ,
    \_ces_2_3_io_outs_down[36] ,
    \_ces_2_3_io_outs_down[35] ,
    \_ces_2_3_io_outs_down[34] ,
    \_ces_2_3_io_outs_down[33] ,
    \_ces_2_3_io_outs_down[32] ,
    \_ces_2_3_io_outs_down[31] ,
    \_ces_2_3_io_outs_down[30] ,
    \_ces_2_3_io_outs_down[29] ,
    \_ces_2_3_io_outs_down[28] ,
    \_ces_2_3_io_outs_down[27] ,
    \_ces_2_3_io_outs_down[26] ,
    \_ces_2_3_io_outs_down[25] ,
    \_ces_2_3_io_outs_down[24] ,
    \_ces_2_3_io_outs_down[23] ,
    \_ces_2_3_io_outs_down[22] ,
    \_ces_2_3_io_outs_down[21] ,
    \_ces_2_3_io_outs_down[20] ,
    \_ces_2_3_io_outs_down[19] ,
    \_ces_2_3_io_outs_down[18] ,
    \_ces_2_3_io_outs_down[17] ,
    \_ces_2_3_io_outs_down[16] ,
    \_ces_2_3_io_outs_down[15] ,
    \_ces_2_3_io_outs_down[14] ,
    \_ces_2_3_io_outs_down[13] ,
    \_ces_2_3_io_outs_down[12] ,
    \_ces_2_3_io_outs_down[11] ,
    \_ces_2_3_io_outs_down[10] ,
    \_ces_2_3_io_outs_down[9] ,
    \_ces_2_3_io_outs_down[8] ,
    \_ces_2_3_io_outs_down[7] ,
    \_ces_2_3_io_outs_down[6] ,
    \_ces_2_3_io_outs_down[5] ,
    \_ces_2_3_io_outs_down[4] ,
    \_ces_2_3_io_outs_down[3] ,
    \_ces_2_3_io_outs_down[2] ,
    \_ces_2_3_io_outs_down[1] ,
    \_ces_2_3_io_outs_down[0] }),
    .io_outs_left({\_ces_2_3_io_outs_left[63] ,
    \_ces_2_3_io_outs_left[62] ,
    \_ces_2_3_io_outs_left[61] ,
    \_ces_2_3_io_outs_left[60] ,
    \_ces_2_3_io_outs_left[59] ,
    \_ces_2_3_io_outs_left[58] ,
    \_ces_2_3_io_outs_left[57] ,
    \_ces_2_3_io_outs_left[56] ,
    \_ces_2_3_io_outs_left[55] ,
    \_ces_2_3_io_outs_left[54] ,
    \_ces_2_3_io_outs_left[53] ,
    \_ces_2_3_io_outs_left[52] ,
    \_ces_2_3_io_outs_left[51] ,
    \_ces_2_3_io_outs_left[50] ,
    \_ces_2_3_io_outs_left[49] ,
    \_ces_2_3_io_outs_left[48] ,
    \_ces_2_3_io_outs_left[47] ,
    \_ces_2_3_io_outs_left[46] ,
    \_ces_2_3_io_outs_left[45] ,
    \_ces_2_3_io_outs_left[44] ,
    \_ces_2_3_io_outs_left[43] ,
    \_ces_2_3_io_outs_left[42] ,
    \_ces_2_3_io_outs_left[41] ,
    \_ces_2_3_io_outs_left[40] ,
    \_ces_2_3_io_outs_left[39] ,
    \_ces_2_3_io_outs_left[38] ,
    \_ces_2_3_io_outs_left[37] ,
    \_ces_2_3_io_outs_left[36] ,
    \_ces_2_3_io_outs_left[35] ,
    \_ces_2_3_io_outs_left[34] ,
    \_ces_2_3_io_outs_left[33] ,
    \_ces_2_3_io_outs_left[32] ,
    \_ces_2_3_io_outs_left[31] ,
    \_ces_2_3_io_outs_left[30] ,
    \_ces_2_3_io_outs_left[29] ,
    \_ces_2_3_io_outs_left[28] ,
    \_ces_2_3_io_outs_left[27] ,
    \_ces_2_3_io_outs_left[26] ,
    \_ces_2_3_io_outs_left[25] ,
    \_ces_2_3_io_outs_left[24] ,
    \_ces_2_3_io_outs_left[23] ,
    \_ces_2_3_io_outs_left[22] ,
    \_ces_2_3_io_outs_left[21] ,
    \_ces_2_3_io_outs_left[20] ,
    \_ces_2_3_io_outs_left[19] ,
    \_ces_2_3_io_outs_left[18] ,
    \_ces_2_3_io_outs_left[17] ,
    \_ces_2_3_io_outs_left[16] ,
    \_ces_2_3_io_outs_left[15] ,
    \_ces_2_3_io_outs_left[14] ,
    \_ces_2_3_io_outs_left[13] ,
    \_ces_2_3_io_outs_left[12] ,
    \_ces_2_3_io_outs_left[11] ,
    \_ces_2_3_io_outs_left[10] ,
    \_ces_2_3_io_outs_left[9] ,
    \_ces_2_3_io_outs_left[8] ,
    \_ces_2_3_io_outs_left[7] ,
    \_ces_2_3_io_outs_left[6] ,
    \_ces_2_3_io_outs_left[5] ,
    \_ces_2_3_io_outs_left[4] ,
    \_ces_2_3_io_outs_left[3] ,
    \_ces_2_3_io_outs_left[2] ,
    \_ces_2_3_io_outs_left[1] ,
    \_ces_2_3_io_outs_left[0] }),
    .io_outs_right({net1751,
    net1750,
    net1749,
    net1748,
    net1746,
    net1745,
    net1744,
    net1743,
    net1742,
    net1741,
    net1740,
    net1739,
    net1738,
    net1737,
    net1735,
    net1734,
    net1733,
    net1732,
    net1731,
    net1730,
    net1729,
    net1728,
    net1727,
    net1726,
    net1724,
    net1723,
    net1722,
    net1721,
    net1720,
    net1719,
    net1718,
    net1717,
    net1716,
    net1715,
    net1713,
    net1712,
    net1711,
    net1710,
    net1709,
    net1708,
    net1707,
    net1706,
    net1705,
    net1704,
    net1702,
    net1701,
    net1700,
    net1699,
    net1698,
    net1697,
    net1696,
    net1695,
    net1694,
    net1693,
    net1755,
    net1754,
    net1753,
    net1752,
    net1747,
    net1736,
    net1725,
    net1714,
    net1703,
    net1692}),
    .io_outs_up({\_ces_2_3_io_outs_up[63] ,
    \_ces_2_3_io_outs_up[62] ,
    \_ces_2_3_io_outs_up[61] ,
    \_ces_2_3_io_outs_up[60] ,
    \_ces_2_3_io_outs_up[59] ,
    \_ces_2_3_io_outs_up[58] ,
    \_ces_2_3_io_outs_up[57] ,
    \_ces_2_3_io_outs_up[56] ,
    \_ces_2_3_io_outs_up[55] ,
    \_ces_2_3_io_outs_up[54] ,
    \_ces_2_3_io_outs_up[53] ,
    \_ces_2_3_io_outs_up[52] ,
    \_ces_2_3_io_outs_up[51] ,
    \_ces_2_3_io_outs_up[50] ,
    \_ces_2_3_io_outs_up[49] ,
    \_ces_2_3_io_outs_up[48] ,
    \_ces_2_3_io_outs_up[47] ,
    \_ces_2_3_io_outs_up[46] ,
    \_ces_2_3_io_outs_up[45] ,
    \_ces_2_3_io_outs_up[44] ,
    \_ces_2_3_io_outs_up[43] ,
    \_ces_2_3_io_outs_up[42] ,
    \_ces_2_3_io_outs_up[41] ,
    \_ces_2_3_io_outs_up[40] ,
    \_ces_2_3_io_outs_up[39] ,
    \_ces_2_3_io_outs_up[38] ,
    \_ces_2_3_io_outs_up[37] ,
    \_ces_2_3_io_outs_up[36] ,
    \_ces_2_3_io_outs_up[35] ,
    \_ces_2_3_io_outs_up[34] ,
    \_ces_2_3_io_outs_up[33] ,
    \_ces_2_3_io_outs_up[32] ,
    \_ces_2_3_io_outs_up[31] ,
    \_ces_2_3_io_outs_up[30] ,
    \_ces_2_3_io_outs_up[29] ,
    \_ces_2_3_io_outs_up[28] ,
    \_ces_2_3_io_outs_up[27] ,
    \_ces_2_3_io_outs_up[26] ,
    \_ces_2_3_io_outs_up[25] ,
    \_ces_2_3_io_outs_up[24] ,
    \_ces_2_3_io_outs_up[23] ,
    \_ces_2_3_io_outs_up[22] ,
    \_ces_2_3_io_outs_up[21] ,
    \_ces_2_3_io_outs_up[20] ,
    \_ces_2_3_io_outs_up[19] ,
    \_ces_2_3_io_outs_up[18] ,
    \_ces_2_3_io_outs_up[17] ,
    \_ces_2_3_io_outs_up[16] ,
    \_ces_2_3_io_outs_up[15] ,
    \_ces_2_3_io_outs_up[14] ,
    \_ces_2_3_io_outs_up[13] ,
    \_ces_2_3_io_outs_up[12] ,
    \_ces_2_3_io_outs_up[11] ,
    \_ces_2_3_io_outs_up[10] ,
    \_ces_2_3_io_outs_up[9] ,
    \_ces_2_3_io_outs_up[8] ,
    \_ces_2_3_io_outs_up[7] ,
    \_ces_2_3_io_outs_up[6] ,
    \_ces_2_3_io_outs_up[5] ,
    \_ces_2_3_io_outs_up[4] ,
    \_ces_2_3_io_outs_up[3] ,
    \_ces_2_3_io_outs_up[2] ,
    \_ces_2_3_io_outs_up[1] ,
    \_ces_2_3_io_outs_up[0] }));
 Element ces_3_0 (.clock(clknet_leaf_0_clock),
    .io_lsbIns_1(net9),
    .io_lsbIns_2(net10),
    .io_lsbIns_3(net11),
    .io_lsbOuts_1(_ces_3_0_io_lsbOuts_1),
    .io_lsbOuts_2(_ces_3_0_io_lsbOuts_2),
    .io_lsbOuts_3(_ces_3_0_io_lsbOuts_3),
    .io_ins_down({net71,
    net70,
    net69,
    net68,
    net66,
    net65,
    net64,
    net63,
    net62,
    net61,
    net60,
    net59,
    net58,
    net57,
    net55,
    net54,
    net53,
    net52,
    net51,
    net50,
    net49,
    net48,
    net47,
    net46,
    net44,
    net43,
    net42,
    net41,
    net40,
    net39,
    net38,
    net37,
    net36,
    net35,
    net33,
    net32,
    net31,
    net30,
    net29,
    net28,
    net27,
    net26,
    net25,
    net24,
    net22,
    net21,
    net20,
    net19,
    net18,
    net17,
    net16,
    net15,
    net14,
    net13,
    net75,
    net74,
    net73,
    net72,
    net67,
    net56,
    net45,
    net34,
    net23,
    net12}),
    .io_ins_left({\_ces_3_1_io_outs_left[63] ,
    \_ces_3_1_io_outs_left[62] ,
    \_ces_3_1_io_outs_left[61] ,
    \_ces_3_1_io_outs_left[60] ,
    \_ces_3_1_io_outs_left[59] ,
    \_ces_3_1_io_outs_left[58] ,
    \_ces_3_1_io_outs_left[57] ,
    \_ces_3_1_io_outs_left[56] ,
    \_ces_3_1_io_outs_left[55] ,
    \_ces_3_1_io_outs_left[54] ,
    \_ces_3_1_io_outs_left[53] ,
    \_ces_3_1_io_outs_left[52] ,
    \_ces_3_1_io_outs_left[51] ,
    \_ces_3_1_io_outs_left[50] ,
    \_ces_3_1_io_outs_left[49] ,
    \_ces_3_1_io_outs_left[48] ,
    \_ces_3_1_io_outs_left[47] ,
    \_ces_3_1_io_outs_left[46] ,
    \_ces_3_1_io_outs_left[45] ,
    \_ces_3_1_io_outs_left[44] ,
    \_ces_3_1_io_outs_left[43] ,
    \_ces_3_1_io_outs_left[42] ,
    \_ces_3_1_io_outs_left[41] ,
    \_ces_3_1_io_outs_left[40] ,
    \_ces_3_1_io_outs_left[39] ,
    \_ces_3_1_io_outs_left[38] ,
    \_ces_3_1_io_outs_left[37] ,
    \_ces_3_1_io_outs_left[36] ,
    \_ces_3_1_io_outs_left[35] ,
    \_ces_3_1_io_outs_left[34] ,
    \_ces_3_1_io_outs_left[33] ,
    \_ces_3_1_io_outs_left[32] ,
    \_ces_3_1_io_outs_left[31] ,
    \_ces_3_1_io_outs_left[30] ,
    \_ces_3_1_io_outs_left[29] ,
    \_ces_3_1_io_outs_left[28] ,
    \_ces_3_1_io_outs_left[27] ,
    \_ces_3_1_io_outs_left[26] ,
    \_ces_3_1_io_outs_left[25] ,
    \_ces_3_1_io_outs_left[24] ,
    \_ces_3_1_io_outs_left[23] ,
    \_ces_3_1_io_outs_left[22] ,
    \_ces_3_1_io_outs_left[21] ,
    \_ces_3_1_io_outs_left[20] ,
    \_ces_3_1_io_outs_left[19] ,
    \_ces_3_1_io_outs_left[18] ,
    \_ces_3_1_io_outs_left[17] ,
    \_ces_3_1_io_outs_left[16] ,
    \_ces_3_1_io_outs_left[15] ,
    \_ces_3_1_io_outs_left[14] ,
    \_ces_3_1_io_outs_left[13] ,
    \_ces_3_1_io_outs_left[12] ,
    \_ces_3_1_io_outs_left[11] ,
    \_ces_3_1_io_outs_left[10] ,
    \_ces_3_1_io_outs_left[9] ,
    \_ces_3_1_io_outs_left[8] ,
    \_ces_3_1_io_outs_left[7] ,
    \_ces_3_1_io_outs_left[6] ,
    \_ces_3_1_io_outs_left[5] ,
    \_ces_3_1_io_outs_left[4] ,
    \_ces_3_1_io_outs_left[3] ,
    \_ces_3_1_io_outs_left[2] ,
    \_ces_3_1_io_outs_left[1] ,
    \_ces_3_1_io_outs_left[0] }),
    .io_ins_right({net775,
    net774,
    net773,
    net772,
    net770,
    net769,
    net768,
    net767,
    net766,
    net765,
    net764,
    net763,
    net762,
    net761,
    net759,
    net758,
    net757,
    net756,
    net755,
    net754,
    net753,
    net752,
    net751,
    net750,
    net748,
    net747,
    net746,
    net745,
    net744,
    net743,
    net742,
    net741,
    net740,
    net739,
    net737,
    net736,
    net735,
    net734,
    net733,
    net732,
    net731,
    net730,
    net729,
    net728,
    net726,
    net725,
    net724,
    net723,
    net722,
    net721,
    net720,
    net719,
    net718,
    net717,
    net779,
    net778,
    net777,
    net776,
    net771,
    net760,
    net749,
    net738,
    net727,
    net716}),
    .io_ins_up({\_ces_2_0_io_outs_up[63] ,
    \_ces_2_0_io_outs_up[62] ,
    \_ces_2_0_io_outs_up[61] ,
    \_ces_2_0_io_outs_up[60] ,
    \_ces_2_0_io_outs_up[59] ,
    \_ces_2_0_io_outs_up[58] ,
    \_ces_2_0_io_outs_up[57] ,
    \_ces_2_0_io_outs_up[56] ,
    \_ces_2_0_io_outs_up[55] ,
    \_ces_2_0_io_outs_up[54] ,
    \_ces_2_0_io_outs_up[53] ,
    \_ces_2_0_io_outs_up[52] ,
    \_ces_2_0_io_outs_up[51] ,
    \_ces_2_0_io_outs_up[50] ,
    \_ces_2_0_io_outs_up[49] ,
    \_ces_2_0_io_outs_up[48] ,
    \_ces_2_0_io_outs_up[47] ,
    \_ces_2_0_io_outs_up[46] ,
    \_ces_2_0_io_outs_up[45] ,
    \_ces_2_0_io_outs_up[44] ,
    \_ces_2_0_io_outs_up[43] ,
    \_ces_2_0_io_outs_up[42] ,
    \_ces_2_0_io_outs_up[41] ,
    \_ces_2_0_io_outs_up[40] ,
    \_ces_2_0_io_outs_up[39] ,
    \_ces_2_0_io_outs_up[38] ,
    \_ces_2_0_io_outs_up[37] ,
    \_ces_2_0_io_outs_up[36] ,
    \_ces_2_0_io_outs_up[35] ,
    \_ces_2_0_io_outs_up[34] ,
    \_ces_2_0_io_outs_up[33] ,
    \_ces_2_0_io_outs_up[32] ,
    \_ces_2_0_io_outs_up[31] ,
    \_ces_2_0_io_outs_up[30] ,
    \_ces_2_0_io_outs_up[29] ,
    \_ces_2_0_io_outs_up[28] ,
    \_ces_2_0_io_outs_up[27] ,
    \_ces_2_0_io_outs_up[26] ,
    \_ces_2_0_io_outs_up[25] ,
    \_ces_2_0_io_outs_up[24] ,
    \_ces_2_0_io_outs_up[23] ,
    \_ces_2_0_io_outs_up[22] ,
    \_ces_2_0_io_outs_up[21] ,
    \_ces_2_0_io_outs_up[20] ,
    \_ces_2_0_io_outs_up[19] ,
    \_ces_2_0_io_outs_up[18] ,
    \_ces_2_0_io_outs_up[17] ,
    \_ces_2_0_io_outs_up[16] ,
    \_ces_2_0_io_outs_up[15] ,
    \_ces_2_0_io_outs_up[14] ,
    \_ces_2_0_io_outs_up[13] ,
    \_ces_2_0_io_outs_up[12] ,
    \_ces_2_0_io_outs_up[11] ,
    \_ces_2_0_io_outs_up[10] ,
    \_ces_2_0_io_outs_up[9] ,
    \_ces_2_0_io_outs_up[8] ,
    \_ces_2_0_io_outs_up[7] ,
    \_ces_2_0_io_outs_up[6] ,
    \_ces_2_0_io_outs_up[5] ,
    \_ces_2_0_io_outs_up[4] ,
    \_ces_2_0_io_outs_up[3] ,
    \_ces_2_0_io_outs_up[2] ,
    \_ces_2_0_io_outs_up[1] ,
    \_ces_2_0_io_outs_up[0] }),
    .io_outs_down({\_ces_3_0_io_outs_down[63] ,
    \_ces_3_0_io_outs_down[62] ,
    \_ces_3_0_io_outs_down[61] ,
    \_ces_3_0_io_outs_down[60] ,
    \_ces_3_0_io_outs_down[59] ,
    \_ces_3_0_io_outs_down[58] ,
    \_ces_3_0_io_outs_down[57] ,
    \_ces_3_0_io_outs_down[56] ,
    \_ces_3_0_io_outs_down[55] ,
    \_ces_3_0_io_outs_down[54] ,
    \_ces_3_0_io_outs_down[53] ,
    \_ces_3_0_io_outs_down[52] ,
    \_ces_3_0_io_outs_down[51] ,
    \_ces_3_0_io_outs_down[50] ,
    \_ces_3_0_io_outs_down[49] ,
    \_ces_3_0_io_outs_down[48] ,
    \_ces_3_0_io_outs_down[47] ,
    \_ces_3_0_io_outs_down[46] ,
    \_ces_3_0_io_outs_down[45] ,
    \_ces_3_0_io_outs_down[44] ,
    \_ces_3_0_io_outs_down[43] ,
    \_ces_3_0_io_outs_down[42] ,
    \_ces_3_0_io_outs_down[41] ,
    \_ces_3_0_io_outs_down[40] ,
    \_ces_3_0_io_outs_down[39] ,
    \_ces_3_0_io_outs_down[38] ,
    \_ces_3_0_io_outs_down[37] ,
    \_ces_3_0_io_outs_down[36] ,
    \_ces_3_0_io_outs_down[35] ,
    \_ces_3_0_io_outs_down[34] ,
    \_ces_3_0_io_outs_down[33] ,
    \_ces_3_0_io_outs_down[32] ,
    \_ces_3_0_io_outs_down[31] ,
    \_ces_3_0_io_outs_down[30] ,
    \_ces_3_0_io_outs_down[29] ,
    \_ces_3_0_io_outs_down[28] ,
    \_ces_3_0_io_outs_down[27] ,
    \_ces_3_0_io_outs_down[26] ,
    \_ces_3_0_io_outs_down[25] ,
    \_ces_3_0_io_outs_down[24] ,
    \_ces_3_0_io_outs_down[23] ,
    \_ces_3_0_io_outs_down[22] ,
    \_ces_3_0_io_outs_down[21] ,
    \_ces_3_0_io_outs_down[20] ,
    \_ces_3_0_io_outs_down[19] ,
    \_ces_3_0_io_outs_down[18] ,
    \_ces_3_0_io_outs_down[17] ,
    \_ces_3_0_io_outs_down[16] ,
    \_ces_3_0_io_outs_down[15] ,
    \_ces_3_0_io_outs_down[14] ,
    \_ces_3_0_io_outs_down[13] ,
    \_ces_3_0_io_outs_down[12] ,
    \_ces_3_0_io_outs_down[11] ,
    \_ces_3_0_io_outs_down[10] ,
    \_ces_3_0_io_outs_down[9] ,
    \_ces_3_0_io_outs_down[8] ,
    \_ces_3_0_io_outs_down[7] ,
    \_ces_3_0_io_outs_down[6] ,
    \_ces_3_0_io_outs_down[5] ,
    \_ces_3_0_io_outs_down[4] ,
    \_ces_3_0_io_outs_down[3] ,
    \_ces_3_0_io_outs_down[2] ,
    \_ces_3_0_io_outs_down[1] ,
    \_ces_3_0_io_outs_down[0] }),
    .io_outs_left({net1559,
    net1558,
    net1557,
    net1556,
    net1554,
    net1553,
    net1552,
    net1551,
    net1550,
    net1549,
    net1548,
    net1547,
    net1546,
    net1545,
    net1543,
    net1542,
    net1541,
    net1540,
    net1539,
    net1538,
    net1537,
    net1536,
    net1535,
    net1534,
    net1532,
    net1531,
    net1530,
    net1529,
    net1528,
    net1527,
    net1526,
    net1525,
    net1524,
    net1523,
    net1521,
    net1520,
    net1519,
    net1518,
    net1517,
    net1516,
    net1515,
    net1514,
    net1513,
    net1512,
    net1510,
    net1509,
    net1508,
    net1507,
    net1506,
    net1505,
    net1504,
    net1503,
    net1502,
    net1501,
    net1563,
    net1562,
    net1561,
    net1560,
    net1555,
    net1544,
    net1533,
    net1522,
    net1511,
    net1500}),
    .io_outs_right({\_ces_3_0_io_outs_right[63] ,
    \_ces_3_0_io_outs_right[62] ,
    \_ces_3_0_io_outs_right[61] ,
    \_ces_3_0_io_outs_right[60] ,
    \_ces_3_0_io_outs_right[59] ,
    \_ces_3_0_io_outs_right[58] ,
    \_ces_3_0_io_outs_right[57] ,
    \_ces_3_0_io_outs_right[56] ,
    \_ces_3_0_io_outs_right[55] ,
    \_ces_3_0_io_outs_right[54] ,
    \_ces_3_0_io_outs_right[53] ,
    \_ces_3_0_io_outs_right[52] ,
    \_ces_3_0_io_outs_right[51] ,
    \_ces_3_0_io_outs_right[50] ,
    \_ces_3_0_io_outs_right[49] ,
    \_ces_3_0_io_outs_right[48] ,
    \_ces_3_0_io_outs_right[47] ,
    \_ces_3_0_io_outs_right[46] ,
    \_ces_3_0_io_outs_right[45] ,
    \_ces_3_0_io_outs_right[44] ,
    \_ces_3_0_io_outs_right[43] ,
    \_ces_3_0_io_outs_right[42] ,
    \_ces_3_0_io_outs_right[41] ,
    \_ces_3_0_io_outs_right[40] ,
    \_ces_3_0_io_outs_right[39] ,
    \_ces_3_0_io_outs_right[38] ,
    \_ces_3_0_io_outs_right[37] ,
    \_ces_3_0_io_outs_right[36] ,
    \_ces_3_0_io_outs_right[35] ,
    \_ces_3_0_io_outs_right[34] ,
    \_ces_3_0_io_outs_right[33] ,
    \_ces_3_0_io_outs_right[32] ,
    \_ces_3_0_io_outs_right[31] ,
    \_ces_3_0_io_outs_right[30] ,
    \_ces_3_0_io_outs_right[29] ,
    \_ces_3_0_io_outs_right[28] ,
    \_ces_3_0_io_outs_right[27] ,
    \_ces_3_0_io_outs_right[26] ,
    \_ces_3_0_io_outs_right[25] ,
    \_ces_3_0_io_outs_right[24] ,
    \_ces_3_0_io_outs_right[23] ,
    \_ces_3_0_io_outs_right[22] ,
    \_ces_3_0_io_outs_right[21] ,
    \_ces_3_0_io_outs_right[20] ,
    \_ces_3_0_io_outs_right[19] ,
    \_ces_3_0_io_outs_right[18] ,
    \_ces_3_0_io_outs_right[17] ,
    \_ces_3_0_io_outs_right[16] ,
    \_ces_3_0_io_outs_right[15] ,
    \_ces_3_0_io_outs_right[14] ,
    \_ces_3_0_io_outs_right[13] ,
    \_ces_3_0_io_outs_right[12] ,
    \_ces_3_0_io_outs_right[11] ,
    \_ces_3_0_io_outs_right[10] ,
    \_ces_3_0_io_outs_right[9] ,
    \_ces_3_0_io_outs_right[8] ,
    \_ces_3_0_io_outs_right[7] ,
    \_ces_3_0_io_outs_right[6] ,
    \_ces_3_0_io_outs_right[5] ,
    \_ces_3_0_io_outs_right[4] ,
    \_ces_3_0_io_outs_right[3] ,
    \_ces_3_0_io_outs_right[2] ,
    \_ces_3_0_io_outs_right[1] ,
    \_ces_3_0_io_outs_right[0] }),
    .io_outs_up({net1879,
    net1878,
    net1877,
    net1876,
    net1874,
    net1873,
    net1872,
    net1871,
    net1870,
    net1869,
    net1868,
    net1867,
    net1866,
    net1865,
    net1863,
    net1862,
    net1861,
    net1860,
    net1859,
    net1858,
    net1857,
    net1856,
    net1855,
    net1854,
    net1852,
    net1851,
    net1850,
    net1849,
    net1848,
    net1847,
    net1846,
    net1845,
    net1844,
    net1843,
    net1841,
    net1840,
    net1839,
    net1838,
    net1837,
    net1836,
    net1835,
    net1834,
    net1833,
    net1832,
    net1830,
    net1829,
    net1828,
    net1827,
    net1826,
    net1825,
    net1824,
    net1823,
    net1822,
    net1821,
    net1883,
    net1882,
    net1881,
    net1880,
    net1875,
    net1864,
    net1853,
    net1842,
    net1831,
    net1820}));
 Element ces_3_1 (.clock(clknet_leaf_0_clock),
    .io_lsbIns_1(_ces_3_0_io_lsbOuts_1),
    .io_lsbIns_2(_ces_3_0_io_lsbOuts_2),
    .io_lsbIns_3(_ces_3_0_io_lsbOuts_3),
    .io_lsbOuts_1(_ces_3_1_io_lsbOuts_1),
    .io_lsbOuts_2(_ces_3_1_io_lsbOuts_2),
    .io_lsbOuts_3(_ces_3_1_io_lsbOuts_3),
    .io_ins_down({net135,
    net134,
    net133,
    net132,
    net130,
    net129,
    net128,
    net127,
    net126,
    net125,
    net124,
    net123,
    net122,
    net121,
    net119,
    net118,
    net117,
    net116,
    net115,
    net114,
    net113,
    net112,
    net111,
    net110,
    net108,
    net107,
    net106,
    net105,
    net104,
    net103,
    net102,
    net101,
    net100,
    net99,
    net97,
    net96,
    net95,
    net94,
    net93,
    net92,
    net91,
    net90,
    net89,
    net88,
    net86,
    net85,
    net84,
    net83,
    net82,
    net81,
    net80,
    net79,
    net78,
    net77,
    net139,
    net138,
    net137,
    net136,
    net131,
    net120,
    net109,
    net98,
    net87,
    net76}),
    .io_ins_left({\_ces_3_2_io_outs_left[63] ,
    \_ces_3_2_io_outs_left[62] ,
    \_ces_3_2_io_outs_left[61] ,
    \_ces_3_2_io_outs_left[60] ,
    \_ces_3_2_io_outs_left[59] ,
    \_ces_3_2_io_outs_left[58] ,
    \_ces_3_2_io_outs_left[57] ,
    \_ces_3_2_io_outs_left[56] ,
    \_ces_3_2_io_outs_left[55] ,
    \_ces_3_2_io_outs_left[54] ,
    \_ces_3_2_io_outs_left[53] ,
    \_ces_3_2_io_outs_left[52] ,
    \_ces_3_2_io_outs_left[51] ,
    \_ces_3_2_io_outs_left[50] ,
    \_ces_3_2_io_outs_left[49] ,
    \_ces_3_2_io_outs_left[48] ,
    \_ces_3_2_io_outs_left[47] ,
    \_ces_3_2_io_outs_left[46] ,
    \_ces_3_2_io_outs_left[45] ,
    \_ces_3_2_io_outs_left[44] ,
    \_ces_3_2_io_outs_left[43] ,
    \_ces_3_2_io_outs_left[42] ,
    \_ces_3_2_io_outs_left[41] ,
    \_ces_3_2_io_outs_left[40] ,
    \_ces_3_2_io_outs_left[39] ,
    \_ces_3_2_io_outs_left[38] ,
    \_ces_3_2_io_outs_left[37] ,
    \_ces_3_2_io_outs_left[36] ,
    \_ces_3_2_io_outs_left[35] ,
    \_ces_3_2_io_outs_left[34] ,
    \_ces_3_2_io_outs_left[33] ,
    \_ces_3_2_io_outs_left[32] ,
    \_ces_3_2_io_outs_left[31] ,
    \_ces_3_2_io_outs_left[30] ,
    \_ces_3_2_io_outs_left[29] ,
    \_ces_3_2_io_outs_left[28] ,
    \_ces_3_2_io_outs_left[27] ,
    \_ces_3_2_io_outs_left[26] ,
    \_ces_3_2_io_outs_left[25] ,
    \_ces_3_2_io_outs_left[24] ,
    \_ces_3_2_io_outs_left[23] ,
    \_ces_3_2_io_outs_left[22] ,
    \_ces_3_2_io_outs_left[21] ,
    \_ces_3_2_io_outs_left[20] ,
    \_ces_3_2_io_outs_left[19] ,
    \_ces_3_2_io_outs_left[18] ,
    \_ces_3_2_io_outs_left[17] ,
    \_ces_3_2_io_outs_left[16] ,
    \_ces_3_2_io_outs_left[15] ,
    \_ces_3_2_io_outs_left[14] ,
    \_ces_3_2_io_outs_left[13] ,
    \_ces_3_2_io_outs_left[12] ,
    \_ces_3_2_io_outs_left[11] ,
    \_ces_3_2_io_outs_left[10] ,
    \_ces_3_2_io_outs_left[9] ,
    \_ces_3_2_io_outs_left[8] ,
    \_ces_3_2_io_outs_left[7] ,
    \_ces_3_2_io_outs_left[6] ,
    \_ces_3_2_io_outs_left[5] ,
    \_ces_3_2_io_outs_left[4] ,
    \_ces_3_2_io_outs_left[3] ,
    \_ces_3_2_io_outs_left[2] ,
    \_ces_3_2_io_outs_left[1] ,
    \_ces_3_2_io_outs_left[0] }),
    .io_ins_right({\_ces_3_0_io_outs_right[63] ,
    \_ces_3_0_io_outs_right[62] ,
    \_ces_3_0_io_outs_right[61] ,
    \_ces_3_0_io_outs_right[60] ,
    \_ces_3_0_io_outs_right[59] ,
    \_ces_3_0_io_outs_right[58] ,
    \_ces_3_0_io_outs_right[57] ,
    \_ces_3_0_io_outs_right[56] ,
    \_ces_3_0_io_outs_right[55] ,
    \_ces_3_0_io_outs_right[54] ,
    \_ces_3_0_io_outs_right[53] ,
    \_ces_3_0_io_outs_right[52] ,
    \_ces_3_0_io_outs_right[51] ,
    \_ces_3_0_io_outs_right[50] ,
    \_ces_3_0_io_outs_right[49] ,
    \_ces_3_0_io_outs_right[48] ,
    \_ces_3_0_io_outs_right[47] ,
    \_ces_3_0_io_outs_right[46] ,
    \_ces_3_0_io_outs_right[45] ,
    \_ces_3_0_io_outs_right[44] ,
    \_ces_3_0_io_outs_right[43] ,
    \_ces_3_0_io_outs_right[42] ,
    \_ces_3_0_io_outs_right[41] ,
    \_ces_3_0_io_outs_right[40] ,
    \_ces_3_0_io_outs_right[39] ,
    \_ces_3_0_io_outs_right[38] ,
    \_ces_3_0_io_outs_right[37] ,
    \_ces_3_0_io_outs_right[36] ,
    \_ces_3_0_io_outs_right[35] ,
    \_ces_3_0_io_outs_right[34] ,
    \_ces_3_0_io_outs_right[33] ,
    \_ces_3_0_io_outs_right[32] ,
    \_ces_3_0_io_outs_right[31] ,
    \_ces_3_0_io_outs_right[30] ,
    \_ces_3_0_io_outs_right[29] ,
    \_ces_3_0_io_outs_right[28] ,
    \_ces_3_0_io_outs_right[27] ,
    \_ces_3_0_io_outs_right[26] ,
    \_ces_3_0_io_outs_right[25] ,
    \_ces_3_0_io_outs_right[24] ,
    \_ces_3_0_io_outs_right[23] ,
    \_ces_3_0_io_outs_right[22] ,
    \_ces_3_0_io_outs_right[21] ,
    \_ces_3_0_io_outs_right[20] ,
    \_ces_3_0_io_outs_right[19] ,
    \_ces_3_0_io_outs_right[18] ,
    \_ces_3_0_io_outs_right[17] ,
    \_ces_3_0_io_outs_right[16] ,
    \_ces_3_0_io_outs_right[15] ,
    \_ces_3_0_io_outs_right[14] ,
    \_ces_3_0_io_outs_right[13] ,
    \_ces_3_0_io_outs_right[12] ,
    \_ces_3_0_io_outs_right[11] ,
    \_ces_3_0_io_outs_right[10] ,
    \_ces_3_0_io_outs_right[9] ,
    \_ces_3_0_io_outs_right[8] ,
    \_ces_3_0_io_outs_right[7] ,
    \_ces_3_0_io_outs_right[6] ,
    \_ces_3_0_io_outs_right[5] ,
    \_ces_3_0_io_outs_right[4] ,
    \_ces_3_0_io_outs_right[3] ,
    \_ces_3_0_io_outs_right[2] ,
    \_ces_3_0_io_outs_right[1] ,
    \_ces_3_0_io_outs_right[0] }),
    .io_ins_up({\_ces_2_1_io_outs_up[63] ,
    \_ces_2_1_io_outs_up[62] ,
    \_ces_2_1_io_outs_up[61] ,
    \_ces_2_1_io_outs_up[60] ,
    \_ces_2_1_io_outs_up[59] ,
    \_ces_2_1_io_outs_up[58] ,
    \_ces_2_1_io_outs_up[57] ,
    \_ces_2_1_io_outs_up[56] ,
    \_ces_2_1_io_outs_up[55] ,
    \_ces_2_1_io_outs_up[54] ,
    \_ces_2_1_io_outs_up[53] ,
    \_ces_2_1_io_outs_up[52] ,
    \_ces_2_1_io_outs_up[51] ,
    \_ces_2_1_io_outs_up[50] ,
    \_ces_2_1_io_outs_up[49] ,
    \_ces_2_1_io_outs_up[48] ,
    \_ces_2_1_io_outs_up[47] ,
    \_ces_2_1_io_outs_up[46] ,
    \_ces_2_1_io_outs_up[45] ,
    \_ces_2_1_io_outs_up[44] ,
    \_ces_2_1_io_outs_up[43] ,
    \_ces_2_1_io_outs_up[42] ,
    \_ces_2_1_io_outs_up[41] ,
    \_ces_2_1_io_outs_up[40] ,
    \_ces_2_1_io_outs_up[39] ,
    \_ces_2_1_io_outs_up[38] ,
    \_ces_2_1_io_outs_up[37] ,
    \_ces_2_1_io_outs_up[36] ,
    \_ces_2_1_io_outs_up[35] ,
    \_ces_2_1_io_outs_up[34] ,
    \_ces_2_1_io_outs_up[33] ,
    \_ces_2_1_io_outs_up[32] ,
    \_ces_2_1_io_outs_up[31] ,
    \_ces_2_1_io_outs_up[30] ,
    \_ces_2_1_io_outs_up[29] ,
    \_ces_2_1_io_outs_up[28] ,
    \_ces_2_1_io_outs_up[27] ,
    \_ces_2_1_io_outs_up[26] ,
    \_ces_2_1_io_outs_up[25] ,
    \_ces_2_1_io_outs_up[24] ,
    \_ces_2_1_io_outs_up[23] ,
    \_ces_2_1_io_outs_up[22] ,
    \_ces_2_1_io_outs_up[21] ,
    \_ces_2_1_io_outs_up[20] ,
    \_ces_2_1_io_outs_up[19] ,
    \_ces_2_1_io_outs_up[18] ,
    \_ces_2_1_io_outs_up[17] ,
    \_ces_2_1_io_outs_up[16] ,
    \_ces_2_1_io_outs_up[15] ,
    \_ces_2_1_io_outs_up[14] ,
    \_ces_2_1_io_outs_up[13] ,
    \_ces_2_1_io_outs_up[12] ,
    \_ces_2_1_io_outs_up[11] ,
    \_ces_2_1_io_outs_up[10] ,
    \_ces_2_1_io_outs_up[9] ,
    \_ces_2_1_io_outs_up[8] ,
    \_ces_2_1_io_outs_up[7] ,
    \_ces_2_1_io_outs_up[6] ,
    \_ces_2_1_io_outs_up[5] ,
    \_ces_2_1_io_outs_up[4] ,
    \_ces_2_1_io_outs_up[3] ,
    \_ces_2_1_io_outs_up[2] ,
    \_ces_2_1_io_outs_up[1] ,
    \_ces_2_1_io_outs_up[0] }),
    .io_outs_down({\_ces_3_1_io_outs_down[63] ,
    \_ces_3_1_io_outs_down[62] ,
    \_ces_3_1_io_outs_down[61] ,
    \_ces_3_1_io_outs_down[60] ,
    \_ces_3_1_io_outs_down[59] ,
    \_ces_3_1_io_outs_down[58] ,
    \_ces_3_1_io_outs_down[57] ,
    \_ces_3_1_io_outs_down[56] ,
    \_ces_3_1_io_outs_down[55] ,
    \_ces_3_1_io_outs_down[54] ,
    \_ces_3_1_io_outs_down[53] ,
    \_ces_3_1_io_outs_down[52] ,
    \_ces_3_1_io_outs_down[51] ,
    \_ces_3_1_io_outs_down[50] ,
    \_ces_3_1_io_outs_down[49] ,
    \_ces_3_1_io_outs_down[48] ,
    \_ces_3_1_io_outs_down[47] ,
    \_ces_3_1_io_outs_down[46] ,
    \_ces_3_1_io_outs_down[45] ,
    \_ces_3_1_io_outs_down[44] ,
    \_ces_3_1_io_outs_down[43] ,
    \_ces_3_1_io_outs_down[42] ,
    \_ces_3_1_io_outs_down[41] ,
    \_ces_3_1_io_outs_down[40] ,
    \_ces_3_1_io_outs_down[39] ,
    \_ces_3_1_io_outs_down[38] ,
    \_ces_3_1_io_outs_down[37] ,
    \_ces_3_1_io_outs_down[36] ,
    \_ces_3_1_io_outs_down[35] ,
    \_ces_3_1_io_outs_down[34] ,
    \_ces_3_1_io_outs_down[33] ,
    \_ces_3_1_io_outs_down[32] ,
    \_ces_3_1_io_outs_down[31] ,
    \_ces_3_1_io_outs_down[30] ,
    \_ces_3_1_io_outs_down[29] ,
    \_ces_3_1_io_outs_down[28] ,
    \_ces_3_1_io_outs_down[27] ,
    \_ces_3_1_io_outs_down[26] ,
    \_ces_3_1_io_outs_down[25] ,
    \_ces_3_1_io_outs_down[24] ,
    \_ces_3_1_io_outs_down[23] ,
    \_ces_3_1_io_outs_down[22] ,
    \_ces_3_1_io_outs_down[21] ,
    \_ces_3_1_io_outs_down[20] ,
    \_ces_3_1_io_outs_down[19] ,
    \_ces_3_1_io_outs_down[18] ,
    \_ces_3_1_io_outs_down[17] ,
    \_ces_3_1_io_outs_down[16] ,
    \_ces_3_1_io_outs_down[15] ,
    \_ces_3_1_io_outs_down[14] ,
    \_ces_3_1_io_outs_down[13] ,
    \_ces_3_1_io_outs_down[12] ,
    \_ces_3_1_io_outs_down[11] ,
    \_ces_3_1_io_outs_down[10] ,
    \_ces_3_1_io_outs_down[9] ,
    \_ces_3_1_io_outs_down[8] ,
    \_ces_3_1_io_outs_down[7] ,
    \_ces_3_1_io_outs_down[6] ,
    \_ces_3_1_io_outs_down[5] ,
    \_ces_3_1_io_outs_down[4] ,
    \_ces_3_1_io_outs_down[3] ,
    \_ces_3_1_io_outs_down[2] ,
    \_ces_3_1_io_outs_down[1] ,
    \_ces_3_1_io_outs_down[0] }),
    .io_outs_left({\_ces_3_1_io_outs_left[63] ,
    \_ces_3_1_io_outs_left[62] ,
    \_ces_3_1_io_outs_left[61] ,
    \_ces_3_1_io_outs_left[60] ,
    \_ces_3_1_io_outs_left[59] ,
    \_ces_3_1_io_outs_left[58] ,
    \_ces_3_1_io_outs_left[57] ,
    \_ces_3_1_io_outs_left[56] ,
    \_ces_3_1_io_outs_left[55] ,
    \_ces_3_1_io_outs_left[54] ,
    \_ces_3_1_io_outs_left[53] ,
    \_ces_3_1_io_outs_left[52] ,
    \_ces_3_1_io_outs_left[51] ,
    \_ces_3_1_io_outs_left[50] ,
    \_ces_3_1_io_outs_left[49] ,
    \_ces_3_1_io_outs_left[48] ,
    \_ces_3_1_io_outs_left[47] ,
    \_ces_3_1_io_outs_left[46] ,
    \_ces_3_1_io_outs_left[45] ,
    \_ces_3_1_io_outs_left[44] ,
    \_ces_3_1_io_outs_left[43] ,
    \_ces_3_1_io_outs_left[42] ,
    \_ces_3_1_io_outs_left[41] ,
    \_ces_3_1_io_outs_left[40] ,
    \_ces_3_1_io_outs_left[39] ,
    \_ces_3_1_io_outs_left[38] ,
    \_ces_3_1_io_outs_left[37] ,
    \_ces_3_1_io_outs_left[36] ,
    \_ces_3_1_io_outs_left[35] ,
    \_ces_3_1_io_outs_left[34] ,
    \_ces_3_1_io_outs_left[33] ,
    \_ces_3_1_io_outs_left[32] ,
    \_ces_3_1_io_outs_left[31] ,
    \_ces_3_1_io_outs_left[30] ,
    \_ces_3_1_io_outs_left[29] ,
    \_ces_3_1_io_outs_left[28] ,
    \_ces_3_1_io_outs_left[27] ,
    \_ces_3_1_io_outs_left[26] ,
    \_ces_3_1_io_outs_left[25] ,
    \_ces_3_1_io_outs_left[24] ,
    \_ces_3_1_io_outs_left[23] ,
    \_ces_3_1_io_outs_left[22] ,
    \_ces_3_1_io_outs_left[21] ,
    \_ces_3_1_io_outs_left[20] ,
    \_ces_3_1_io_outs_left[19] ,
    \_ces_3_1_io_outs_left[18] ,
    \_ces_3_1_io_outs_left[17] ,
    \_ces_3_1_io_outs_left[16] ,
    \_ces_3_1_io_outs_left[15] ,
    \_ces_3_1_io_outs_left[14] ,
    \_ces_3_1_io_outs_left[13] ,
    \_ces_3_1_io_outs_left[12] ,
    \_ces_3_1_io_outs_left[11] ,
    \_ces_3_1_io_outs_left[10] ,
    \_ces_3_1_io_outs_left[9] ,
    \_ces_3_1_io_outs_left[8] ,
    \_ces_3_1_io_outs_left[7] ,
    \_ces_3_1_io_outs_left[6] ,
    \_ces_3_1_io_outs_left[5] ,
    \_ces_3_1_io_outs_left[4] ,
    \_ces_3_1_io_outs_left[3] ,
    \_ces_3_1_io_outs_left[2] ,
    \_ces_3_1_io_outs_left[1] ,
    \_ces_3_1_io_outs_left[0] }),
    .io_outs_right({\_ces_3_1_io_outs_right[63] ,
    \_ces_3_1_io_outs_right[62] ,
    \_ces_3_1_io_outs_right[61] ,
    \_ces_3_1_io_outs_right[60] ,
    \_ces_3_1_io_outs_right[59] ,
    \_ces_3_1_io_outs_right[58] ,
    \_ces_3_1_io_outs_right[57] ,
    \_ces_3_1_io_outs_right[56] ,
    \_ces_3_1_io_outs_right[55] ,
    \_ces_3_1_io_outs_right[54] ,
    \_ces_3_1_io_outs_right[53] ,
    \_ces_3_1_io_outs_right[52] ,
    \_ces_3_1_io_outs_right[51] ,
    \_ces_3_1_io_outs_right[50] ,
    \_ces_3_1_io_outs_right[49] ,
    \_ces_3_1_io_outs_right[48] ,
    \_ces_3_1_io_outs_right[47] ,
    \_ces_3_1_io_outs_right[46] ,
    \_ces_3_1_io_outs_right[45] ,
    \_ces_3_1_io_outs_right[44] ,
    \_ces_3_1_io_outs_right[43] ,
    \_ces_3_1_io_outs_right[42] ,
    \_ces_3_1_io_outs_right[41] ,
    \_ces_3_1_io_outs_right[40] ,
    \_ces_3_1_io_outs_right[39] ,
    \_ces_3_1_io_outs_right[38] ,
    \_ces_3_1_io_outs_right[37] ,
    \_ces_3_1_io_outs_right[36] ,
    \_ces_3_1_io_outs_right[35] ,
    \_ces_3_1_io_outs_right[34] ,
    \_ces_3_1_io_outs_right[33] ,
    \_ces_3_1_io_outs_right[32] ,
    \_ces_3_1_io_outs_right[31] ,
    \_ces_3_1_io_outs_right[30] ,
    \_ces_3_1_io_outs_right[29] ,
    \_ces_3_1_io_outs_right[28] ,
    \_ces_3_1_io_outs_right[27] ,
    \_ces_3_1_io_outs_right[26] ,
    \_ces_3_1_io_outs_right[25] ,
    \_ces_3_1_io_outs_right[24] ,
    \_ces_3_1_io_outs_right[23] ,
    \_ces_3_1_io_outs_right[22] ,
    \_ces_3_1_io_outs_right[21] ,
    \_ces_3_1_io_outs_right[20] ,
    \_ces_3_1_io_outs_right[19] ,
    \_ces_3_1_io_outs_right[18] ,
    \_ces_3_1_io_outs_right[17] ,
    \_ces_3_1_io_outs_right[16] ,
    \_ces_3_1_io_outs_right[15] ,
    \_ces_3_1_io_outs_right[14] ,
    \_ces_3_1_io_outs_right[13] ,
    \_ces_3_1_io_outs_right[12] ,
    \_ces_3_1_io_outs_right[11] ,
    \_ces_3_1_io_outs_right[10] ,
    \_ces_3_1_io_outs_right[9] ,
    \_ces_3_1_io_outs_right[8] ,
    \_ces_3_1_io_outs_right[7] ,
    \_ces_3_1_io_outs_right[6] ,
    \_ces_3_1_io_outs_right[5] ,
    \_ces_3_1_io_outs_right[4] ,
    \_ces_3_1_io_outs_right[3] ,
    \_ces_3_1_io_outs_right[2] ,
    \_ces_3_1_io_outs_right[1] ,
    \_ces_3_1_io_outs_right[0] }),
    .io_outs_up({net1943,
    net1942,
    net1941,
    net1940,
    net1938,
    net1937,
    net1936,
    net1935,
    net1934,
    net1933,
    net1932,
    net1931,
    net1930,
    net1929,
    net1927,
    net1926,
    net1925,
    net1924,
    net1923,
    net1922,
    net1921,
    net1920,
    net1919,
    net1918,
    net1916,
    net1915,
    net1914,
    net1913,
    net1912,
    net1911,
    net1910,
    net1909,
    net1908,
    net1907,
    net1905,
    net1904,
    net1903,
    net1902,
    net1901,
    net1900,
    net1899,
    net1898,
    net1897,
    net1896,
    net1894,
    net1893,
    net1892,
    net1891,
    net1890,
    net1889,
    net1888,
    net1887,
    net1886,
    net1885,
    net1947,
    net1946,
    net1945,
    net1944,
    net1939,
    net1928,
    net1917,
    net1906,
    net1895,
    net1884}));
 Element ces_3_2 (.clock(clknet_leaf_1_clock),
    .io_lsbIns_1(_ces_3_1_io_lsbOuts_1),
    .io_lsbIns_2(_ces_3_1_io_lsbOuts_2),
    .io_lsbIns_3(_ces_3_1_io_lsbOuts_3),
    .io_lsbOuts_1(_ces_3_2_io_lsbOuts_1),
    .io_lsbOuts_2(_ces_3_2_io_lsbOuts_2),
    .io_lsbOuts_3(_ces_3_2_io_lsbOuts_3),
    .io_ins_down({net199,
    net198,
    net197,
    net196,
    net194,
    net193,
    net192,
    net191,
    net190,
    net189,
    net188,
    net187,
    net186,
    net185,
    net183,
    net182,
    net181,
    net180,
    net179,
    net178,
    net177,
    net176,
    net175,
    net174,
    net172,
    net171,
    net170,
    net169,
    net168,
    net167,
    net166,
    net165,
    net164,
    net163,
    net161,
    net160,
    net159,
    net158,
    net157,
    net156,
    net155,
    net154,
    net153,
    net152,
    net150,
    net149,
    net148,
    net147,
    net146,
    net145,
    net144,
    net143,
    net142,
    net141,
    net203,
    net202,
    net201,
    net200,
    net195,
    net184,
    net173,
    net162,
    net151,
    net140}),
    .io_ins_left({\_ces_3_3_io_outs_left[63] ,
    \_ces_3_3_io_outs_left[62] ,
    \_ces_3_3_io_outs_left[61] ,
    \_ces_3_3_io_outs_left[60] ,
    \_ces_3_3_io_outs_left[59] ,
    \_ces_3_3_io_outs_left[58] ,
    \_ces_3_3_io_outs_left[57] ,
    \_ces_3_3_io_outs_left[56] ,
    \_ces_3_3_io_outs_left[55] ,
    \_ces_3_3_io_outs_left[54] ,
    \_ces_3_3_io_outs_left[53] ,
    \_ces_3_3_io_outs_left[52] ,
    \_ces_3_3_io_outs_left[51] ,
    \_ces_3_3_io_outs_left[50] ,
    \_ces_3_3_io_outs_left[49] ,
    \_ces_3_3_io_outs_left[48] ,
    \_ces_3_3_io_outs_left[47] ,
    \_ces_3_3_io_outs_left[46] ,
    \_ces_3_3_io_outs_left[45] ,
    \_ces_3_3_io_outs_left[44] ,
    \_ces_3_3_io_outs_left[43] ,
    \_ces_3_3_io_outs_left[42] ,
    \_ces_3_3_io_outs_left[41] ,
    \_ces_3_3_io_outs_left[40] ,
    \_ces_3_3_io_outs_left[39] ,
    \_ces_3_3_io_outs_left[38] ,
    \_ces_3_3_io_outs_left[37] ,
    \_ces_3_3_io_outs_left[36] ,
    \_ces_3_3_io_outs_left[35] ,
    \_ces_3_3_io_outs_left[34] ,
    \_ces_3_3_io_outs_left[33] ,
    \_ces_3_3_io_outs_left[32] ,
    \_ces_3_3_io_outs_left[31] ,
    \_ces_3_3_io_outs_left[30] ,
    \_ces_3_3_io_outs_left[29] ,
    \_ces_3_3_io_outs_left[28] ,
    \_ces_3_3_io_outs_left[27] ,
    \_ces_3_3_io_outs_left[26] ,
    \_ces_3_3_io_outs_left[25] ,
    \_ces_3_3_io_outs_left[24] ,
    \_ces_3_3_io_outs_left[23] ,
    \_ces_3_3_io_outs_left[22] ,
    \_ces_3_3_io_outs_left[21] ,
    \_ces_3_3_io_outs_left[20] ,
    \_ces_3_3_io_outs_left[19] ,
    \_ces_3_3_io_outs_left[18] ,
    \_ces_3_3_io_outs_left[17] ,
    \_ces_3_3_io_outs_left[16] ,
    \_ces_3_3_io_outs_left[15] ,
    \_ces_3_3_io_outs_left[14] ,
    \_ces_3_3_io_outs_left[13] ,
    \_ces_3_3_io_outs_left[12] ,
    \_ces_3_3_io_outs_left[11] ,
    \_ces_3_3_io_outs_left[10] ,
    \_ces_3_3_io_outs_left[9] ,
    \_ces_3_3_io_outs_left[8] ,
    \_ces_3_3_io_outs_left[7] ,
    \_ces_3_3_io_outs_left[6] ,
    \_ces_3_3_io_outs_left[5] ,
    \_ces_3_3_io_outs_left[4] ,
    \_ces_3_3_io_outs_left[3] ,
    \_ces_3_3_io_outs_left[2] ,
    \_ces_3_3_io_outs_left[1] ,
    \_ces_3_3_io_outs_left[0] }),
    .io_ins_right({\_ces_3_1_io_outs_right[63] ,
    \_ces_3_1_io_outs_right[62] ,
    \_ces_3_1_io_outs_right[61] ,
    \_ces_3_1_io_outs_right[60] ,
    \_ces_3_1_io_outs_right[59] ,
    \_ces_3_1_io_outs_right[58] ,
    \_ces_3_1_io_outs_right[57] ,
    \_ces_3_1_io_outs_right[56] ,
    \_ces_3_1_io_outs_right[55] ,
    \_ces_3_1_io_outs_right[54] ,
    \_ces_3_1_io_outs_right[53] ,
    \_ces_3_1_io_outs_right[52] ,
    \_ces_3_1_io_outs_right[51] ,
    \_ces_3_1_io_outs_right[50] ,
    \_ces_3_1_io_outs_right[49] ,
    \_ces_3_1_io_outs_right[48] ,
    \_ces_3_1_io_outs_right[47] ,
    \_ces_3_1_io_outs_right[46] ,
    \_ces_3_1_io_outs_right[45] ,
    \_ces_3_1_io_outs_right[44] ,
    \_ces_3_1_io_outs_right[43] ,
    \_ces_3_1_io_outs_right[42] ,
    \_ces_3_1_io_outs_right[41] ,
    \_ces_3_1_io_outs_right[40] ,
    \_ces_3_1_io_outs_right[39] ,
    \_ces_3_1_io_outs_right[38] ,
    \_ces_3_1_io_outs_right[37] ,
    \_ces_3_1_io_outs_right[36] ,
    \_ces_3_1_io_outs_right[35] ,
    \_ces_3_1_io_outs_right[34] ,
    \_ces_3_1_io_outs_right[33] ,
    \_ces_3_1_io_outs_right[32] ,
    \_ces_3_1_io_outs_right[31] ,
    \_ces_3_1_io_outs_right[30] ,
    \_ces_3_1_io_outs_right[29] ,
    \_ces_3_1_io_outs_right[28] ,
    \_ces_3_1_io_outs_right[27] ,
    \_ces_3_1_io_outs_right[26] ,
    \_ces_3_1_io_outs_right[25] ,
    \_ces_3_1_io_outs_right[24] ,
    \_ces_3_1_io_outs_right[23] ,
    \_ces_3_1_io_outs_right[22] ,
    \_ces_3_1_io_outs_right[21] ,
    \_ces_3_1_io_outs_right[20] ,
    \_ces_3_1_io_outs_right[19] ,
    \_ces_3_1_io_outs_right[18] ,
    \_ces_3_1_io_outs_right[17] ,
    \_ces_3_1_io_outs_right[16] ,
    \_ces_3_1_io_outs_right[15] ,
    \_ces_3_1_io_outs_right[14] ,
    \_ces_3_1_io_outs_right[13] ,
    \_ces_3_1_io_outs_right[12] ,
    \_ces_3_1_io_outs_right[11] ,
    \_ces_3_1_io_outs_right[10] ,
    \_ces_3_1_io_outs_right[9] ,
    \_ces_3_1_io_outs_right[8] ,
    \_ces_3_1_io_outs_right[7] ,
    \_ces_3_1_io_outs_right[6] ,
    \_ces_3_1_io_outs_right[5] ,
    \_ces_3_1_io_outs_right[4] ,
    \_ces_3_1_io_outs_right[3] ,
    \_ces_3_1_io_outs_right[2] ,
    \_ces_3_1_io_outs_right[1] ,
    \_ces_3_1_io_outs_right[0] }),
    .io_ins_up({\_ces_2_2_io_outs_up[63] ,
    \_ces_2_2_io_outs_up[62] ,
    \_ces_2_2_io_outs_up[61] ,
    \_ces_2_2_io_outs_up[60] ,
    \_ces_2_2_io_outs_up[59] ,
    \_ces_2_2_io_outs_up[58] ,
    \_ces_2_2_io_outs_up[57] ,
    \_ces_2_2_io_outs_up[56] ,
    \_ces_2_2_io_outs_up[55] ,
    \_ces_2_2_io_outs_up[54] ,
    \_ces_2_2_io_outs_up[53] ,
    \_ces_2_2_io_outs_up[52] ,
    \_ces_2_2_io_outs_up[51] ,
    \_ces_2_2_io_outs_up[50] ,
    \_ces_2_2_io_outs_up[49] ,
    \_ces_2_2_io_outs_up[48] ,
    \_ces_2_2_io_outs_up[47] ,
    \_ces_2_2_io_outs_up[46] ,
    \_ces_2_2_io_outs_up[45] ,
    \_ces_2_2_io_outs_up[44] ,
    \_ces_2_2_io_outs_up[43] ,
    \_ces_2_2_io_outs_up[42] ,
    \_ces_2_2_io_outs_up[41] ,
    \_ces_2_2_io_outs_up[40] ,
    \_ces_2_2_io_outs_up[39] ,
    \_ces_2_2_io_outs_up[38] ,
    \_ces_2_2_io_outs_up[37] ,
    \_ces_2_2_io_outs_up[36] ,
    \_ces_2_2_io_outs_up[35] ,
    \_ces_2_2_io_outs_up[34] ,
    \_ces_2_2_io_outs_up[33] ,
    \_ces_2_2_io_outs_up[32] ,
    \_ces_2_2_io_outs_up[31] ,
    \_ces_2_2_io_outs_up[30] ,
    \_ces_2_2_io_outs_up[29] ,
    \_ces_2_2_io_outs_up[28] ,
    \_ces_2_2_io_outs_up[27] ,
    \_ces_2_2_io_outs_up[26] ,
    \_ces_2_2_io_outs_up[25] ,
    \_ces_2_2_io_outs_up[24] ,
    \_ces_2_2_io_outs_up[23] ,
    \_ces_2_2_io_outs_up[22] ,
    \_ces_2_2_io_outs_up[21] ,
    \_ces_2_2_io_outs_up[20] ,
    \_ces_2_2_io_outs_up[19] ,
    \_ces_2_2_io_outs_up[18] ,
    \_ces_2_2_io_outs_up[17] ,
    \_ces_2_2_io_outs_up[16] ,
    \_ces_2_2_io_outs_up[15] ,
    \_ces_2_2_io_outs_up[14] ,
    \_ces_2_2_io_outs_up[13] ,
    \_ces_2_2_io_outs_up[12] ,
    \_ces_2_2_io_outs_up[11] ,
    \_ces_2_2_io_outs_up[10] ,
    \_ces_2_2_io_outs_up[9] ,
    \_ces_2_2_io_outs_up[8] ,
    \_ces_2_2_io_outs_up[7] ,
    \_ces_2_2_io_outs_up[6] ,
    \_ces_2_2_io_outs_up[5] ,
    \_ces_2_2_io_outs_up[4] ,
    \_ces_2_2_io_outs_up[3] ,
    \_ces_2_2_io_outs_up[2] ,
    \_ces_2_2_io_outs_up[1] ,
    \_ces_2_2_io_outs_up[0] }),
    .io_outs_down({\_ces_3_2_io_outs_down[63] ,
    \_ces_3_2_io_outs_down[62] ,
    \_ces_3_2_io_outs_down[61] ,
    \_ces_3_2_io_outs_down[60] ,
    \_ces_3_2_io_outs_down[59] ,
    \_ces_3_2_io_outs_down[58] ,
    \_ces_3_2_io_outs_down[57] ,
    \_ces_3_2_io_outs_down[56] ,
    \_ces_3_2_io_outs_down[55] ,
    \_ces_3_2_io_outs_down[54] ,
    \_ces_3_2_io_outs_down[53] ,
    \_ces_3_2_io_outs_down[52] ,
    \_ces_3_2_io_outs_down[51] ,
    \_ces_3_2_io_outs_down[50] ,
    \_ces_3_2_io_outs_down[49] ,
    \_ces_3_2_io_outs_down[48] ,
    \_ces_3_2_io_outs_down[47] ,
    \_ces_3_2_io_outs_down[46] ,
    \_ces_3_2_io_outs_down[45] ,
    \_ces_3_2_io_outs_down[44] ,
    \_ces_3_2_io_outs_down[43] ,
    \_ces_3_2_io_outs_down[42] ,
    \_ces_3_2_io_outs_down[41] ,
    \_ces_3_2_io_outs_down[40] ,
    \_ces_3_2_io_outs_down[39] ,
    \_ces_3_2_io_outs_down[38] ,
    \_ces_3_2_io_outs_down[37] ,
    \_ces_3_2_io_outs_down[36] ,
    \_ces_3_2_io_outs_down[35] ,
    \_ces_3_2_io_outs_down[34] ,
    \_ces_3_2_io_outs_down[33] ,
    \_ces_3_2_io_outs_down[32] ,
    \_ces_3_2_io_outs_down[31] ,
    \_ces_3_2_io_outs_down[30] ,
    \_ces_3_2_io_outs_down[29] ,
    \_ces_3_2_io_outs_down[28] ,
    \_ces_3_2_io_outs_down[27] ,
    \_ces_3_2_io_outs_down[26] ,
    \_ces_3_2_io_outs_down[25] ,
    \_ces_3_2_io_outs_down[24] ,
    \_ces_3_2_io_outs_down[23] ,
    \_ces_3_2_io_outs_down[22] ,
    \_ces_3_2_io_outs_down[21] ,
    \_ces_3_2_io_outs_down[20] ,
    \_ces_3_2_io_outs_down[19] ,
    \_ces_3_2_io_outs_down[18] ,
    \_ces_3_2_io_outs_down[17] ,
    \_ces_3_2_io_outs_down[16] ,
    \_ces_3_2_io_outs_down[15] ,
    \_ces_3_2_io_outs_down[14] ,
    \_ces_3_2_io_outs_down[13] ,
    \_ces_3_2_io_outs_down[12] ,
    \_ces_3_2_io_outs_down[11] ,
    \_ces_3_2_io_outs_down[10] ,
    \_ces_3_2_io_outs_down[9] ,
    \_ces_3_2_io_outs_down[8] ,
    \_ces_3_2_io_outs_down[7] ,
    \_ces_3_2_io_outs_down[6] ,
    \_ces_3_2_io_outs_down[5] ,
    \_ces_3_2_io_outs_down[4] ,
    \_ces_3_2_io_outs_down[3] ,
    \_ces_3_2_io_outs_down[2] ,
    \_ces_3_2_io_outs_down[1] ,
    \_ces_3_2_io_outs_down[0] }),
    .io_outs_left({\_ces_3_2_io_outs_left[63] ,
    \_ces_3_2_io_outs_left[62] ,
    \_ces_3_2_io_outs_left[61] ,
    \_ces_3_2_io_outs_left[60] ,
    \_ces_3_2_io_outs_left[59] ,
    \_ces_3_2_io_outs_left[58] ,
    \_ces_3_2_io_outs_left[57] ,
    \_ces_3_2_io_outs_left[56] ,
    \_ces_3_2_io_outs_left[55] ,
    \_ces_3_2_io_outs_left[54] ,
    \_ces_3_2_io_outs_left[53] ,
    \_ces_3_2_io_outs_left[52] ,
    \_ces_3_2_io_outs_left[51] ,
    \_ces_3_2_io_outs_left[50] ,
    \_ces_3_2_io_outs_left[49] ,
    \_ces_3_2_io_outs_left[48] ,
    \_ces_3_2_io_outs_left[47] ,
    \_ces_3_2_io_outs_left[46] ,
    \_ces_3_2_io_outs_left[45] ,
    \_ces_3_2_io_outs_left[44] ,
    \_ces_3_2_io_outs_left[43] ,
    \_ces_3_2_io_outs_left[42] ,
    \_ces_3_2_io_outs_left[41] ,
    \_ces_3_2_io_outs_left[40] ,
    \_ces_3_2_io_outs_left[39] ,
    \_ces_3_2_io_outs_left[38] ,
    \_ces_3_2_io_outs_left[37] ,
    \_ces_3_2_io_outs_left[36] ,
    \_ces_3_2_io_outs_left[35] ,
    \_ces_3_2_io_outs_left[34] ,
    \_ces_3_2_io_outs_left[33] ,
    \_ces_3_2_io_outs_left[32] ,
    \_ces_3_2_io_outs_left[31] ,
    \_ces_3_2_io_outs_left[30] ,
    \_ces_3_2_io_outs_left[29] ,
    \_ces_3_2_io_outs_left[28] ,
    \_ces_3_2_io_outs_left[27] ,
    \_ces_3_2_io_outs_left[26] ,
    \_ces_3_2_io_outs_left[25] ,
    \_ces_3_2_io_outs_left[24] ,
    \_ces_3_2_io_outs_left[23] ,
    \_ces_3_2_io_outs_left[22] ,
    \_ces_3_2_io_outs_left[21] ,
    \_ces_3_2_io_outs_left[20] ,
    \_ces_3_2_io_outs_left[19] ,
    \_ces_3_2_io_outs_left[18] ,
    \_ces_3_2_io_outs_left[17] ,
    \_ces_3_2_io_outs_left[16] ,
    \_ces_3_2_io_outs_left[15] ,
    \_ces_3_2_io_outs_left[14] ,
    \_ces_3_2_io_outs_left[13] ,
    \_ces_3_2_io_outs_left[12] ,
    \_ces_3_2_io_outs_left[11] ,
    \_ces_3_2_io_outs_left[10] ,
    \_ces_3_2_io_outs_left[9] ,
    \_ces_3_2_io_outs_left[8] ,
    \_ces_3_2_io_outs_left[7] ,
    \_ces_3_2_io_outs_left[6] ,
    \_ces_3_2_io_outs_left[5] ,
    \_ces_3_2_io_outs_left[4] ,
    \_ces_3_2_io_outs_left[3] ,
    \_ces_3_2_io_outs_left[2] ,
    \_ces_3_2_io_outs_left[1] ,
    \_ces_3_2_io_outs_left[0] }),
    .io_outs_right({\_ces_3_2_io_outs_right[63] ,
    \_ces_3_2_io_outs_right[62] ,
    \_ces_3_2_io_outs_right[61] ,
    \_ces_3_2_io_outs_right[60] ,
    \_ces_3_2_io_outs_right[59] ,
    \_ces_3_2_io_outs_right[58] ,
    \_ces_3_2_io_outs_right[57] ,
    \_ces_3_2_io_outs_right[56] ,
    \_ces_3_2_io_outs_right[55] ,
    \_ces_3_2_io_outs_right[54] ,
    \_ces_3_2_io_outs_right[53] ,
    \_ces_3_2_io_outs_right[52] ,
    \_ces_3_2_io_outs_right[51] ,
    \_ces_3_2_io_outs_right[50] ,
    \_ces_3_2_io_outs_right[49] ,
    \_ces_3_2_io_outs_right[48] ,
    \_ces_3_2_io_outs_right[47] ,
    \_ces_3_2_io_outs_right[46] ,
    \_ces_3_2_io_outs_right[45] ,
    \_ces_3_2_io_outs_right[44] ,
    \_ces_3_2_io_outs_right[43] ,
    \_ces_3_2_io_outs_right[42] ,
    \_ces_3_2_io_outs_right[41] ,
    \_ces_3_2_io_outs_right[40] ,
    \_ces_3_2_io_outs_right[39] ,
    \_ces_3_2_io_outs_right[38] ,
    \_ces_3_2_io_outs_right[37] ,
    \_ces_3_2_io_outs_right[36] ,
    \_ces_3_2_io_outs_right[35] ,
    \_ces_3_2_io_outs_right[34] ,
    \_ces_3_2_io_outs_right[33] ,
    \_ces_3_2_io_outs_right[32] ,
    \_ces_3_2_io_outs_right[31] ,
    \_ces_3_2_io_outs_right[30] ,
    \_ces_3_2_io_outs_right[29] ,
    \_ces_3_2_io_outs_right[28] ,
    \_ces_3_2_io_outs_right[27] ,
    \_ces_3_2_io_outs_right[26] ,
    \_ces_3_2_io_outs_right[25] ,
    \_ces_3_2_io_outs_right[24] ,
    \_ces_3_2_io_outs_right[23] ,
    \_ces_3_2_io_outs_right[22] ,
    \_ces_3_2_io_outs_right[21] ,
    \_ces_3_2_io_outs_right[20] ,
    \_ces_3_2_io_outs_right[19] ,
    \_ces_3_2_io_outs_right[18] ,
    \_ces_3_2_io_outs_right[17] ,
    \_ces_3_2_io_outs_right[16] ,
    \_ces_3_2_io_outs_right[15] ,
    \_ces_3_2_io_outs_right[14] ,
    \_ces_3_2_io_outs_right[13] ,
    \_ces_3_2_io_outs_right[12] ,
    \_ces_3_2_io_outs_right[11] ,
    \_ces_3_2_io_outs_right[10] ,
    \_ces_3_2_io_outs_right[9] ,
    \_ces_3_2_io_outs_right[8] ,
    \_ces_3_2_io_outs_right[7] ,
    \_ces_3_2_io_outs_right[6] ,
    \_ces_3_2_io_outs_right[5] ,
    \_ces_3_2_io_outs_right[4] ,
    \_ces_3_2_io_outs_right[3] ,
    \_ces_3_2_io_outs_right[2] ,
    \_ces_3_2_io_outs_right[1] ,
    \_ces_3_2_io_outs_right[0] }),
    .io_outs_up({net2007,
    net2006,
    net2005,
    net2004,
    net2002,
    net2001,
    net2000,
    net1999,
    net1998,
    net1997,
    net1996,
    net1995,
    net1994,
    net1993,
    net1991,
    net1990,
    net1989,
    net1988,
    net1987,
    net1986,
    net1985,
    net1984,
    net1983,
    net1982,
    net1980,
    net1979,
    net1978,
    net1977,
    net1976,
    net1975,
    net1974,
    net1973,
    net1972,
    net1971,
    net1969,
    net1968,
    net1967,
    net1966,
    net1965,
    net1964,
    net1963,
    net1962,
    net1961,
    net1960,
    net1958,
    net1957,
    net1956,
    net1955,
    net1954,
    net1953,
    net1952,
    net1951,
    net1950,
    net1949,
    net2011,
    net2010,
    net2009,
    net2008,
    net2003,
    net1992,
    net1981,
    net1970,
    net1959,
    net1948}));
 Element ces_3_3 (.clock(clknet_leaf_1_clock),
    .io_lsbIns_1(_ces_3_2_io_lsbOuts_1),
    .io_lsbIns_2(_ces_3_2_io_lsbOuts_2),
    .io_lsbIns_3(_ces_3_2_io_lsbOuts_3),
    .io_lsbOuts_0(_ces_3_3_io_lsbOuts_0),
    .io_lsbOuts_1(_ces_3_3_io_lsbOuts_1),
    .io_lsbOuts_2(_ces_3_3_io_lsbOuts_2),
    .io_lsbOuts_3(_ces_3_3_io_lsbOuts_3),
    .io_ins_down({net263,
    net262,
    net261,
    net260,
    net258,
    net257,
    net256,
    net255,
    net254,
    net253,
    net252,
    net251,
    net250,
    net249,
    net247,
    net246,
    net245,
    net244,
    net243,
    net242,
    net241,
    net240,
    net239,
    net238,
    net236,
    net235,
    net234,
    net233,
    net232,
    net231,
    net230,
    net229,
    net228,
    net227,
    net225,
    net224,
    net223,
    net222,
    net221,
    net220,
    net219,
    net218,
    net217,
    net216,
    net214,
    net213,
    net212,
    net211,
    net210,
    net209,
    net208,
    net207,
    net206,
    net205,
    net267,
    net266,
    net265,
    net264,
    net259,
    net248,
    net237,
    net226,
    net215,
    net204}),
    .io_ins_left({net519,
    net518,
    net517,
    net516,
    net514,
    net513,
    net512,
    net511,
    net510,
    net509,
    net508,
    net507,
    net506,
    net505,
    net503,
    net502,
    net501,
    net500,
    net499,
    net498,
    net497,
    net496,
    net495,
    net494,
    net492,
    net491,
    net490,
    net489,
    net488,
    net487,
    net486,
    net485,
    net484,
    net483,
    net481,
    net480,
    net479,
    net478,
    net477,
    net476,
    net475,
    net474,
    net473,
    net472,
    net470,
    net469,
    net468,
    net467,
    net466,
    net465,
    net464,
    net463,
    net462,
    net461,
    net523,
    net522,
    net521,
    net520,
    net515,
    net504,
    net493,
    net482,
    net471,
    net460}),
    .io_ins_right({\_ces_3_2_io_outs_right[63] ,
    \_ces_3_2_io_outs_right[62] ,
    \_ces_3_2_io_outs_right[61] ,
    \_ces_3_2_io_outs_right[60] ,
    \_ces_3_2_io_outs_right[59] ,
    \_ces_3_2_io_outs_right[58] ,
    \_ces_3_2_io_outs_right[57] ,
    \_ces_3_2_io_outs_right[56] ,
    \_ces_3_2_io_outs_right[55] ,
    \_ces_3_2_io_outs_right[54] ,
    \_ces_3_2_io_outs_right[53] ,
    \_ces_3_2_io_outs_right[52] ,
    \_ces_3_2_io_outs_right[51] ,
    \_ces_3_2_io_outs_right[50] ,
    \_ces_3_2_io_outs_right[49] ,
    \_ces_3_2_io_outs_right[48] ,
    \_ces_3_2_io_outs_right[47] ,
    \_ces_3_2_io_outs_right[46] ,
    \_ces_3_2_io_outs_right[45] ,
    \_ces_3_2_io_outs_right[44] ,
    \_ces_3_2_io_outs_right[43] ,
    \_ces_3_2_io_outs_right[42] ,
    \_ces_3_2_io_outs_right[41] ,
    \_ces_3_2_io_outs_right[40] ,
    \_ces_3_2_io_outs_right[39] ,
    \_ces_3_2_io_outs_right[38] ,
    \_ces_3_2_io_outs_right[37] ,
    \_ces_3_2_io_outs_right[36] ,
    \_ces_3_2_io_outs_right[35] ,
    \_ces_3_2_io_outs_right[34] ,
    \_ces_3_2_io_outs_right[33] ,
    \_ces_3_2_io_outs_right[32] ,
    \_ces_3_2_io_outs_right[31] ,
    \_ces_3_2_io_outs_right[30] ,
    \_ces_3_2_io_outs_right[29] ,
    \_ces_3_2_io_outs_right[28] ,
    \_ces_3_2_io_outs_right[27] ,
    \_ces_3_2_io_outs_right[26] ,
    \_ces_3_2_io_outs_right[25] ,
    \_ces_3_2_io_outs_right[24] ,
    \_ces_3_2_io_outs_right[23] ,
    \_ces_3_2_io_outs_right[22] ,
    \_ces_3_2_io_outs_right[21] ,
    \_ces_3_2_io_outs_right[20] ,
    \_ces_3_2_io_outs_right[19] ,
    \_ces_3_2_io_outs_right[18] ,
    \_ces_3_2_io_outs_right[17] ,
    \_ces_3_2_io_outs_right[16] ,
    \_ces_3_2_io_outs_right[15] ,
    \_ces_3_2_io_outs_right[14] ,
    \_ces_3_2_io_outs_right[13] ,
    \_ces_3_2_io_outs_right[12] ,
    \_ces_3_2_io_outs_right[11] ,
    \_ces_3_2_io_outs_right[10] ,
    \_ces_3_2_io_outs_right[9] ,
    \_ces_3_2_io_outs_right[8] ,
    \_ces_3_2_io_outs_right[7] ,
    \_ces_3_2_io_outs_right[6] ,
    \_ces_3_2_io_outs_right[5] ,
    \_ces_3_2_io_outs_right[4] ,
    \_ces_3_2_io_outs_right[3] ,
    \_ces_3_2_io_outs_right[2] ,
    \_ces_3_2_io_outs_right[1] ,
    \_ces_3_2_io_outs_right[0] }),
    .io_ins_up({\_ces_2_3_io_outs_up[63] ,
    \_ces_2_3_io_outs_up[62] ,
    \_ces_2_3_io_outs_up[61] ,
    \_ces_2_3_io_outs_up[60] ,
    \_ces_2_3_io_outs_up[59] ,
    \_ces_2_3_io_outs_up[58] ,
    \_ces_2_3_io_outs_up[57] ,
    \_ces_2_3_io_outs_up[56] ,
    \_ces_2_3_io_outs_up[55] ,
    \_ces_2_3_io_outs_up[54] ,
    \_ces_2_3_io_outs_up[53] ,
    \_ces_2_3_io_outs_up[52] ,
    \_ces_2_3_io_outs_up[51] ,
    \_ces_2_3_io_outs_up[50] ,
    \_ces_2_3_io_outs_up[49] ,
    \_ces_2_3_io_outs_up[48] ,
    \_ces_2_3_io_outs_up[47] ,
    \_ces_2_3_io_outs_up[46] ,
    \_ces_2_3_io_outs_up[45] ,
    \_ces_2_3_io_outs_up[44] ,
    \_ces_2_3_io_outs_up[43] ,
    \_ces_2_3_io_outs_up[42] ,
    \_ces_2_3_io_outs_up[41] ,
    \_ces_2_3_io_outs_up[40] ,
    \_ces_2_3_io_outs_up[39] ,
    \_ces_2_3_io_outs_up[38] ,
    \_ces_2_3_io_outs_up[37] ,
    \_ces_2_3_io_outs_up[36] ,
    \_ces_2_3_io_outs_up[35] ,
    \_ces_2_3_io_outs_up[34] ,
    \_ces_2_3_io_outs_up[33] ,
    \_ces_2_3_io_outs_up[32] ,
    \_ces_2_3_io_outs_up[31] ,
    \_ces_2_3_io_outs_up[30] ,
    \_ces_2_3_io_outs_up[29] ,
    \_ces_2_3_io_outs_up[28] ,
    \_ces_2_3_io_outs_up[27] ,
    \_ces_2_3_io_outs_up[26] ,
    \_ces_2_3_io_outs_up[25] ,
    \_ces_2_3_io_outs_up[24] ,
    \_ces_2_3_io_outs_up[23] ,
    \_ces_2_3_io_outs_up[22] ,
    \_ces_2_3_io_outs_up[21] ,
    \_ces_2_3_io_outs_up[20] ,
    \_ces_2_3_io_outs_up[19] ,
    \_ces_2_3_io_outs_up[18] ,
    \_ces_2_3_io_outs_up[17] ,
    \_ces_2_3_io_outs_up[16] ,
    \_ces_2_3_io_outs_up[15] ,
    \_ces_2_3_io_outs_up[14] ,
    \_ces_2_3_io_outs_up[13] ,
    \_ces_2_3_io_outs_up[12] ,
    \_ces_2_3_io_outs_up[11] ,
    \_ces_2_3_io_outs_up[10] ,
    \_ces_2_3_io_outs_up[9] ,
    \_ces_2_3_io_outs_up[8] ,
    \_ces_2_3_io_outs_up[7] ,
    \_ces_2_3_io_outs_up[6] ,
    \_ces_2_3_io_outs_up[5] ,
    \_ces_2_3_io_outs_up[4] ,
    \_ces_2_3_io_outs_up[3] ,
    \_ces_2_3_io_outs_up[2] ,
    \_ces_2_3_io_outs_up[1] ,
    \_ces_2_3_io_outs_up[0] }),
    .io_outs_down({\_ces_3_3_io_outs_down[63] ,
    \_ces_3_3_io_outs_down[62] ,
    \_ces_3_3_io_outs_down[61] ,
    \_ces_3_3_io_outs_down[60] ,
    \_ces_3_3_io_outs_down[59] ,
    \_ces_3_3_io_outs_down[58] ,
    \_ces_3_3_io_outs_down[57] ,
    \_ces_3_3_io_outs_down[56] ,
    \_ces_3_3_io_outs_down[55] ,
    \_ces_3_3_io_outs_down[54] ,
    \_ces_3_3_io_outs_down[53] ,
    \_ces_3_3_io_outs_down[52] ,
    \_ces_3_3_io_outs_down[51] ,
    \_ces_3_3_io_outs_down[50] ,
    \_ces_3_3_io_outs_down[49] ,
    \_ces_3_3_io_outs_down[48] ,
    \_ces_3_3_io_outs_down[47] ,
    \_ces_3_3_io_outs_down[46] ,
    \_ces_3_3_io_outs_down[45] ,
    \_ces_3_3_io_outs_down[44] ,
    \_ces_3_3_io_outs_down[43] ,
    \_ces_3_3_io_outs_down[42] ,
    \_ces_3_3_io_outs_down[41] ,
    \_ces_3_3_io_outs_down[40] ,
    \_ces_3_3_io_outs_down[39] ,
    \_ces_3_3_io_outs_down[38] ,
    \_ces_3_3_io_outs_down[37] ,
    \_ces_3_3_io_outs_down[36] ,
    \_ces_3_3_io_outs_down[35] ,
    \_ces_3_3_io_outs_down[34] ,
    \_ces_3_3_io_outs_down[33] ,
    \_ces_3_3_io_outs_down[32] ,
    \_ces_3_3_io_outs_down[31] ,
    \_ces_3_3_io_outs_down[30] ,
    \_ces_3_3_io_outs_down[29] ,
    \_ces_3_3_io_outs_down[28] ,
    \_ces_3_3_io_outs_down[27] ,
    \_ces_3_3_io_outs_down[26] ,
    \_ces_3_3_io_outs_down[25] ,
    \_ces_3_3_io_outs_down[24] ,
    \_ces_3_3_io_outs_down[23] ,
    \_ces_3_3_io_outs_down[22] ,
    \_ces_3_3_io_outs_down[21] ,
    \_ces_3_3_io_outs_down[20] ,
    \_ces_3_3_io_outs_down[19] ,
    \_ces_3_3_io_outs_down[18] ,
    \_ces_3_3_io_outs_down[17] ,
    \_ces_3_3_io_outs_down[16] ,
    \_ces_3_3_io_outs_down[15] ,
    \_ces_3_3_io_outs_down[14] ,
    \_ces_3_3_io_outs_down[13] ,
    \_ces_3_3_io_outs_down[12] ,
    \_ces_3_3_io_outs_down[11] ,
    \_ces_3_3_io_outs_down[10] ,
    \_ces_3_3_io_outs_down[9] ,
    \_ces_3_3_io_outs_down[8] ,
    \_ces_3_3_io_outs_down[7] ,
    \_ces_3_3_io_outs_down[6] ,
    \_ces_3_3_io_outs_down[5] ,
    \_ces_3_3_io_outs_down[4] ,
    \_ces_3_3_io_outs_down[3] ,
    \_ces_3_3_io_outs_down[2] ,
    \_ces_3_3_io_outs_down[1] ,
    \_ces_3_3_io_outs_down[0] }),
    .io_outs_left({\_ces_3_3_io_outs_left[63] ,
    \_ces_3_3_io_outs_left[62] ,
    \_ces_3_3_io_outs_left[61] ,
    \_ces_3_3_io_outs_left[60] ,
    \_ces_3_3_io_outs_left[59] ,
    \_ces_3_3_io_outs_left[58] ,
    \_ces_3_3_io_outs_left[57] ,
    \_ces_3_3_io_outs_left[56] ,
    \_ces_3_3_io_outs_left[55] ,
    \_ces_3_3_io_outs_left[54] ,
    \_ces_3_3_io_outs_left[53] ,
    \_ces_3_3_io_outs_left[52] ,
    \_ces_3_3_io_outs_left[51] ,
    \_ces_3_3_io_outs_left[50] ,
    \_ces_3_3_io_outs_left[49] ,
    \_ces_3_3_io_outs_left[48] ,
    \_ces_3_3_io_outs_left[47] ,
    \_ces_3_3_io_outs_left[46] ,
    \_ces_3_3_io_outs_left[45] ,
    \_ces_3_3_io_outs_left[44] ,
    \_ces_3_3_io_outs_left[43] ,
    \_ces_3_3_io_outs_left[42] ,
    \_ces_3_3_io_outs_left[41] ,
    \_ces_3_3_io_outs_left[40] ,
    \_ces_3_3_io_outs_left[39] ,
    \_ces_3_3_io_outs_left[38] ,
    \_ces_3_3_io_outs_left[37] ,
    \_ces_3_3_io_outs_left[36] ,
    \_ces_3_3_io_outs_left[35] ,
    \_ces_3_3_io_outs_left[34] ,
    \_ces_3_3_io_outs_left[33] ,
    \_ces_3_3_io_outs_left[32] ,
    \_ces_3_3_io_outs_left[31] ,
    \_ces_3_3_io_outs_left[30] ,
    \_ces_3_3_io_outs_left[29] ,
    \_ces_3_3_io_outs_left[28] ,
    \_ces_3_3_io_outs_left[27] ,
    \_ces_3_3_io_outs_left[26] ,
    \_ces_3_3_io_outs_left[25] ,
    \_ces_3_3_io_outs_left[24] ,
    \_ces_3_3_io_outs_left[23] ,
    \_ces_3_3_io_outs_left[22] ,
    \_ces_3_3_io_outs_left[21] ,
    \_ces_3_3_io_outs_left[20] ,
    \_ces_3_3_io_outs_left[19] ,
    \_ces_3_3_io_outs_left[18] ,
    \_ces_3_3_io_outs_left[17] ,
    \_ces_3_3_io_outs_left[16] ,
    \_ces_3_3_io_outs_left[15] ,
    \_ces_3_3_io_outs_left[14] ,
    \_ces_3_3_io_outs_left[13] ,
    \_ces_3_3_io_outs_left[12] ,
    \_ces_3_3_io_outs_left[11] ,
    \_ces_3_3_io_outs_left[10] ,
    \_ces_3_3_io_outs_left[9] ,
    \_ces_3_3_io_outs_left[8] ,
    \_ces_3_3_io_outs_left[7] ,
    \_ces_3_3_io_outs_left[6] ,
    \_ces_3_3_io_outs_left[5] ,
    \_ces_3_3_io_outs_left[4] ,
    \_ces_3_3_io_outs_left[3] ,
    \_ces_3_3_io_outs_left[2] ,
    \_ces_3_3_io_outs_left[1] ,
    \_ces_3_3_io_outs_left[0] }),
    .io_outs_right({net1815,
    net1814,
    net1813,
    net1812,
    net1810,
    net1809,
    net1808,
    net1807,
    net1806,
    net1805,
    net1804,
    net1803,
    net1802,
    net1801,
    net1799,
    net1798,
    net1797,
    net1796,
    net1795,
    net1794,
    net1793,
    net1792,
    net1791,
    net1790,
    net1788,
    net1787,
    net1786,
    net1785,
    net1784,
    net1783,
    net1782,
    net1781,
    net1780,
    net1779,
    net1777,
    net1776,
    net1775,
    net1774,
    net1773,
    net1772,
    net1771,
    net1770,
    net1769,
    net1768,
    net1766,
    net1765,
    net1764,
    net1763,
    net1762,
    net1761,
    net1760,
    net1759,
    net1758,
    net1757,
    net1819,
    net1818,
    net1817,
    net1816,
    net1811,
    net1800,
    net1789,
    net1778,
    net1767,
    net1756}),
    .io_outs_up({net2071,
    net2070,
    net2069,
    net2068,
    net2066,
    net2065,
    net2064,
    net2063,
    net2062,
    net2061,
    net2060,
    net2059,
    net2058,
    net2057,
    net2055,
    net2054,
    net2053,
    net2052,
    net2051,
    net2050,
    net2049,
    net2048,
    net2047,
    net2046,
    net2044,
    net2043,
    net2042,
    net2041,
    net2040,
    net2039,
    net2038,
    net2037,
    net2036,
    net2035,
    net2033,
    net2032,
    net2031,
    net2030,
    net2029,
    net2028,
    net2027,
    net2026,
    net2025,
    net2024,
    net2022,
    net2021,
    net2020,
    net2019,
    net2018,
    net2017,
    net2016,
    net2015,
    net2014,
    net2013,
    net2075,
    net2074,
    net2073,
    net2072,
    net2067,
    net2056,
    net2045,
    net2034,
    net2023,
    net2012}));
endmodule
