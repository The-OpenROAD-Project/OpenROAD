VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 2000 ;
END UNITS

MACRO ENDCAP_X4_LEFTBOTTOMCORNER_Y
  PROPERTY LEF58_CLASS " CLASS ENDCAP LEFTBOTTOMCORNER ; " ;
  ORIGIN 0 0 ;
  FOREIGN ENDCAP_X4 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.76 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.76 0.085 ;
    END
  END VSS
END ENDCAP_X4_LEFTBOTTOMCORNER_Y

MACRO ENDCAP_X4_LEFTTOPCORNER_Y
  PROPERTY LEF58_CLASS " CLASS ENDCAP LEFTTOPCORNER ; " ;
  ORIGIN 0 0 ;
  FOREIGN ENDCAP_X4 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.76 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.76 0.085 ;
    END
  END VSS
END ENDCAP_X4_LEFTTOPCORNER_Y

MACRO ENDCAP_X4_LEFTBOTTOMEDGE_Y
  PROPERTY LEF58_CLASS " CLASS ENDCAP LEFTBOTTOMEDGE ; " ;
  ORIGIN 0 0 ;
  FOREIGN ENDCAP_X4 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.76 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.76 0.085 ;
    END
  END VSS
END ENDCAP_X4_LEFTBOTTOMEDGE_Y

MACRO ENDCAP_X4_LEFTTOPEDGE_Y
  PROPERTY LEF58_CLASS " CLASS ENDCAP LEFTTOPEDGE ; " ;
  ORIGIN 0 0 ;
  FOREIGN ENDCAP_X4 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.76 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.76 0.085 ;
    END
  END VSS
END ENDCAP_X4_LEFTTOPEDGE_Y

MACRO ENDCAP_X4_RIGHTEDGE_Y
  PROPERTY LEF58_CLASS " CLASS ENDCAP RIGHTEDGE ; " ;
  ORIGIN 0 0 ;
  FOREIGN ENDCAP_X4 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.76 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.76 0.085 ;
    END
  END VSS
END ENDCAP_X4_RIGHTEDGE_Y

END LIBRARY
#
# End of file
#
