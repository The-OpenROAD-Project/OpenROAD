VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO SLC
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SLC 0 0 ;
  SIZE 13.34 BY 2.72 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.95 0.85 2.12 1.18 ;
    END
  END IN
  PIN INB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.28 1.225 9.71 1.395 ;
    END
  END INB
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 13.34 0.24 ;
      LAYER li1 ;
        RECT 0 -0.085 13.34 0.085 ;
        RECT 11.595 -0.085 11.845 0.635 ;
        RECT 10.715 -0.085 10.965 0.635 ;
        RECT 9.835 -0.085 10.085 0.635 ;
        RECT 8.955 -0.085 9.205 0.635 ;
        RECT 8.075 -0.085 8.325 0.635 ;
        RECT 7.195 -0.085 7.445 0.635 ;
        RECT 6.565 -0.085 6.815 0.635 ;
        RECT 5.685 -0.085 5.935 0.635 ;
        RECT 4.805 -0.085 5.055 0.635 ;
        RECT 3.925 -0.085 4.175 0.635 ;
        RECT 3.045 -0.085 3.295 0.635 ;
        RECT 2.165 -0.085 2.415 0.635 ;
        RECT 1.53 -0.085 1.78 0.635 ;
      LAYER mcon ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 12.505 0.265 12.795 0.81 ;
        RECT 0.545 0.265 0.835 0.81 ;
    END
  END VNB
  PIN VOUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.32 1.835 2.57 2.4 ;
        RECT 1.01 1.835 2.57 2.005 ;
        RECT 1.01 0.305 1.26 1.195 ;
        RECT 1.01 0.305 1.18 2.005 ;
    END
  END VOUT
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 12.505 1.47 12.795 2.455 ;
        RECT 0.545 1.47 0.835 2.455 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 13.34 2.96 ;
      LAYER li1 ;
        RECT 0 2.635 13.34 2.805 ;
        RECT 5.715 2.085 5.965 2.805 ;
        RECT 4.805 2.085 5.055 2.805 ;
        RECT 2.76 2.175 3.01 2.805 ;
        RECT 1.88 2.175 2.13 2.805 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
    END
  END VPWR
  OBS
    LAYER mcon ;
      RECT 3.345 1.165 3.515 1.335 ;
      RECT 3.345 2.085 3.515 2.255 ;
    LAYER met1 ;
      RECT 3.285 2.055 3.575 2.285 ;
      RECT 3.36 1.135 3.5 2.285 ;
      RECT 3.285 1.135 3.575 1.365 ;
    LAYER li1 ;
      RECT 6.675 1.665 6.885 2.425 ;
      RECT 4.67 1.665 7.84 1.835 ;
      RECT 7.635 0.305 7.84 1.835 ;
      RECT 7.42 1.505 7.84 1.835 ;
      RECT 4.67 1.505 4.92 1.835 ;
      RECT 7.635 0.805 11.855 0.975 ;
      RECT 11.155 0.305 11.405 0.975 ;
      RECT 10.275 0.305 10.525 0.975 ;
      RECT 9.395 0.305 9.645 0.975 ;
      RECT 8.515 0.305 8.765 0.975 ;
      RECT 7.635 0.305 7.885 0.975 ;
      RECT 1.35 1.415 2.46 1.585 ;
      RECT 2.29 1.165 2.46 1.585 ;
      RECT 5.825 1.165 6.175 1.46 ;
      RECT 3.975 1.165 4.305 1.46 ;
      RECT 2.29 1.165 6.175 1.335 ;
      RECT 3.345 0.805 3.515 1.335 ;
      RECT 2.605 0.805 6.955 0.975 ;
      RECT 6.125 0.305 6.375 0.975 ;
      RECT 5.245 0.305 5.495 0.975 ;
      RECT 4.365 0.305 4.615 0.975 ;
      RECT 3.485 0.305 3.735 0.975 ;
      RECT 2.605 0.305 2.855 0.975 ;
      RECT 4.285 2.085 4.535 2.425 ;
      RECT 4.285 1.745 4.455 2.425 ;
      RECT 3.01 1.745 4.455 1.915 ;
      RECT 3.01 1.515 3.18 1.915 ;
      RECT 2.74 1.515 3.18 1.685 ;
      RECT 3.845 2.085 4.095 2.425 ;
      RECT 3.285 2.085 4.095 2.255 ;
  END
END SLC

END LIBRARY
