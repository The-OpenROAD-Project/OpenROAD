module multi_sink (clk);
 input clk;

 wire gclk1;
 wire gclk3;
 wire gclk4;


 CLKGATE_X1 gclk1 (.CK(clk), .GCK(gclk1));
   DFF_X1 ff278 (.CK(gclk1));
   DFF_X1 ff277 (.CK(gclk1));
   DFF_X1 ff276 (.CK(gclk1));
   DFF_X1 ff275 (.CK(gclk1));
   DFF_X1 ff274 (.CK(gclk1));
   DFF_X1 ff273 (.CK(gclk1));
   DFF_X1 ff272 (.CK(gclk1));
   DFF_X1 ff271 (.CK(gclk1));
   DFF_X1 ff270 (.CK(gclk1));
   DFF_X1 ff260 (.CK(gclk1));
   DFF_X1 ff259 (.CK(gclk1));
   DFF_X1 ff258 (.CK(gclk1));
   DFF_X1 ff257 (.CK(gclk1));
   DFF_X1 ff256 (.CK(gclk1));
   DFF_X1 ff255 (.CK(gclk1));
   DFF_X1 ff254 (.CK(gclk1));
   DFF_X1 ff253 (.CK(gclk1));
   DFF_X1 ff252 (.CK(gclk1));
   DFF_X1 ff242 (.CK(gclk1));
   DFF_X1 ff241 (.CK(gclk1));
   DFF_X1 ff240 (.CK(gclk1));
   DFF_X1 ff239 (.CK(gclk1));
   DFF_X1 ff238 (.CK(gclk1));
   DFF_X1 ff237 (.CK(gclk1));
   DFF_X1 ff236 (.CK(gclk1));
   DFF_X1 ff235 (.CK(gclk1));
   DFF_X1 ff234 (.CK(gclk1));
   DFF_X1 ff224 (.CK(gclk1));
   DFF_X1 ff223 (.CK(gclk1));
   DFF_X1 ff222 (.CK(gclk1));
   DFF_X1 ff221 (.CK(gclk1));
   DFF_X1 ff220 (.CK(gclk1));
   DFF_X1 ff219 (.CK(gclk1));
   DFF_X1 ff218 (.CK(gclk1));
   DFF_X1 ff217 (.CK(gclk1));
   DFF_X1 ff216 (.CK(gclk1));
 CLKGATE_X1 gclk3 (.CK(gclk4), .GCK(gclk3));
 DFF_X1 ff287 (.CK(gclk3));
 DFF_X1 ff286 (.CK(gclk3));
 DFF_X1 ff285 (.CK(gclk3));
 DFF_X1 ff284 (.CK(gclk3));
 DFF_X1 ff283 (.CK(gclk3));
 DFF_X1 ff282 (.CK(gclk3));
 DFF_X1 ff281 (.CK(gclk3));
 DFF_X1 ff280 (.CK(gclk3));
 DFF_X1 ff279 (.CK(gclk3));
 DFF_X1 ff269 (.CK(gclk3));
 DFF_X1 ff268 (.CK(gclk3));
 DFF_X1 ff267 (.CK(gclk3));
 DFF_X1 ff266 (.CK(gclk3));
 DFF_X1 ff265 (.CK(gclk3));
 DFF_X1 ff264 (.CK(gclk3));
 DFF_X1 ff263 (.CK(gclk3));
 DFF_X1 ff262 (.CK(gclk3));
 DFF_X1 ff261 (.CK(gclk3));
 DFF_X1 ff251 (.CK(gclk3));
 DFF_X1 ff250 (.CK(gclk3));
 DFF_X1 ff249 (.CK(gclk3));
 DFF_X1 ff248 (.CK(gclk3));
 DFF_X1 ff247 (.CK(gclk3));
 DFF_X1 ff246 (.CK(gclk3));
 DFF_X1 ff245 (.CK(gclk3));
 DFF_X1 ff244 (.CK(gclk3));
 DFF_X1 ff243 (.CK(gclk3));
 DFF_X1 ff233 (.CK(gclk3));
 DFF_X1 ff232 (.CK(gclk3));
 DFF_X1 ff231 (.CK(gclk3));
 DFF_X1 ff230 (.CK(gclk3));
 DFF_X1 ff229 (.CK(gclk3));
 DFF_X1 ff228 (.CK(gclk3));
 DFF_X1 ff227 (.CK(gclk3));
 DFF_X1 ff226 (.CK(gclk3));
 DFF_X1 ff225 (.CK(gclk3));
 CLKGATE_X1 gclk4 (.CK(clk), .GCK(gclk4));
 DFF_X1 ff197 (.CK(gclk4));
 DFF_X1 ff196 (.CK(gclk4));
 DFF_X1 ff195 (.CK(gclk4));
 DFF_X1 ff194 (.CK(gclk4));
 DFF_X1 ff193 (.CK(gclk4));
 DFF_X1 ff192 (.CK(gclk4));
 DFF_X1 ff191 (.CK(gclk4));
 DFF_X1 ff190 (.CK(gclk4));
 DFF_X1 ff189 (.CK(gclk4));
 DFF_X1 ff179 (.CK(gclk4));
 DFF_X1 ff178 (.CK(gclk4));
 DFF_X1 ff177 (.CK(gclk4));
 DFF_X1 ff176 (.CK(gclk4));
 DFF_X1 ff175 (.CK(gclk4));
 DFF_X1 ff174 (.CK(gclk4));
 DFF_X1 ff173 (.CK(gclk4));
 DFF_X1 ff172 (.CK(gclk4));
 DFF_X1 ff171 (.CK(gclk4));
 DFF_X1 ff161 (.CK(gclk4));
 DFF_X1 ff160 (.CK(gclk4));
 DFF_X1 ff159 (.CK(gclk4));
 DFF_X1 ff158 (.CK(gclk4));
 DFF_X1 ff157 (.CK(gclk4));
 DFF_X1 ff156 (.CK(gclk4));
 DFF_X1 ff155 (.CK(gclk4));
 DFF_X1 ff154 (.CK(gclk4));
 DFF_X1 ff153 (.CK(gclk4));
 DFF_X1 ff215 (.CK(gclk4));
 DFF_X1 ff214 (.CK(gclk4));
 DFF_X1 ff213 (.CK(gclk4));
 DFF_X1 ff212 (.CK(gclk4));
 DFF_X1 ff211 (.CK(gclk4));
 DFF_X1 ff210 (.CK(gclk4));
 DFF_X1 ff209 (.CK(gclk4));
 DFF_X1 ff208 (.CK(gclk4));
 DFF_X1 ff207 (.CK(gclk4));

 wire hi_gclk2;
 wire hi_gclk5;

 CLKGATE_X1 \hi_inst/gclk2_inst (.CK(clk), .GCK(hi_gclk2));
 DFF_X1 \h1/ff152 (.CK(hi_gclk2));
 DFF_X1 \h1/ff151 (.CK(hi_gclk2));
 DFF_X1 \h1/ff150 (.CK(hi_gclk2));
 DFF_X1 \h1/ff149 (.CK(hi_gclk2));
 DFF_X1 \h1/ff148 (.CK(hi_gclk2));
 DFF_X1 \h1/ff147 (.CK(hi_gclk2));
 DFF_X1 \h1/ff146 (.CK(hi_gclk2));
 DFF_X1 \h1/ff145 (.CK(hi_gclk2));
 DFF_X1 \h1/ff144 (.CK(hi_gclk2));
 DFF_X1 \h1/ff170 (.CK(hi_gclk2));
 DFF_X1 \h1/ff169 (.CK(hi_gclk2));
 DFF_X1 \h1/ff168 (.CK(hi_gclk2));
 DFF_X1 \h1/ff167 (.CK(hi_gclk2));
 DFF_X1 \h1/ff166 (.CK(hi_gclk2));
 DFF_X1 \h1/ff165 (.CK(hi_gclk2));
 DFF_X1 \h1/ff164 (.CK(hi_gclk2));
 DFF_X1 \h1/ff163 (.CK(hi_gclk2));
 DFF_X1 \h1/ff162 (.CK(hi_gclk2));
 DFF_X1 \h1/ff188 (.CK(hi_gclk2));
 DFF_X1 \h1/ff187 (.CK(hi_gclk2));
 DFF_X1 \h1/ff186 (.CK(hi_gclk2));
 DFF_X1 \h1/ff185 (.CK(hi_gclk2));
 DFF_X1 \h1/ff184 (.CK(hi_gclk2));
 DFF_X1 \h1/ff183 (.CK(hi_gclk2));
 DFF_X1 \h1/ff182 (.CK(hi_gclk2));
 DFF_X1 \h1/ff181 (.CK(hi_gclk2));
 DFF_X1 \h1/ff180 (.CK(hi_gclk2));
 DFF_X1 \h1/ff206 (.CK(hi_gclk2));
 DFF_X1 \h1/ff205 (.CK(hi_gclk2));
 DFF_X1 \h1/ff204 (.CK(hi_gclk2));
 DFF_X1 \h1/ff203 (.CK(hi_gclk2));
 DFF_X1 \h1/ff202 (.CK(hi_gclk2));
 DFF_X1 \h1/ff201 (.CK(hi_gclk2));
 DFF_X1 \h1/ff200 (.CK(hi_gclk2));
 DFF_X1 \h1/ff199 (.CK(hi_gclk2));
 DFF_X1 \h1/ff198 (.CK(hi_gclk2));
 CLKGATE_X1 hi_gclk5 (.CK(clk), .GCK(hi_gclk5));
 DFF_X1 \h1/ff143 (.CK(hi_gclk5));
 DFF_X1 \h1/ff142 (.CK(hi_gclk5));
 DFF_X1 \h1/ff141 (.CK(hi_gclk5));
 DFF_X1 \h1/ff140 (.CK(hi_gclk5));
 DFF_X1 \h1/ff139 (.CK(hi_gclk5));
 DFF_X1 \h1/ff138 (.CK(hi_gclk5));
 DFF_X1 \h1/ff137 (.CK(hi_gclk5));
 DFF_X1 \h1/ff136 (.CK(hi_gclk5));
 DFF_X1 \h1/ff135 (.CK(hi_gclk5));
 DFF_X1 \h1/ff134 (.CK(hi_gclk5));
 DFF_X1 \h1/ff133 (.CK(hi_gclk5));
 DFF_X1 \h1/ff132 (.CK(hi_gclk5));
 DFF_X1 \h1/ff131 (.CK(hi_gclk5));
 DFF_X1 \h1/ff130 (.CK(hi_gclk5));
 DFF_X1 \h1/ff129 (.CK(hi_gclk5));
 DFF_X1 \h1/ff125 (.CK(hi_gclk5));
 DFF_X1 \h1/ff124 (.CK(hi_gclk5));
 DFF_X1 \h1/ff123 (.CK(hi_gclk5));
 DFF_X1 \h1/ff122 (.CK(hi_gclk5));
 DFF_X1 \h1/ff121 (.CK(hi_gclk5));
 DFF_X1 \h1/ff120 (.CK(hi_gclk5));
 DFF_X1 \h1/ff119 (.CK(hi_gclk5));
 DFF_X1 \h1/ff118 (.CK(hi_gclk5));
 DFF_X1 \h1/ff117 (.CK(hi_gclk5));
 DFF_X1 \h1/ff116 (.CK(hi_gclk5));
 DFF_X1 \h1/ff115 (.CK(hi_gclk5));
 DFF_X1 \h1/ff114 (.CK(hi_gclk5));
 DFF_X1 \h1/ff113 (.CK(hi_gclk5));
 DFF_X1 \h1/ff112 (.CK(hi_gclk5));
 DFF_X1 \h1/ff111 (.CK(hi_gclk5));
 DFF_X1 \h1/ff107 (.CK(hi_gclk5));
 DFF_X1 \h1/ff106 (.CK(hi_gclk5));
 DFF_X1 \h1/ff105 (.CK(hi_gclk5));
 DFF_X1 \h1/ff104 (.CK(hi_gclk5));
 DFF_X1 \h1/ff103 (.CK(hi_gclk5));
 DFF_X1 \h1/ff102 (.CK(hi_gclk5));
 DFF_X1 \h1/ff101 (.CK(hi_gclk5));
 DFF_X1 \h1/ff100 (.CK(hi_gclk5));
 DFF_X1 \h1/ff99 (.CK(hi_gclk5));
 DFF_X1 \h1/ff98 (.CK(hi_gclk5));
 DFF_X1 \h1/ff97 (.CK(hi_gclk5));
 DFF_X1 \h1/ff96 (.CK(hi_gclk5));
 DFF_X1 \h1/ff95 (.CK(hi_gclk5));
 DFF_X1 \h1/ff94 (.CK(hi_gclk5));
 DFF_X1 \h1/ff93 (.CK(hi_gclk5));
 DFF_X1 \h1/ff92 (.CK(hi_gclk5));
 DFF_X1 \h1/ff89 (.CK(hi_gclk5));
 DFF_X1 \h1/ff88 (.CK(hi_gclk5));
 DFF_X1 \h1/ff87 (.CK(hi_gclk5));
 DFF_X1 \h1/ff86 (.CK(hi_gclk5));
 DFF_X1 \h1/ff85 (.CK(hi_gclk5));
 DFF_X1 \h1/ff84 (.CK(hi_gclk5));
 DFF_X1 \h1/ff83 (.CK(hi_gclk5));
 DFF_X1 \h1/ff82 (.CK(hi_gclk5));
 DFF_X1 \h1/ff81 (.CK(hi_gclk5));
 DFF_X1 \h1/ff80 (.CK(hi_gclk5));
 DFF_X1 \h1/ff79 (.CK(hi_gclk5));
 DFF_X1 \h1/ff78 (.CK(hi_gclk5));
 DFF_X1 \h1/ff77 (.CK(hi_gclk5));
 DFF_X1 \h1/ff76 (.CK(hi_gclk5));
 DFF_X1 \h1/ff75 (.CK(hi_gclk5));
 DFF_X1 \h1/ff74 (.CK(hi_gclk5));
 DFF_X1 \h1/ff71 (.CK(hi_gclk5));
 DFF_X1 \h1/ff70 (.CK(hi_gclk5));
 DFF_X1 \h1/ff69 (.CK(hi_gclk5));
 DFF_X1 \h1/ff68 (.CK(hi_gclk5));
 DFF_X1 \h1/ff67 (.CK(hi_gclk5));
 DFF_X1 \h1/ff66 (.CK(hi_gclk5));
 DFF_X1 \h1/ff65 (.CK(hi_gclk5));
 DFF_X1 \h1/ff64 (.CK(hi_gclk5));
 DFF_X1 \h1/ff63 (.CK(hi_gclk5));
 DFF_X1 \h1/ff62 (.CK(hi_gclk5));
 DFF_X1 \h1/ff61 (.CK(hi_gclk5));
 DFF_X1 \h1/ff60 (.CK(hi_gclk5));
 DFF_X1 \h1/ff59 (.CK(hi_gclk5));
 DFF_X1 \h1/ff58 (.CK(hi_gclk5));
 DFF_X1 \h1/ff57 (.CK(hi_gclk5));
 DFF_X1 \h1/ff56 (.CK(hi_gclk5));
 DFF_X1 \h1/ff55 (.CK(hi_gclk5));
 DFF_X1 \h1/ff54 (.CK(hi_gclk5));
 DFF_X1 \h1/ff53 (.CK(hi_gclk5));
 DFF_X1 \h1/ff52 (.CK(hi_gclk5));
 DFF_X1 \h1/ff51 (.CK(hi_gclk5));
 DFF_X1 \h1/ff50 (.CK(hi_gclk5));
 DFF_X1 \h1/ff49 (.CK(hi_gclk5));
 DFF_X1 \h1/ff48 (.CK(hi_gclk5));
 DFF_X1 \h1/ff47 (.CK(hi_gclk5));
 DFF_X1 \h1/ff46 (.CK(hi_gclk5));
 DFF_X1 \h1/ff45 (.CK(hi_gclk5));
 DFF_X1 \h1/ff44 (.CK(hi_gclk5));
 DFF_X1 \h1/ff43 (.CK(hi_gclk5));
 DFF_X1 \h1/ff42 (.CK(hi_gclk5));
 DFF_X1 \h1/ff41 (.CK(hi_gclk5));
 DFF_X1 \h1/ff40 (.CK(hi_gclk5));
 DFF_X1 \h1/ff39 (.CK(hi_gclk5));
 DFF_X1 \h1/ff38 (.CK(hi_gclk5));
 DFF_X1 \h1/ff37 (.CK(hi_gclk5));
 DFF_X1 \h1/ff36 (.CK(hi_gclk5));
 DFF_X1 \h1/ff35 (.CK(hi_gclk5));
 DFF_X1 \h1/ff34 (.CK(hi_gclk5));
 DFF_X1 \h1/ff33 (.CK(hi_gclk5));
 DFF_X1 \h1/ff32 (.CK(hi_gclk5));
 DFF_X1 \h1/ff31 (.CK(hi_gclk5));
 DFF_X1 \h1/ff30 (.CK(hi_gclk5));
 DFF_X1 \h1/ff29 (.CK(hi_gclk5));
 DFF_X1 \h1/ff28 (.CK(hi_gclk5));
 DFF_X1 \h1/ff27 (.CK(hi_gclk5));
 DFF_X1 \h1/ff26 (.CK(hi_gclk5));
 DFF_X1 \h1/ff25 (.CK(hi_gclk5));
 DFF_X1 \h1/ff24 (.CK(hi_gclk5));
 DFF_X1 \h1/ff23 (.CK(hi_gclk5));
 DFF_X1 \h1/ff22 (.CK(hi_gclk5));
 DFF_X1 \h1/ff21 (.CK(hi_gclk5));
 DFF_X1 \h1/ff20 (.CK(hi_gclk5));
 DFF_X1 \h1/ff19 (.CK(hi_gclk5));
 DFF_X1 \h1/ff18 (.CK(hi_gclk5));
 DFF_X1 \h1/ff17 (.CK(hi_gclk5));
 DFF_X1 \h1/ff16 (.CK(hi_gclk5));
 DFF_X1 \h1/ff15 (.CK(hi_gclk5));
 DFF_X1 \h1/ff14 (.CK(hi_gclk5));
 DFF_X1 \h1/ff13 (.CK(hi_gclk5));
 DFF_X1 \h1/ff12 (.CK(hi_gclk5));
 DFF_X1 \h1/ff11 (.CK(hi_gclk5));
 DFF_X1 \h1/ff10 (.CK(hi_gclk5));
 DFF_X1 \h1/ff9 (.CK(hi_gclk5));
 DFF_X1 \h1/ff8 (.CK(hi_gclk5));
 DFF_X1 \h1/ff7 (.CK(hi_gclk5));
 DFF_X1 \h1/ff6 (.CK(hi_gclk5));
 DFF_X1 \h1/ff5 (.CK(hi_gclk5));
 DFF_X1 \h1/ff4 (.CK(hi_gclk5));
 DFF_X1 \h1/ff3 (.CK(hi_gclk5));
 DFF_X1 \h1/ff2 (.CK(hi_gclk5));
 DFF_X1 \h1/ff1 (.CK(hi_gclk5));
 DFF_X1 \ff0/name (.CK(hi_gclk5));
 
endmodule // multi_sink
