VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MACRO snl_1nsdel
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_1nsdel

MACRO snl_2nsdel
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_2nsdel

MACRO snl_4nsdel
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_4nsdel

MACRO snl_add05x1
 SIZE 50 BY 20 ;
 PIN S DIRECTION OUTPUT ; END S
 PIN CO DIRECTION OUTPUT ; END CO
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_add05x1

MACRO snl_add05x2
 SIZE 50 BY 20 ;
 PIN S DIRECTION OUTPUT ; END S
 PIN CO DIRECTION OUTPUT ; END CO
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_add05x2

MACRO snl_add1x1
 SIZE 50 BY 20 ;
 PIN S DIRECTION OUTPUT ; END S
 PIN CO DIRECTION OUTPUT ; END CO
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN CI DIRECTION INPUT ; END CI
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_add1x1

MACRO snl_add1x2
 SIZE 50 BY 20 ;
 PIN S DIRECTION OUTPUT ; END S
 PIN CO DIRECTION OUTPUT ; END CO
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN CI DIRECTION INPUT ; END CI
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_add1x2

MACRO snl_addprop1x1
 SIZE 50 BY 20 ;
 PIN S DIRECTION OUTPUT ; END S
 PIN P DIRECTION OUTPUT ; END P
 PIN CO DIRECTION OUTPUT ; END CO
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN CI DIRECTION INPUT ; END CI
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_addprop1x1

MACRO snl_addprop1x2
 SIZE 50 BY 20 ;
 PIN S DIRECTION OUTPUT ; END S
 PIN P DIRECTION OUTPUT ; END P
 PIN CO DIRECTION OUTPUT ; END CO
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN CI DIRECTION INPUT ; END CI
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_addprop1x2

MACRO snl_and02x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and02x1

MACRO snl_and02x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and02x2

MACRO snl_and02x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and02x4

MACRO snl_and02x8
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and02x8

MACRO snl_and03x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and03x1

MACRO snl_and03x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and03x2

MACRO snl_and03x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and03x4

MACRO snl_and03x8
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and03x8

MACRO snl_and04x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and04x1

MACRO snl_and04x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and04x2

MACRO snl_and04x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and04x4

MACRO snl_and04x8
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and04x8

MACRO snl_and05x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and05x1

MACRO snl_and05x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and05x2

MACRO snl_and05x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and05x4

MACRO snl_and05x8
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and05x8

MACRO snl_and06x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and06x1

MACRO snl_and06x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and06x2

MACRO snl_and06x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and06x4

MACRO snl_and06x8
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and06x8

MACRO snl_and08x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and08x1

MACRO snl_and08x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and08x2

MACRO snl_and08x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and08x4

MACRO snl_and08x8
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and08x8

MACRO snl_and12x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and12x1

MACRO snl_and12x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and12x2

MACRO snl_and12x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and12x4

MACRO snl_and12x8
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and12x8

MACRO snl_and13x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and13x1

MACRO snl_and13x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and13x2

MACRO snl_and13x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and13x4

MACRO snl_and13x8
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and13x8

MACRO snl_and14x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and14x1

MACRO snl_and14x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and14x2

MACRO snl_and14x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and14x4

MACRO snl_and14x8
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and14x8

MACRO snl_and23x0
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and23x0

MACRO snl_and23x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and23x1

MACRO snl_and23x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and23x2

MACRO snl_and23x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and23x4

MACRO snl_and23x8
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and23x8

MACRO snl_and24x0
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and24x0

MACRO snl_and24x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and24x1

MACRO snl_and24x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and24x2

MACRO snl_and24x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and24x4

MACRO snl_and24x8
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and24x8

MACRO snl_and34x0
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and34x0

MACRO snl_and34x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and34x1

MACRO snl_and34x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and34x2

MACRO snl_and34x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and34x4

MACRO snl_and34x8
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and34x8

MACRO snl_ao012x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao012x1

MACRO snl_ao012x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao012x2

MACRO snl_ao012x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao012x4

MACRO snl_ao013x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao013x1

MACRO snl_ao013x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao013x2

MACRO snl_ao013x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao013x4

MACRO snl_ao01b2x0
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao01b2x0

MACRO snl_ao01b2x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao01b2x1

MACRO snl_ao01b2x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao01b2x2

MACRO snl_ao01b2x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao01b2x4

MACRO snl_ao01b3x0
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao01b3x0

MACRO snl_ao01b3x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao01b3x1

MACRO snl_ao01b3x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao01b3x2

MACRO snl_ao01b3x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao01b3x4

MACRO snl_ao022x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao022x1

MACRO snl_ao022x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao022x2

MACRO snl_ao022x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao022x4

MACRO snl_ao023x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao023x1

MACRO snl_ao023x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao023x2

MACRO snl_ao023x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao023x4

MACRO snl_ao02b2x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao02b2x1

MACRO snl_ao02b2x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao02b2x2

MACRO snl_ao02b2x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao02b2x4

MACRO snl_ao02b3x0
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao02b3x0

MACRO snl_ao02b3x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao02b3x1

MACRO snl_ao02b3x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao02b3x2

MACRO snl_ao02b3x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao02b3x4

MACRO snl_ao033x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao033x1

MACRO snl_ao033x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao033x2

MACRO snl_ao033x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao033x4

MACRO snl_ao03b3x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao03b3x1

MACRO snl_ao03b3x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao03b3x2

MACRO snl_ao03b3x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao03b3x4

MACRO snl_ao0b12x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao0b12x1

MACRO snl_ao0b12x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao0b12x2

MACRO snl_ao0b12x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao0b12x4

MACRO snl_ao0b13x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao0b13x1

MACRO snl_ao0b13x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao0b13x2

MACRO snl_ao0b13x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao0b13x4

MACRO snl_ao0b23x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao0b23x1

MACRO snl_ao0b23x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao0b23x2

MACRO snl_ao0b23x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao0b23x4

MACRO snl_ao112x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao112x1

MACRO snl_ao112x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao112x2

MACRO snl_ao112x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao112x4

MACRO snl_ao113x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao113x1

MACRO snl_ao113x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao113x2

MACRO snl_ao113x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao113x4

MACRO snl_ao11b2x0
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao11b2x0

MACRO snl_ao11b2x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao11b2x1

MACRO snl_ao11b2x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao11b2x2

MACRO snl_ao11b2x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao11b2x4

MACRO snl_ao11b3x0
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao11b3x0

MACRO snl_ao11b3x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao11b3x1

MACRO snl_ao11b3x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao11b3x2

MACRO snl_ao11b3x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao11b3x4

MACRO snl_ao122x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao122x1

MACRO snl_ao122x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao122x2

MACRO snl_ao122x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao122x4

MACRO snl_ao123x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao123x1

MACRO snl_ao123x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao123x2

MACRO snl_ao123x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao123x4

MACRO snl_ao12b2x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao12b2x1

MACRO snl_ao12b2x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao12b2x2

MACRO snl_ao12b2x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao12b2x4

MACRO snl_ao12b3x0
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao12b3x0

MACRO snl_ao12b3x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao12b3x1

MACRO snl_ao12b3x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao12b3x2

MACRO snl_ao12b3x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao12b3x4

MACRO snl_ao133x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao133x1

MACRO snl_ao133x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao133x2

MACRO snl_ao133x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao133x4

MACRO snl_ao13b3x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao13b3x1

MACRO snl_ao13b3x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao13b3x2

MACRO snl_ao13b3x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao13b3x4

MACRO snl_ao1b12x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao1b12x1

MACRO snl_ao1b12x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao1b12x2

MACRO snl_ao1b12x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao1b12x4

MACRO snl_ao1b13x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao1b13x1

MACRO snl_ao1b13x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao1b13x2

MACRO snl_ao1b13x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao1b13x4

MACRO snl_ao1b1b2x0
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao1b1b2x0

MACRO snl_ao1b1b2x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao1b1b2x1

MACRO snl_ao1b1b2x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao1b1b2x2

MACRO snl_ao1b1b2x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao1b1b2x4

MACRO snl_ao1b1b3x0
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao1b1b3x0

MACRO snl_ao1b1b3x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao1b1b3x1

MACRO snl_ao1b1b3x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao1b1b3x2

MACRO snl_ao1b1b3x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao1b1b3x4

MACRO snl_ao1b23x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao1b23x1

MACRO snl_ao1b23x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao1b23x2

MACRO snl_ao1b23x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao1b23x4

MACRO snl_ao1b2b2x0
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao1b2b2x0

MACRO snl_ao1b2b2x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao1b2b2x1

MACRO snl_ao1b2b2x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao1b2b2x2

MACRO snl_ao1b2b2x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao1b2b2x4

MACRO snl_ao1b2b3x0
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao1b2b3x0

MACRO snl_ao1b2b3x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao1b2b3x1

MACRO snl_ao1b2b3x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao1b2b3x2

MACRO snl_ao1b2b3x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao1b2b3x4

MACRO snl_ao1b3b3x0
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao1b3b3x0

MACRO snl_ao1b3b3x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao1b3b3x1

MACRO snl_ao1b3b3x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao1b3b3x2

MACRO snl_ao1b3b3x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao1b3b3x4

MACRO snl_ao2222x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao2222x1

MACRO snl_ao2222x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao2222x2

MACRO snl_ao2222x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao2222x4

MACRO snl_ao222x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao222x1

MACRO snl_ao222x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao222x2

MACRO snl_ao222x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao222x4

MACRO snl_ao223x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao223x1

MACRO snl_ao223x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao223x2

MACRO snl_ao223x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao223x4

MACRO snl_ao22b2x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao22b2x1

MACRO snl_ao22b2x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao22b2x2

MACRO snl_ao22b2x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao22b2x4

MACRO snl_ao22b3x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao22b3x1

MACRO snl_ao22b3x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao22b3x2

MACRO snl_ao22b3x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao22b3x4

MACRO snl_ao233x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao233x1

MACRO snl_ao233x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao233x2

MACRO snl_ao233x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao233x4

MACRO snl_ao23b3x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao23b3x1

MACRO snl_ao23b3x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao23b3x2

MACRO snl_ao23b3x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao23b3x4

MACRO snl_ao2b23x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao2b23x1

MACRO snl_ao2b23x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao2b23x2

MACRO snl_ao2b23x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao2b23x4

MACRO snl_ao2b2b2x0
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao2b2b2x0

MACRO snl_ao2b2b2x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao2b2b2x1

MACRO snl_ao2b2b2x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao2b2b2x2

MACRO snl_ao2b2b2x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao2b2b2x4

MACRO snl_ao2b2b3x0
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao2b2b3x0

MACRO snl_ao2b2b3x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao2b2b3x1

MACRO snl_ao2b2b3x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao2b2b3x2

MACRO snl_ao2b2b3x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao2b2b3x4

MACRO snl_ao2b3b3x0
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao2b3b3x0

MACRO snl_ao2b3b3x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao2b3b3x1

MACRO snl_ao2b3b3x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao2b3b3x2

MACRO snl_ao2b3b3x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao2b3b3x4

MACRO snl_ao333x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN I DIRECTION INPUT ; END I
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao333x1

MACRO snl_ao333x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN I DIRECTION INPUT ; END I
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao333x2

MACRO snl_ao333x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN I DIRECTION INPUT ; END I
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao333x4

MACRO snl_ao33b3x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN I DIRECTION INPUT ; END I
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao33b3x1

MACRO snl_ao33b3x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN I DIRECTION INPUT ; END I
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao33b3x2

MACRO snl_ao33b3x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN I DIRECTION INPUT ; END I
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao33b3x4

MACRO snl_ao3b3b3x0
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN I DIRECTION INPUT ; END I
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao3b3b3x0

MACRO snl_ao3b3b3x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN I DIRECTION INPUT ; END I
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao3b3b3x1

MACRO snl_ao3b3b3x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN I DIRECTION INPUT ; END I
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao3b3b3x2

MACRO snl_ao3b3b3x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN I DIRECTION INPUT ; END I
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ao3b3b3x4

MACRO snl_aob122x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob122x1

MACRO snl_aob122x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob122x2

MACRO snl_aob122x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob122x4

MACRO snl_aob123x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob123x1

MACRO snl_aob123x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob123x2

MACRO snl_aob123x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob123x4

MACRO snl_aob12b2x0
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob12b2x0

MACRO snl_aob12b2x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob12b2x1

MACRO snl_aob12b2x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob12b2x2

MACRO snl_aob12b2x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob12b2x4

MACRO snl_aob12b3x0
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob12b3x0

MACRO snl_aob12b3x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob12b3x1

MACRO snl_aob12b3x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob12b3x2

MACRO snl_aob12b3x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob12b3x4

MACRO snl_aob133x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob133x1

MACRO snl_aob133x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob133x2

MACRO snl_aob133x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob133x4

MACRO snl_aob13b3x0
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob13b3x0

MACRO snl_aob13b3x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob13b3x1

MACRO snl_aob13b3x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob13b3x2

MACRO snl_aob13b3x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob13b3x4

MACRO snl_aob1b12x0
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob1b12x0

MACRO snl_aob1b12x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob1b12x1

MACRO snl_aob1b12x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob1b12x2

MACRO snl_aob1b12x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob1b12x4

MACRO snl_aob1b13x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob1b13x1

MACRO snl_aob1b13x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob1b13x2

MACRO snl_aob1b13x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob1b13x4

MACRO snl_aob1b23x0
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob1b23x0

MACRO snl_aob1b23x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob1b23x1

MACRO snl_aob1b23x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob1b23x2

MACRO snl_aob1b23x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob1b23x4

MACRO snl_aob233x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob233x1

MACRO snl_aob233x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob233x2

MACRO snl_aob233x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob233x4

MACRO snl_aob23b3x0
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob23b3x0

MACRO snl_aob23b3x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob23b3x1

MACRO snl_aob23b3x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob23b3x2

MACRO snl_aob23b3x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob23b3x4

MACRO snl_aob2b23x0
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob2b23x0

MACRO snl_aob2b23x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob2b23x1

MACRO snl_aob2b23x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob2b23x2

MACRO snl_aob2b23x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aob2b23x4

MACRO snl_aoi012x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi012x1

MACRO snl_aoi012x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi012x2

MACRO snl_aoi012x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi012x4

MACRO snl_aoi013x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi013x0

MACRO snl_aoi013x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi013x1

MACRO snl_aoi013x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi013x2

MACRO snl_aoi013x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi013x4

MACRO snl_aoi01b2x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi01b2x1

MACRO snl_aoi01b2x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi01b2x2

MACRO snl_aoi01b2x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi01b2x4

MACRO snl_aoi01b3x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi01b3x1

MACRO snl_aoi01b3x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi01b3x2

MACRO snl_aoi01b3x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi01b3x4

MACRO snl_aoi022x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi022x1

MACRO snl_aoi022x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi022x2

MACRO snl_aoi022x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi022x4

MACRO snl_aoi023x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi023x0

MACRO snl_aoi023x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi023x1

MACRO snl_aoi023x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi023x2

MACRO snl_aoi023x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi023x4

MACRO snl_aoi02b2x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi02b2x0

MACRO snl_aoi02b2x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi02b2x1

MACRO snl_aoi02b2x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi02b2x2

MACRO snl_aoi02b2x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi02b2x4

MACRO snl_aoi02b3x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi02b3x1

MACRO snl_aoi02b3x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi02b3x2

MACRO snl_aoi02b3x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi02b3x4

MACRO snl_aoi033x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi033x0

MACRO snl_aoi033x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi033x1

MACRO snl_aoi033x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi033x2

MACRO snl_aoi033x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi033x4

MACRO snl_aoi03b3x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi03b3x0

MACRO snl_aoi03b3x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi03b3x1

MACRO snl_aoi03b3x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi03b3x2

MACRO snl_aoi03b3x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi03b3x4

MACRO snl_aoi0b12x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi0b12x0

MACRO snl_aoi0b12x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi0b12x1

MACRO snl_aoi0b12x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi0b12x2

MACRO snl_aoi0b12x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi0b12x4

MACRO snl_aoi0b13x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi0b13x0

MACRO snl_aoi0b13x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi0b13x1

MACRO snl_aoi0b13x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi0b13x2

MACRO snl_aoi0b13x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi0b13x4

MACRO snl_aoi0b23x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi0b23x0

MACRO snl_aoi0b23x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi0b23x1

MACRO snl_aoi0b23x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi0b23x2

MACRO snl_aoi0b23x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi0b23x4

MACRO snl_aoi112x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi112x0

MACRO snl_aoi112x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi112x1

MACRO snl_aoi112x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi112x2

MACRO snl_aoi112x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi112x4

MACRO snl_aoi113x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi113x0

MACRO snl_aoi113x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi113x1

MACRO snl_aoi113x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi113x2

MACRO snl_aoi113x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi113x4

MACRO snl_aoi11b2x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi11b2x0

MACRO snl_aoi11b2x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi11b2x1

MACRO snl_aoi11b2x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi11b2x2

MACRO snl_aoi11b2x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi11b2x4

MACRO snl_aoi11b3x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi11b3x1

MACRO snl_aoi11b3x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi11b3x2

MACRO snl_aoi11b3x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi11b3x4

MACRO snl_aoi122x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi122x0

MACRO snl_aoi122x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi122x1

MACRO snl_aoi122x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi122x2

MACRO snl_aoi122x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi122x4

MACRO snl_aoi123x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi123x0

MACRO snl_aoi123x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi123x1

MACRO snl_aoi123x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi123x2

MACRO snl_aoi123x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi123x4

MACRO snl_aoi12b2x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi12b2x0

MACRO snl_aoi12b2x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi12b2x1

MACRO snl_aoi12b2x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi12b2x2

MACRO snl_aoi12b2x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi12b2x4

MACRO snl_aoi12b3x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi12b3x0

MACRO snl_aoi12b3x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi12b3x1

MACRO snl_aoi12b3x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi12b3x2

MACRO snl_aoi12b3x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi12b3x4

MACRO snl_aoi133x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi133x0

MACRO snl_aoi133x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi133x1

MACRO snl_aoi133x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi133x2

MACRO snl_aoi133x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi133x4

MACRO snl_aoi13b3x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi13b3x0

MACRO snl_aoi13b3x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi13b3x1

MACRO snl_aoi13b3x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi13b3x2

MACRO snl_aoi13b3x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi13b3x4

MACRO snl_aoi1b12x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi1b12x0

MACRO snl_aoi1b12x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi1b12x1

MACRO snl_aoi1b12x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi1b12x2

MACRO snl_aoi1b12x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi1b12x4

MACRO snl_aoi1b13x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi1b13x0

MACRO snl_aoi1b13x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi1b13x1

MACRO snl_aoi1b13x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi1b13x2

MACRO snl_aoi1b13x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi1b13x4

MACRO snl_aoi1b1b2x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi1b1b2x1

MACRO snl_aoi1b1b2x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi1b1b2x2

MACRO snl_aoi1b1b2x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi1b1b2x4

MACRO snl_aoi1b1b3x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi1b1b3x1

MACRO snl_aoi1b1b3x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi1b1b3x2

MACRO snl_aoi1b1b3x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi1b1b3x4

MACRO snl_aoi1b23x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi1b23x0

MACRO snl_aoi1b23x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi1b23x1

MACRO snl_aoi1b23x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi1b23x2

MACRO snl_aoi1b23x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi1b23x4

MACRO snl_aoi1b2b2x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi1b2b2x1

MACRO snl_aoi1b2b2x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi1b2b2x2

MACRO snl_aoi1b2b2x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi1b2b2x4

MACRO snl_aoi1b2b3x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi1b2b3x1

MACRO snl_aoi1b2b3x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi1b2b3x2

MACRO snl_aoi1b2b3x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi1b2b3x4

MACRO snl_aoi1b3b3x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi1b3b3x1

MACRO snl_aoi1b3b3x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi1b3b3x2

MACRO snl_aoi1b3b3x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi1b3b3x4

MACRO snl_aoi2222x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi2222x0

MACRO snl_aoi2222x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi2222x1

MACRO snl_aoi2222x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi2222x2

MACRO snl_aoi2222x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi2222x4

MACRO snl_aoi222x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi222x0

MACRO snl_aoi222x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi222x1

MACRO snl_aoi222x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi222x2

MACRO snl_aoi222x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi222x4

MACRO snl_aoi223x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi223x0

MACRO snl_aoi223x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi223x1

MACRO snl_aoi223x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi223x2

MACRO snl_aoi223x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi223x4

MACRO snl_aoi22b2x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi22b2x0

MACRO snl_aoi22b2x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi22b2x1

MACRO snl_aoi22b2x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi22b2x2

MACRO snl_aoi22b2x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi22b2x4

MACRO snl_aoi22b3x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi22b3x0

MACRO snl_aoi22b3x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi22b3x1

MACRO snl_aoi22b3x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi22b3x2

MACRO snl_aoi22b3x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi22b3x4

MACRO snl_aoi233x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi233x0

MACRO snl_aoi233x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi233x1

MACRO snl_aoi233x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi233x2

MACRO snl_aoi233x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi233x4

MACRO snl_aoi23b3x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi23b3x0

MACRO snl_aoi23b3x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi23b3x1

MACRO snl_aoi23b3x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi23b3x2

MACRO snl_aoi23b3x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi23b3x4

MACRO snl_aoi2b23x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi2b23x0

MACRO snl_aoi2b23x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi2b23x1

MACRO snl_aoi2b23x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi2b23x2

MACRO snl_aoi2b23x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi2b23x4

MACRO snl_aoi2b2b2x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi2b2b2x1

MACRO snl_aoi2b2b2x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi2b2b2x2

MACRO snl_aoi2b2b2x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi2b2b2x4

MACRO snl_aoi2b2b3x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi2b2b3x1

MACRO snl_aoi2b2b3x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi2b2b3x2

MACRO snl_aoi2b2b3x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi2b2b3x4

MACRO snl_aoi2b3b3x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi2b3b3x1

MACRO snl_aoi2b3b3x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi2b3b3x2

MACRO snl_aoi2b3b3x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi2b3b3x4

MACRO snl_aoi333x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN I DIRECTION INPUT ; END I
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi333x0

MACRO snl_aoi333x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN I DIRECTION INPUT ; END I
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi333x1

MACRO snl_aoi333x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN I DIRECTION INPUT ; END I
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi333x2

MACRO snl_aoi333x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN I DIRECTION INPUT ; END I
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi333x4

MACRO snl_aoi33b3x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN I DIRECTION INPUT ; END I
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi33b3x0

MACRO snl_aoi33b3x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN I DIRECTION INPUT ; END I
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi33b3x1

MACRO snl_aoi33b3x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN I DIRECTION INPUT ; END I
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi33b3x2

MACRO snl_aoi33b3x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN I DIRECTION INPUT ; END I
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi33b3x4

MACRO snl_aoi3b3b3x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN I DIRECTION INPUT ; END I
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi3b3b3x1

MACRO snl_aoi3b3b3x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN I DIRECTION INPUT ; END I
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi3b3b3x2

MACRO snl_aoi3b3b3x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN I DIRECTION INPUT ; END I
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoi3b3b3x4

MACRO snl_aoib122x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib122x0

MACRO snl_aoib122x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib122x1

MACRO snl_aoib122x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib122x2

MACRO snl_aoib122x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib122x4

MACRO snl_aoib123x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib123x0

MACRO snl_aoib123x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib123x1

MACRO snl_aoib123x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib123x2

MACRO snl_aoib123x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib123x4

MACRO snl_aoib12b2x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib12b2x1

MACRO snl_aoib12b2x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib12b2x2

MACRO snl_aoib12b2x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib12b2x4

MACRO snl_aoib12b3x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib12b3x1

MACRO snl_aoib12b3x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib12b3x2

MACRO snl_aoib12b3x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib12b3x4

MACRO snl_aoib133x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib133x0

MACRO snl_aoib133x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib133x1

MACRO snl_aoib133x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib133x2

MACRO snl_aoib133x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib133x4

MACRO snl_aoib13b3x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib13b3x1

MACRO snl_aoib13b3x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib13b3x2

MACRO snl_aoib13b3x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib13b3x4

MACRO snl_aoib1b12x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib1b12x0

MACRO snl_aoib1b12x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib1b12x1

MACRO snl_aoib1b12x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib1b12x2

MACRO snl_aoib1b12x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib1b12x4

MACRO snl_aoib1b13x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib1b13x0

MACRO snl_aoib1b13x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib1b13x1

MACRO snl_aoib1b13x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib1b13x2

MACRO snl_aoib1b13x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib1b13x4

MACRO snl_aoib1b23x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib1b23x0

MACRO snl_aoib1b23x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib1b23x1

MACRO snl_aoib1b23x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib1b23x2

MACRO snl_aoib1b23x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib1b23x4

MACRO snl_aoib233x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib233x0

MACRO snl_aoib233x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib233x1

MACRO snl_aoib233x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib233x2

MACRO snl_aoib233x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib233x4

MACRO snl_aoib23b3x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib23b3x1

MACRO snl_aoib23b3x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib23b3x2

MACRO snl_aoib23b3x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib23b3x4

MACRO snl_aoib2b23x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib2b23x1

MACRO snl_aoib2b23x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib2b23x2

MACRO snl_aoib2b23x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_aoib2b23x4

MACRO snl_bufx1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_bufx1

MACRO snl_bufx12
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_bufx12

MACRO snl_bufx16
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_bufx16

MACRO snl_bufx2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_bufx2

MACRO snl_bufx20
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_bufx20

MACRO snl_bufx24
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_bufx24

MACRO snl_bufx4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_bufx4

MACRO snl_bufx8
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_bufx8

MACRO snl_clkbufx1
 SIZE 50 BY 20 ;
 PIN CP DIRECTION OUTPUT ; END CP
 PIN CN DIRECTION OUTPUT ; END CN
 PIN CLK DIRECTION INPUT ; END CLK
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_clkbufx1

MACRO snl_clkbufx12
 SIZE 50 BY 20 ;
 PIN CP DIRECTION OUTPUT ; END CP
 PIN CN DIRECTION OUTPUT ; END CN
 PIN CLK DIRECTION INPUT ; END CLK
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_clkbufx12

MACRO snl_clkbufx16
 SIZE 50 BY 20 ;
 PIN CP DIRECTION OUTPUT ; END CP
 PIN CN DIRECTION OUTPUT ; END CN
 PIN CLK DIRECTION INPUT ; END CLK
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_clkbufx16

MACRO snl_clkbufx2
 SIZE 50 BY 20 ;
 PIN CP DIRECTION OUTPUT ; END CP
 PIN CN DIRECTION OUTPUT ; END CN
 PIN CLK DIRECTION INPUT ; END CLK
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_clkbufx2

MACRO snl_clkbufx20
 SIZE 50 BY 20 ;
 PIN CP DIRECTION OUTPUT ; END CP
 PIN CN DIRECTION OUTPUT ; END CN
 PIN CLK DIRECTION INPUT ; END CLK
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_clkbufx20

MACRO snl_clkbufx24
 SIZE 50 BY 20 ;
 PIN CP DIRECTION OUTPUT ; END CP
 PIN CN DIRECTION OUTPUT ; END CN
 PIN CLK DIRECTION INPUT ; END CLK
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_clkbufx24

MACRO snl_clkbufx4
 SIZE 50 BY 20 ;
 PIN CP DIRECTION OUTPUT ; END CP
 PIN CN DIRECTION OUTPUT ; END CN
 PIN CLK DIRECTION INPUT ; END CLK
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_clkbufx4

MACRO snl_clkbufx8
 SIZE 50 BY 20 ;
 PIN CP DIRECTION OUTPUT ; END CP
 PIN CN DIRECTION OUTPUT ; END CN
 PIN CLK DIRECTION INPUT ; END CLK
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_clkbufx8

MACRO snl_dec24x1
 SIZE 50 BY 20 ;
 PIN Z1 DIRECTION OUTPUT ; END Z1
 PIN Z2 DIRECTION OUTPUT ; END Z2
 PIN Z3 DIRECTION OUTPUT ; END Z3
 PIN Z4 DIRECTION OUTPUT ; END Z4
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_dec24x1

MACRO snl_dec24x2
 SIZE 50 BY 20 ;
 PIN Z1 DIRECTION OUTPUT ; END Z1
 PIN Z2 DIRECTION OUTPUT ; END Z2
 PIN Z3 DIRECTION OUTPUT ; END Z3
 PIN Z4 DIRECTION OUTPUT ; END Z4
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_dec24x2

MACRO snl_deci24x1
 SIZE 50 BY 20 ;
 PIN ZN1 DIRECTION OUTPUT ; END ZN1
 PIN ZN2 DIRECTION OUTPUT ; END ZN2
 PIN ZN3 DIRECTION OUTPUT ; END ZN3
 PIN ZN4 DIRECTION OUTPUT ; END ZN4
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_deci24x1

MACRO snl_deci24x2
 SIZE 50 BY 20 ;
 PIN ZN1 DIRECTION OUTPUT ; END ZN1
 PIN ZN2 DIRECTION OUTPUT ; END ZN2
 PIN ZN3 DIRECTION OUTPUT ; END ZN3
 PIN ZN4 DIRECTION OUTPUT ; END ZN4
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_deci24x2

MACRO snl_ffandnorx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffandnorx1

MACRO snl_ffandnorx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffandnorx2

MACRO snl_ffandnorx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffandnorx4

MACRO snl_ffandorx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffandorx1

MACRO snl_ffandorx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffandorx2

MACRO snl_ffandorx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffandorx4

MACRO snl_ffandx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffandx1

MACRO snl_ffandx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffandx2

MACRO snl_ffandx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffandx4

MACRO snl_ffmu2x1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN S DIRECTION INPUT ; END S
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffmu2x1

MACRO snl_ffmu2x2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN S DIRECTION INPUT ; END S
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffmu2x2

MACRO snl_ffmu2x4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN S DIRECTION INPUT ; END S
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffmu2x4

MACRO snl_ffnandx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffnandx1

MACRO snl_ffnandx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffnandx2

MACRO snl_ffnandx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffnandx4

MACRO snl_ffnorx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffnorx1

MACRO snl_ffnorx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffnorx2

MACRO snl_ffnorx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffnorx4

MACRO snl_fforandx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_fforandx1

MACRO snl_fforandx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_fforandx2

MACRO snl_fforandx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_fforandx4

MACRO snl_ffornandx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffornandx1

MACRO snl_ffornandx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffornandx2

MACRO snl_ffornandx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffornandx4

MACRO snl_fforx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_fforx1

MACRO snl_fforx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_fforx2

MACRO snl_fforx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_fforx4

MACRO snl_ffqenrnx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN RN DIRECTION INPUT ; END RN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqenrnx1

MACRO snl_ffqenrnx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN RN DIRECTION INPUT ; END RN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqenrnx2

MACRO snl_ffqenrnx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN RN DIRECTION INPUT ; END RN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqenrnx4

MACRO snl_ffqensnx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN SN DIRECTION INPUT ; END SN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqensnx1

MACRO snl_ffqensnx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN SN DIRECTION INPUT ; END SN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqensnx2

MACRO snl_ffqensnx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN SN DIRECTION INPUT ; END SN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqensnx4

MACRO snl_ffqenx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqenx1

MACRO snl_ffqenx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqenx2

MACRO snl_ffqenx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqenx4

MACRO snl_ffqnenrnx1
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN RN DIRECTION INPUT ; END RN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqnenrnx1

MACRO snl_ffqnenrnx2
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN RN DIRECTION INPUT ; END RN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqnenrnx2

MACRO snl_ffqnenrnx4
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN RN DIRECTION INPUT ; END RN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqnenrnx4

MACRO snl_ffqnensnx1
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN SN DIRECTION INPUT ; END SN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqnensnx1

MACRO snl_ffqnensnx2
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN SN DIRECTION INPUT ; END SN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqnensnx2

MACRO snl_ffqnensnx4
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN SN DIRECTION INPUT ; END SN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqnensnx4

MACRO snl_ffqnenx1
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqnenx1

MACRO snl_ffqnenx2
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqnenx2

MACRO snl_ffqnenx4
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqnenx4

MACRO snl_ffqnrnx1
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqnrnx1

MACRO snl_ffqnrnx2
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqnrnx2

MACRO snl_ffqnrnx4
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqnrnx4

MACRO snl_ffqnsnx1
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN SN DIRECTION INPUT ; END SN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqnsnx1

MACRO snl_ffqnsnx2
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN SN DIRECTION INPUT ; END SN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqnsnx2

MACRO snl_ffqnsnx4
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN SN DIRECTION INPUT ; END SN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqnsnx4

MACRO snl_ffqnx1
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqnx1

MACRO snl_ffqnx2
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqnx2

MACRO snl_ffqnx4
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqnx4

MACRO snl_ffqqnenrnx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN RN DIRECTION INPUT ; END RN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqqnenrnx1

MACRO snl_ffqqnenrnx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN RN DIRECTION INPUT ; END RN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqqnenrnx2

MACRO snl_ffqqnensnx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN SN DIRECTION INPUT ; END SN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqqnensnx1

MACRO snl_ffqqnensnx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN SN DIRECTION INPUT ; END SN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqqnensnx2

MACRO snl_ffqqnenx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqqnenx1

MACRO snl_ffqqnenx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqqnenx2

MACRO snl_ffqqnrnsnx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqqnrnsnx1

MACRO snl_ffqqnrnsnx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqqnrnsnx2

MACRO snl_ffqqnrnx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqqnrnx1

MACRO snl_ffqqnrnx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqqnrnx2

MACRO snl_ffqqnsnx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN SN DIRECTION INPUT ; END SN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqqnsnx1

MACRO snl_ffqqnsnx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN SN DIRECTION INPUT ; END SN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqqnsnx2

MACRO snl_ffqqnx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqqnx1

MACRO snl_ffqqnx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqqnx2

MACRO snl_ffqrnx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqrnx1

MACRO snl_ffqrnx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqrnx2

MACRO snl_ffqrnx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqrnx4

MACRO snl_ffqsnx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN SN DIRECTION INPUT ; END SN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqsnx1

MACRO snl_ffqsnx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN SN DIRECTION INPUT ; END SN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqsnx2

MACRO snl_ffqsnx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN SN DIRECTION INPUT ; END SN
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqsnx4

MACRO snl_ffqx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqx1

MACRO snl_ffqx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqx2

MACRO snl_ffqx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqx4

MACRO snl_invx05
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_invx05

MACRO snl_invx1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_invx1

MACRO snl_invx12
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_invx12

MACRO snl_invx16
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_invx16

MACRO snl_invx2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_invx2

MACRO snl_invx20
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_invx20

MACRO snl_invx24
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_invx24

MACRO snl_invx3
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_invx3

MACRO snl_invx4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_invx4

MACRO snl_invx5
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_invx5

MACRO snl_invx6
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_invx6

MACRO snl_invx7
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_invx7

MACRO snl_invx8
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_invx8

MACRO snl_landnorx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_landnorx1

MACRO snl_landnorx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_landnorx2

MACRO snl_landnorx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_landnorx4

MACRO snl_landorx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_landorx1

MACRO snl_landorx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_landorx2

MACRO snl_landorx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_landorx4

MACRO snl_landx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_landx1

MACRO snl_landx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_landx2

MACRO snl_landx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_landx4

MACRO snl_lenqnrnsnx1
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqnrnsnx1

MACRO snl_lenqnrnsnx2
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqnrnsnx2

MACRO snl_lenqnrnsnx4
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqnrnsnx4

MACRO snl_lenqnrnx1
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqnrnx1

MACRO snl_lenqnrnx2
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqnrnx2

MACRO snl_lenqnrnx4
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqnrnx4

MACRO snl_lenqnsnrnx1
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqnsnrnx1

MACRO snl_lenqnsnrnx2
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqnsnrnx2

MACRO snl_lenqnsnrnx4
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqnsnrnx4

MACRO snl_lenqnsnx1
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN SN DIRECTION INPUT ; END SN
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqnsnx1

MACRO snl_lenqnsnx2
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN SN DIRECTION INPUT ; END SN
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqnsnx2

MACRO snl_lenqnsnx4
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN SN DIRECTION INPUT ; END SN
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqnsnx4

MACRO snl_lenqnx1
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqnx1

MACRO snl_lenqnx2
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqnx2

MACRO snl_lenqnx4
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqnx4

MACRO snl_lenqqnrnsnx1
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqqnrnsnx1

MACRO snl_lenqqnrnsnx2
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqqnrnsnx2

MACRO snl_lenqqnrnx1
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqqnrnx1

MACRO snl_lenqqnrnx2
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqqnrnx2

MACRO snl_lenqqnsnrnx1
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqqnsnrnx1

MACRO snl_lenqqnsnrnx2
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqqnsnrnx2

MACRO snl_lenqqnsnx1
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN SN DIRECTION INPUT ; END SN
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqqnsnx1

MACRO snl_lenqqnsnx2
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN SN DIRECTION INPUT ; END SN
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqqnsnx2

MACRO snl_lenqqnx1
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqqnx1

MACRO snl_lenqqnx2
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqqnx2

MACRO snl_lenqrnsnx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqrnsnx1

MACRO snl_lenqrnsnx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqrnsnx2

MACRO snl_lenqrnsnx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqrnsnx4

MACRO snl_lenqrnx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqrnx1

MACRO snl_lenqrnx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqrnx2

MACRO snl_lenqrnx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqrnx4

MACRO snl_lenqsnrnx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqsnrnx1

MACRO snl_lenqsnrnx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqsnrnx2

MACRO snl_lenqsnrnx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqsnrnx4

MACRO snl_lenqsnx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN SN DIRECTION INPUT ; END SN
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqsnx1

MACRO snl_lenqsnx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN SN DIRECTION INPUT ; END SN
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqsnx2

MACRO snl_lenqsnx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN SN DIRECTION INPUT ; END SN
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqsnx4

MACRO snl_lenqx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqx1

MACRO snl_lenqx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqx2

MACRO snl_lenqx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lenqx4

MACRO snl_lmu2x1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN S DIRECTION INPUT ; END S
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lmu2x1

MACRO snl_lmu2x2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN S DIRECTION INPUT ; END S
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lmu2x2

MACRO snl_lmu2x4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN S DIRECTION INPUT ; END S
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lmu2x4

MACRO snl_lnandx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lnandx1

MACRO snl_lnandx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lnandx2

MACRO snl_lnandx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lnandx4

MACRO snl_lnorx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lnorx1

MACRO snl_lnorx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lnorx2

MACRO snl_lnorx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lnorx4

MACRO snl_lorandx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lorandx1

MACRO snl_lorandx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lorandx2

MACRO snl_lorandx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lorandx4

MACRO snl_lornandx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lornandx1

MACRO snl_lornandx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lornandx2

MACRO snl_lornandx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lornandx4

MACRO snl_lorx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lorx1

MACRO snl_lorx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lorx2

MACRO snl_lorx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lorx4

MACRO snl_lqnrnsnx1
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqnrnsnx1

MACRO snl_lqnrnsnx2
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqnrnsnx2

MACRO snl_lqnrnsnx4
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqnrnsnx4

MACRO snl_lqnrnx1
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqnrnx1

MACRO snl_lqnrnx2
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqnrnx2

MACRO snl_lqnrnx4
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqnrnx4

MACRO snl_lqnsnrnx1
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqnsnrnx1

MACRO snl_lqnsnrnx2
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqnsnrnx2

MACRO snl_lqnsnrnx4
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqnsnrnx4

MACRO snl_lqnsnx1
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN SN DIRECTION INPUT ; END SN
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqnsnx1

MACRO snl_lqnsnx2
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN SN DIRECTION INPUT ; END SN
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqnsnx2

MACRO snl_lqnsnx4
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN SN DIRECTION INPUT ; END SN
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqnsnx4

MACRO snl_lqnx1
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqnx1

MACRO snl_lqnx2
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqnx2

MACRO snl_lqnx4
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqnx4

MACRO snl_lqqnrnsnx1
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqqnrnsnx1

MACRO snl_lqqnrnsnx2
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqqnrnsnx2

MACRO snl_lqqnrnx1
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqqnrnx1

MACRO snl_lqqnrnx2
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqqnrnx2

MACRO snl_lqqnsnrnx1
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqqnsnrnx1

MACRO snl_lqqnsnrnx2
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqqnsnrnx2

MACRO snl_lqqnsnx1
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN SN DIRECTION INPUT ; END SN
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqqnsnx1

MACRO snl_lqqnsnx2
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN SN DIRECTION INPUT ; END SN
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqqnsnx2

MACRO snl_lqqnx1
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqqnx1

MACRO snl_lqqnx2
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqqnx2

MACRO snl_lqrnsnx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqrnsnx1

MACRO snl_lqrnsnx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqrnsnx2

MACRO snl_lqrnsnx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqrnsnx4

MACRO snl_lqrnx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqrnx1

MACRO snl_lqrnx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqrnx2

MACRO snl_lqrnx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqrnx4

MACRO snl_lqsnrnx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqsnrnx1

MACRO snl_lqsnrnx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqsnrnx2

MACRO snl_lqsnrnx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqsnrnx4

MACRO snl_lqsnx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN SN DIRECTION INPUT ; END SN
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqsnx1

MACRO snl_lqsnx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN SN DIRECTION INPUT ; END SN
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqsnx2

MACRO snl_lqsnx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN SN DIRECTION INPUT ; END SN
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqsnx4

MACRO snl_lqx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqx1

MACRO snl_lqx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqx2

MACRO snl_lqx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_lqx4

MACRO snl_mux21x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN S DIRECTION INPUT ; END S
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_mux21x1

MACRO snl_mux21x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN S DIRECTION INPUT ; END S
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_mux21x2

MACRO snl_mux21x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN S DIRECTION INPUT ; END S
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_mux21x4

MACRO snl_mux21x8
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN S DIRECTION INPUT ; END S
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_mux21x8

MACRO snl_mux42x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN S1 DIRECTION INPUT ; END S1
 PIN S2 DIRECTION INPUT ; END S2
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_mux42x1

MACRO snl_mux42x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN S1 DIRECTION INPUT ; END S1
 PIN S2 DIRECTION INPUT ; END S2
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_mux42x2

MACRO snl_mux42x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN S1 DIRECTION INPUT ; END S1
 PIN S2 DIRECTION INPUT ; END S2
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_mux42x4

MACRO snl_mux42x8
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN S1 DIRECTION INPUT ; END S1
 PIN S2 DIRECTION INPUT ; END S2
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_mux42x8

MACRO snl_muxi21x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN S DIRECTION INPUT ; END S
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_muxi21x1

MACRO snl_muxi21x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN S DIRECTION INPUT ; END S
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_muxi21x2

MACRO snl_muxi21x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN S DIRECTION INPUT ; END S
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_muxi21x4

MACRO snl_muxi21x8
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN S DIRECTION INPUT ; END S
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_muxi21x8

MACRO snl_muxi42x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN S1 DIRECTION INPUT ; END S1
 PIN S2 DIRECTION INPUT ; END S2
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_muxi42x0

MACRO snl_muxi42x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN S1 DIRECTION INPUT ; END S1
 PIN S2 DIRECTION INPUT ; END S2
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_muxi42x1

MACRO snl_muxi42x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN S1 DIRECTION INPUT ; END S1
 PIN S2 DIRECTION INPUT ; END S2
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_muxi42x2

MACRO snl_muxi42x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN S1 DIRECTION INPUT ; END S1
 PIN S2 DIRECTION INPUT ; END S2
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_muxi42x4

MACRO snl_muxi42x8
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN S1 DIRECTION INPUT ; END S1
 PIN S2 DIRECTION INPUT ; END S2
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_muxi42x8

MACRO snl_nand02x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand02x1

MACRO snl_nand02x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand02x2

MACRO snl_nand02x3
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand02x3

MACRO snl_nand02x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand02x4

MACRO snl_nand02x8
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand02x8

MACRO snl_nand03x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand03x0

MACRO snl_nand03x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand03x1

MACRO snl_nand03x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand03x2

MACRO snl_nand03x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand03x4

MACRO snl_nand03x8
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand03x8

MACRO snl_nand04x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand04x0

MACRO snl_nand04x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand04x1

MACRO snl_nand04x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand04x2

MACRO snl_nand04x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand04x4

MACRO snl_nand04x8
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand04x8

MACRO snl_nand05x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand05x1

MACRO snl_nand05x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand05x2

MACRO snl_nand05x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand05x4

MACRO snl_nand05x8
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand05x8

MACRO snl_nand06x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand06x1

MACRO snl_nand06x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand06x2

MACRO snl_nand06x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand06x4

MACRO snl_nand06x8
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand06x8

MACRO snl_nand08x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand08x1

MACRO snl_nand08x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand08x2

MACRO snl_nand08x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand08x4

MACRO snl_nand08x8
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand08x8

MACRO snl_nand12x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand12x1

MACRO snl_nand12x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand12x2

MACRO snl_nand12x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand12x4

MACRO snl_nand12x8
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand12x8

MACRO snl_nand13x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand13x1

MACRO snl_nand13x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand13x2

MACRO snl_nand13x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand13x4

MACRO snl_nand13x8
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand13x8

MACRO snl_nand14x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand14x0

MACRO snl_nand14x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand14x1

MACRO snl_nand14x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand14x2

MACRO snl_nand14x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand14x4

MACRO snl_nand14x8
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand14x8

MACRO snl_nand23x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand23x1

MACRO snl_nand23x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand23x2

MACRO snl_nand23x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand23x4

MACRO snl_nand23x8
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand23x8

MACRO snl_nand24x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand24x0

MACRO snl_nand24x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand24x1

MACRO snl_nand24x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand24x2

MACRO snl_nand24x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand24x4

MACRO snl_nand24x8
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand24x8

MACRO snl_nand34x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand34x1

MACRO snl_nand34x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand34x2

MACRO snl_nand34x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand34x4

MACRO snl_nand34x8
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nand34x8

MACRO snl_nor02x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nor02x1

MACRO snl_nor02x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nor02x2

MACRO snl_nor02x3
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nor02x3

MACRO snl_nor02x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nor02x4

MACRO snl_nor02x8
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nor02x8

MACRO snl_nor03x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nor03x0

MACRO snl_nor03x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nor03x1

MACRO snl_nor03x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nor03x2

MACRO snl_nor03x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nor03x4

MACRO snl_nor03x8
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nor03x8

MACRO snl_nor04x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nor04x0

MACRO snl_nor04x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nor04x1

MACRO snl_nor04x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nor04x2

MACRO snl_nor04x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nor04x4

MACRO snl_nor04x8
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nor04x8

MACRO snl_nor05x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nor05x1

MACRO snl_nor05x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nor05x2

MACRO snl_nor05x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nor05x4

MACRO snl_nor05x8
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nor05x8

MACRO snl_nor06x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nor06x1

MACRO snl_nor06x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nor06x2

MACRO snl_nor06x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nor06x4

MACRO snl_nor06x8
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nor06x8

MACRO snl_nor08x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nor08x1

MACRO snl_nor08x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nor08x2

MACRO snl_nor08x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nor08x4

MACRO snl_nor08x8
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nor08x8

MACRO snl_oa012x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa012x1

MACRO snl_oa012x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa012x2

MACRO snl_oa012x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa012x4

MACRO snl_oa013x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa013x1

MACRO snl_oa013x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa013x2

MACRO snl_oa013x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa013x4

MACRO snl_oa022x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa022x1

MACRO snl_oa022x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa022x2

MACRO snl_oa022x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa022x4

MACRO snl_oa023x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa023x1

MACRO snl_oa023x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa023x2

MACRO snl_oa023x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa023x4

MACRO snl_oa033x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa033x1

MACRO snl_oa033x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa033x2

MACRO snl_oa033x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa033x4

MACRO snl_oa112x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa112x1

MACRO snl_oa112x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa112x2

MACRO snl_oa112x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa112x4

MACRO snl_oa113x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa113x1

MACRO snl_oa113x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa113x2

MACRO snl_oa113x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa113x4

MACRO snl_oa122x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa122x1

MACRO snl_oa122x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa122x2

MACRO snl_oa122x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa122x4

MACRO snl_oa123x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa123x1

MACRO snl_oa123x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa123x2

MACRO snl_oa123x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa123x4

MACRO snl_oa133x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa133x1

MACRO snl_oa133x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa133x2

MACRO snl_oa133x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa133x4

MACRO snl_oa2222x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa2222x1

MACRO snl_oa2222x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa2222x2

MACRO snl_oa2222x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa2222x4

MACRO snl_oa222x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa222x1

MACRO snl_oa222x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa222x2

MACRO snl_oa222x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa222x4

MACRO snl_oa223x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa223x1

MACRO snl_oa223x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa223x2

MACRO snl_oa223x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa223x4

MACRO snl_oa233x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa233x1

MACRO snl_oa233x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa233x2

MACRO snl_oa233x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa233x4

MACRO snl_oa333x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN I DIRECTION INPUT ; END I
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa333x1

MACRO snl_oa333x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN I DIRECTION INPUT ; END I
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa333x2

MACRO snl_oa333x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN I DIRECTION INPUT ; END I
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oa333x4

MACRO snl_oai012x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai012x1

MACRO snl_oai012x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai012x2

MACRO snl_oai012x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai012x4

MACRO snl_oai013x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai013x0

MACRO snl_oai013x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai013x1

MACRO snl_oai013x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai013x2

MACRO snl_oai013x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai013x4

MACRO snl_oai022x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai022x1

MACRO snl_oai022x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai022x2

MACRO snl_oai022x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai022x4

MACRO snl_oai023x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai023x0

MACRO snl_oai023x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai023x1

MACRO snl_oai023x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai023x2

MACRO snl_oai023x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai023x4

MACRO snl_oai033x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai033x0

MACRO snl_oai033x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai033x1

MACRO snl_oai033x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai033x2

MACRO snl_oai033x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai033x4

MACRO snl_oai112x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai112x0

MACRO snl_oai112x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai112x1

MACRO snl_oai112x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai112x2

MACRO snl_oai112x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai112x4

MACRO snl_oai113x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai113x0

MACRO snl_oai113x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai113x1

MACRO snl_oai113x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai113x2

MACRO snl_oai113x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai113x4

MACRO snl_oai122x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai122x0

MACRO snl_oai122x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai122x1

MACRO snl_oai122x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai122x2

MACRO snl_oai122x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai122x4

MACRO snl_oai123x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai123x0

MACRO snl_oai123x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai123x1

MACRO snl_oai123x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai123x2

MACRO snl_oai123x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai123x4

MACRO snl_oai133x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai133x0

MACRO snl_oai133x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai133x1

MACRO snl_oai133x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai133x2

MACRO snl_oai133x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai133x4

MACRO snl_oai2222x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai2222x0

MACRO snl_oai2222x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai2222x1

MACRO snl_oai2222x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai2222x2

MACRO snl_oai2222x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai2222x4

MACRO snl_oai222x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai222x0

MACRO snl_oai222x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai222x1

MACRO snl_oai222x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai222x2

MACRO snl_oai222x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai222x4

MACRO snl_oai223x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai223x0

MACRO snl_oai223x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai223x1

MACRO snl_oai223x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai223x2

MACRO snl_oai223x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai223x4

MACRO snl_oai233x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai233x0

MACRO snl_oai233x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai233x1

MACRO snl_oai233x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai233x2

MACRO snl_oai233x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai233x4

MACRO snl_oai333x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN I DIRECTION INPUT ; END I
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai333x0

MACRO snl_oai333x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN I DIRECTION INPUT ; END I
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai333x1

MACRO snl_oai333x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN I DIRECTION INPUT ; END I
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai333x2

MACRO snl_oai333x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN I DIRECTION INPUT ; END I
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_oai333x4

MACRO snl_or02x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_or02x1

MACRO snl_or02x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_or02x2

MACRO snl_or02x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_or02x4

MACRO snl_or02x8
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_or02x8

MACRO snl_or03x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_or03x1

MACRO snl_or03x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_or03x2

MACRO snl_or03x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_or03x4

MACRO snl_or03x8
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_or03x8

MACRO snl_or04x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_or04x1

MACRO snl_or04x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_or04x2

MACRO snl_or04x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_or04x4

MACRO snl_or04x8
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_or04x8

MACRO snl_or05x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_or05x1

MACRO snl_or05x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_or05x2

MACRO snl_or05x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_or05x4

MACRO snl_or05x8
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_or05x8

MACRO snl_or06x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_or06x1

MACRO snl_or06x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_or06x2

MACRO snl_or06x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_or06x4

MACRO snl_or06x8
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_or06x8

MACRO snl_or08x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_or08x1

MACRO snl_or08x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_or08x2

MACRO snl_or08x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_or08x4

MACRO snl_or08x8
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN D DIRECTION INPUT ; END D
 PIN E DIRECTION INPUT ; END E
 PIN F DIRECTION INPUT ; END F
 PIN G DIRECTION INPUT ; END G
 PIN H DIRECTION INPUT ; END H
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_or08x8

MACRO snl_rep
 SIZE 50 BY 20 ;
 PIN I DIRECTION INOUT ; END I
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_rep

MACRO snl_sffandnorx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffandnorx1

MACRO snl_sffandnorx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffandnorx2

MACRO snl_sffandnorx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffandnorx4

MACRO snl_sffandorx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffandorx1

MACRO snl_sffandorx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffandorx2

MACRO snl_sffandorx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffandorx4

MACRO snl_sffandx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffandx1

MACRO snl_sffandx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffandx2

MACRO snl_sffandx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffandx4

MACRO snl_sffmu2x1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN S DIRECTION INPUT ; END S
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffmu2x1

MACRO snl_sffmu2x2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN S DIRECTION INPUT ; END S
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffmu2x2

MACRO snl_sffmu2x4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN S DIRECTION INPUT ; END S
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffmu2x4

MACRO snl_sffnandx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffnandx1

MACRO snl_sffnandx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffnandx2

MACRO snl_sffnandx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffnandx4

MACRO snl_sffnorx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffnorx1

MACRO snl_sffnorx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffnorx2

MACRO snl_sffnorx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffnorx4

MACRO snl_sfforandx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sfforandx1

MACRO snl_sfforandx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sfforandx2

MACRO snl_sfforandx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sfforandx4

MACRO snl_sffornandx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffornandx1

MACRO snl_sffornandx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffornandx2

MACRO snl_sffornandx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffornandx4

MACRO snl_sfforx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sfforx1

MACRO snl_sfforx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sfforx2

MACRO snl_sfforx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sfforx4

MACRO snl_sffqenrnx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN RN DIRECTION INPUT ; END RN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqenrnx1

MACRO snl_sffqenrnx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN RN DIRECTION INPUT ; END RN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqenrnx2

MACRO snl_sffqenrnx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN RN DIRECTION INPUT ; END RN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqenrnx4

MACRO snl_sffqensnx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN SN DIRECTION INPUT ; END SN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqensnx1

MACRO snl_sffqensnx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN SN DIRECTION INPUT ; END SN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqensnx2

MACRO snl_sffqensnx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN SN DIRECTION INPUT ; END SN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqensnx4

MACRO snl_sffqenx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqenx1

MACRO snl_sffqenx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqenx2

MACRO snl_sffqenx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqenx4

MACRO snl_sffqnenrnx1
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN RN DIRECTION INPUT ; END RN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqnenrnx1

MACRO snl_sffqnenrnx2
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN RN DIRECTION INPUT ; END RN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqnenrnx2

MACRO snl_sffqnenrnx4
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN RN DIRECTION INPUT ; END RN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqnenrnx4

MACRO snl_sffqnensnx1
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN SN DIRECTION INPUT ; END SN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqnensnx1

MACRO snl_sffqnensnx2
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN SN DIRECTION INPUT ; END SN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqnensnx2

MACRO snl_sffqnensnx4
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN SN DIRECTION INPUT ; END SN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqnensnx4

MACRO snl_sffqnenx1
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqnenx1

MACRO snl_sffqnenx2
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqnenx2

MACRO snl_sffqnenx4
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqnenx4

MACRO snl_sffqnrnx1
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqnrnx1

MACRO snl_sffqnrnx2
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqnrnx2

MACRO snl_sffqnrnx4
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqnrnx4

MACRO snl_sffqnsnx1
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN SN DIRECTION INPUT ; END SN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqnsnx1

MACRO snl_sffqnsnx2
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN SN DIRECTION INPUT ; END SN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqnsnx2

MACRO snl_sffqnsnx4
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN SN DIRECTION INPUT ; END SN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqnsnx4

MACRO snl_sffqnx1
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqnx1

MACRO snl_sffqnx2
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqnx2

MACRO snl_sffqnx4
 SIZE 50 BY 20 ;
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqnx4

MACRO snl_sffqqnenrnx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN RN DIRECTION INPUT ; END RN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqqnenrnx1

MACRO snl_sffqqnenrnx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN RN DIRECTION INPUT ; END RN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqqnenrnx2

MACRO snl_sffqqnensnx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN SN DIRECTION INPUT ; END SN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqqnensnx1

MACRO snl_sffqqnensnx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN SN DIRECTION INPUT ; END SN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqqnensnx2

MACRO snl_sffqqnenx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqqnenx1

MACRO snl_sffqqnenx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN EN DIRECTION INPUT ; END EN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqqnenx2

MACRO snl_sffqqnrnsnx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqqnrnsnx1

MACRO snl_sffqqnrnsnx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SN DIRECTION INPUT ; END SN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqqnrnsnx2

MACRO snl_sffqqnrnx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqqnrnx1

MACRO snl_sffqqnrnx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqqnrnx2

MACRO snl_sffqqnsnx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN SN DIRECTION INPUT ; END SN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqqnsnx1

MACRO snl_sffqqnsnx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN SN DIRECTION INPUT ; END SN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqqnsnx2

MACRO snl_sffqqnx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqqnx1

MACRO snl_sffqqnx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN QN DIRECTION OUTPUT ; END QN
 PIN D DIRECTION INPUT ; END D
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqqnx2

MACRO snl_sffqrnx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqrnx1

MACRO snl_sffqrnx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqrnx2

MACRO snl_sffqrnx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN RN DIRECTION INPUT ; END RN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqrnx4

MACRO snl_sffqsnx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN SN DIRECTION INPUT ; END SN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqsnx1

MACRO snl_sffqsnx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN SN DIRECTION INPUT ; END SN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqsnx2

MACRO snl_sffqsnx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN SN DIRECTION INPUT ; END SN
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqsnx4

MACRO snl_sffqx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqx1

MACRO snl_sffqx2
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqx2

MACRO snl_sffqx4
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN SD DIRECTION INPUT ; END SD
 PIN SE DIRECTION INPUT ; END SE
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_sffqx4

MACRO snl_tbufx1
 SIZE 50 BY 20 ;
 PIN A DIRECTION INPUT ; END A
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_tbufx1

MACRO snl_tbufx12
 SIZE 50 BY 20 ;
 PIN A DIRECTION INPUT ; END A
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_tbufx12

MACRO snl_tbufx2
 SIZE 50 BY 20 ;
 PIN A DIRECTION INPUT ; END A
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_tbufx2

MACRO snl_tbufx4
 SIZE 50 BY 20 ;
 PIN A DIRECTION INPUT ; END A
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_tbufx4

MACRO snl_tbufx8
 SIZE 50 BY 20 ;
 PIN A DIRECTION INPUT ; END A
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_tbufx8

MACRO snl_tinvx1
 SIZE 50 BY 20 ;
 PIN A DIRECTION INPUT ; END A
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_tinvx1

MACRO snl_tinvx12
 SIZE 50 BY 20 ;
 PIN A DIRECTION INPUT ; END A
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_tinvx12

MACRO snl_tinvx2
 SIZE 50 BY 20 ;
 PIN A DIRECTION INPUT ; END A
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_tinvx2

MACRO snl_tinvx4
 SIZE 50 BY 20 ;
 PIN A DIRECTION INPUT ; END A
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_tinvx4

MACRO snl_tinvx8
 SIZE 50 BY 20 ;
 PIN A DIRECTION INPUT ; END A
 PIN E DIRECTION INPUT ; END E
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_tinvx8

MACRO snl_xnor2x0
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_xnor2x0

MACRO snl_xnor2x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_xnor2x1

MACRO snl_xnor2x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_xnor2x2

MACRO snl_xnor2x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_xnor2x4

MACRO snl_xnor2x8
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_xnor2x8

MACRO snl_xnor3x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_xnor3x1

MACRO snl_xnor3x2
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_xnor3x2

MACRO snl_xnor3x4
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_xnor3x4

MACRO snl_xnor3x8
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_xnor3x8

MACRO snl_xor2x0
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_xor2x0

MACRO snl_xor2x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_xor2x1

MACRO snl_xor2x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_xor2x2

MACRO snl_xor2x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_xor2x4

MACRO snl_xor2x8
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_xor2x8

MACRO snl_xor3x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_xor3x1

MACRO snl_xor3x2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_xor3x2

MACRO snl_xor3x4
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_xor3x4

MACRO snl_xor3x8
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN C DIRECTION INPUT ; END C
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_xor3x8

END LIBRARY
