module test (
  sig1,
  sig2,
  sig3,
  sig4,
  sig5,
  sig6,
  sig7,
  sig8,
  sig9,
  sig10,
  sig11,
  sig12,
  sig13,
  sig14,
  sig15,
  sig16,
  sig17,
  sig18,
  sig19,
  sig20,
  sig21,
  sig22,
  sig23,
  sig24,
  sig25,
  sig26,
  sig27,
  sig28,
  sig29,
  sig30,
  sig31,
  sig32,
  sig33,
  sig34,
  sig35,
  sig36,
  sig37,
  sig38,
  sig39,
  sig40,
  sig41,
  sig42,
  sig43,
  sig44,
  sig45,
  sig46,
  sig47,
  sig48,
  sig49,
  sig50,
  sig51,
  sig52,
  sig53,
  sig54,
  sig55,
  sig56,
  sig57,
  sig58,
  sig59,
  sig60,
  sig61,
  sig62,
  sig63,
  sig64,
  sig65,
  sig66,
  sig67,
  sig68,
  sig69,
  sig70,
  sig71,
  sig72,
  sig73,
  sig74,
  sig75,
  sig76,
  sig77,
  sig78,
  sig79,
  sig80,
  sig81,
  sig82,
  sig83,
  sig84,
  sig85,
  sig86,
  sig87,
  sig88,
  sig89,
  sig90,
  sig91,
  sig92,
  sig93,
  sig94,
  sig95,
  sig96,
  sig97,
  sig98,
  sig99,
  sig100,
  sig101,
  sig102,
  sig103,
  sig104,
  sig105,
  sig106,
  sig107,
  sig108,
  sig109,
  sig110,
  sig111,
  sig112,
  sig113,
  sig114,
  sig115,
  sig116,
  sig117,
  sig118,
  sig119,
  sig120,
  sig121,
  sig122,
  sig123,
  sig124,
  sig125,
  sig126,
  sig127,
  sig128,
  sig129,
  sig130,
  sig131,
  sig132,
  sig133,
  sig134,
  sig135,
  sig136,
  sig137,
  sig138,
  sig139,
  sig140,
  sig141,
  sig142,
  sig143,
  sig144,
  sig145,
  sig146,
  sig147,
  sig148,
  sig149,
  sig150,
  sig151,
  sig152,
  sig153,
  sig154,
  sig155,
  sig156,
  sig157,
  sig158,
  sig159,
  sig160,
  sig161,
  sig162,
  sig163,
  sig164,
  sig165,
  sig166,
  sig167,
  sig168,
  sig169,
  sig170,
  sig171,
  sig172,
  sig173,
  sig174,
  sig175,
  sig176,
  sig177,
  sig178,
  sig179,
  sig180,
  sig181,
  sig182,
  sig183,
  sig184,
  sig185,
  sig186,
  sig187,
  sig188,
  sig189,
  sig190,
  sig191,
  sig192,
  sig193,
  sig194,
  sig195,
  sig196,
  sig197,
  sig198,
  sig199,
  sig200,
  sig201,
  sig202,
  sig203,
  sig204,
  sig205,
  sig206,
  sig207,
  sig208,
  sig209,
  sig210,
  sig211,
  sig212,
  sig213,
  sig214,
  sig215,
  sig216,
  sig217,
  sig218,
  sig219,
  sig220,
  sig221,
  sig222,
  sig223,
  sig224,
  sig225,
  sig226,
  sig227,
  sig228,
  sig229,
  sig230,
  sig231,
  sig232,
  sig233,
  sig234,
  sig235,
  sig236,
  sig237,
  sig238,
  sig239,
  sig240,
  sig241,
  sig242,
  sig243,
  sig244,
  sig245,
  sig246,
  sig247,
  sig248,
  sig249,
  sig250,
  sig251,
  sig252
) ;
  output sig1 ;
  input  sig2 ;
  output sig3 ;
  input  sig4 ;
  output sig5 ;
  input  sig6 ;
  output sig7 ;
  input  sig8 ;
  output sig9 ;
  input  sig10 ;
  output sig11 ;
  input  sig12 ;
  output sig13 ;
  input  sig14 ;
  output sig15 ;
  input  sig16 ;
  output sig17 ;
  input  sig18 ;
  output sig19 ;
  input  sig20 ;
  output sig21 ;
  input  sig22 ;
  output sig23 ;
  input  sig24 ;
  output sig25 ;
  input  sig26 ;
  output sig27 ;
  input  sig28 ;
  output sig29 ;
  input  sig30 ;
  output sig31 ;
  input  sig32 ;
  output sig33 ;
  input  sig34 ;
  output sig35 ;
  input  sig36 ;
  output sig37 ;
  input  sig38 ;
  output sig39 ;
  input  sig40 ;
  output sig41 ;
  input  sig42 ;
  output sig43 ;
  input  sig44 ;
  output sig45 ;
  input  sig46 ;
  output sig47 ;
  input  sig48 ;
  output sig49 ;
  input  sig50 ;
  output sig51 ;
  input  sig52 ;
  output sig53 ;
  input  sig54 ;
  output sig55 ;
  input  sig56 ;
  output sig57 ;
  input  sig58 ;
  output sig59 ;
  input  sig60 ;
  output sig61 ;
  input  sig62 ;
  output sig63 ;
  input  sig64 ;
  output sig65 ;
  input  sig66 ;
  output sig67 ;
  input  sig68 ;
  output sig69 ;
  input  sig70 ;
  output sig71 ;
  input  sig72 ;
  output sig73 ;
  input  sig74 ;
  output sig75 ;
  input  sig76 ;
  output sig77 ;
  input  sig78 ;
  output sig79 ;
  input  sig80 ;
  output sig81 ;
  input  sig82 ;
  output sig83 ;
  input  sig84 ;
  output sig85 ;
  input  sig86 ;
  output sig87 ;
  input  sig88 ;
  output sig89 ;
  input  sig90 ;
  output sig91 ;
  input  sig92 ;
  output sig93 ;
  input  sig94 ;
  output sig95 ;
  input  sig96 ;
  output sig97 ;
  input  sig98 ;
  output sig99 ;
  input  sig100 ;
  output sig101 ;
  input  sig102 ;
  output sig103 ;
  input  sig104 ;
  output sig105 ;
  input  sig106 ;
  output sig107 ;
  input  sig108 ;
  output sig109 ;
  input  sig110 ;
  output sig111 ;
  input  sig112 ;
  output sig113 ;
  input  sig114 ;
  output sig115 ;
  input  sig116 ;
  output sig117 ;
  input  sig118 ;
  output sig119 ;
  input  sig120 ;
  output sig121 ;
  input  sig122 ;
  output sig123 ;
  input  sig124 ;
  output sig125 ;
  input  sig126 ;
  output sig127 ;
  input  sig128 ;
  output sig129 ;
  input  sig130 ;
  output sig131 ;
  input  sig132 ;
  output sig133 ;
  input  sig134 ;
  output sig135 ;
  input  sig136 ;
  output sig137 ;
  input  sig138 ;
  output sig139 ;
  input  sig140 ;
  output sig141 ;
  input  sig142 ;
  output sig143 ;
  input  sig144 ;
  output sig145 ;
  input  sig146 ;
  output sig147 ;
  input  sig148 ;
  output sig149 ;
  input  sig150 ;
  output sig151 ;
  input  sig152 ;
  output sig153 ;
  input  sig154 ;
  output sig155 ;
  input  sig156 ;
  output sig157 ;
  input  sig158 ;
  output sig159 ;
  input  sig160 ;
  output sig161 ;
  input  sig162 ;
  output sig163 ;
  input  sig164 ;
  output sig165 ;
  input  sig166 ;
  output sig167 ;
  input  sig168 ;
  output sig169 ;
  input  sig170 ;
  output sig171 ;
  input  sig172 ;
  output sig173 ;
  input  sig174 ;
  output sig175 ;
  input  sig176 ;
  output sig177 ;
  input  sig178 ;
  output sig179 ;
  input  sig180 ;
  output sig181 ;
  input  sig182 ;
  output sig183 ;
  input  sig184 ;
  output sig185 ;
  input  sig186 ;
  output sig187 ;
  input  sig188 ;
  output sig189 ;
  input  sig190 ;
  output sig191 ;
  input  sig192 ;
  output sig193 ;
  input  sig194 ;
  output sig195 ;
  input  sig196 ;
  output sig197 ;
  input  sig198 ;
  output sig199 ;
  input  sig200 ;
  output sig201 ;
  input  sig202 ;
  output sig203 ;
  input  sig204 ;
  output sig205 ;
  input  sig206 ;
  output sig207 ;
  input  sig208 ;
  output sig209 ;
  input  sig210 ;
  output sig211 ;
  input  sig212 ;
  output sig213 ;
  input  sig214 ;
  output sig215 ;
  input  sig216 ;
  output sig217 ;
  input  sig218 ;
  output sig219 ;
  input  sig220 ;
  output sig221 ;
  input  sig222 ;
  output sig223 ;
  input  sig224 ;
  output sig225 ;
  input  sig226 ;
  output sig227 ;
  input  sig228 ;
  output sig229 ;
  input  sig230 ;
  output sig231 ;
  input  sig232 ;
  output sig233 ;
  input  sig234 ;
  output sig235 ;
  input  sig236 ;
  output sig237 ;
  input  sig238 ;
  output sig239 ;
  input  sig240 ;
  output sig241 ;
  input  sig242 ;
  output sig243 ;
  input  sig244 ;
  output sig245 ;
  input  sig246 ;
  output sig247 ;
  input  sig248 ;
  output sig249 ;
  input  sig250 ;
  output sig251 ;
  input  sig252 ;
  PADCELL_SIG_V u_sig1 (.PAD(sig1), .A(core_sig1));
  PADCELL_SIG_V u_sig2 (.PAD(sig2), .Y(core_sig2));
  PADCELL_SIG_V u_sig3 (.PAD(sig3), .A(core_sig3));
  PADCELL_SIG_V u_sig4 (.PAD(sig4), .Y(core_sig4));
  PADCELL_SIG_V u_sig5 (.PAD(sig5), .A(core_sig5));
  PADCELL_SIG_V u_sig6 (.PAD(sig6), .Y(core_sig6));
  PADCELL_SIG_V u_sig7 (.PAD(sig7), .A(core_sig7));
  PADCELL_SIG_V u_sig8 (.PAD(sig8), .Y(core_sig8));
  PADCELL_SIG_V u_sig9 (.PAD(sig9), .A(core_sig9));
  PADCELL_SIG_V u_sig10 (.PAD(sig10), .Y(core_sig10));
  PADCELL_SIG_V u_sig11 (.PAD(sig11), .A(core_sig11));
  PADCELL_SIG_V u_sig12 (.PAD(sig12), .Y(core_sig12));
  PADCELL_SIG_V u_sig13 (.PAD(sig13), .A(core_sig13));
  PADCELL_SIG_V u_sig14 (.PAD(sig14), .Y(core_sig14));
  PADCELL_SIG_V u_sig15 (.PAD(sig15), .A(core_sig15));
  PADCELL_SIG_V u_sig16 (.PAD(sig16), .Y(core_sig16));
  PADCELL_SIG_V u_sig17 (.PAD(sig17), .A(core_sig17));
  PADCELL_SIG_V u_sig18 (.PAD(sig18), .Y(core_sig18));
  PADCELL_SIG_V u_sig19 (.PAD(sig19), .A(core_sig19));
  PADCELL_SIG_V u_sig20 (.PAD(sig20), .Y(core_sig20));
  PADCELL_SIG_V u_sig21 (.PAD(sig21), .A(core_sig21));
  PADCELL_SIG_V u_sig22 (.PAD(sig22), .Y(core_sig22));
  PADCELL_SIG_V u_sig23 (.PAD(sig23), .A(core_sig23));
  PADCELL_SIG_V u_sig24 (.PAD(sig24), .Y(core_sig24));
  PADCELL_SIG_V u_sig25 (.PAD(sig25), .A(core_sig25));
  PADCELL_SIG_V u_sig26 (.PAD(sig26), .Y(core_sig26));
  PADCELL_SIG_V u_sig27 (.PAD(sig27), .A(core_sig27));
  PADCELL_SIG_V u_sig28 (.PAD(sig28), .Y(core_sig28));
  PADCELL_SIG_V u_sig29 (.PAD(sig29), .A(core_sig29));
  PADCELL_SIG_V u_sig30 (.PAD(sig30), .Y(core_sig30));
  PADCELL_SIG_V u_sig31 (.PAD(sig31), .A(core_sig31));
  PADCELL_SIG_V u_sig32 (.PAD(sig32), .Y(core_sig32));
  PADCELL_SIG_V u_sig33 (.PAD(sig33), .A(core_sig33));
  PADCELL_SIG_V u_sig34 (.PAD(sig34), .Y(core_sig34));
  PADCELL_SIG_V u_sig35 (.PAD(sig35), .A(core_sig35));
  PADCELL_SIG_V u_sig36 (.PAD(sig36), .Y(core_sig36));
  PADCELL_SIG_V u_sig37 (.PAD(sig37), .A(core_sig37));
  PADCELL_SIG_V u_sig38 (.PAD(sig38), .Y(core_sig38));
  PADCELL_SIG_V u_sig39 (.PAD(sig39), .A(core_sig39));
  PADCELL_SIG_V u_sig40 (.PAD(sig40), .Y(core_sig40));
  PADCELL_SIG_V u_sig41 (.PAD(sig41), .A(core_sig41));
  PADCELL_SIG_V u_sig42 (.PAD(sig42), .Y(core_sig42));
  PADCELL_SIG_V u_sig43 (.PAD(sig43), .A(core_sig43));
  PADCELL_SIG_V u_sig44 (.PAD(sig44), .Y(core_sig44));
  PADCELL_SIG_V u_sig45 (.PAD(sig45), .A(core_sig45));
  PADCELL_SIG_V u_sig46 (.PAD(sig46), .Y(core_sig46));
  PADCELL_SIG_V u_sig47 (.PAD(sig47), .A(core_sig47));
  PADCELL_SIG_V u_sig48 (.PAD(sig48), .Y(core_sig48));
  PADCELL_SIG_V u_sig49 (.PAD(sig49), .A(core_sig49));
  PADCELL_SIG_V u_sig50 (.PAD(sig50), .Y(core_sig50));
  PADCELL_SIG_V u_sig51 (.PAD(sig51), .A(core_sig51));
  PADCELL_SIG_V u_sig52 (.PAD(sig52), .Y(core_sig52));
  PADCELL_SIG_V u_sig53 (.PAD(sig53), .A(core_sig53));
  PADCELL_SIG_V u_sig54 (.PAD(sig54), .Y(core_sig54));
  PADCELL_SIG_V u_sig55 (.PAD(sig55), .A(core_sig55));
  PADCELL_SIG_V u_sig56 (.PAD(sig56), .Y(core_sig56));
  PADCELL_SIG_V u_sig57 (.PAD(sig57), .A(core_sig57));
  PADCELL_SIG_V u_sig58 (.PAD(sig58), .Y(core_sig58));
  PADCELL_SIG_V u_sig59 (.PAD(sig59), .A(core_sig59));
  PADCELL_SIG_V u_sig60 (.PAD(sig60), .Y(core_sig60));
  PADCELL_SIG_V u_sig61 (.PAD(sig61), .A(core_sig61));
  PADCELL_SIG_V u_sig62 (.PAD(sig62), .Y(core_sig62));
  PADCELL_SIG_V u_sig63 (.PAD(sig63), .A(core_sig63));
  PADCELL_SIG_H u_sig64 (.PAD(sig64), .Y(core_sig64));
  PADCELL_SIG_H u_sig65 (.PAD(sig65), .A(core_sig65));
  PADCELL_SIG_H u_sig66 (.PAD(sig66), .Y(core_sig66));
  PADCELL_SIG_H u_sig67 (.PAD(sig67), .A(core_sig67));
  PADCELL_SIG_H u_sig68 (.PAD(sig68), .Y(core_sig68));
  PADCELL_SIG_H u_sig69 (.PAD(sig69), .A(core_sig69));
  PADCELL_SIG_H u_sig70 (.PAD(sig70), .Y(core_sig70));
  PADCELL_SIG_H u_sig71 (.PAD(sig71), .A(core_sig71));
  PADCELL_SIG_H u_sig72 (.PAD(sig72), .Y(core_sig72));
  PADCELL_SIG_H u_sig73 (.PAD(sig73), .A(core_sig73));
  PADCELL_SIG_H u_sig74 (.PAD(sig74), .Y(core_sig74));
  PADCELL_SIG_H u_sig75 (.PAD(sig75), .A(core_sig75));
  PADCELL_SIG_H u_sig76 (.PAD(sig76), .Y(core_sig76));
  PADCELL_SIG_H u_sig77 (.PAD(sig77), .A(core_sig77));
  PADCELL_SIG_H u_sig78 (.PAD(sig78), .Y(core_sig78));
  PADCELL_SIG_H u_sig79 (.PAD(sig79), .A(core_sig79));
  PADCELL_SIG_H u_sig80 (.PAD(sig80), .Y(core_sig80));
  PADCELL_SIG_H u_sig81 (.PAD(sig81), .A(core_sig81));
  PADCELL_SIG_H u_sig82 (.PAD(sig82), .Y(core_sig82));
  PADCELL_SIG_H u_sig83 (.PAD(sig83), .A(core_sig83));
  PADCELL_SIG_H u_sig84 (.PAD(sig84), .Y(core_sig84));
  PADCELL_SIG_H u_sig85 (.PAD(sig85), .A(core_sig85));
  PADCELL_SIG_H u_sig86 (.PAD(sig86), .Y(core_sig86));
  PADCELL_SIG_H u_sig87 (.PAD(sig87), .A(core_sig87));
  PADCELL_SIG_H u_sig88 (.PAD(sig88), .Y(core_sig88));
  PADCELL_SIG_H u_sig89 (.PAD(sig89), .A(core_sig89));
  PADCELL_SIG_H u_sig90 (.PAD(sig90), .Y(core_sig90));
  PADCELL_SIG_H u_sig91 (.PAD(sig91), .A(core_sig91));
  PADCELL_SIG_H u_sig92 (.PAD(sig92), .Y(core_sig92));
  PADCELL_SIG_H u_sig93 (.PAD(sig93), .A(core_sig93));
  PADCELL_SIG_H u_sig94 (.PAD(sig94), .Y(core_sig94));
  PADCELL_SIG_H u_sig95 (.PAD(sig95), .A(core_sig95));
  PADCELL_SIG_H u_sig96 (.PAD(sig96), .Y(core_sig96));
  PADCELL_SIG_H u_sig97 (.PAD(sig97), .A(core_sig97));
  PADCELL_SIG_H u_sig98 (.PAD(sig98), .Y(core_sig98));
  PADCELL_SIG_H u_sig99 (.PAD(sig99), .A(core_sig99));
  PADCELL_SIG_H u_sig100 (.PAD(sig100), .Y(core_sig100));
  PADCELL_SIG_H u_sig101 (.PAD(sig101), .A(core_sig101));
  PADCELL_SIG_H u_sig102 (.PAD(sig102), .Y(core_sig102));
  PADCELL_SIG_H u_sig103 (.PAD(sig103), .A(core_sig103));
  PADCELL_SIG_H u_sig104 (.PAD(sig104), .Y(core_sig104));
  PADCELL_SIG_H u_sig105 (.PAD(sig105), .A(core_sig105));
  PADCELL_SIG_H u_sig106 (.PAD(sig106), .Y(core_sig106));
  PADCELL_SIG_H u_sig107 (.PAD(sig107), .A(core_sig107));
  PADCELL_SIG_H u_sig108 (.PAD(sig108), .Y(core_sig108));
  PADCELL_SIG_H u_sig109 (.PAD(sig109), .A(core_sig109));
  PADCELL_SIG_H u_sig110 (.PAD(sig110), .Y(core_sig110));
  PADCELL_SIG_H u_sig111 (.PAD(sig111), .A(core_sig111));
  PADCELL_SIG_H u_sig112 (.PAD(sig112), .Y(core_sig112));
  PADCELL_SIG_H u_sig113 (.PAD(sig113), .A(core_sig113));
  PADCELL_SIG_H u_sig114 (.PAD(sig114), .Y(core_sig114));
  PADCELL_SIG_H u_sig115 (.PAD(sig115), .A(core_sig115));
  PADCELL_SIG_H u_sig116 (.PAD(sig116), .Y(core_sig116));
  PADCELL_SIG_H u_sig117 (.PAD(sig117), .A(core_sig117));
  PADCELL_SIG_H u_sig118 (.PAD(sig118), .Y(core_sig118));
  PADCELL_SIG_H u_sig119 (.PAD(sig119), .A(core_sig119));
  PADCELL_SIG_H u_sig120 (.PAD(sig120), .Y(core_sig120));
  PADCELL_SIG_H u_sig121 (.PAD(sig121), .A(core_sig121));
  PADCELL_SIG_H u_sig122 (.PAD(sig122), .Y(core_sig122));
  PADCELL_SIG_H u_sig123 (.PAD(sig123), .A(core_sig123));
  PADCELL_SIG_H u_sig124 (.PAD(sig124), .Y(core_sig124));
  PADCELL_SIG_H u_sig125 (.PAD(sig125), .A(core_sig125));
  PADCELL_SIG_H u_sig126 (.PAD(sig126), .Y(core_sig126));
  PADCELL_SIG_V u_sig127 (.PAD(sig127), .A(core_sig127));
  PADCELL_SIG_V u_sig128 (.PAD(sig128), .Y(core_sig128));
  PADCELL_SIG_V u_sig129 (.PAD(sig129), .A(core_sig129));
  PADCELL_SIG_V u_sig130 (.PAD(sig130), .Y(core_sig130));
  PADCELL_SIG_V u_sig131 (.PAD(sig131), .A(core_sig131));
  PADCELL_SIG_V u_sig132 (.PAD(sig132), .Y(core_sig132));
  PADCELL_SIG_V u_sig133 (.PAD(sig133), .A(core_sig133));
  PADCELL_SIG_V u_sig134 (.PAD(sig134), .Y(core_sig134));
  PADCELL_SIG_V u_sig135 (.PAD(sig135), .A(core_sig135));
  PADCELL_SIG_V u_sig136 (.PAD(sig136), .Y(core_sig136));
  PADCELL_SIG_V u_sig137 (.PAD(sig137), .A(core_sig137));
  PADCELL_SIG_V u_sig138 (.PAD(sig138), .Y(core_sig138));
  PADCELL_SIG_V u_sig139 (.PAD(sig139), .A(core_sig139));
  PADCELL_SIG_V u_sig140 (.PAD(sig140), .Y(core_sig140));
  PADCELL_SIG_V u_sig141 (.PAD(sig141), .A(core_sig141));
  PADCELL_SIG_V u_sig142 (.PAD(sig142), .Y(core_sig142));
  PADCELL_SIG_V u_sig143 (.PAD(sig143), .A(core_sig143));
  PADCELL_SIG_V u_sig144 (.PAD(sig144), .Y(core_sig144));
  PADCELL_SIG_V u_sig145 (.PAD(sig145), .A(core_sig145));
  PADCELL_SIG_V u_sig146 (.PAD(sig146), .Y(core_sig146));
  PADCELL_SIG_V u_sig147 (.PAD(sig147), .A(core_sig147));
  PADCELL_SIG_V u_sig148 (.PAD(sig148), .Y(core_sig148));
  PADCELL_SIG_V u_sig149 (.PAD(sig149), .A(core_sig149));
  PADCELL_SIG_V u_sig150 (.PAD(sig150), .Y(core_sig150));
  PADCELL_SIG_V u_sig151 (.PAD(sig151), .A(core_sig151));
  PADCELL_SIG_V u_sig152 (.PAD(sig152), .Y(core_sig152));
  PADCELL_SIG_V u_sig153 (.PAD(sig153), .A(core_sig153));
  PADCELL_SIG_V u_sig154 (.PAD(sig154), .Y(core_sig154));
  PADCELL_SIG_V u_sig155 (.PAD(sig155), .A(core_sig155));
  PADCELL_SIG_V u_sig156 (.PAD(sig156), .Y(core_sig156));
  PADCELL_SIG_V u_sig157 (.PAD(sig157), .A(core_sig157));
  PADCELL_SIG_V u_sig158 (.PAD(sig158), .Y(core_sig158));
  PADCELL_SIG_V u_sig159 (.PAD(sig159), .A(core_sig159));
  PADCELL_SIG_V u_sig160 (.PAD(sig160), .Y(core_sig160));
  PADCELL_SIG_V u_sig161 (.PAD(sig161), .A(core_sig161));
  PADCELL_SIG_V u_sig162 (.PAD(sig162), .Y(core_sig162));
  PADCELL_SIG_V u_sig163 (.PAD(sig163), .A(core_sig163));
  PADCELL_SIG_V u_sig164 (.PAD(sig164), .Y(core_sig164));
  PADCELL_SIG_V u_sig165 (.PAD(sig165), .A(core_sig165));
  PADCELL_SIG_V u_sig166 (.PAD(sig166), .Y(core_sig166));
  PADCELL_SIG_V u_sig167 (.PAD(sig167), .A(core_sig167));
  PADCELL_SIG_V u_sig168 (.PAD(sig168), .Y(core_sig168));
  PADCELL_SIG_V u_sig169 (.PAD(sig169), .A(core_sig169));
  PADCELL_SIG_V u_sig170 (.PAD(sig170), .Y(core_sig170));
  PADCELL_SIG_V u_sig171 (.PAD(sig171), .A(core_sig171));
  PADCELL_SIG_V u_sig172 (.PAD(sig172), .Y(core_sig172));
  PADCELL_SIG_V u_sig173 (.PAD(sig173), .A(core_sig173));
  PADCELL_SIG_V u_sig174 (.PAD(sig174), .Y(core_sig174));
  PADCELL_SIG_V u_sig175 (.PAD(sig175), .A(core_sig175));
  PADCELL_SIG_V u_sig176 (.PAD(sig176), .Y(core_sig176));
  PADCELL_SIG_V u_sig177 (.PAD(sig177), .A(core_sig177));
  PADCELL_SIG_V u_sig178 (.PAD(sig178), .Y(core_sig178));
  PADCELL_SIG_V u_sig179 (.PAD(sig179), .A(core_sig179));
  PADCELL_SIG_V u_sig180 (.PAD(sig180), .Y(core_sig180));
  PADCELL_SIG_V u_sig181 (.PAD(sig181), .A(core_sig181));
  PADCELL_SIG_V u_sig182 (.PAD(sig182), .Y(core_sig182));
  PADCELL_SIG_V u_sig183 (.PAD(sig183), .A(core_sig183));
  PADCELL_SIG_V u_sig184 (.PAD(sig184), .Y(core_sig184));
  PADCELL_SIG_V u_sig185 (.PAD(sig185), .A(core_sig185));
  PADCELL_SIG_V u_sig186 (.PAD(sig186), .Y(core_sig186));
  PADCELL_SIG_V u_sig187 (.PAD(sig187), .A(core_sig187));
  PADCELL_SIG_V u_sig188 (.PAD(sig188), .Y(core_sig188));
  PADCELL_SIG_V u_sig189 (.PAD(sig189), .A(core_sig189));
  PADCELL_SIG_H u_sig190 (.PAD(sig190), .Y(core_sig190));
  PADCELL_SIG_H u_sig191 (.PAD(sig191), .A(core_sig191));
  PADCELL_SIG_H u_sig192 (.PAD(sig192), .Y(core_sig192));
  PADCELL_SIG_H u_sig193 (.PAD(sig193), .A(core_sig193));
  PADCELL_SIG_H u_sig194 (.PAD(sig194), .Y(core_sig194));
  PADCELL_SIG_H u_sig195 (.PAD(sig195), .A(core_sig195));
  PADCELL_SIG_H u_sig196 (.PAD(sig196), .Y(core_sig196));
  PADCELL_SIG_H u_sig197 (.PAD(sig197), .A(core_sig197));
  PADCELL_SIG_H u_sig198 (.PAD(sig198), .Y(core_sig198));
  PADCELL_SIG_H u_sig199 (.PAD(sig199), .A(core_sig199));
  PADCELL_SIG_H u_sig200 (.PAD(sig200), .Y(core_sig200));
  PADCELL_SIG_H u_sig201 (.PAD(sig201), .A(core_sig201));
  PADCELL_SIG_H u_sig202 (.PAD(sig202), .Y(core_sig202));
  PADCELL_SIG_H u_sig203 (.PAD(sig203), .A(core_sig203));
  PADCELL_SIG_H u_sig204 (.PAD(sig204), .Y(core_sig204));
  PADCELL_SIG_H u_sig205 (.PAD(sig205), .A(core_sig205));
  PADCELL_SIG_H u_sig206 (.PAD(sig206), .Y(core_sig206));
  PADCELL_SIG_H u_sig207 (.PAD(sig207), .A(core_sig207));
  PADCELL_SIG_H u_sig208 (.PAD(sig208), .Y(core_sig208));
  PADCELL_SIG_H u_sig209 (.PAD(sig209), .A(core_sig209));
  PADCELL_SIG_H u_sig210 (.PAD(sig210), .Y(core_sig210));
  PADCELL_SIG_H u_sig211 (.PAD(sig211), .A(core_sig211));
  PADCELL_SIG_H u_sig212 (.PAD(sig212), .Y(core_sig212));
  PADCELL_SIG_H u_sig213 (.PAD(sig213), .A(core_sig213));
  PADCELL_SIG_H u_sig214 (.PAD(sig214), .Y(core_sig214));
  PADCELL_SIG_H u_sig215 (.PAD(sig215), .A(core_sig215));
  PADCELL_SIG_H u_sig216 (.PAD(sig216), .Y(core_sig216));
  PADCELL_SIG_H u_sig217 (.PAD(sig217), .A(core_sig217));
  PADCELL_SIG_H u_sig218 (.PAD(sig218), .Y(core_sig218));
  PADCELL_SIG_H u_sig219 (.PAD(sig219), .A(core_sig219));
  PADCELL_SIG_H u_sig220 (.PAD(sig220), .Y(core_sig220));
  PADCELL_SIG_H u_sig221 (.PAD(sig221), .A(core_sig221));
  PADCELL_SIG_H u_sig222 (.PAD(sig222), .Y(core_sig222));
  PADCELL_SIG_H u_sig223 (.PAD(sig223), .A(core_sig223));
  PADCELL_SIG_H u_sig224 (.PAD(sig224), .Y(core_sig224));
  PADCELL_SIG_H u_sig225 (.PAD(sig225), .A(core_sig225));
  PADCELL_SIG_H u_sig226 (.PAD(sig226), .Y(core_sig226));
  PADCELL_SIG_H u_sig227 (.PAD(sig227), .A(core_sig227));
  PADCELL_SIG_H u_sig228 (.PAD(sig228), .Y(core_sig228));
  PADCELL_SIG_H u_sig229 (.PAD(sig229), .A(core_sig229));
  PADCELL_SIG_H u_sig230 (.PAD(sig230), .Y(core_sig230));
  PADCELL_SIG_H u_sig231 (.PAD(sig231), .A(core_sig231));
  PADCELL_SIG_H u_sig232 (.PAD(sig232), .Y(core_sig232));
  PADCELL_SIG_H u_sig233 (.PAD(sig233), .A(core_sig233));
  PADCELL_SIG_H u_sig234 (.PAD(sig234), .Y(core_sig234));
  PADCELL_SIG_H u_sig235 (.PAD(sig235), .A(core_sig235));
  PADCELL_SIG_H u_sig236 (.PAD(sig236), .Y(core_sig236));
  PADCELL_SIG_H u_sig237 (.PAD(sig237), .A(core_sig237));
  PADCELL_SIG_H u_sig238 (.PAD(sig238), .Y(core_sig238));
  PADCELL_SIG_H u_sig239 (.PAD(sig239), .A(core_sig239));
  PADCELL_SIG_H u_sig240 (.PAD(sig240), .Y(core_sig240));
  PADCELL_SIG_H u_sig241 (.PAD(sig241), .A(core_sig241));
  PADCELL_SIG_H u_sig242 (.PAD(sig242), .Y(core_sig242));
  PADCELL_SIG_H u_sig243 (.PAD(sig243), .A(core_sig243));
  PADCELL_SIG_H u_sig244 (.PAD(sig244), .Y(core_sig244));
  PADCELL_SIG_H u_sig245 (.PAD(sig245), .A(core_sig245));
  PADCELL_SIG_H u_sig246 (.PAD(sig246), .Y(core_sig246));
  PADCELL_SIG_H u_sig247 (.PAD(sig247), .A(core_sig247));
  PADCELL_SIG_H u_sig248 (.PAD(sig248), .Y(core_sig248));
  PADCELL_SIG_H u_sig249 (.PAD(sig249), .A(core_sig249));
  PADCELL_SIG_H u_sig250 (.PAD(sig250), .Y(core_sig250));
  PADCELL_SIG_H u_sig251 (.PAD(sig251), .A(core_sig251));
  PADCELL_SIG_H u_sig252 (.PAD(sig252), .Y(core_sig252));
endmodule
