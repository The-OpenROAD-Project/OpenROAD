# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_io__overlay_vccd_hvc
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 200 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 1.270000 56.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 53.125000 75.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 1.270000 51.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 48.365000 75.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.495000 8.890000 24.395000 13.530000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390000 8.890000 74.290000 13.530000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 8.885000 24.370000 13.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.415000 8.885000 75.000000 13.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 8.985000 1.270000 13.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 8.985000 75.000000 13.435000 ;
    END
    PORT
      LAYER via3 ;
        RECT  0.585000  8.960000  0.785000  9.160000 ;
        RECT  0.585000  9.390000  0.785000  9.590000 ;
        RECT  0.585000  9.820000  0.785000 10.020000 ;
        RECT  0.585000 10.250000  0.785000 10.450000 ;
        RECT  0.585000 10.680000  0.785000 10.880000 ;
        RECT  0.585000 11.110000  0.785000 11.310000 ;
        RECT  0.585000 11.540000  0.785000 11.740000 ;
        RECT  0.585000 11.970000  0.785000 12.170000 ;
        RECT  0.585000 12.400000  0.785000 12.600000 ;
        RECT  0.585000 12.830000  0.785000 13.030000 ;
        RECT  0.585000 13.260000  0.785000 13.460000 ;
        RECT  0.995000  8.960000  1.195000  9.160000 ;
        RECT  0.995000  9.390000  1.195000  9.590000 ;
        RECT  0.995000  9.820000  1.195000 10.020000 ;
        RECT  0.995000 10.250000  1.195000 10.450000 ;
        RECT  0.995000 10.680000  1.195000 10.880000 ;
        RECT  0.995000 11.110000  1.195000 11.310000 ;
        RECT  0.995000 11.540000  1.195000 11.740000 ;
        RECT  0.995000 11.970000  1.195000 12.170000 ;
        RECT  0.995000 12.400000  1.195000 12.600000 ;
        RECT  0.995000 12.830000  1.195000 13.030000 ;
        RECT  0.995000 13.260000  1.195000 13.460000 ;
        RECT  1.405000  8.960000  1.605000  9.160000 ;
        RECT  1.405000  9.390000  1.605000  9.590000 ;
        RECT  1.405000  9.820000  1.605000 10.020000 ;
        RECT  1.405000 10.250000  1.605000 10.450000 ;
        RECT  1.405000 10.680000  1.605000 10.880000 ;
        RECT  1.405000 11.110000  1.605000 11.310000 ;
        RECT  1.405000 11.540000  1.605000 11.740000 ;
        RECT  1.405000 11.970000  1.605000 12.170000 ;
        RECT  1.405000 12.400000  1.605000 12.600000 ;
        RECT  1.405000 12.830000  1.605000 13.030000 ;
        RECT  1.405000 13.260000  1.605000 13.460000 ;
        RECT  1.815000  8.960000  2.015000  9.160000 ;
        RECT  1.815000  9.390000  2.015000  9.590000 ;
        RECT  1.815000  9.820000  2.015000 10.020000 ;
        RECT  1.815000 10.250000  2.015000 10.450000 ;
        RECT  1.815000 10.680000  2.015000 10.880000 ;
        RECT  1.815000 11.110000  2.015000 11.310000 ;
        RECT  1.815000 11.540000  2.015000 11.740000 ;
        RECT  1.815000 11.970000  2.015000 12.170000 ;
        RECT  1.815000 12.400000  2.015000 12.600000 ;
        RECT  1.815000 12.830000  2.015000 13.030000 ;
        RECT  1.815000 13.260000  2.015000 13.460000 ;
        RECT  2.225000  8.960000  2.425000  9.160000 ;
        RECT  2.225000  9.390000  2.425000  9.590000 ;
        RECT  2.225000  9.820000  2.425000 10.020000 ;
        RECT  2.225000 10.250000  2.425000 10.450000 ;
        RECT  2.225000 10.680000  2.425000 10.880000 ;
        RECT  2.225000 11.110000  2.425000 11.310000 ;
        RECT  2.225000 11.540000  2.425000 11.740000 ;
        RECT  2.225000 11.970000  2.425000 12.170000 ;
        RECT  2.225000 12.400000  2.425000 12.600000 ;
        RECT  2.225000 12.830000  2.425000 13.030000 ;
        RECT  2.225000 13.260000  2.425000 13.460000 ;
        RECT  2.635000  8.960000  2.835000  9.160000 ;
        RECT  2.635000  9.390000  2.835000  9.590000 ;
        RECT  2.635000  9.820000  2.835000 10.020000 ;
        RECT  2.635000 10.250000  2.835000 10.450000 ;
        RECT  2.635000 10.680000  2.835000 10.880000 ;
        RECT  2.635000 11.110000  2.835000 11.310000 ;
        RECT  2.635000 11.540000  2.835000 11.740000 ;
        RECT  2.635000 11.970000  2.835000 12.170000 ;
        RECT  2.635000 12.400000  2.835000 12.600000 ;
        RECT  2.635000 12.830000  2.835000 13.030000 ;
        RECT  2.635000 13.260000  2.835000 13.460000 ;
        RECT  3.045000  8.960000  3.245000  9.160000 ;
        RECT  3.045000  9.390000  3.245000  9.590000 ;
        RECT  3.045000  9.820000  3.245000 10.020000 ;
        RECT  3.045000 10.250000  3.245000 10.450000 ;
        RECT  3.045000 10.680000  3.245000 10.880000 ;
        RECT  3.045000 11.110000  3.245000 11.310000 ;
        RECT  3.045000 11.540000  3.245000 11.740000 ;
        RECT  3.045000 11.970000  3.245000 12.170000 ;
        RECT  3.045000 12.400000  3.245000 12.600000 ;
        RECT  3.045000 12.830000  3.245000 13.030000 ;
        RECT  3.045000 13.260000  3.245000 13.460000 ;
        RECT  3.450000  8.960000  3.650000  9.160000 ;
        RECT  3.450000  9.390000  3.650000  9.590000 ;
        RECT  3.450000  9.820000  3.650000 10.020000 ;
        RECT  3.450000 10.250000  3.650000 10.450000 ;
        RECT  3.450000 10.680000  3.650000 10.880000 ;
        RECT  3.450000 11.110000  3.650000 11.310000 ;
        RECT  3.450000 11.540000  3.650000 11.740000 ;
        RECT  3.450000 11.970000  3.650000 12.170000 ;
        RECT  3.450000 12.400000  3.650000 12.600000 ;
        RECT  3.450000 12.830000  3.650000 13.030000 ;
        RECT  3.450000 13.260000  3.650000 13.460000 ;
        RECT  3.855000  8.960000  4.055000  9.160000 ;
        RECT  3.855000  9.390000  4.055000  9.590000 ;
        RECT  3.855000  9.820000  4.055000 10.020000 ;
        RECT  3.855000 10.250000  4.055000 10.450000 ;
        RECT  3.855000 10.680000  4.055000 10.880000 ;
        RECT  3.855000 11.110000  4.055000 11.310000 ;
        RECT  3.855000 11.540000  4.055000 11.740000 ;
        RECT  3.855000 11.970000  4.055000 12.170000 ;
        RECT  3.855000 12.400000  4.055000 12.600000 ;
        RECT  3.855000 12.830000  4.055000 13.030000 ;
        RECT  3.855000 13.260000  4.055000 13.460000 ;
        RECT  4.260000  8.960000  4.460000  9.160000 ;
        RECT  4.260000  9.390000  4.460000  9.590000 ;
        RECT  4.260000  9.820000  4.460000 10.020000 ;
        RECT  4.260000 10.250000  4.460000 10.450000 ;
        RECT  4.260000 10.680000  4.460000 10.880000 ;
        RECT  4.260000 11.110000  4.460000 11.310000 ;
        RECT  4.260000 11.540000  4.460000 11.740000 ;
        RECT  4.260000 11.970000  4.460000 12.170000 ;
        RECT  4.260000 12.400000  4.460000 12.600000 ;
        RECT  4.260000 12.830000  4.460000 13.030000 ;
        RECT  4.260000 13.260000  4.460000 13.460000 ;
        RECT  4.665000  8.960000  4.865000  9.160000 ;
        RECT  4.665000  9.390000  4.865000  9.590000 ;
        RECT  4.665000  9.820000  4.865000 10.020000 ;
        RECT  4.665000 10.250000  4.865000 10.450000 ;
        RECT  4.665000 10.680000  4.865000 10.880000 ;
        RECT  4.665000 11.110000  4.865000 11.310000 ;
        RECT  4.665000 11.540000  4.865000 11.740000 ;
        RECT  4.665000 11.970000  4.865000 12.170000 ;
        RECT  4.665000 12.400000  4.865000 12.600000 ;
        RECT  4.665000 12.830000  4.865000 13.030000 ;
        RECT  4.665000 13.260000  4.865000 13.460000 ;
        RECT  5.070000  8.960000  5.270000  9.160000 ;
        RECT  5.070000  9.390000  5.270000  9.590000 ;
        RECT  5.070000  9.820000  5.270000 10.020000 ;
        RECT  5.070000 10.250000  5.270000 10.450000 ;
        RECT  5.070000 10.680000  5.270000 10.880000 ;
        RECT  5.070000 11.110000  5.270000 11.310000 ;
        RECT  5.070000 11.540000  5.270000 11.740000 ;
        RECT  5.070000 11.970000  5.270000 12.170000 ;
        RECT  5.070000 12.400000  5.270000 12.600000 ;
        RECT  5.070000 12.830000  5.270000 13.030000 ;
        RECT  5.070000 13.260000  5.270000 13.460000 ;
        RECT  5.475000  8.960000  5.675000  9.160000 ;
        RECT  5.475000  9.390000  5.675000  9.590000 ;
        RECT  5.475000  9.820000  5.675000 10.020000 ;
        RECT  5.475000 10.250000  5.675000 10.450000 ;
        RECT  5.475000 10.680000  5.675000 10.880000 ;
        RECT  5.475000 11.110000  5.675000 11.310000 ;
        RECT  5.475000 11.540000  5.675000 11.740000 ;
        RECT  5.475000 11.970000  5.675000 12.170000 ;
        RECT  5.475000 12.400000  5.675000 12.600000 ;
        RECT  5.475000 12.830000  5.675000 13.030000 ;
        RECT  5.475000 13.260000  5.675000 13.460000 ;
        RECT  5.880000  8.960000  6.080000  9.160000 ;
        RECT  5.880000  9.390000  6.080000  9.590000 ;
        RECT  5.880000  9.820000  6.080000 10.020000 ;
        RECT  5.880000 10.250000  6.080000 10.450000 ;
        RECT  5.880000 10.680000  6.080000 10.880000 ;
        RECT  5.880000 11.110000  6.080000 11.310000 ;
        RECT  5.880000 11.540000  6.080000 11.740000 ;
        RECT  5.880000 11.970000  6.080000 12.170000 ;
        RECT  5.880000 12.400000  6.080000 12.600000 ;
        RECT  5.880000 12.830000  6.080000 13.030000 ;
        RECT  5.880000 13.260000  6.080000 13.460000 ;
        RECT  6.285000  8.960000  6.485000  9.160000 ;
        RECT  6.285000  9.390000  6.485000  9.590000 ;
        RECT  6.285000  9.820000  6.485000 10.020000 ;
        RECT  6.285000 10.250000  6.485000 10.450000 ;
        RECT  6.285000 10.680000  6.485000 10.880000 ;
        RECT  6.285000 11.110000  6.485000 11.310000 ;
        RECT  6.285000 11.540000  6.485000 11.740000 ;
        RECT  6.285000 11.970000  6.485000 12.170000 ;
        RECT  6.285000 12.400000  6.485000 12.600000 ;
        RECT  6.285000 12.830000  6.485000 13.030000 ;
        RECT  6.285000 13.260000  6.485000 13.460000 ;
        RECT  6.690000  8.960000  6.890000  9.160000 ;
        RECT  6.690000  9.390000  6.890000  9.590000 ;
        RECT  6.690000  9.820000  6.890000 10.020000 ;
        RECT  6.690000 10.250000  6.890000 10.450000 ;
        RECT  6.690000 10.680000  6.890000 10.880000 ;
        RECT  6.690000 11.110000  6.890000 11.310000 ;
        RECT  6.690000 11.540000  6.890000 11.740000 ;
        RECT  6.690000 11.970000  6.890000 12.170000 ;
        RECT  6.690000 12.400000  6.890000 12.600000 ;
        RECT  6.690000 12.830000  6.890000 13.030000 ;
        RECT  6.690000 13.260000  6.890000 13.460000 ;
        RECT  7.095000  8.960000  7.295000  9.160000 ;
        RECT  7.095000  9.390000  7.295000  9.590000 ;
        RECT  7.095000  9.820000  7.295000 10.020000 ;
        RECT  7.095000 10.250000  7.295000 10.450000 ;
        RECT  7.095000 10.680000  7.295000 10.880000 ;
        RECT  7.095000 11.110000  7.295000 11.310000 ;
        RECT  7.095000 11.540000  7.295000 11.740000 ;
        RECT  7.095000 11.970000  7.295000 12.170000 ;
        RECT  7.095000 12.400000  7.295000 12.600000 ;
        RECT  7.095000 12.830000  7.295000 13.030000 ;
        RECT  7.095000 13.260000  7.295000 13.460000 ;
        RECT  7.500000  8.960000  7.700000  9.160000 ;
        RECT  7.500000  9.390000  7.700000  9.590000 ;
        RECT  7.500000  9.820000  7.700000 10.020000 ;
        RECT  7.500000 10.250000  7.700000 10.450000 ;
        RECT  7.500000 10.680000  7.700000 10.880000 ;
        RECT  7.500000 11.110000  7.700000 11.310000 ;
        RECT  7.500000 11.540000  7.700000 11.740000 ;
        RECT  7.500000 11.970000  7.700000 12.170000 ;
        RECT  7.500000 12.400000  7.700000 12.600000 ;
        RECT  7.500000 12.830000  7.700000 13.030000 ;
        RECT  7.500000 13.260000  7.700000 13.460000 ;
        RECT  7.905000  8.960000  8.105000  9.160000 ;
        RECT  7.905000  9.390000  8.105000  9.590000 ;
        RECT  7.905000  9.820000  8.105000 10.020000 ;
        RECT  7.905000 10.250000  8.105000 10.450000 ;
        RECT  7.905000 10.680000  8.105000 10.880000 ;
        RECT  7.905000 11.110000  8.105000 11.310000 ;
        RECT  7.905000 11.540000  8.105000 11.740000 ;
        RECT  7.905000 11.970000  8.105000 12.170000 ;
        RECT  7.905000 12.400000  8.105000 12.600000 ;
        RECT  7.905000 12.830000  8.105000 13.030000 ;
        RECT  7.905000 13.260000  8.105000 13.460000 ;
        RECT  8.310000  8.960000  8.510000  9.160000 ;
        RECT  8.310000  9.390000  8.510000  9.590000 ;
        RECT  8.310000  9.820000  8.510000 10.020000 ;
        RECT  8.310000 10.250000  8.510000 10.450000 ;
        RECT  8.310000 10.680000  8.510000 10.880000 ;
        RECT  8.310000 11.110000  8.510000 11.310000 ;
        RECT  8.310000 11.540000  8.510000 11.740000 ;
        RECT  8.310000 11.970000  8.510000 12.170000 ;
        RECT  8.310000 12.400000  8.510000 12.600000 ;
        RECT  8.310000 12.830000  8.510000 13.030000 ;
        RECT  8.310000 13.260000  8.510000 13.460000 ;
        RECT  8.715000  8.960000  8.915000  9.160000 ;
        RECT  8.715000  9.390000  8.915000  9.590000 ;
        RECT  8.715000  9.820000  8.915000 10.020000 ;
        RECT  8.715000 10.250000  8.915000 10.450000 ;
        RECT  8.715000 10.680000  8.915000 10.880000 ;
        RECT  8.715000 11.110000  8.915000 11.310000 ;
        RECT  8.715000 11.540000  8.915000 11.740000 ;
        RECT  8.715000 11.970000  8.915000 12.170000 ;
        RECT  8.715000 12.400000  8.915000 12.600000 ;
        RECT  8.715000 12.830000  8.915000 13.030000 ;
        RECT  8.715000 13.260000  8.915000 13.460000 ;
        RECT  9.120000  8.960000  9.320000  9.160000 ;
        RECT  9.120000  9.390000  9.320000  9.590000 ;
        RECT  9.120000  9.820000  9.320000 10.020000 ;
        RECT  9.120000 10.250000  9.320000 10.450000 ;
        RECT  9.120000 10.680000  9.320000 10.880000 ;
        RECT  9.120000 11.110000  9.320000 11.310000 ;
        RECT  9.120000 11.540000  9.320000 11.740000 ;
        RECT  9.120000 11.970000  9.320000 12.170000 ;
        RECT  9.120000 12.400000  9.320000 12.600000 ;
        RECT  9.120000 12.830000  9.320000 13.030000 ;
        RECT  9.120000 13.260000  9.320000 13.460000 ;
        RECT  9.525000  8.960000  9.725000  9.160000 ;
        RECT  9.525000  9.390000  9.725000  9.590000 ;
        RECT  9.525000  9.820000  9.725000 10.020000 ;
        RECT  9.525000 10.250000  9.725000 10.450000 ;
        RECT  9.525000 10.680000  9.725000 10.880000 ;
        RECT  9.525000 11.110000  9.725000 11.310000 ;
        RECT  9.525000 11.540000  9.725000 11.740000 ;
        RECT  9.525000 11.970000  9.725000 12.170000 ;
        RECT  9.525000 12.400000  9.725000 12.600000 ;
        RECT  9.525000 12.830000  9.725000 13.030000 ;
        RECT  9.525000 13.260000  9.725000 13.460000 ;
        RECT  9.930000  8.960000 10.130000  9.160000 ;
        RECT  9.930000  9.390000 10.130000  9.590000 ;
        RECT  9.930000  9.820000 10.130000 10.020000 ;
        RECT  9.930000 10.250000 10.130000 10.450000 ;
        RECT  9.930000 10.680000 10.130000 10.880000 ;
        RECT  9.930000 11.110000 10.130000 11.310000 ;
        RECT  9.930000 11.540000 10.130000 11.740000 ;
        RECT  9.930000 11.970000 10.130000 12.170000 ;
        RECT  9.930000 12.400000 10.130000 12.600000 ;
        RECT  9.930000 12.830000 10.130000 13.030000 ;
        RECT  9.930000 13.260000 10.130000 13.460000 ;
        RECT 10.335000  8.960000 10.535000  9.160000 ;
        RECT 10.335000  9.390000 10.535000  9.590000 ;
        RECT 10.335000  9.820000 10.535000 10.020000 ;
        RECT 10.335000 10.250000 10.535000 10.450000 ;
        RECT 10.335000 10.680000 10.535000 10.880000 ;
        RECT 10.335000 11.110000 10.535000 11.310000 ;
        RECT 10.335000 11.540000 10.535000 11.740000 ;
        RECT 10.335000 11.970000 10.535000 12.170000 ;
        RECT 10.335000 12.400000 10.535000 12.600000 ;
        RECT 10.335000 12.830000 10.535000 13.030000 ;
        RECT 10.335000 13.260000 10.535000 13.460000 ;
        RECT 10.740000  8.960000 10.940000  9.160000 ;
        RECT 10.740000  9.390000 10.940000  9.590000 ;
        RECT 10.740000  9.820000 10.940000 10.020000 ;
        RECT 10.740000 10.250000 10.940000 10.450000 ;
        RECT 10.740000 10.680000 10.940000 10.880000 ;
        RECT 10.740000 11.110000 10.940000 11.310000 ;
        RECT 10.740000 11.540000 10.940000 11.740000 ;
        RECT 10.740000 11.970000 10.940000 12.170000 ;
        RECT 10.740000 12.400000 10.940000 12.600000 ;
        RECT 10.740000 12.830000 10.940000 13.030000 ;
        RECT 10.740000 13.260000 10.940000 13.460000 ;
        RECT 11.145000  8.960000 11.345000  9.160000 ;
        RECT 11.145000  9.390000 11.345000  9.590000 ;
        RECT 11.145000  9.820000 11.345000 10.020000 ;
        RECT 11.145000 10.250000 11.345000 10.450000 ;
        RECT 11.145000 10.680000 11.345000 10.880000 ;
        RECT 11.145000 11.110000 11.345000 11.310000 ;
        RECT 11.145000 11.540000 11.345000 11.740000 ;
        RECT 11.145000 11.970000 11.345000 12.170000 ;
        RECT 11.145000 12.400000 11.345000 12.600000 ;
        RECT 11.145000 12.830000 11.345000 13.030000 ;
        RECT 11.145000 13.260000 11.345000 13.460000 ;
        RECT 11.550000  8.960000 11.750000  9.160000 ;
        RECT 11.550000  9.390000 11.750000  9.590000 ;
        RECT 11.550000  9.820000 11.750000 10.020000 ;
        RECT 11.550000 10.250000 11.750000 10.450000 ;
        RECT 11.550000 10.680000 11.750000 10.880000 ;
        RECT 11.550000 11.110000 11.750000 11.310000 ;
        RECT 11.550000 11.540000 11.750000 11.740000 ;
        RECT 11.550000 11.970000 11.750000 12.170000 ;
        RECT 11.550000 12.400000 11.750000 12.600000 ;
        RECT 11.550000 12.830000 11.750000 13.030000 ;
        RECT 11.550000 13.260000 11.750000 13.460000 ;
        RECT 11.955000  8.960000 12.155000  9.160000 ;
        RECT 11.955000  9.390000 12.155000  9.590000 ;
        RECT 11.955000  9.820000 12.155000 10.020000 ;
        RECT 11.955000 10.250000 12.155000 10.450000 ;
        RECT 11.955000 10.680000 12.155000 10.880000 ;
        RECT 11.955000 11.110000 12.155000 11.310000 ;
        RECT 11.955000 11.540000 12.155000 11.740000 ;
        RECT 11.955000 11.970000 12.155000 12.170000 ;
        RECT 11.955000 12.400000 12.155000 12.600000 ;
        RECT 11.955000 12.830000 12.155000 13.030000 ;
        RECT 11.955000 13.260000 12.155000 13.460000 ;
        RECT 12.360000  8.960000 12.560000  9.160000 ;
        RECT 12.360000  9.390000 12.560000  9.590000 ;
        RECT 12.360000  9.820000 12.560000 10.020000 ;
        RECT 12.360000 10.250000 12.560000 10.450000 ;
        RECT 12.360000 10.680000 12.560000 10.880000 ;
        RECT 12.360000 11.110000 12.560000 11.310000 ;
        RECT 12.360000 11.540000 12.560000 11.740000 ;
        RECT 12.360000 11.970000 12.560000 12.170000 ;
        RECT 12.360000 12.400000 12.560000 12.600000 ;
        RECT 12.360000 12.830000 12.560000 13.030000 ;
        RECT 12.360000 13.260000 12.560000 13.460000 ;
        RECT 12.765000  8.960000 12.965000  9.160000 ;
        RECT 12.765000  9.390000 12.965000  9.590000 ;
        RECT 12.765000  9.820000 12.965000 10.020000 ;
        RECT 12.765000 10.250000 12.965000 10.450000 ;
        RECT 12.765000 10.680000 12.965000 10.880000 ;
        RECT 12.765000 11.110000 12.965000 11.310000 ;
        RECT 12.765000 11.540000 12.965000 11.740000 ;
        RECT 12.765000 11.970000 12.965000 12.170000 ;
        RECT 12.765000 12.400000 12.965000 12.600000 ;
        RECT 12.765000 12.830000 12.965000 13.030000 ;
        RECT 12.765000 13.260000 12.965000 13.460000 ;
        RECT 13.170000  8.960000 13.370000  9.160000 ;
        RECT 13.170000  9.390000 13.370000  9.590000 ;
        RECT 13.170000  9.820000 13.370000 10.020000 ;
        RECT 13.170000 10.250000 13.370000 10.450000 ;
        RECT 13.170000 10.680000 13.370000 10.880000 ;
        RECT 13.170000 11.110000 13.370000 11.310000 ;
        RECT 13.170000 11.540000 13.370000 11.740000 ;
        RECT 13.170000 11.970000 13.370000 12.170000 ;
        RECT 13.170000 12.400000 13.370000 12.600000 ;
        RECT 13.170000 12.830000 13.370000 13.030000 ;
        RECT 13.170000 13.260000 13.370000 13.460000 ;
        RECT 13.575000  8.960000 13.775000  9.160000 ;
        RECT 13.575000  9.390000 13.775000  9.590000 ;
        RECT 13.575000  9.820000 13.775000 10.020000 ;
        RECT 13.575000 10.250000 13.775000 10.450000 ;
        RECT 13.575000 10.680000 13.775000 10.880000 ;
        RECT 13.575000 11.110000 13.775000 11.310000 ;
        RECT 13.575000 11.540000 13.775000 11.740000 ;
        RECT 13.575000 11.970000 13.775000 12.170000 ;
        RECT 13.575000 12.400000 13.775000 12.600000 ;
        RECT 13.575000 12.830000 13.775000 13.030000 ;
        RECT 13.575000 13.260000 13.775000 13.460000 ;
        RECT 13.980000  8.960000 14.180000  9.160000 ;
        RECT 13.980000  9.390000 14.180000  9.590000 ;
        RECT 13.980000  9.820000 14.180000 10.020000 ;
        RECT 13.980000 10.250000 14.180000 10.450000 ;
        RECT 13.980000 10.680000 14.180000 10.880000 ;
        RECT 13.980000 11.110000 14.180000 11.310000 ;
        RECT 13.980000 11.540000 14.180000 11.740000 ;
        RECT 13.980000 11.970000 14.180000 12.170000 ;
        RECT 13.980000 12.400000 14.180000 12.600000 ;
        RECT 13.980000 12.830000 14.180000 13.030000 ;
        RECT 13.980000 13.260000 14.180000 13.460000 ;
        RECT 14.385000  8.960000 14.585000  9.160000 ;
        RECT 14.385000  9.390000 14.585000  9.590000 ;
        RECT 14.385000  9.820000 14.585000 10.020000 ;
        RECT 14.385000 10.250000 14.585000 10.450000 ;
        RECT 14.385000 10.680000 14.585000 10.880000 ;
        RECT 14.385000 11.110000 14.585000 11.310000 ;
        RECT 14.385000 11.540000 14.585000 11.740000 ;
        RECT 14.385000 11.970000 14.585000 12.170000 ;
        RECT 14.385000 12.400000 14.585000 12.600000 ;
        RECT 14.385000 12.830000 14.585000 13.030000 ;
        RECT 14.385000 13.260000 14.585000 13.460000 ;
        RECT 14.790000  8.960000 14.990000  9.160000 ;
        RECT 14.790000  9.390000 14.990000  9.590000 ;
        RECT 14.790000  9.820000 14.990000 10.020000 ;
        RECT 14.790000 10.250000 14.990000 10.450000 ;
        RECT 14.790000 10.680000 14.990000 10.880000 ;
        RECT 14.790000 11.110000 14.990000 11.310000 ;
        RECT 14.790000 11.540000 14.990000 11.740000 ;
        RECT 14.790000 11.970000 14.990000 12.170000 ;
        RECT 14.790000 12.400000 14.990000 12.600000 ;
        RECT 14.790000 12.830000 14.990000 13.030000 ;
        RECT 14.790000 13.260000 14.990000 13.460000 ;
        RECT 15.195000  8.960000 15.395000  9.160000 ;
        RECT 15.195000  9.390000 15.395000  9.590000 ;
        RECT 15.195000  9.820000 15.395000 10.020000 ;
        RECT 15.195000 10.250000 15.395000 10.450000 ;
        RECT 15.195000 10.680000 15.395000 10.880000 ;
        RECT 15.195000 11.110000 15.395000 11.310000 ;
        RECT 15.195000 11.540000 15.395000 11.740000 ;
        RECT 15.195000 11.970000 15.395000 12.170000 ;
        RECT 15.195000 12.400000 15.395000 12.600000 ;
        RECT 15.195000 12.830000 15.395000 13.030000 ;
        RECT 15.195000 13.260000 15.395000 13.460000 ;
        RECT 15.600000  8.960000 15.800000  9.160000 ;
        RECT 15.600000  9.390000 15.800000  9.590000 ;
        RECT 15.600000  9.820000 15.800000 10.020000 ;
        RECT 15.600000 10.250000 15.800000 10.450000 ;
        RECT 15.600000 10.680000 15.800000 10.880000 ;
        RECT 15.600000 11.110000 15.800000 11.310000 ;
        RECT 15.600000 11.540000 15.800000 11.740000 ;
        RECT 15.600000 11.970000 15.800000 12.170000 ;
        RECT 15.600000 12.400000 15.800000 12.600000 ;
        RECT 15.600000 12.830000 15.800000 13.030000 ;
        RECT 15.600000 13.260000 15.800000 13.460000 ;
        RECT 16.005000  8.960000 16.205000  9.160000 ;
        RECT 16.005000  9.390000 16.205000  9.590000 ;
        RECT 16.005000  9.820000 16.205000 10.020000 ;
        RECT 16.005000 10.250000 16.205000 10.450000 ;
        RECT 16.005000 10.680000 16.205000 10.880000 ;
        RECT 16.005000 11.110000 16.205000 11.310000 ;
        RECT 16.005000 11.540000 16.205000 11.740000 ;
        RECT 16.005000 11.970000 16.205000 12.170000 ;
        RECT 16.005000 12.400000 16.205000 12.600000 ;
        RECT 16.005000 12.830000 16.205000 13.030000 ;
        RECT 16.005000 13.260000 16.205000 13.460000 ;
        RECT 16.410000  8.960000 16.610000  9.160000 ;
        RECT 16.410000  9.390000 16.610000  9.590000 ;
        RECT 16.410000  9.820000 16.610000 10.020000 ;
        RECT 16.410000 10.250000 16.610000 10.450000 ;
        RECT 16.410000 10.680000 16.610000 10.880000 ;
        RECT 16.410000 11.110000 16.610000 11.310000 ;
        RECT 16.410000 11.540000 16.610000 11.740000 ;
        RECT 16.410000 11.970000 16.610000 12.170000 ;
        RECT 16.410000 12.400000 16.610000 12.600000 ;
        RECT 16.410000 12.830000 16.610000 13.030000 ;
        RECT 16.410000 13.260000 16.610000 13.460000 ;
        RECT 16.815000  8.960000 17.015000  9.160000 ;
        RECT 16.815000  9.390000 17.015000  9.590000 ;
        RECT 16.815000  9.820000 17.015000 10.020000 ;
        RECT 16.815000 10.250000 17.015000 10.450000 ;
        RECT 16.815000 10.680000 17.015000 10.880000 ;
        RECT 16.815000 11.110000 17.015000 11.310000 ;
        RECT 16.815000 11.540000 17.015000 11.740000 ;
        RECT 16.815000 11.970000 17.015000 12.170000 ;
        RECT 16.815000 12.400000 17.015000 12.600000 ;
        RECT 16.815000 12.830000 17.015000 13.030000 ;
        RECT 16.815000 13.260000 17.015000 13.460000 ;
        RECT 17.220000  8.960000 17.420000  9.160000 ;
        RECT 17.220000  9.390000 17.420000  9.590000 ;
        RECT 17.220000  9.820000 17.420000 10.020000 ;
        RECT 17.220000 10.250000 17.420000 10.450000 ;
        RECT 17.220000 10.680000 17.420000 10.880000 ;
        RECT 17.220000 11.110000 17.420000 11.310000 ;
        RECT 17.220000 11.540000 17.420000 11.740000 ;
        RECT 17.220000 11.970000 17.420000 12.170000 ;
        RECT 17.220000 12.400000 17.420000 12.600000 ;
        RECT 17.220000 12.830000 17.420000 13.030000 ;
        RECT 17.220000 13.260000 17.420000 13.460000 ;
        RECT 17.625000  8.960000 17.825000  9.160000 ;
        RECT 17.625000  9.390000 17.825000  9.590000 ;
        RECT 17.625000  9.820000 17.825000 10.020000 ;
        RECT 17.625000 10.250000 17.825000 10.450000 ;
        RECT 17.625000 10.680000 17.825000 10.880000 ;
        RECT 17.625000 11.110000 17.825000 11.310000 ;
        RECT 17.625000 11.540000 17.825000 11.740000 ;
        RECT 17.625000 11.970000 17.825000 12.170000 ;
        RECT 17.625000 12.400000 17.825000 12.600000 ;
        RECT 17.625000 12.830000 17.825000 13.030000 ;
        RECT 17.625000 13.260000 17.825000 13.460000 ;
        RECT 18.030000  8.960000 18.230000  9.160000 ;
        RECT 18.030000  9.390000 18.230000  9.590000 ;
        RECT 18.030000  9.820000 18.230000 10.020000 ;
        RECT 18.030000 10.250000 18.230000 10.450000 ;
        RECT 18.030000 10.680000 18.230000 10.880000 ;
        RECT 18.030000 11.110000 18.230000 11.310000 ;
        RECT 18.030000 11.540000 18.230000 11.740000 ;
        RECT 18.030000 11.970000 18.230000 12.170000 ;
        RECT 18.030000 12.400000 18.230000 12.600000 ;
        RECT 18.030000 12.830000 18.230000 13.030000 ;
        RECT 18.030000 13.260000 18.230000 13.460000 ;
        RECT 18.435000  8.960000 18.635000  9.160000 ;
        RECT 18.435000  9.390000 18.635000  9.590000 ;
        RECT 18.435000  9.820000 18.635000 10.020000 ;
        RECT 18.435000 10.250000 18.635000 10.450000 ;
        RECT 18.435000 10.680000 18.635000 10.880000 ;
        RECT 18.435000 11.110000 18.635000 11.310000 ;
        RECT 18.435000 11.540000 18.635000 11.740000 ;
        RECT 18.435000 11.970000 18.635000 12.170000 ;
        RECT 18.435000 12.400000 18.635000 12.600000 ;
        RECT 18.435000 12.830000 18.635000 13.030000 ;
        RECT 18.435000 13.260000 18.635000 13.460000 ;
        RECT 18.840000  8.960000 19.040000  9.160000 ;
        RECT 18.840000  9.390000 19.040000  9.590000 ;
        RECT 18.840000  9.820000 19.040000 10.020000 ;
        RECT 18.840000 10.250000 19.040000 10.450000 ;
        RECT 18.840000 10.680000 19.040000 10.880000 ;
        RECT 18.840000 11.110000 19.040000 11.310000 ;
        RECT 18.840000 11.540000 19.040000 11.740000 ;
        RECT 18.840000 11.970000 19.040000 12.170000 ;
        RECT 18.840000 12.400000 19.040000 12.600000 ;
        RECT 18.840000 12.830000 19.040000 13.030000 ;
        RECT 18.840000 13.260000 19.040000 13.460000 ;
        RECT 19.245000  8.960000 19.445000  9.160000 ;
        RECT 19.245000  9.390000 19.445000  9.590000 ;
        RECT 19.245000  9.820000 19.445000 10.020000 ;
        RECT 19.245000 10.250000 19.445000 10.450000 ;
        RECT 19.245000 10.680000 19.445000 10.880000 ;
        RECT 19.245000 11.110000 19.445000 11.310000 ;
        RECT 19.245000 11.540000 19.445000 11.740000 ;
        RECT 19.245000 11.970000 19.445000 12.170000 ;
        RECT 19.245000 12.400000 19.445000 12.600000 ;
        RECT 19.245000 12.830000 19.445000 13.030000 ;
        RECT 19.245000 13.260000 19.445000 13.460000 ;
        RECT 19.650000  8.960000 19.850000  9.160000 ;
        RECT 19.650000  9.390000 19.850000  9.590000 ;
        RECT 19.650000  9.820000 19.850000 10.020000 ;
        RECT 19.650000 10.250000 19.850000 10.450000 ;
        RECT 19.650000 10.680000 19.850000 10.880000 ;
        RECT 19.650000 11.110000 19.850000 11.310000 ;
        RECT 19.650000 11.540000 19.850000 11.740000 ;
        RECT 19.650000 11.970000 19.850000 12.170000 ;
        RECT 19.650000 12.400000 19.850000 12.600000 ;
        RECT 19.650000 12.830000 19.850000 13.030000 ;
        RECT 19.650000 13.260000 19.850000 13.460000 ;
        RECT 20.055000  8.960000 20.255000  9.160000 ;
        RECT 20.055000  9.390000 20.255000  9.590000 ;
        RECT 20.055000  9.820000 20.255000 10.020000 ;
        RECT 20.055000 10.250000 20.255000 10.450000 ;
        RECT 20.055000 10.680000 20.255000 10.880000 ;
        RECT 20.055000 11.110000 20.255000 11.310000 ;
        RECT 20.055000 11.540000 20.255000 11.740000 ;
        RECT 20.055000 11.970000 20.255000 12.170000 ;
        RECT 20.055000 12.400000 20.255000 12.600000 ;
        RECT 20.055000 12.830000 20.255000 13.030000 ;
        RECT 20.055000 13.260000 20.255000 13.460000 ;
        RECT 20.460000  8.960000 20.660000  9.160000 ;
        RECT 20.460000  9.390000 20.660000  9.590000 ;
        RECT 20.460000  9.820000 20.660000 10.020000 ;
        RECT 20.460000 10.250000 20.660000 10.450000 ;
        RECT 20.460000 10.680000 20.660000 10.880000 ;
        RECT 20.460000 11.110000 20.660000 11.310000 ;
        RECT 20.460000 11.540000 20.660000 11.740000 ;
        RECT 20.460000 11.970000 20.660000 12.170000 ;
        RECT 20.460000 12.400000 20.660000 12.600000 ;
        RECT 20.460000 12.830000 20.660000 13.030000 ;
        RECT 20.460000 13.260000 20.660000 13.460000 ;
        RECT 20.865000  8.960000 21.065000  9.160000 ;
        RECT 20.865000  9.390000 21.065000  9.590000 ;
        RECT 20.865000  9.820000 21.065000 10.020000 ;
        RECT 20.865000 10.250000 21.065000 10.450000 ;
        RECT 20.865000 10.680000 21.065000 10.880000 ;
        RECT 20.865000 11.110000 21.065000 11.310000 ;
        RECT 20.865000 11.540000 21.065000 11.740000 ;
        RECT 20.865000 11.970000 21.065000 12.170000 ;
        RECT 20.865000 12.400000 21.065000 12.600000 ;
        RECT 20.865000 12.830000 21.065000 13.030000 ;
        RECT 20.865000 13.260000 21.065000 13.460000 ;
        RECT 21.270000  8.960000 21.470000  9.160000 ;
        RECT 21.270000  9.390000 21.470000  9.590000 ;
        RECT 21.270000  9.820000 21.470000 10.020000 ;
        RECT 21.270000 10.250000 21.470000 10.450000 ;
        RECT 21.270000 10.680000 21.470000 10.880000 ;
        RECT 21.270000 11.110000 21.470000 11.310000 ;
        RECT 21.270000 11.540000 21.470000 11.740000 ;
        RECT 21.270000 11.970000 21.470000 12.170000 ;
        RECT 21.270000 12.400000 21.470000 12.600000 ;
        RECT 21.270000 12.830000 21.470000 13.030000 ;
        RECT 21.270000 13.260000 21.470000 13.460000 ;
        RECT 21.675000  8.960000 21.875000  9.160000 ;
        RECT 21.675000  9.390000 21.875000  9.590000 ;
        RECT 21.675000  9.820000 21.875000 10.020000 ;
        RECT 21.675000 10.250000 21.875000 10.450000 ;
        RECT 21.675000 10.680000 21.875000 10.880000 ;
        RECT 21.675000 11.110000 21.875000 11.310000 ;
        RECT 21.675000 11.540000 21.875000 11.740000 ;
        RECT 21.675000 11.970000 21.875000 12.170000 ;
        RECT 21.675000 12.400000 21.875000 12.600000 ;
        RECT 21.675000 12.830000 21.875000 13.030000 ;
        RECT 21.675000 13.260000 21.875000 13.460000 ;
        RECT 22.080000  8.960000 22.280000  9.160000 ;
        RECT 22.080000  9.390000 22.280000  9.590000 ;
        RECT 22.080000  9.820000 22.280000 10.020000 ;
        RECT 22.080000 10.250000 22.280000 10.450000 ;
        RECT 22.080000 10.680000 22.280000 10.880000 ;
        RECT 22.080000 11.110000 22.280000 11.310000 ;
        RECT 22.080000 11.540000 22.280000 11.740000 ;
        RECT 22.080000 11.970000 22.280000 12.170000 ;
        RECT 22.080000 12.400000 22.280000 12.600000 ;
        RECT 22.080000 12.830000 22.280000 13.030000 ;
        RECT 22.080000 13.260000 22.280000 13.460000 ;
        RECT 22.485000  8.960000 22.685000  9.160000 ;
        RECT 22.485000  9.390000 22.685000  9.590000 ;
        RECT 22.485000  9.820000 22.685000 10.020000 ;
        RECT 22.485000 10.250000 22.685000 10.450000 ;
        RECT 22.485000 10.680000 22.685000 10.880000 ;
        RECT 22.485000 11.110000 22.685000 11.310000 ;
        RECT 22.485000 11.540000 22.685000 11.740000 ;
        RECT 22.485000 11.970000 22.685000 12.170000 ;
        RECT 22.485000 12.400000 22.685000 12.600000 ;
        RECT 22.485000 12.830000 22.685000 13.030000 ;
        RECT 22.485000 13.260000 22.685000 13.460000 ;
        RECT 22.890000  8.960000 23.090000  9.160000 ;
        RECT 22.890000  9.390000 23.090000  9.590000 ;
        RECT 22.890000  9.820000 23.090000 10.020000 ;
        RECT 22.890000 10.250000 23.090000 10.450000 ;
        RECT 22.890000 10.680000 23.090000 10.880000 ;
        RECT 22.890000 11.110000 23.090000 11.310000 ;
        RECT 22.890000 11.540000 23.090000 11.740000 ;
        RECT 22.890000 11.970000 23.090000 12.170000 ;
        RECT 22.890000 12.400000 23.090000 12.600000 ;
        RECT 22.890000 12.830000 23.090000 13.030000 ;
        RECT 22.890000 13.260000 23.090000 13.460000 ;
        RECT 23.295000  8.960000 23.495000  9.160000 ;
        RECT 23.295000  9.390000 23.495000  9.590000 ;
        RECT 23.295000  9.820000 23.495000 10.020000 ;
        RECT 23.295000 10.250000 23.495000 10.450000 ;
        RECT 23.295000 10.680000 23.495000 10.880000 ;
        RECT 23.295000 11.110000 23.495000 11.310000 ;
        RECT 23.295000 11.540000 23.495000 11.740000 ;
        RECT 23.295000 11.970000 23.495000 12.170000 ;
        RECT 23.295000 12.400000 23.495000 12.600000 ;
        RECT 23.295000 12.830000 23.495000 13.030000 ;
        RECT 23.295000 13.260000 23.495000 13.460000 ;
        RECT 23.700000  8.960000 23.900000  9.160000 ;
        RECT 23.700000  9.390000 23.900000  9.590000 ;
        RECT 23.700000  9.820000 23.900000 10.020000 ;
        RECT 23.700000 10.250000 23.900000 10.450000 ;
        RECT 23.700000 10.680000 23.900000 10.880000 ;
        RECT 23.700000 11.110000 23.900000 11.310000 ;
        RECT 23.700000 11.540000 23.900000 11.740000 ;
        RECT 23.700000 11.970000 23.900000 12.170000 ;
        RECT 23.700000 12.400000 23.900000 12.600000 ;
        RECT 23.700000 12.830000 23.900000 13.030000 ;
        RECT 23.700000 13.260000 23.900000 13.460000 ;
        RECT 24.105000  8.960000 24.305000  9.160000 ;
        RECT 24.105000  9.390000 24.305000  9.590000 ;
        RECT 24.105000  9.820000 24.305000 10.020000 ;
        RECT 24.105000 10.250000 24.305000 10.450000 ;
        RECT 24.105000 10.680000 24.305000 10.880000 ;
        RECT 24.105000 11.110000 24.305000 11.310000 ;
        RECT 24.105000 11.540000 24.305000 11.740000 ;
        RECT 24.105000 11.970000 24.305000 12.170000 ;
        RECT 24.105000 12.400000 24.305000 12.600000 ;
        RECT 24.105000 12.830000 24.305000 13.030000 ;
        RECT 24.105000 13.260000 24.305000 13.460000 ;
        RECT 50.480000  8.960000 50.680000  9.160000 ;
        RECT 50.480000  9.390000 50.680000  9.590000 ;
        RECT 50.480000  9.820000 50.680000 10.020000 ;
        RECT 50.480000 10.250000 50.680000 10.450000 ;
        RECT 50.480000 10.680000 50.680000 10.880000 ;
        RECT 50.480000 11.110000 50.680000 11.310000 ;
        RECT 50.480000 11.540000 50.680000 11.740000 ;
        RECT 50.480000 11.970000 50.680000 12.170000 ;
        RECT 50.480000 12.400000 50.680000 12.600000 ;
        RECT 50.480000 12.830000 50.680000 13.030000 ;
        RECT 50.480000 13.260000 50.680000 13.460000 ;
        RECT 50.890000  8.960000 51.090000  9.160000 ;
        RECT 50.890000  9.390000 51.090000  9.590000 ;
        RECT 50.890000  9.820000 51.090000 10.020000 ;
        RECT 50.890000 10.250000 51.090000 10.450000 ;
        RECT 50.890000 10.680000 51.090000 10.880000 ;
        RECT 50.890000 11.110000 51.090000 11.310000 ;
        RECT 50.890000 11.540000 51.090000 11.740000 ;
        RECT 50.890000 11.970000 51.090000 12.170000 ;
        RECT 50.890000 12.400000 51.090000 12.600000 ;
        RECT 50.890000 12.830000 51.090000 13.030000 ;
        RECT 50.890000 13.260000 51.090000 13.460000 ;
        RECT 51.300000  8.960000 51.500000  9.160000 ;
        RECT 51.300000  9.390000 51.500000  9.590000 ;
        RECT 51.300000  9.820000 51.500000 10.020000 ;
        RECT 51.300000 10.250000 51.500000 10.450000 ;
        RECT 51.300000 10.680000 51.500000 10.880000 ;
        RECT 51.300000 11.110000 51.500000 11.310000 ;
        RECT 51.300000 11.540000 51.500000 11.740000 ;
        RECT 51.300000 11.970000 51.500000 12.170000 ;
        RECT 51.300000 12.400000 51.500000 12.600000 ;
        RECT 51.300000 12.830000 51.500000 13.030000 ;
        RECT 51.300000 13.260000 51.500000 13.460000 ;
        RECT 51.710000  8.960000 51.910000  9.160000 ;
        RECT 51.710000  9.390000 51.910000  9.590000 ;
        RECT 51.710000  9.820000 51.910000 10.020000 ;
        RECT 51.710000 10.250000 51.910000 10.450000 ;
        RECT 51.710000 10.680000 51.910000 10.880000 ;
        RECT 51.710000 11.110000 51.910000 11.310000 ;
        RECT 51.710000 11.540000 51.910000 11.740000 ;
        RECT 51.710000 11.970000 51.910000 12.170000 ;
        RECT 51.710000 12.400000 51.910000 12.600000 ;
        RECT 51.710000 12.830000 51.910000 13.030000 ;
        RECT 51.710000 13.260000 51.910000 13.460000 ;
        RECT 52.120000  8.960000 52.320000  9.160000 ;
        RECT 52.120000  9.390000 52.320000  9.590000 ;
        RECT 52.120000  9.820000 52.320000 10.020000 ;
        RECT 52.120000 10.250000 52.320000 10.450000 ;
        RECT 52.120000 10.680000 52.320000 10.880000 ;
        RECT 52.120000 11.110000 52.320000 11.310000 ;
        RECT 52.120000 11.540000 52.320000 11.740000 ;
        RECT 52.120000 11.970000 52.320000 12.170000 ;
        RECT 52.120000 12.400000 52.320000 12.600000 ;
        RECT 52.120000 12.830000 52.320000 13.030000 ;
        RECT 52.120000 13.260000 52.320000 13.460000 ;
        RECT 52.530000  8.960000 52.730000  9.160000 ;
        RECT 52.530000  9.390000 52.730000  9.590000 ;
        RECT 52.530000  9.820000 52.730000 10.020000 ;
        RECT 52.530000 10.250000 52.730000 10.450000 ;
        RECT 52.530000 10.680000 52.730000 10.880000 ;
        RECT 52.530000 11.110000 52.730000 11.310000 ;
        RECT 52.530000 11.540000 52.730000 11.740000 ;
        RECT 52.530000 11.970000 52.730000 12.170000 ;
        RECT 52.530000 12.400000 52.730000 12.600000 ;
        RECT 52.530000 12.830000 52.730000 13.030000 ;
        RECT 52.530000 13.260000 52.730000 13.460000 ;
        RECT 52.940000  8.960000 53.140000  9.160000 ;
        RECT 52.940000  9.390000 53.140000  9.590000 ;
        RECT 52.940000  9.820000 53.140000 10.020000 ;
        RECT 52.940000 10.250000 53.140000 10.450000 ;
        RECT 52.940000 10.680000 53.140000 10.880000 ;
        RECT 52.940000 11.110000 53.140000 11.310000 ;
        RECT 52.940000 11.540000 53.140000 11.740000 ;
        RECT 52.940000 11.970000 53.140000 12.170000 ;
        RECT 52.940000 12.400000 53.140000 12.600000 ;
        RECT 52.940000 12.830000 53.140000 13.030000 ;
        RECT 52.940000 13.260000 53.140000 13.460000 ;
        RECT 53.345000  8.960000 53.545000  9.160000 ;
        RECT 53.345000  9.390000 53.545000  9.590000 ;
        RECT 53.345000  9.820000 53.545000 10.020000 ;
        RECT 53.345000 10.250000 53.545000 10.450000 ;
        RECT 53.345000 10.680000 53.545000 10.880000 ;
        RECT 53.345000 11.110000 53.545000 11.310000 ;
        RECT 53.345000 11.540000 53.545000 11.740000 ;
        RECT 53.345000 11.970000 53.545000 12.170000 ;
        RECT 53.345000 12.400000 53.545000 12.600000 ;
        RECT 53.345000 12.830000 53.545000 13.030000 ;
        RECT 53.345000 13.260000 53.545000 13.460000 ;
        RECT 53.750000  8.960000 53.950000  9.160000 ;
        RECT 53.750000  9.390000 53.950000  9.590000 ;
        RECT 53.750000  9.820000 53.950000 10.020000 ;
        RECT 53.750000 10.250000 53.950000 10.450000 ;
        RECT 53.750000 10.680000 53.950000 10.880000 ;
        RECT 53.750000 11.110000 53.950000 11.310000 ;
        RECT 53.750000 11.540000 53.950000 11.740000 ;
        RECT 53.750000 11.970000 53.950000 12.170000 ;
        RECT 53.750000 12.400000 53.950000 12.600000 ;
        RECT 53.750000 12.830000 53.950000 13.030000 ;
        RECT 53.750000 13.260000 53.950000 13.460000 ;
        RECT 54.155000  8.960000 54.355000  9.160000 ;
        RECT 54.155000  9.390000 54.355000  9.590000 ;
        RECT 54.155000  9.820000 54.355000 10.020000 ;
        RECT 54.155000 10.250000 54.355000 10.450000 ;
        RECT 54.155000 10.680000 54.355000 10.880000 ;
        RECT 54.155000 11.110000 54.355000 11.310000 ;
        RECT 54.155000 11.540000 54.355000 11.740000 ;
        RECT 54.155000 11.970000 54.355000 12.170000 ;
        RECT 54.155000 12.400000 54.355000 12.600000 ;
        RECT 54.155000 12.830000 54.355000 13.030000 ;
        RECT 54.155000 13.260000 54.355000 13.460000 ;
        RECT 54.560000  8.960000 54.760000  9.160000 ;
        RECT 54.560000  9.390000 54.760000  9.590000 ;
        RECT 54.560000  9.820000 54.760000 10.020000 ;
        RECT 54.560000 10.250000 54.760000 10.450000 ;
        RECT 54.560000 10.680000 54.760000 10.880000 ;
        RECT 54.560000 11.110000 54.760000 11.310000 ;
        RECT 54.560000 11.540000 54.760000 11.740000 ;
        RECT 54.560000 11.970000 54.760000 12.170000 ;
        RECT 54.560000 12.400000 54.760000 12.600000 ;
        RECT 54.560000 12.830000 54.760000 13.030000 ;
        RECT 54.560000 13.260000 54.760000 13.460000 ;
        RECT 54.965000  8.960000 55.165000  9.160000 ;
        RECT 54.965000  9.390000 55.165000  9.590000 ;
        RECT 54.965000  9.820000 55.165000 10.020000 ;
        RECT 54.965000 10.250000 55.165000 10.450000 ;
        RECT 54.965000 10.680000 55.165000 10.880000 ;
        RECT 54.965000 11.110000 55.165000 11.310000 ;
        RECT 54.965000 11.540000 55.165000 11.740000 ;
        RECT 54.965000 11.970000 55.165000 12.170000 ;
        RECT 54.965000 12.400000 55.165000 12.600000 ;
        RECT 54.965000 12.830000 55.165000 13.030000 ;
        RECT 54.965000 13.260000 55.165000 13.460000 ;
        RECT 55.370000  8.960000 55.570000  9.160000 ;
        RECT 55.370000  9.390000 55.570000  9.590000 ;
        RECT 55.370000  9.820000 55.570000 10.020000 ;
        RECT 55.370000 10.250000 55.570000 10.450000 ;
        RECT 55.370000 10.680000 55.570000 10.880000 ;
        RECT 55.370000 11.110000 55.570000 11.310000 ;
        RECT 55.370000 11.540000 55.570000 11.740000 ;
        RECT 55.370000 11.970000 55.570000 12.170000 ;
        RECT 55.370000 12.400000 55.570000 12.600000 ;
        RECT 55.370000 12.830000 55.570000 13.030000 ;
        RECT 55.370000 13.260000 55.570000 13.460000 ;
        RECT 55.775000  8.960000 55.975000  9.160000 ;
        RECT 55.775000  9.390000 55.975000  9.590000 ;
        RECT 55.775000  9.820000 55.975000 10.020000 ;
        RECT 55.775000 10.250000 55.975000 10.450000 ;
        RECT 55.775000 10.680000 55.975000 10.880000 ;
        RECT 55.775000 11.110000 55.975000 11.310000 ;
        RECT 55.775000 11.540000 55.975000 11.740000 ;
        RECT 55.775000 11.970000 55.975000 12.170000 ;
        RECT 55.775000 12.400000 55.975000 12.600000 ;
        RECT 55.775000 12.830000 55.975000 13.030000 ;
        RECT 55.775000 13.260000 55.975000 13.460000 ;
        RECT 56.180000  8.960000 56.380000  9.160000 ;
        RECT 56.180000  9.390000 56.380000  9.590000 ;
        RECT 56.180000  9.820000 56.380000 10.020000 ;
        RECT 56.180000 10.250000 56.380000 10.450000 ;
        RECT 56.180000 10.680000 56.380000 10.880000 ;
        RECT 56.180000 11.110000 56.380000 11.310000 ;
        RECT 56.180000 11.540000 56.380000 11.740000 ;
        RECT 56.180000 11.970000 56.380000 12.170000 ;
        RECT 56.180000 12.400000 56.380000 12.600000 ;
        RECT 56.180000 12.830000 56.380000 13.030000 ;
        RECT 56.180000 13.260000 56.380000 13.460000 ;
        RECT 56.585000  8.960000 56.785000  9.160000 ;
        RECT 56.585000  9.390000 56.785000  9.590000 ;
        RECT 56.585000  9.820000 56.785000 10.020000 ;
        RECT 56.585000 10.250000 56.785000 10.450000 ;
        RECT 56.585000 10.680000 56.785000 10.880000 ;
        RECT 56.585000 11.110000 56.785000 11.310000 ;
        RECT 56.585000 11.540000 56.785000 11.740000 ;
        RECT 56.585000 11.970000 56.785000 12.170000 ;
        RECT 56.585000 12.400000 56.785000 12.600000 ;
        RECT 56.585000 12.830000 56.785000 13.030000 ;
        RECT 56.585000 13.260000 56.785000 13.460000 ;
        RECT 56.990000  8.960000 57.190000  9.160000 ;
        RECT 56.990000  9.390000 57.190000  9.590000 ;
        RECT 56.990000  9.820000 57.190000 10.020000 ;
        RECT 56.990000 10.250000 57.190000 10.450000 ;
        RECT 56.990000 10.680000 57.190000 10.880000 ;
        RECT 56.990000 11.110000 57.190000 11.310000 ;
        RECT 56.990000 11.540000 57.190000 11.740000 ;
        RECT 56.990000 11.970000 57.190000 12.170000 ;
        RECT 56.990000 12.400000 57.190000 12.600000 ;
        RECT 56.990000 12.830000 57.190000 13.030000 ;
        RECT 56.990000 13.260000 57.190000 13.460000 ;
        RECT 57.395000  8.960000 57.595000  9.160000 ;
        RECT 57.395000  9.390000 57.595000  9.590000 ;
        RECT 57.395000  9.820000 57.595000 10.020000 ;
        RECT 57.395000 10.250000 57.595000 10.450000 ;
        RECT 57.395000 10.680000 57.595000 10.880000 ;
        RECT 57.395000 11.110000 57.595000 11.310000 ;
        RECT 57.395000 11.540000 57.595000 11.740000 ;
        RECT 57.395000 11.970000 57.595000 12.170000 ;
        RECT 57.395000 12.400000 57.595000 12.600000 ;
        RECT 57.395000 12.830000 57.595000 13.030000 ;
        RECT 57.395000 13.260000 57.595000 13.460000 ;
        RECT 57.800000  8.960000 58.000000  9.160000 ;
        RECT 57.800000  9.390000 58.000000  9.590000 ;
        RECT 57.800000  9.820000 58.000000 10.020000 ;
        RECT 57.800000 10.250000 58.000000 10.450000 ;
        RECT 57.800000 10.680000 58.000000 10.880000 ;
        RECT 57.800000 11.110000 58.000000 11.310000 ;
        RECT 57.800000 11.540000 58.000000 11.740000 ;
        RECT 57.800000 11.970000 58.000000 12.170000 ;
        RECT 57.800000 12.400000 58.000000 12.600000 ;
        RECT 57.800000 12.830000 58.000000 13.030000 ;
        RECT 57.800000 13.260000 58.000000 13.460000 ;
        RECT 58.205000  8.960000 58.405000  9.160000 ;
        RECT 58.205000  9.390000 58.405000  9.590000 ;
        RECT 58.205000  9.820000 58.405000 10.020000 ;
        RECT 58.205000 10.250000 58.405000 10.450000 ;
        RECT 58.205000 10.680000 58.405000 10.880000 ;
        RECT 58.205000 11.110000 58.405000 11.310000 ;
        RECT 58.205000 11.540000 58.405000 11.740000 ;
        RECT 58.205000 11.970000 58.405000 12.170000 ;
        RECT 58.205000 12.400000 58.405000 12.600000 ;
        RECT 58.205000 12.830000 58.405000 13.030000 ;
        RECT 58.205000 13.260000 58.405000 13.460000 ;
        RECT 58.610000  8.960000 58.810000  9.160000 ;
        RECT 58.610000  9.390000 58.810000  9.590000 ;
        RECT 58.610000  9.820000 58.810000 10.020000 ;
        RECT 58.610000 10.250000 58.810000 10.450000 ;
        RECT 58.610000 10.680000 58.810000 10.880000 ;
        RECT 58.610000 11.110000 58.810000 11.310000 ;
        RECT 58.610000 11.540000 58.810000 11.740000 ;
        RECT 58.610000 11.970000 58.810000 12.170000 ;
        RECT 58.610000 12.400000 58.810000 12.600000 ;
        RECT 58.610000 12.830000 58.810000 13.030000 ;
        RECT 58.610000 13.260000 58.810000 13.460000 ;
        RECT 59.015000  8.960000 59.215000  9.160000 ;
        RECT 59.015000  9.390000 59.215000  9.590000 ;
        RECT 59.015000  9.820000 59.215000 10.020000 ;
        RECT 59.015000 10.250000 59.215000 10.450000 ;
        RECT 59.015000 10.680000 59.215000 10.880000 ;
        RECT 59.015000 11.110000 59.215000 11.310000 ;
        RECT 59.015000 11.540000 59.215000 11.740000 ;
        RECT 59.015000 11.970000 59.215000 12.170000 ;
        RECT 59.015000 12.400000 59.215000 12.600000 ;
        RECT 59.015000 12.830000 59.215000 13.030000 ;
        RECT 59.015000 13.260000 59.215000 13.460000 ;
        RECT 59.420000  8.960000 59.620000  9.160000 ;
        RECT 59.420000  9.390000 59.620000  9.590000 ;
        RECT 59.420000  9.820000 59.620000 10.020000 ;
        RECT 59.420000 10.250000 59.620000 10.450000 ;
        RECT 59.420000 10.680000 59.620000 10.880000 ;
        RECT 59.420000 11.110000 59.620000 11.310000 ;
        RECT 59.420000 11.540000 59.620000 11.740000 ;
        RECT 59.420000 11.970000 59.620000 12.170000 ;
        RECT 59.420000 12.400000 59.620000 12.600000 ;
        RECT 59.420000 12.830000 59.620000 13.030000 ;
        RECT 59.420000 13.260000 59.620000 13.460000 ;
        RECT 59.825000  8.960000 60.025000  9.160000 ;
        RECT 59.825000  9.390000 60.025000  9.590000 ;
        RECT 59.825000  9.820000 60.025000 10.020000 ;
        RECT 59.825000 10.250000 60.025000 10.450000 ;
        RECT 59.825000 10.680000 60.025000 10.880000 ;
        RECT 59.825000 11.110000 60.025000 11.310000 ;
        RECT 59.825000 11.540000 60.025000 11.740000 ;
        RECT 59.825000 11.970000 60.025000 12.170000 ;
        RECT 59.825000 12.400000 60.025000 12.600000 ;
        RECT 59.825000 12.830000 60.025000 13.030000 ;
        RECT 59.825000 13.260000 60.025000 13.460000 ;
        RECT 60.230000  8.960000 60.430000  9.160000 ;
        RECT 60.230000  9.390000 60.430000  9.590000 ;
        RECT 60.230000  9.820000 60.430000 10.020000 ;
        RECT 60.230000 10.250000 60.430000 10.450000 ;
        RECT 60.230000 10.680000 60.430000 10.880000 ;
        RECT 60.230000 11.110000 60.430000 11.310000 ;
        RECT 60.230000 11.540000 60.430000 11.740000 ;
        RECT 60.230000 11.970000 60.430000 12.170000 ;
        RECT 60.230000 12.400000 60.430000 12.600000 ;
        RECT 60.230000 12.830000 60.430000 13.030000 ;
        RECT 60.230000 13.260000 60.430000 13.460000 ;
        RECT 60.635000  8.960000 60.835000  9.160000 ;
        RECT 60.635000  9.390000 60.835000  9.590000 ;
        RECT 60.635000  9.820000 60.835000 10.020000 ;
        RECT 60.635000 10.250000 60.835000 10.450000 ;
        RECT 60.635000 10.680000 60.835000 10.880000 ;
        RECT 60.635000 11.110000 60.835000 11.310000 ;
        RECT 60.635000 11.540000 60.835000 11.740000 ;
        RECT 60.635000 11.970000 60.835000 12.170000 ;
        RECT 60.635000 12.400000 60.835000 12.600000 ;
        RECT 60.635000 12.830000 60.835000 13.030000 ;
        RECT 60.635000 13.260000 60.835000 13.460000 ;
        RECT 61.040000  8.960000 61.240000  9.160000 ;
        RECT 61.040000  9.390000 61.240000  9.590000 ;
        RECT 61.040000  9.820000 61.240000 10.020000 ;
        RECT 61.040000 10.250000 61.240000 10.450000 ;
        RECT 61.040000 10.680000 61.240000 10.880000 ;
        RECT 61.040000 11.110000 61.240000 11.310000 ;
        RECT 61.040000 11.540000 61.240000 11.740000 ;
        RECT 61.040000 11.970000 61.240000 12.170000 ;
        RECT 61.040000 12.400000 61.240000 12.600000 ;
        RECT 61.040000 12.830000 61.240000 13.030000 ;
        RECT 61.040000 13.260000 61.240000 13.460000 ;
        RECT 61.445000  8.960000 61.645000  9.160000 ;
        RECT 61.445000  9.390000 61.645000  9.590000 ;
        RECT 61.445000  9.820000 61.645000 10.020000 ;
        RECT 61.445000 10.250000 61.645000 10.450000 ;
        RECT 61.445000 10.680000 61.645000 10.880000 ;
        RECT 61.445000 11.110000 61.645000 11.310000 ;
        RECT 61.445000 11.540000 61.645000 11.740000 ;
        RECT 61.445000 11.970000 61.645000 12.170000 ;
        RECT 61.445000 12.400000 61.645000 12.600000 ;
        RECT 61.445000 12.830000 61.645000 13.030000 ;
        RECT 61.445000 13.260000 61.645000 13.460000 ;
        RECT 61.850000  8.960000 62.050000  9.160000 ;
        RECT 61.850000  9.390000 62.050000  9.590000 ;
        RECT 61.850000  9.820000 62.050000 10.020000 ;
        RECT 61.850000 10.250000 62.050000 10.450000 ;
        RECT 61.850000 10.680000 62.050000 10.880000 ;
        RECT 61.850000 11.110000 62.050000 11.310000 ;
        RECT 61.850000 11.540000 62.050000 11.740000 ;
        RECT 61.850000 11.970000 62.050000 12.170000 ;
        RECT 61.850000 12.400000 62.050000 12.600000 ;
        RECT 61.850000 12.830000 62.050000 13.030000 ;
        RECT 61.850000 13.260000 62.050000 13.460000 ;
        RECT 62.255000  8.960000 62.455000  9.160000 ;
        RECT 62.255000  9.390000 62.455000  9.590000 ;
        RECT 62.255000  9.820000 62.455000 10.020000 ;
        RECT 62.255000 10.250000 62.455000 10.450000 ;
        RECT 62.255000 10.680000 62.455000 10.880000 ;
        RECT 62.255000 11.110000 62.455000 11.310000 ;
        RECT 62.255000 11.540000 62.455000 11.740000 ;
        RECT 62.255000 11.970000 62.455000 12.170000 ;
        RECT 62.255000 12.400000 62.455000 12.600000 ;
        RECT 62.255000 12.830000 62.455000 13.030000 ;
        RECT 62.255000 13.260000 62.455000 13.460000 ;
        RECT 62.660000  8.960000 62.860000  9.160000 ;
        RECT 62.660000  9.390000 62.860000  9.590000 ;
        RECT 62.660000  9.820000 62.860000 10.020000 ;
        RECT 62.660000 10.250000 62.860000 10.450000 ;
        RECT 62.660000 10.680000 62.860000 10.880000 ;
        RECT 62.660000 11.110000 62.860000 11.310000 ;
        RECT 62.660000 11.540000 62.860000 11.740000 ;
        RECT 62.660000 11.970000 62.860000 12.170000 ;
        RECT 62.660000 12.400000 62.860000 12.600000 ;
        RECT 62.660000 12.830000 62.860000 13.030000 ;
        RECT 62.660000 13.260000 62.860000 13.460000 ;
        RECT 63.065000  8.960000 63.265000  9.160000 ;
        RECT 63.065000  9.390000 63.265000  9.590000 ;
        RECT 63.065000  9.820000 63.265000 10.020000 ;
        RECT 63.065000 10.250000 63.265000 10.450000 ;
        RECT 63.065000 10.680000 63.265000 10.880000 ;
        RECT 63.065000 11.110000 63.265000 11.310000 ;
        RECT 63.065000 11.540000 63.265000 11.740000 ;
        RECT 63.065000 11.970000 63.265000 12.170000 ;
        RECT 63.065000 12.400000 63.265000 12.600000 ;
        RECT 63.065000 12.830000 63.265000 13.030000 ;
        RECT 63.065000 13.260000 63.265000 13.460000 ;
        RECT 63.470000  8.960000 63.670000  9.160000 ;
        RECT 63.470000  9.390000 63.670000  9.590000 ;
        RECT 63.470000  9.820000 63.670000 10.020000 ;
        RECT 63.470000 10.250000 63.670000 10.450000 ;
        RECT 63.470000 10.680000 63.670000 10.880000 ;
        RECT 63.470000 11.110000 63.670000 11.310000 ;
        RECT 63.470000 11.540000 63.670000 11.740000 ;
        RECT 63.470000 11.970000 63.670000 12.170000 ;
        RECT 63.470000 12.400000 63.670000 12.600000 ;
        RECT 63.470000 12.830000 63.670000 13.030000 ;
        RECT 63.470000 13.260000 63.670000 13.460000 ;
        RECT 63.875000  8.960000 64.075000  9.160000 ;
        RECT 63.875000  9.390000 64.075000  9.590000 ;
        RECT 63.875000  9.820000 64.075000 10.020000 ;
        RECT 63.875000 10.250000 64.075000 10.450000 ;
        RECT 63.875000 10.680000 64.075000 10.880000 ;
        RECT 63.875000 11.110000 64.075000 11.310000 ;
        RECT 63.875000 11.540000 64.075000 11.740000 ;
        RECT 63.875000 11.970000 64.075000 12.170000 ;
        RECT 63.875000 12.400000 64.075000 12.600000 ;
        RECT 63.875000 12.830000 64.075000 13.030000 ;
        RECT 63.875000 13.260000 64.075000 13.460000 ;
        RECT 64.280000  8.960000 64.480000  9.160000 ;
        RECT 64.280000  9.390000 64.480000  9.590000 ;
        RECT 64.280000  9.820000 64.480000 10.020000 ;
        RECT 64.280000 10.250000 64.480000 10.450000 ;
        RECT 64.280000 10.680000 64.480000 10.880000 ;
        RECT 64.280000 11.110000 64.480000 11.310000 ;
        RECT 64.280000 11.540000 64.480000 11.740000 ;
        RECT 64.280000 11.970000 64.480000 12.170000 ;
        RECT 64.280000 12.400000 64.480000 12.600000 ;
        RECT 64.280000 12.830000 64.480000 13.030000 ;
        RECT 64.280000 13.260000 64.480000 13.460000 ;
        RECT 64.685000  8.960000 64.885000  9.160000 ;
        RECT 64.685000  9.390000 64.885000  9.590000 ;
        RECT 64.685000  9.820000 64.885000 10.020000 ;
        RECT 64.685000 10.250000 64.885000 10.450000 ;
        RECT 64.685000 10.680000 64.885000 10.880000 ;
        RECT 64.685000 11.110000 64.885000 11.310000 ;
        RECT 64.685000 11.540000 64.885000 11.740000 ;
        RECT 64.685000 11.970000 64.885000 12.170000 ;
        RECT 64.685000 12.400000 64.885000 12.600000 ;
        RECT 64.685000 12.830000 64.885000 13.030000 ;
        RECT 64.685000 13.260000 64.885000 13.460000 ;
        RECT 65.090000  8.960000 65.290000  9.160000 ;
        RECT 65.090000  9.390000 65.290000  9.590000 ;
        RECT 65.090000  9.820000 65.290000 10.020000 ;
        RECT 65.090000 10.250000 65.290000 10.450000 ;
        RECT 65.090000 10.680000 65.290000 10.880000 ;
        RECT 65.090000 11.110000 65.290000 11.310000 ;
        RECT 65.090000 11.540000 65.290000 11.740000 ;
        RECT 65.090000 11.970000 65.290000 12.170000 ;
        RECT 65.090000 12.400000 65.290000 12.600000 ;
        RECT 65.090000 12.830000 65.290000 13.030000 ;
        RECT 65.090000 13.260000 65.290000 13.460000 ;
        RECT 65.495000  8.960000 65.695000  9.160000 ;
        RECT 65.495000  9.390000 65.695000  9.590000 ;
        RECT 65.495000  9.820000 65.695000 10.020000 ;
        RECT 65.495000 10.250000 65.695000 10.450000 ;
        RECT 65.495000 10.680000 65.695000 10.880000 ;
        RECT 65.495000 11.110000 65.695000 11.310000 ;
        RECT 65.495000 11.540000 65.695000 11.740000 ;
        RECT 65.495000 11.970000 65.695000 12.170000 ;
        RECT 65.495000 12.400000 65.695000 12.600000 ;
        RECT 65.495000 12.830000 65.695000 13.030000 ;
        RECT 65.495000 13.260000 65.695000 13.460000 ;
        RECT 65.900000  8.960000 66.100000  9.160000 ;
        RECT 65.900000  9.390000 66.100000  9.590000 ;
        RECT 65.900000  9.820000 66.100000 10.020000 ;
        RECT 65.900000 10.250000 66.100000 10.450000 ;
        RECT 65.900000 10.680000 66.100000 10.880000 ;
        RECT 65.900000 11.110000 66.100000 11.310000 ;
        RECT 65.900000 11.540000 66.100000 11.740000 ;
        RECT 65.900000 11.970000 66.100000 12.170000 ;
        RECT 65.900000 12.400000 66.100000 12.600000 ;
        RECT 65.900000 12.830000 66.100000 13.030000 ;
        RECT 65.900000 13.260000 66.100000 13.460000 ;
        RECT 66.305000  8.960000 66.505000  9.160000 ;
        RECT 66.305000  9.390000 66.505000  9.590000 ;
        RECT 66.305000  9.820000 66.505000 10.020000 ;
        RECT 66.305000 10.250000 66.505000 10.450000 ;
        RECT 66.305000 10.680000 66.505000 10.880000 ;
        RECT 66.305000 11.110000 66.505000 11.310000 ;
        RECT 66.305000 11.540000 66.505000 11.740000 ;
        RECT 66.305000 11.970000 66.505000 12.170000 ;
        RECT 66.305000 12.400000 66.505000 12.600000 ;
        RECT 66.305000 12.830000 66.505000 13.030000 ;
        RECT 66.305000 13.260000 66.505000 13.460000 ;
        RECT 66.710000  8.960000 66.910000  9.160000 ;
        RECT 66.710000  9.390000 66.910000  9.590000 ;
        RECT 66.710000  9.820000 66.910000 10.020000 ;
        RECT 66.710000 10.250000 66.910000 10.450000 ;
        RECT 66.710000 10.680000 66.910000 10.880000 ;
        RECT 66.710000 11.110000 66.910000 11.310000 ;
        RECT 66.710000 11.540000 66.910000 11.740000 ;
        RECT 66.710000 11.970000 66.910000 12.170000 ;
        RECT 66.710000 12.400000 66.910000 12.600000 ;
        RECT 66.710000 12.830000 66.910000 13.030000 ;
        RECT 66.710000 13.260000 66.910000 13.460000 ;
        RECT 67.115000  8.960000 67.315000  9.160000 ;
        RECT 67.115000  9.390000 67.315000  9.590000 ;
        RECT 67.115000  9.820000 67.315000 10.020000 ;
        RECT 67.115000 10.250000 67.315000 10.450000 ;
        RECT 67.115000 10.680000 67.315000 10.880000 ;
        RECT 67.115000 11.110000 67.315000 11.310000 ;
        RECT 67.115000 11.540000 67.315000 11.740000 ;
        RECT 67.115000 11.970000 67.315000 12.170000 ;
        RECT 67.115000 12.400000 67.315000 12.600000 ;
        RECT 67.115000 12.830000 67.315000 13.030000 ;
        RECT 67.115000 13.260000 67.315000 13.460000 ;
        RECT 67.520000  8.960000 67.720000  9.160000 ;
        RECT 67.520000  9.390000 67.720000  9.590000 ;
        RECT 67.520000  9.820000 67.720000 10.020000 ;
        RECT 67.520000 10.250000 67.720000 10.450000 ;
        RECT 67.520000 10.680000 67.720000 10.880000 ;
        RECT 67.520000 11.110000 67.720000 11.310000 ;
        RECT 67.520000 11.540000 67.720000 11.740000 ;
        RECT 67.520000 11.970000 67.720000 12.170000 ;
        RECT 67.520000 12.400000 67.720000 12.600000 ;
        RECT 67.520000 12.830000 67.720000 13.030000 ;
        RECT 67.520000 13.260000 67.720000 13.460000 ;
        RECT 67.925000  8.960000 68.125000  9.160000 ;
        RECT 67.925000  9.390000 68.125000  9.590000 ;
        RECT 67.925000  9.820000 68.125000 10.020000 ;
        RECT 67.925000 10.250000 68.125000 10.450000 ;
        RECT 67.925000 10.680000 68.125000 10.880000 ;
        RECT 67.925000 11.110000 68.125000 11.310000 ;
        RECT 67.925000 11.540000 68.125000 11.740000 ;
        RECT 67.925000 11.970000 68.125000 12.170000 ;
        RECT 67.925000 12.400000 68.125000 12.600000 ;
        RECT 67.925000 12.830000 68.125000 13.030000 ;
        RECT 67.925000 13.260000 68.125000 13.460000 ;
        RECT 68.330000  8.960000 68.530000  9.160000 ;
        RECT 68.330000  9.390000 68.530000  9.590000 ;
        RECT 68.330000  9.820000 68.530000 10.020000 ;
        RECT 68.330000 10.250000 68.530000 10.450000 ;
        RECT 68.330000 10.680000 68.530000 10.880000 ;
        RECT 68.330000 11.110000 68.530000 11.310000 ;
        RECT 68.330000 11.540000 68.530000 11.740000 ;
        RECT 68.330000 11.970000 68.530000 12.170000 ;
        RECT 68.330000 12.400000 68.530000 12.600000 ;
        RECT 68.330000 12.830000 68.530000 13.030000 ;
        RECT 68.330000 13.260000 68.530000 13.460000 ;
        RECT 68.735000  8.960000 68.935000  9.160000 ;
        RECT 68.735000  9.390000 68.935000  9.590000 ;
        RECT 68.735000  9.820000 68.935000 10.020000 ;
        RECT 68.735000 10.250000 68.935000 10.450000 ;
        RECT 68.735000 10.680000 68.935000 10.880000 ;
        RECT 68.735000 11.110000 68.935000 11.310000 ;
        RECT 68.735000 11.540000 68.935000 11.740000 ;
        RECT 68.735000 11.970000 68.935000 12.170000 ;
        RECT 68.735000 12.400000 68.935000 12.600000 ;
        RECT 68.735000 12.830000 68.935000 13.030000 ;
        RECT 68.735000 13.260000 68.935000 13.460000 ;
        RECT 69.140000  8.960000 69.340000  9.160000 ;
        RECT 69.140000  9.390000 69.340000  9.590000 ;
        RECT 69.140000  9.820000 69.340000 10.020000 ;
        RECT 69.140000 10.250000 69.340000 10.450000 ;
        RECT 69.140000 10.680000 69.340000 10.880000 ;
        RECT 69.140000 11.110000 69.340000 11.310000 ;
        RECT 69.140000 11.540000 69.340000 11.740000 ;
        RECT 69.140000 11.970000 69.340000 12.170000 ;
        RECT 69.140000 12.400000 69.340000 12.600000 ;
        RECT 69.140000 12.830000 69.340000 13.030000 ;
        RECT 69.140000 13.260000 69.340000 13.460000 ;
        RECT 69.545000  8.960000 69.745000  9.160000 ;
        RECT 69.545000  9.390000 69.745000  9.590000 ;
        RECT 69.545000  9.820000 69.745000 10.020000 ;
        RECT 69.545000 10.250000 69.745000 10.450000 ;
        RECT 69.545000 10.680000 69.745000 10.880000 ;
        RECT 69.545000 11.110000 69.745000 11.310000 ;
        RECT 69.545000 11.540000 69.745000 11.740000 ;
        RECT 69.545000 11.970000 69.745000 12.170000 ;
        RECT 69.545000 12.400000 69.745000 12.600000 ;
        RECT 69.545000 12.830000 69.745000 13.030000 ;
        RECT 69.545000 13.260000 69.745000 13.460000 ;
        RECT 69.950000  8.960000 70.150000  9.160000 ;
        RECT 69.950000  9.390000 70.150000  9.590000 ;
        RECT 69.950000  9.820000 70.150000 10.020000 ;
        RECT 69.950000 10.250000 70.150000 10.450000 ;
        RECT 69.950000 10.680000 70.150000 10.880000 ;
        RECT 69.950000 11.110000 70.150000 11.310000 ;
        RECT 69.950000 11.540000 70.150000 11.740000 ;
        RECT 69.950000 11.970000 70.150000 12.170000 ;
        RECT 69.950000 12.400000 70.150000 12.600000 ;
        RECT 69.950000 12.830000 70.150000 13.030000 ;
        RECT 69.950000 13.260000 70.150000 13.460000 ;
        RECT 70.355000  8.960000 70.555000  9.160000 ;
        RECT 70.355000  9.390000 70.555000  9.590000 ;
        RECT 70.355000  9.820000 70.555000 10.020000 ;
        RECT 70.355000 10.250000 70.555000 10.450000 ;
        RECT 70.355000 10.680000 70.555000 10.880000 ;
        RECT 70.355000 11.110000 70.555000 11.310000 ;
        RECT 70.355000 11.540000 70.555000 11.740000 ;
        RECT 70.355000 11.970000 70.555000 12.170000 ;
        RECT 70.355000 12.400000 70.555000 12.600000 ;
        RECT 70.355000 12.830000 70.555000 13.030000 ;
        RECT 70.355000 13.260000 70.555000 13.460000 ;
        RECT 70.760000  8.960000 70.960000  9.160000 ;
        RECT 70.760000  9.390000 70.960000  9.590000 ;
        RECT 70.760000  9.820000 70.960000 10.020000 ;
        RECT 70.760000 10.250000 70.960000 10.450000 ;
        RECT 70.760000 10.680000 70.960000 10.880000 ;
        RECT 70.760000 11.110000 70.960000 11.310000 ;
        RECT 70.760000 11.540000 70.960000 11.740000 ;
        RECT 70.760000 11.970000 70.960000 12.170000 ;
        RECT 70.760000 12.400000 70.960000 12.600000 ;
        RECT 70.760000 12.830000 70.960000 13.030000 ;
        RECT 70.760000 13.260000 70.960000 13.460000 ;
        RECT 71.165000  8.960000 71.365000  9.160000 ;
        RECT 71.165000  9.390000 71.365000  9.590000 ;
        RECT 71.165000  9.820000 71.365000 10.020000 ;
        RECT 71.165000 10.250000 71.365000 10.450000 ;
        RECT 71.165000 10.680000 71.365000 10.880000 ;
        RECT 71.165000 11.110000 71.365000 11.310000 ;
        RECT 71.165000 11.540000 71.365000 11.740000 ;
        RECT 71.165000 11.970000 71.365000 12.170000 ;
        RECT 71.165000 12.400000 71.365000 12.600000 ;
        RECT 71.165000 12.830000 71.365000 13.030000 ;
        RECT 71.165000 13.260000 71.365000 13.460000 ;
        RECT 71.570000  8.960000 71.770000  9.160000 ;
        RECT 71.570000  9.390000 71.770000  9.590000 ;
        RECT 71.570000  9.820000 71.770000 10.020000 ;
        RECT 71.570000 10.250000 71.770000 10.450000 ;
        RECT 71.570000 10.680000 71.770000 10.880000 ;
        RECT 71.570000 11.110000 71.770000 11.310000 ;
        RECT 71.570000 11.540000 71.770000 11.740000 ;
        RECT 71.570000 11.970000 71.770000 12.170000 ;
        RECT 71.570000 12.400000 71.770000 12.600000 ;
        RECT 71.570000 12.830000 71.770000 13.030000 ;
        RECT 71.570000 13.260000 71.770000 13.460000 ;
        RECT 71.975000  8.960000 72.175000  9.160000 ;
        RECT 71.975000  9.390000 72.175000  9.590000 ;
        RECT 71.975000  9.820000 72.175000 10.020000 ;
        RECT 71.975000 10.250000 72.175000 10.450000 ;
        RECT 71.975000 10.680000 72.175000 10.880000 ;
        RECT 71.975000 11.110000 72.175000 11.310000 ;
        RECT 71.975000 11.540000 72.175000 11.740000 ;
        RECT 71.975000 11.970000 72.175000 12.170000 ;
        RECT 71.975000 12.400000 72.175000 12.600000 ;
        RECT 71.975000 12.830000 72.175000 13.030000 ;
        RECT 71.975000 13.260000 72.175000 13.460000 ;
        RECT 72.380000  8.960000 72.580000  9.160000 ;
        RECT 72.380000  9.390000 72.580000  9.590000 ;
        RECT 72.380000  9.820000 72.580000 10.020000 ;
        RECT 72.380000 10.250000 72.580000 10.450000 ;
        RECT 72.380000 10.680000 72.580000 10.880000 ;
        RECT 72.380000 11.110000 72.580000 11.310000 ;
        RECT 72.380000 11.540000 72.580000 11.740000 ;
        RECT 72.380000 11.970000 72.580000 12.170000 ;
        RECT 72.380000 12.400000 72.580000 12.600000 ;
        RECT 72.380000 12.830000 72.580000 13.030000 ;
        RECT 72.380000 13.260000 72.580000 13.460000 ;
        RECT 72.785000  8.960000 72.985000  9.160000 ;
        RECT 72.785000  9.390000 72.985000  9.590000 ;
        RECT 72.785000  9.820000 72.985000 10.020000 ;
        RECT 72.785000 10.250000 72.985000 10.450000 ;
        RECT 72.785000 10.680000 72.985000 10.880000 ;
        RECT 72.785000 11.110000 72.985000 11.310000 ;
        RECT 72.785000 11.540000 72.985000 11.740000 ;
        RECT 72.785000 11.970000 72.985000 12.170000 ;
        RECT 72.785000 12.400000 72.985000 12.600000 ;
        RECT 72.785000 12.830000 72.985000 13.030000 ;
        RECT 72.785000 13.260000 72.985000 13.460000 ;
        RECT 73.190000  8.960000 73.390000  9.160000 ;
        RECT 73.190000  9.390000 73.390000  9.590000 ;
        RECT 73.190000  9.820000 73.390000 10.020000 ;
        RECT 73.190000 10.250000 73.390000 10.450000 ;
        RECT 73.190000 10.680000 73.390000 10.880000 ;
        RECT 73.190000 11.110000 73.390000 11.310000 ;
        RECT 73.190000 11.540000 73.390000 11.740000 ;
        RECT 73.190000 11.970000 73.390000 12.170000 ;
        RECT 73.190000 12.400000 73.390000 12.600000 ;
        RECT 73.190000 12.830000 73.390000 13.030000 ;
        RECT 73.190000 13.260000 73.390000 13.460000 ;
        RECT 73.595000  8.960000 73.795000  9.160000 ;
        RECT 73.595000  9.390000 73.795000  9.590000 ;
        RECT 73.595000  9.820000 73.795000 10.020000 ;
        RECT 73.595000 10.250000 73.795000 10.450000 ;
        RECT 73.595000 10.680000 73.795000 10.880000 ;
        RECT 73.595000 11.110000 73.795000 11.310000 ;
        RECT 73.595000 11.540000 73.795000 11.740000 ;
        RECT 73.595000 11.970000 73.795000 12.170000 ;
        RECT 73.595000 12.400000 73.795000 12.600000 ;
        RECT 73.595000 12.830000 73.795000 13.030000 ;
        RECT 73.595000 13.260000 73.795000 13.460000 ;
        RECT 74.000000  8.960000 74.200000  9.160000 ;
        RECT 74.000000  9.390000 74.200000  9.590000 ;
        RECT 74.000000  9.820000 74.200000 10.020000 ;
        RECT 74.000000 10.250000 74.200000 10.450000 ;
        RECT 74.000000 10.680000 74.200000 10.880000 ;
        RECT 74.000000 11.110000 74.200000 11.310000 ;
        RECT 74.000000 11.540000 74.200000 11.740000 ;
        RECT 74.000000 11.970000 74.200000 12.170000 ;
        RECT 74.000000 12.400000 74.200000 12.600000 ;
        RECT 74.000000 12.830000 74.200000 13.030000 ;
        RECT 74.000000 13.260000 74.200000 13.460000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2.035000 1.270000 7.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 2.035000 75.000000 7.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 2.135000 1.270000 7.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 2.135000 75.000000 7.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 14.935000 0.965000 18.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035000 14.935000 75.000000 18.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 15.035000 0.965000 18.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 15.035000 75.000000 18.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 19.785000 1.270000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 70.035000 1.270000 95.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 19.785000 75.000000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 70.035000 75.000000 95.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 19.885000 1.270000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 70.035000 1.270000 94.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 19.885000 75.000000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 70.035000 75.000000 94.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 64.085000 1.270000 68.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 64.085000 75.000000 68.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 64.185000 1.270000 68.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 64.185000 75.000000 68.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 36.735000 1.270000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 47.735000 1.270000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 51.645000 1.270000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 56.405000 1.270000 56.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 36.735000 75.000000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 47.735000 75.000000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.645000 75.000000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 56.405000 75.000000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 36.840000 1.270000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 47.735000 1.270000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 36.840000 75.000000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 47.735000 75.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 41.585000 1.270000 46.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 41.585000 75.000000 46.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 41.685000 1.270000 46.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 41.685000 75.000000 46.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 25.835000 1.270000 30.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 25.835000 75.000000 30.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 25.935000 1.270000 30.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 25.935000 75.000000 30.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 58.235000 1.270000 62.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 58.235000 75.000000 62.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 58.335000 1.270000 62.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 58.335000 75.000000 62.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 31.885000 1.270000 35.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 31.885000 75.000000 35.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 31.985000 1.270000 35.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 31.985000 75.000000 35.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met1 ;
      RECT 0.000000 0.000000 75.000000 200.000000 ;
  END
END sky130_fd_io__overlay_vccd_hvc
END LIBRARY
