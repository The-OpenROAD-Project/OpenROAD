module gcd (clk,
    req_rdy,
    req_val,
    reset,
    resp_rdy,
    resp_val,
    req_msg,
    resp_msg);
 input clk;
 output req_rdy;
 input req_val;
 input reset;
 input resp_rdy;
 output resp_val;
 input [31:0] req_msg;
 output [15:0] resp_msg;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire net2;
 wire net1;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire clknet_2_3__leaf_clk;
 wire _171_;
 wire _172_;
 wire clknet_2_2__leaf_clk;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire clknet_2_1__leaf_clk;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire clknet_2_0__leaf_clk;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire clknet_0_clk;
 wire _205_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire \ctrl.state.out[1] ;
 wire \ctrl.state.out[2] ;
 wire \dpath.a_lt_b$in0[0] ;
 wire \dpath.a_lt_b$in0[10] ;
 wire \dpath.a_lt_b$in0[11] ;
 wire \dpath.a_lt_b$in0[12] ;
 wire \dpath.a_lt_b$in0[13] ;
 wire \dpath.a_lt_b$in0[14] ;
 wire \dpath.a_lt_b$in0[15] ;
 wire \dpath.a_lt_b$in0[1] ;
 wire \dpath.a_lt_b$in0[2] ;
 wire \dpath.a_lt_b$in0[3] ;
 wire \dpath.a_lt_b$in0[4] ;
 wire \dpath.a_lt_b$in0[5] ;
 wire \dpath.a_lt_b$in0[6] ;
 wire \dpath.a_lt_b$in0[7] ;
 wire \dpath.a_lt_b$in0[8] ;
 wire \dpath.a_lt_b$in0[9] ;
 wire \dpath.a_lt_b$in1[0] ;
 wire \dpath.a_lt_b$in1[10] ;
 wire \dpath.a_lt_b$in1[11] ;
 wire \dpath.a_lt_b$in1[12] ;
 wire \dpath.a_lt_b$in1[13] ;
 wire \dpath.a_lt_b$in1[14] ;
 wire \dpath.a_lt_b$in1[15] ;
 wire \dpath.a_lt_b$in1[1] ;
 wire \dpath.a_lt_b$in1[2] ;
 wire \dpath.a_lt_b$in1[3] ;
 wire \dpath.a_lt_b$in1[4] ;
 wire \dpath.a_lt_b$in1[5] ;
 wire \dpath.a_lt_b$in1[6] ;
 wire \dpath.a_lt_b$in1[7] ;
 wire \dpath.a_lt_b$in1[8] ;
 wire \dpath.a_lt_b$in1[9] ;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;

 sky130_fd_sc_hs__nor2b_4 _252_ (.A(\dpath.a_lt_b$in0[0] ),
    .B_N(\dpath.a_lt_b$in1[0] ),
    .Y(_035_));
 sky130_fd_sc_hs__nor2b_2 _253_ (.A(\dpath.a_lt_b$in0[1] ),
    .B_N(\dpath.a_lt_b$in1[1] ),
    .Y(_036_));
 sky130_fd_sc_hs__inv_2 _254_ (.A(\dpath.a_lt_b$in1[1] ),
    .Y(_037_));
 sky130_fd_sc_hs__nand2_1 _255_ (.A(_037_),
    .B(\dpath.a_lt_b$in0[1] ),
    .Y(_038_));
 sky130_fd_sc_hs__o21ai_4 _256_ (.A1(_035_),
    .A2(_036_),
    .B1(_038_),
    .Y(_039_));
 sky130_fd_sc_hs__nand2b_1 _257_ (.A_N(\dpath.a_lt_b$in1[3] ),
    .B(\dpath.a_lt_b$in0[3] ),
    .Y(_040_));
 sky130_fd_sc_hs__nand2b_1 _258_ (.A_N(\dpath.a_lt_b$in0[3] ),
    .B(\dpath.a_lt_b$in1[3] ),
    .Y(_041_));
 sky130_fd_sc_hs__nand2_2 _259_ (.A(_040_),
    .B(_041_),
    .Y(_042_));
 sky130_fd_sc_hs__nand2b_2 _260_ (.A_N(\dpath.a_lt_b$in1[2] ),
    .B(\dpath.a_lt_b$in0[2] ),
    .Y(_043_));
 sky130_fd_sc_hs__nand2b_2 _261_ (.A_N(\dpath.a_lt_b$in0[2] ),
    .B(\dpath.a_lt_b$in1[2] ),
    .Y(_044_));
 sky130_fd_sc_hs__nand2_2 _262_ (.A(_043_),
    .B(_044_),
    .Y(_045_));
 sky130_fd_sc_hs__nor2_2 _263_ (.A(_042_),
    .B(_045_),
    .Y(_046_));
 sky130_fd_sc_hs__nand2_2 _264_ (.A(_039_),
    .B(_046_),
    .Y(_047_));
 sky130_fd_sc_hs__inv_1 _265_ (.A(\dpath.a_lt_b$in1[3] ),
    .Y(_048_));
 sky130_fd_sc_hs__nor2_1 _266_ (.A(\dpath.a_lt_b$in0[3] ),
    .B(_048_),
    .Y(_049_));
 sky130_fd_sc_hs__o21a_1 _267_ (.A1(_043_),
    .A2(_049_),
    .B1(_040_),
    .X(_050_));
 sky130_fd_sc_hs__nand2_8 _268_ (.A(_047_),
    .B(_050_),
    .Y(_051_));
 sky130_fd_sc_hs__inv_1 _269_ (.A(\dpath.a_lt_b$in1[7] ),
    .Y(_052_));
 sky130_fd_sc_hs__nand2_1 _270_ (.A(_052_),
    .B(\dpath.a_lt_b$in0[7] ),
    .Y(_053_));
 sky130_fd_sc_hs__nand2b_1 _271_ (.A_N(\dpath.a_lt_b$in0[7] ),
    .B(\dpath.a_lt_b$in1[7] ),
    .Y(_054_));
 sky130_fd_sc_hs__and2_2 _272_ (.A(_053_),
    .B(_054_),
    .X(_055_));
 sky130_fd_sc_hs__xnor2_4 _273_ (.A(\dpath.a_lt_b$in1[6] ),
    .B(\dpath.a_lt_b$in0[6] ),
    .Y(_056_));
 sky130_fd_sc_hs__nand2_2 _274_ (.A(_055_),
    .B(_056_),
    .Y(_057_));
 sky130_fd_sc_hs__inv_1 _275_ (.A(\dpath.a_lt_b$in1[5] ),
    .Y(_058_));
 sky130_fd_sc_hs__nand2_2 _276_ (.A(_058_),
    .B(\dpath.a_lt_b$in0[5] ),
    .Y(_059_));
 sky130_fd_sc_hs__nand2b_2 _277_ (.A_N(\dpath.a_lt_b$in0[5] ),
    .B(\dpath.a_lt_b$in1[5] ),
    .Y(_060_));
 sky130_fd_sc_hs__and2_4 _278_ (.A(_059_),
    .B(_060_),
    .X(_061_));
 sky130_fd_sc_hs__xnor2_4 _279_ (.A(\dpath.a_lt_b$in1[4] ),
    .B(\dpath.a_lt_b$in0[4] ),
    .Y(_062_));
 sky130_fd_sc_hs__nand2_1 _280_ (.A(_061_),
    .B(_062_),
    .Y(_063_));
 sky130_fd_sc_hs__nor2_4 _281_ (.A(_057_),
    .B(_063_),
    .Y(_064_));
 sky130_fd_sc_hs__nand2_2 _282_ (.A(_051_),
    .B(_064_),
    .Y(_065_));
 sky130_fd_sc_hs__inv_2 _283_ (.A(\dpath.a_lt_b$in1[6] ),
    .Y(_066_));
 sky130_fd_sc_hs__nand2_1 _284_ (.A(_066_),
    .B(\dpath.a_lt_b$in0[6] ),
    .Y(_067_));
 sky130_fd_sc_hs__a21boi_1 _285_ (.A1(_053_),
    .A2(_067_),
    .B1_N(_054_),
    .Y(_068_));
 sky130_fd_sc_hs__inv_2 _286_ (.A(\dpath.a_lt_b$in1[4] ),
    .Y(_069_));
 sky130_fd_sc_hs__nand2_1 _287_ (.A(_069_),
    .B(\dpath.a_lt_b$in0[4] ),
    .Y(_070_));
 sky130_fd_sc_hs__nand2_1 _288_ (.A(_059_),
    .B(_070_),
    .Y(_071_));
 sky130_fd_sc_hs__nand2_1 _289_ (.A(_071_),
    .B(_060_),
    .Y(_072_));
 sky130_fd_sc_hs__nor2_2 _290_ (.A(_072_),
    .B(_057_),
    .Y(_073_));
 sky130_fd_sc_hs__nor2_2 _291_ (.A(_068_),
    .B(_073_),
    .Y(_074_));
 sky130_fd_sc_hs__nand2_8 _292_ (.A(_065_),
    .B(_074_),
    .Y(_075_));
 sky130_fd_sc_hs__inv_2 _293_ (.A(\dpath.a_lt_b$in0[9] ),
    .Y(_076_));
 sky130_fd_sc_hs__xnor2_4 _294_ (.A(\dpath.a_lt_b$in1[9] ),
    .B(_076_),
    .Y(_077_));
 sky130_fd_sc_hs__inv_2 _295_ (.A(\dpath.a_lt_b$in1[8] ),
    .Y(_078_));
 sky130_fd_sc_hs__nand2_4 _296_ (.A(_078_),
    .B(\dpath.a_lt_b$in0[8] ),
    .Y(_079_));
 sky130_fd_sc_hs__inv_2 _297_ (.A(\dpath.a_lt_b$in0[8] ),
    .Y(_080_));
 sky130_fd_sc_hs__nand2_1 _298_ (.A(_080_),
    .B(\dpath.a_lt_b$in1[8] ),
    .Y(_081_));
 sky130_fd_sc_hs__nand2_4 _299_ (.A(_079_),
    .B(_081_),
    .Y(_082_));
 sky130_fd_sc_hs__xnor2_4 _300_ (.A(\dpath.a_lt_b$in1[10] ),
    .B(\dpath.a_lt_b$in0[10] ),
    .Y(_083_));
 sky130_fd_sc_hs__inv_1 _301_ (.A(\dpath.a_lt_b$in1[11] ),
    .Y(_084_));
 sky130_fd_sc_hs__nand2_2 _302_ (.A(_084_),
    .B(\dpath.a_lt_b$in0[11] ),
    .Y(_085_));
 sky130_fd_sc_hs__inv_1 _303_ (.A(\dpath.a_lt_b$in0[11] ),
    .Y(_086_));
 sky130_fd_sc_hs__nand2_1 _304_ (.A(_086_),
    .B(\dpath.a_lt_b$in1[11] ),
    .Y(_087_));
 sky130_fd_sc_hs__nand3_4 _305_ (.A(_083_),
    .B(_085_),
    .C(_087_),
    .Y(_088_));
 sky130_fd_sc_hs__nor3_4 _306_ (.A(_077_),
    .B(_082_),
    .C(_088_),
    .Y(_089_));
 sky130_fd_sc_hs__nand2_2 _307_ (.A(_075_),
    .B(_089_),
    .Y(_090_));
 sky130_fd_sc_hs__inv_1 _308_ (.A(\dpath.a_lt_b$in1[10] ),
    .Y(_091_));
 sky130_fd_sc_hs__nand2_1 _309_ (.A(_091_),
    .B(\dpath.a_lt_b$in0[10] ),
    .Y(_092_));
 sky130_fd_sc_hs__nand2_2 _310_ (.A(_085_),
    .B(_087_),
    .Y(_093_));
 sky130_fd_sc_hs__o21ai_1 _311_ (.A1(_092_),
    .A2(_093_),
    .B1(_085_),
    .Y(_094_));
 sky130_fd_sc_hs__maj3_1 _312_ (.A(\dpath.a_lt_b$in1[9] ),
    .B(_079_),
    .C(_076_),
    .X(_095_));
 sky130_fd_sc_hs__nor2_1 _313_ (.A(_088_),
    .B(_095_),
    .Y(_096_));
 sky130_fd_sc_hs__nor2_1 _314_ (.A(_094_),
    .B(_096_),
    .Y(_097_));
 sky130_fd_sc_hs__nand2_2 _315_ (.A(_090_),
    .B(_097_),
    .Y(_098_));
 sky130_fd_sc_hs__inv_2 _316_ (.A(\dpath.a_lt_b$in0[12] ),
    .Y(_099_));
 sky130_fd_sc_hs__nor2_2 _317_ (.A(\dpath.a_lt_b$in1[12] ),
    .B(_099_),
    .Y(_100_));
 sky130_fd_sc_hs__clkinv_2 _318_ (.A(_100_),
    .Y(_101_));
 sky130_fd_sc_hs__nand2_1 _319_ (.A(_099_),
    .B(\dpath.a_lt_b$in1[12] ),
    .Y(_102_));
 sky130_fd_sc_hs__nand2_8 _320_ (.A(_101_),
    .B(_102_),
    .Y(_103_));
 sky130_fd_sc_hs__inv_2 _321_ (.A(\dpath.a_lt_b$in1[13] ),
    .Y(_104_));
 sky130_fd_sc_hs__nor2_1 _322_ (.A(\dpath.a_lt_b$in0[13] ),
    .B(_104_),
    .Y(_105_));
 sky130_fd_sc_hs__and2_1 _323_ (.A(_104_),
    .B(\dpath.a_lt_b$in0[13] ),
    .X(_106_));
 sky130_fd_sc_hs__nor2_2 _324_ (.A(_105_),
    .B(_106_),
    .Y(_107_));
 sky130_fd_sc_hs__inv_2 _325_ (.A(_107_),
    .Y(_108_));
 sky130_fd_sc_hs__nor2_1 _326_ (.A(_103_),
    .B(_108_),
    .Y(_109_));
 sky130_fd_sc_hs__nand2_2 _327_ (.A(_098_),
    .B(_109_),
    .Y(_110_));
 sky130_fd_sc_hs__a21oi_2 _328_ (.A1(_107_),
    .A2(_100_),
    .B1(_106_),
    .Y(_111_));
 sky130_fd_sc_hs__nand2_2 _329_ (.A(_110_),
    .B(_111_),
    .Y(_112_));
 sky130_fd_sc_hs__xnor2_4 _330_ (.A(\dpath.a_lt_b$in1[14] ),
    .B(\dpath.a_lt_b$in0[14] ),
    .Y(_113_));
 sky130_fd_sc_hs__nand2_2 _331_ (.A(_112_),
    .B(_113_),
    .Y(_114_));
 sky130_fd_sc_hs__inv_1 _332_ (.A(\dpath.a_lt_b$in0[14] ),
    .Y(_115_));
 sky130_fd_sc_hs__nor2_1 _333_ (.A(\dpath.a_lt_b$in1[14] ),
    .B(_115_),
    .Y(_116_));
 sky130_fd_sc_hs__inv_1 _334_ (.A(_116_),
    .Y(_117_));
 sky130_fd_sc_hs__nand2_1 _335_ (.A(_114_),
    .B(_117_),
    .Y(_118_));
 sky130_fd_sc_hs__inv_2 _336_ (.A(\dpath.a_lt_b$in1[15] ),
    .Y(_119_));
 sky130_fd_sc_hs__nor2_1 _337_ (.A(\dpath.a_lt_b$in0[15] ),
    .B(_119_),
    .Y(_120_));
 sky130_fd_sc_hs__and2_1 _338_ (.A(_119_),
    .B(\dpath.a_lt_b$in0[15] ),
    .X(_121_));
 sky130_fd_sc_hs__nor2_4 _339_ (.A(_120_),
    .B(_121_),
    .Y(_122_));
 sky130_fd_sc_hs__nand2_1 _340_ (.A(_118_),
    .B(_122_),
    .Y(_123_));
 sky130_fd_sc_hs__inv_1 _341_ (.A(_122_),
    .Y(_124_));
 sky130_fd_sc_hs__nand3_1 _342_ (.A(_114_),
    .B(_117_),
    .C(_124_),
    .Y(_125_));
 sky130_fd_sc_hs__and2_2 _343_ (.A(_123_),
    .B(_125_),
    .X(resp_msg[15]));
 sky130_fd_sc_hs__xnor2_4 _344_ (.A(\dpath.a_lt_b$in1[1] ),
    .B(\dpath.a_lt_b$in0[1] ),
    .Y(_126_));
 sky130_fd_sc_hs__xnor2_4 _345_ (.A(_035_),
    .B(_126_),
    .Y(resp_msg[1]));
 sky130_fd_sc_hs__xnor2_4 _346_ (.A(_045_),
    .B(net2),
    .Y(resp_msg[2]));
 sky130_fd_sc_hs__a21boi_2 _347_ (.A1(_039_),
    .A2(_044_),
    .B1_N(_043_),
    .Y(_127_));
 sky130_fd_sc_hs__xor2_4 _348_ (.A(net11),
    .B(_127_),
    .X(resp_msg[3]));
 sky130_fd_sc_hs__xor2_4 _349_ (.A(_062_),
    .B(net7),
    .X(resp_msg[4]));
 sky130_fd_sc_hs__nand2_1 _350_ (.A(_051_),
    .B(_062_),
    .Y(_128_));
 sky130_fd_sc_hs__nand2_2 _351_ (.A(_128_),
    .B(_070_),
    .Y(_129_));
 sky130_fd_sc_hs__xor2_4 _352_ (.A(_061_),
    .B(_129_),
    .X(resp_msg[5]));
 sky130_fd_sc_hs__nand3_1 _353_ (.A(_051_),
    .B(_061_),
    .C(_062_),
    .Y(_130_));
 sky130_fd_sc_hs__nand2_2 _354_ (.A(_130_),
    .B(_072_),
    .Y(_131_));
 sky130_fd_sc_hs__xor2_4 _355_ (.A(_056_),
    .B(_131_),
    .X(resp_msg[6]));
 sky130_fd_sc_hs__nand2_1 _356_ (.A(_131_),
    .B(net8),
    .Y(_132_));
 sky130_fd_sc_hs__nand2_2 _357_ (.A(_132_),
    .B(_067_),
    .Y(_133_));
 sky130_fd_sc_hs__xor2_4 _358_ (.A(_055_),
    .B(_133_),
    .X(resp_msg[7]));
 sky130_fd_sc_hs__xnor2_4 _359_ (.A(_082_),
    .B(_075_),
    .Y(resp_msg[8]));
 sky130_fd_sc_hs__nand3_1 _360_ (.A(_075_),
    .B(_079_),
    .C(_081_),
    .Y(_134_));
 sky130_fd_sc_hs__nand2_1 _361_ (.A(_134_),
    .B(_079_),
    .Y(_135_));
 sky130_fd_sc_hs__xnor2_4 _362_ (.A(_077_),
    .B(_135_),
    .Y(resp_msg[9]));
 sky130_fd_sc_hs__nor2_1 _363_ (.A(_082_),
    .B(_077_),
    .Y(_136_));
 sky130_fd_sc_hs__nand2_1 _364_ (.A(_075_),
    .B(_136_),
    .Y(_137_));
 sky130_fd_sc_hs__nand2_4 _365_ (.A(_137_),
    .B(_095_),
    .Y(_138_));
 sky130_fd_sc_hs__xor2_4 _366_ (.A(_083_),
    .B(_138_),
    .X(resp_msg[10]));
 sky130_fd_sc_hs__nand2_1 _367_ (.A(_138_),
    .B(_083_),
    .Y(_139_));
 sky130_fd_sc_hs__nand2_2 _368_ (.A(_139_),
    .B(_092_),
    .Y(_140_));
 sky130_fd_sc_hs__xnor2_4 _369_ (.A(_093_),
    .B(_140_),
    .Y(resp_msg[11]));
 sky130_fd_sc_hs__xnor2_4 _370_ (.A(_103_),
    .B(_098_),
    .Y(resp_msg[12]));
 sky130_fd_sc_hs__inv_1 _371_ (.A(_103_),
    .Y(_141_));
 sky130_fd_sc_hs__nand2_1 _372_ (.A(net5),
    .B(_141_),
    .Y(_142_));
 sky130_fd_sc_hs__nand2_2 _373_ (.A(_142_),
    .B(_101_),
    .Y(_143_));
 sky130_fd_sc_hs__xnor2_4 _374_ (.A(_108_),
    .B(_143_),
    .Y(resp_msg[13]));
 sky130_fd_sc_hs__xor2_4 _375_ (.A(_113_),
    .B(net10),
    .X(resp_msg[14]));
 sky130_fd_sc_hs__inv_2 _376_ (.A(\dpath.a_lt_b$in1[0] ),
    .Y(_144_));
 sky130_fd_sc_hs__xnor2_4 _377_ (.A(\dpath.a_lt_b$in0[0] ),
    .B(_144_),
    .Y(resp_msg[0]));
 sky130_fd_sc_hs__clkinv_1 _378_ (.A(\ctrl.state.out[2] ),
    .Y(_145_));
 sky130_fd_sc_hs__nor2_1 _379_ (.A(reset),
    .B(_145_),
    .Y(_146_));
 sky130_fd_sc_hs__nor4_4 _380_ (.A(\dpath.a_lt_b$in1[12] ),
    .B(\dpath.a_lt_b$in1[13] ),
    .C(\dpath.a_lt_b$in1[14] ),
    .D(\dpath.a_lt_b$in1[15] ),
    .Y(_147_));
 sky130_fd_sc_hs__nor4_4 _381_ (.A(\dpath.a_lt_b$in1[8] ),
    .B(\dpath.a_lt_b$in1[9] ),
    .C(\dpath.a_lt_b$in1[10] ),
    .D(\dpath.a_lt_b$in1[11] ),
    .Y(_148_));
 sky130_fd_sc_hs__nor4_4 _382_ (.A(\dpath.a_lt_b$in1[4] ),
    .B(net9),
    .C(\dpath.a_lt_b$in1[6] ),
    .D(net6),
    .Y(_149_));
 sky130_fd_sc_hs__nor4_4 _383_ (.A(net3),
    .B(net1),
    .C(\dpath.a_lt_b$in1[0] ),
    .D(\dpath.a_lt_b$in1[1] ),
    .Y(_150_));
 sky130_fd_sc_hs__nand4_4 _384_ (.A(_147_),
    .B(_148_),
    .C(_149_),
    .D(_150_),
    .Y(_151_));
 sky130_fd_sc_hs__tap_1 TAP_8 ();
 sky130_fd_sc_hs__tap_1 TAP_7 ();
 sky130_fd_sc_hs__nand2_1 _387_ (.A(req_rdy),
    .B(req_val),
    .Y(_154_));
 sky130_fd_sc_hs__o2bb2ai_1 _388_ (.A1_N(_146_),
    .A2_N(_151_),
    .B1(reset),
    .B2(_154_),
    .Y(_002_));
 sky130_fd_sc_hs__nor2_8 _389_ (.A(\ctrl.state.out[2] ),
    .B(req_rdy),
    .Y(_155_));
 sky130_fd_sc_hs__and2_1 _390_ (.A(_155_),
    .B(\ctrl.state.out[1] ),
    .X(resp_val));
 sky130_fd_sc_hs__clkinv_4 _391_ (.A(req_rdy),
    .Y(_156_));
 sky130_fd_sc_hs__a21oi_1 _392_ (.A1(resp_val),
    .A2(resp_rdy),
    .B1(reset),
    .Y(_157_));
 sky130_fd_sc_hs__o21ai_1 _393_ (.A1(_156_),
    .A2(req_val),
    .B1(_157_),
    .Y(_000_));
 sky130_fd_sc_hs__nand2_1 _394_ (.A(_157_),
    .B(\ctrl.state.out[1] ),
    .Y(_158_));
 sky130_fd_sc_hs__o31ai_1 _395_ (.A1(_145_),
    .A2(reset),
    .A3(_151_),
    .B1(_158_),
    .Y(_001_));
 sky130_fd_sc_hs__or2_1 _396_ (.A(_094_),
    .B(_096_),
    .X(_159_));
 sky130_fd_sc_hs__nand2_2 _397_ (.A(_122_),
    .B(_113_),
    .Y(_160_));
 sky130_fd_sc_hs__nor3_4 _398_ (.A(_103_),
    .B(_160_),
    .C(_108_),
    .Y(_161_));
 sky130_fd_sc_hs__a21oi_1 _399_ (.A1(_122_),
    .A2(_116_),
    .B1(_121_),
    .Y(_162_));
 sky130_fd_sc_hs__o21ai_1 _400_ (.A1(_160_),
    .A2(_111_),
    .B1(_162_),
    .Y(_163_));
 sky130_fd_sc_hs__a21oi_4 _401_ (.A1(_159_),
    .A2(_161_),
    .B1(_163_),
    .Y(_164_));
 sky130_fd_sc_hs__nand3_4 _402_ (.A(net4),
    .B(_161_),
    .C(_089_),
    .Y(_165_));
 sky130_fd_sc_hs__nand2_4 _403_ (.A(_164_),
    .B(_165_),
    .Y(_166_));
 sky130_fd_sc_hs__nor2_2 _404_ (.A(_145_),
    .B(_166_),
    .Y(_167_));
 sky130_fd_sc_hs__nor2_8 _405_ (.A(req_rdy),
    .B(_167_),
    .Y(_168_));
 sky130_fd_sc_hs__inv_8 _406_ (.A(_168_),
    .Y(_169_));
 sky130_fd_sc_hs__tap_1 TAP_6 ();
 sky130_fd_sc_hs__nand2_4 _408_ (.A(_156_),
    .B(\ctrl.state.out[2] ),
    .Y(_171_));
 sky130_fd_sc_hs__nor2_8 _409_ (.A(_171_),
    .B(_166_),
    .Y(_172_));
 sky130_fd_sc_hs__tap_1 TAP_5 ();
 sky130_fd_sc_hs__a22oi_1 _411_ (.A1(req_rdy),
    .A2(req_msg[0]),
    .B1(_172_),
    .B2(\dpath.a_lt_b$in0[0] ),
    .Y(_174_));
 sky130_fd_sc_hs__o21ai_1 _412_ (.A1(_144_),
    .A2(_169_),
    .B1(_174_),
    .Y(_003_));
 sky130_fd_sc_hs__a22oi_1 _413_ (.A1(req_rdy),
    .A2(req_msg[1]),
    .B1(_172_),
    .B2(\dpath.a_lt_b$in0[1] ),
    .Y(_175_));
 sky130_fd_sc_hs__o21ai_1 _414_ (.A1(_037_),
    .A2(_169_),
    .B1(_175_),
    .Y(_004_));
 sky130_fd_sc_hs__inv_1 _415_ (.A(\dpath.a_lt_b$in1[2] ),
    .Y(_176_));
 sky130_fd_sc_hs__a22oi_1 _416_ (.A1(req_rdy),
    .A2(req_msg[2]),
    .B1(_172_),
    .B2(\dpath.a_lt_b$in0[2] ),
    .Y(_177_));
 sky130_fd_sc_hs__o21ai_1 _417_ (.A1(_176_),
    .A2(_169_),
    .B1(_177_),
    .Y(_005_));
 sky130_fd_sc_hs__tap_1 TAP_4 ();
 sky130_fd_sc_hs__a22oi_1 _419_ (.A1(req_rdy),
    .A2(req_msg[3]),
    .B1(_172_),
    .B2(\dpath.a_lt_b$in0[3] ),
    .Y(_179_));
 sky130_fd_sc_hs__o21ai_1 _420_ (.A1(_048_),
    .A2(_169_),
    .B1(_179_),
    .Y(_006_));
 sky130_fd_sc_hs__a22oi_1 _421_ (.A1(req_rdy),
    .A2(req_msg[4]),
    .B1(_172_),
    .B2(\dpath.a_lt_b$in0[4] ),
    .Y(_180_));
 sky130_fd_sc_hs__o21ai_1 _422_ (.A1(_069_),
    .A2(_169_),
    .B1(_180_),
    .Y(_007_));
 sky130_fd_sc_hs__a22oi_1 _423_ (.A1(req_rdy),
    .A2(req_msg[5]),
    .B1(_172_),
    .B2(\dpath.a_lt_b$in0[5] ),
    .Y(_181_));
 sky130_fd_sc_hs__o21ai_1 _424_ (.A1(_058_),
    .A2(_169_),
    .B1(_181_),
    .Y(_008_));
 sky130_fd_sc_hs__a22oi_1 _425_ (.A1(req_rdy),
    .A2(req_msg[6]),
    .B1(_172_),
    .B2(\dpath.a_lt_b$in0[6] ),
    .Y(_182_));
 sky130_fd_sc_hs__o21ai_1 _426_ (.A1(_066_),
    .A2(_169_),
    .B1(_182_),
    .Y(_009_));
 sky130_fd_sc_hs__a22oi_1 _427_ (.A1(req_rdy),
    .A2(req_msg[7]),
    .B1(_172_),
    .B2(\dpath.a_lt_b$in0[7] ),
    .Y(_183_));
 sky130_fd_sc_hs__o21ai_1 _428_ (.A1(_052_),
    .A2(_169_),
    .B1(_183_),
    .Y(_010_));
 sky130_fd_sc_hs__nor2_1 _429_ (.A(req_msg[8]),
    .B(_156_),
    .Y(_184_));
 sky130_fd_sc_hs__a21oi_1 _430_ (.A1(_156_),
    .A2(_080_),
    .B1(_184_),
    .Y(_185_));
 sky130_fd_sc_hs__nor2_1 _431_ (.A(_185_),
    .B(_168_),
    .Y(_186_));
 sky130_fd_sc_hs__a21oi_1 _432_ (.A1(_078_),
    .A2(_168_),
    .B1(_186_),
    .Y(_011_));
 sky130_fd_sc_hs__nand2_1 _433_ (.A(_168_),
    .B(\dpath.a_lt_b$in1[9] ),
    .Y(_187_));
 sky130_fd_sc_hs__nor2_1 _434_ (.A(req_msg[9]),
    .B(_156_),
    .Y(_188_));
 sky130_fd_sc_hs__a21oi_1 _435_ (.A1(_156_),
    .A2(_076_),
    .B1(_188_),
    .Y(_189_));
 sky130_fd_sc_hs__nand2_1 _436_ (.A(_169_),
    .B(_189_),
    .Y(_190_));
 sky130_fd_sc_hs__nand2_1 _437_ (.A(_187_),
    .B(_190_),
    .Y(_012_));
 sky130_fd_sc_hs__a22oi_1 _438_ (.A1(req_rdy),
    .A2(req_msg[10]),
    .B1(_172_),
    .B2(\dpath.a_lt_b$in0[10] ),
    .Y(_191_));
 sky130_fd_sc_hs__o21ai_1 _439_ (.A1(_091_),
    .A2(_169_),
    .B1(_191_),
    .Y(_013_));
 sky130_fd_sc_hs__nor2_1 _440_ (.A(req_msg[11]),
    .B(_156_),
    .Y(_192_));
 sky130_fd_sc_hs__a21oi_1 _441_ (.A1(_156_),
    .A2(_086_),
    .B1(_192_),
    .Y(_193_));
 sky130_fd_sc_hs__nor2_1 _442_ (.A(_193_),
    .B(_168_),
    .Y(_194_));
 sky130_fd_sc_hs__a21oi_1 _443_ (.A1(_084_),
    .A2(_168_),
    .B1(_194_),
    .Y(_014_));
 sky130_fd_sc_hs__tap_1 TAP_3 ();
 sky130_fd_sc_hs__a22oi_1 _445_ (.A1(req_rdy),
    .A2(req_msg[12]),
    .B1(_172_),
    .B2(\dpath.a_lt_b$in0[12] ),
    .Y(_196_));
 sky130_fd_sc_hs__nand2_1 _446_ (.A(_168_),
    .B(\dpath.a_lt_b$in1[12] ),
    .Y(_197_));
 sky130_fd_sc_hs__nand2_1 _447_ (.A(_196_),
    .B(_197_),
    .Y(_015_));
 sky130_fd_sc_hs__a22oi_1 _448_ (.A1(req_rdy),
    .A2(req_msg[13]),
    .B1(_172_),
    .B2(\dpath.a_lt_b$in0[13] ),
    .Y(_198_));
 sky130_fd_sc_hs__o21ai_1 _449_ (.A1(_104_),
    .A2(_169_),
    .B1(_198_),
    .Y(_016_));
 sky130_fd_sc_hs__a22oi_1 _450_ (.A1(req_rdy),
    .A2(req_msg[14]),
    .B1(_172_),
    .B2(\dpath.a_lt_b$in0[14] ),
    .Y(_199_));
 sky130_fd_sc_hs__nand2_1 _451_ (.A(_168_),
    .B(\dpath.a_lt_b$in1[14] ),
    .Y(_200_));
 sky130_fd_sc_hs__nand2_1 _452_ (.A(_199_),
    .B(_200_),
    .Y(_017_));
 sky130_fd_sc_hs__a22oi_1 _453_ (.A1(req_rdy),
    .A2(req_msg[15]),
    .B1(_172_),
    .B2(\dpath.a_lt_b$in0[15] ),
    .Y(_201_));
 sky130_fd_sc_hs__o21ai_1 _454_ (.A1(_119_),
    .A2(_169_),
    .B1(_201_),
    .Y(_018_));
 sky130_fd_sc_hs__inv_4 _455_ (.A(_172_),
    .Y(_202_));
 sky130_fd_sc_hs__a21oi_4 _456_ (.A1(_164_),
    .A2(_165_),
    .B1(_171_),
    .Y(_203_));
 sky130_fd_sc_hs__tap_1 TAP_2 ();
 sky130_fd_sc_hs__nand2_1 _458_ (.A(_203_),
    .B(resp_msg[0]),
    .Y(_205_));
 sky130_fd_sc_hs__tap_1 TAP_1 ();
 sky130_fd_sc_hs__a22oi_1 _460_ (.A1(req_rdy),
    .A2(req_msg[16]),
    .B1(_155_),
    .B2(\dpath.a_lt_b$in0[0] ),
    .Y(_207_));
 sky130_fd_sc_hs__o211ai_1 _461_ (.A1(_144_),
    .A2(_202_),
    .B1(_205_),
    .C1(_207_),
    .Y(_019_));
 sky130_fd_sc_hs__nand2_1 _462_ (.A(_203_),
    .B(resp_msg[1]),
    .Y(_208_));
 sky130_fd_sc_hs__nand2_1 _463_ (.A(_172_),
    .B(\dpath.a_lt_b$in1[1] ),
    .Y(_209_));
 sky130_fd_sc_hs__nand2_1 _464_ (.A(_155_),
    .B(\dpath.a_lt_b$in0[1] ),
    .Y(_210_));
 sky130_fd_sc_hs__nand2_1 _465_ (.A(req_rdy),
    .B(req_msg[17]),
    .Y(_211_));
 sky130_fd_sc_hs__nand4_1 _466_ (.A(_208_),
    .B(_209_),
    .C(_210_),
    .D(_211_),
    .Y(_020_));
 sky130_fd_sc_hs__nand2_1 _467_ (.A(_203_),
    .B(resp_msg[2]),
    .Y(_212_));
 sky130_fd_sc_hs__tap_1 TAP_0 ();
 sky130_fd_sc_hs__a22oi_1 _469_ (.A1(req_msg[18]),
    .A2(req_rdy),
    .B1(_155_),
    .B2(\dpath.a_lt_b$in0[2] ),
    .Y(_214_));
 sky130_fd_sc_hs__o211ai_1 _470_ (.A1(_176_),
    .A2(_202_),
    .B1(_212_),
    .C1(_214_),
    .Y(_021_));
 sky130_fd_sc_hs__nand2_1 _471_ (.A(_203_),
    .B(resp_msg[3]),
    .Y(_215_));
 sky130_fd_sc_hs__a22oi_1 _472_ (.A1(req_msg[19]),
    .A2(req_rdy),
    .B1(_155_),
    .B2(\dpath.a_lt_b$in0[3] ),
    .Y(_216_));
 sky130_fd_sc_hs__o211ai_1 _473_ (.A1(_048_),
    .A2(_202_),
    .B1(_215_),
    .C1(_216_),
    .Y(_022_));
 sky130_fd_sc_hs__nand2_1 _474_ (.A(_203_),
    .B(resp_msg[4]),
    .Y(_217_));
 sky130_fd_sc_hs__a22oi_1 _475_ (.A1(req_msg[20]),
    .A2(req_rdy),
    .B1(_155_),
    .B2(\dpath.a_lt_b$in0[4] ),
    .Y(_218_));
 sky130_fd_sc_hs__o211ai_1 _476_ (.A1(_069_),
    .A2(_202_),
    .B1(_217_),
    .C1(_218_),
    .Y(_023_));
 sky130_fd_sc_hs__nand2_1 _477_ (.A(_203_),
    .B(resp_msg[5]),
    .Y(_219_));
 sky130_fd_sc_hs__a22oi_1 _478_ (.A1(req_msg[21]),
    .A2(req_rdy),
    .B1(_155_),
    .B2(\dpath.a_lt_b$in0[5] ),
    .Y(_220_));
 sky130_fd_sc_hs__o211ai_1 _479_ (.A1(_058_),
    .A2(_202_),
    .B1(_219_),
    .C1(_220_),
    .Y(_024_));
 sky130_fd_sc_hs__nand2_1 _480_ (.A(_203_),
    .B(resp_msg[6]),
    .Y(_221_));
 sky130_fd_sc_hs__a22oi_1 _481_ (.A1(req_msg[22]),
    .A2(req_rdy),
    .B1(_155_),
    .B2(\dpath.a_lt_b$in0[6] ),
    .Y(_222_));
 sky130_fd_sc_hs__o211ai_1 _482_ (.A1(_066_),
    .A2(_202_),
    .B1(_221_),
    .C1(_222_),
    .Y(_025_));
 sky130_fd_sc_hs__a22oi_1 _483_ (.A1(req_msg[23]),
    .A2(req_rdy),
    .B1(_155_),
    .B2(\dpath.a_lt_b$in0[7] ),
    .Y(_223_));
 sky130_fd_sc_hs__nand2_1 _484_ (.A(resp_msg[7]),
    .B(_203_),
    .Y(_224_));
 sky130_fd_sc_hs__o211ai_1 _485_ (.A1(_052_),
    .A2(_202_),
    .B1(_223_),
    .C1(_224_),
    .Y(_026_));
 sky130_fd_sc_hs__nand2_1 _486_ (.A(_203_),
    .B(resp_msg[8]),
    .Y(_225_));
 sky130_fd_sc_hs__nand2_1 _487_ (.A(_172_),
    .B(\dpath.a_lt_b$in1[8] ),
    .Y(_226_));
 sky130_fd_sc_hs__nand2_4 _488_ (.A(req_msg[24]),
    .B(req_rdy),
    .Y(_227_));
 sky130_fd_sc_hs__nand2_1 _489_ (.A(_155_),
    .B(\dpath.a_lt_b$in0[8] ),
    .Y(_228_));
 sky130_fd_sc_hs__nand4_1 _490_ (.A(_225_),
    .B(_226_),
    .C(_227_),
    .D(_228_),
    .Y(_027_));
 sky130_fd_sc_hs__nand2_1 _491_ (.A(resp_msg[9]),
    .B(_203_),
    .Y(_229_));
 sky130_fd_sc_hs__nand2_1 _492_ (.A(_172_),
    .B(\dpath.a_lt_b$in1[9] ),
    .Y(_230_));
 sky130_fd_sc_hs__nand2_1 _493_ (.A(req_msg[25]),
    .B(req_rdy),
    .Y(_231_));
 sky130_fd_sc_hs__nand2_1 _494_ (.A(_155_),
    .B(\dpath.a_lt_b$in0[9] ),
    .Y(_232_));
 sky130_fd_sc_hs__nand4_1 _495_ (.A(_229_),
    .B(_230_),
    .C(_231_),
    .D(_232_),
    .Y(_028_));
 sky130_fd_sc_hs__nand2_1 _496_ (.A(_203_),
    .B(resp_msg[10]),
    .Y(_233_));
 sky130_fd_sc_hs__a22oi_1 _497_ (.A1(req_msg[26]),
    .A2(req_rdy),
    .B1(_155_),
    .B2(\dpath.a_lt_b$in0[10] ),
    .Y(_234_));
 sky130_fd_sc_hs__o211ai_1 _498_ (.A1(_091_),
    .A2(_202_),
    .B1(_233_),
    .C1(_234_),
    .Y(_029_));
 sky130_fd_sc_hs__nand2_1 _499_ (.A(resp_msg[11]),
    .B(_203_),
    .Y(_235_));
 sky130_fd_sc_hs__nand2_1 _500_ (.A(_172_),
    .B(\dpath.a_lt_b$in1[11] ),
    .Y(_236_));
 sky130_fd_sc_hs__nor3_1 _501_ (.A(\ctrl.state.out[2] ),
    .B(req_rdy),
    .C(_086_),
    .Y(_237_));
 sky130_fd_sc_hs__a21oi_1 _502_ (.A1(req_msg[27]),
    .A2(req_rdy),
    .B1(_237_),
    .Y(_238_));
 sky130_fd_sc_hs__nand3_1 _503_ (.A(_235_),
    .B(_236_),
    .C(_238_),
    .Y(_030_));
 sky130_fd_sc_hs__nand2_1 _504_ (.A(_203_),
    .B(resp_msg[12]),
    .Y(_239_));
 sky130_fd_sc_hs__nand2_1 _505_ (.A(_172_),
    .B(\dpath.a_lt_b$in1[12] ),
    .Y(_240_));
 sky130_fd_sc_hs__nand2_1 _506_ (.A(_155_),
    .B(\dpath.a_lt_b$in0[12] ),
    .Y(_241_));
 sky130_fd_sc_hs__nand2_2 _507_ (.A(req_msg[28]),
    .B(req_rdy),
    .Y(_242_));
 sky130_fd_sc_hs__nand4_1 _508_ (.A(_239_),
    .B(_240_),
    .C(_241_),
    .D(_242_),
    .Y(_031_));
 sky130_fd_sc_hs__nand2_1 _509_ (.A(resp_msg[13]),
    .B(_203_),
    .Y(_243_));
 sky130_fd_sc_hs__nand2_1 _510_ (.A(_172_),
    .B(\dpath.a_lt_b$in1[13] ),
    .Y(_244_));
 sky130_fd_sc_hs__a22oi_1 _511_ (.A1(req_msg[29]),
    .A2(req_rdy),
    .B1(_155_),
    .B2(\dpath.a_lt_b$in0[13] ),
    .Y(_245_));
 sky130_fd_sc_hs__nand3_1 _512_ (.A(_243_),
    .B(_244_),
    .C(_245_),
    .Y(_032_));
 sky130_fd_sc_hs__nand2_1 _513_ (.A(resp_msg[14]),
    .B(_203_),
    .Y(_246_));
 sky130_fd_sc_hs__nand2_1 _514_ (.A(_172_),
    .B(\dpath.a_lt_b$in1[14] ),
    .Y(_247_));
 sky130_fd_sc_hs__a22oi_1 _515_ (.A1(req_msg[30]),
    .A2(req_rdy),
    .B1(_155_),
    .B2(\dpath.a_lt_b$in0[14] ),
    .Y(_248_));
 sky130_fd_sc_hs__nand3_1 _516_ (.A(_246_),
    .B(_247_),
    .C(_248_),
    .Y(_033_));
 sky130_fd_sc_hs__nand3_1 _517_ (.A(net12),
    .B(_125_),
    .C(_203_),
    .Y(_249_));
 sky130_fd_sc_hs__a22o_1 _518_ (.A1(req_msg[31]),
    .A2(req_rdy),
    .B1(_155_),
    .B2(\dpath.a_lt_b$in0[15] ),
    .X(_250_));
 sky130_fd_sc_hs__a21oi_1 _519_ (.A1(_172_),
    .A2(\dpath.a_lt_b$in1[15] ),
    .B1(_250_),
    .Y(_251_));
 sky130_fd_sc_hs__nand2_1 _520_ (.A(_249_),
    .B(_251_),
    .Y(_034_));
 sky130_fd_sc_hs__dfxtp_4 _521_ (.D(_000_),
    .Q(req_rdy),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hs__dfxtp_1 _522_ (.D(_001_),
    .Q(\ctrl.state.out[1] ),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hs__dfxtp_4 _523_ (.D(_002_),
    .Q(\ctrl.state.out[2] ),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _524_ (.D(_003_),
    .Q(\dpath.a_lt_b$in1[0] ),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hs__dfxtp_4 _525_ (.D(_004_),
    .Q(\dpath.a_lt_b$in1[1] ),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _526_ (.D(_005_),
    .Q(\dpath.a_lt_b$in1[2] ),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _527_ (.D(_006_),
    .Q(\dpath.a_lt_b$in1[3] ),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hs__dfxtp_4 _528_ (.D(_007_),
    .Q(\dpath.a_lt_b$in1[4] ),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _529_ (.D(_008_),
    .Q(\dpath.a_lt_b$in1[5] ),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _530_ (.D(_009_),
    .Q(\dpath.a_lt_b$in1[6] ),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _531_ (.D(_010_),
    .Q(\dpath.a_lt_b$in1[7] ),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _532_ (.D(_011_),
    .Q(\dpath.a_lt_b$in1[8] ),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _533_ (.D(_012_),
    .Q(\dpath.a_lt_b$in1[9] ),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _534_ (.D(_013_),
    .Q(\dpath.a_lt_b$in1[10] ),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _535_ (.D(_014_),
    .Q(\dpath.a_lt_b$in1[11] ),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _536_ (.D(_015_),
    .Q(\dpath.a_lt_b$in1[12] ),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hs__dfxtp_1 _537_ (.D(_016_),
    .Q(\dpath.a_lt_b$in1[13] ),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _538_ (.D(_017_),
    .Q(\dpath.a_lt_b$in1[14] ),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _539_ (.D(_018_),
    .Q(\dpath.a_lt_b$in1[15] ),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _540_ (.D(_019_),
    .Q(\dpath.a_lt_b$in0[0] ),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _541_ (.D(_020_),
    .Q(\dpath.a_lt_b$in0[1] ),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _542_ (.D(_021_),
    .Q(\dpath.a_lt_b$in0[2] ),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _543_ (.D(_022_),
    .Q(\dpath.a_lt_b$in0[3] ),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _544_ (.D(_023_),
    .Q(\dpath.a_lt_b$in0[4] ),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _545_ (.D(_024_),
    .Q(\dpath.a_lt_b$in0[5] ),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _546_ (.D(_025_),
    .Q(\dpath.a_lt_b$in0[6] ),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hs__dfxtp_1 _547_ (.D(_026_),
    .Q(\dpath.a_lt_b$in0[7] ),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hs__dfxtp_1 _548_ (.D(_027_),
    .Q(\dpath.a_lt_b$in0[8] ),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hs__dfxtp_1 _549_ (.D(_028_),
    .Q(\dpath.a_lt_b$in0[9] ),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _550_ (.D(_029_),
    .Q(\dpath.a_lt_b$in0[10] ),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hs__dfxtp_1 _551_ (.D(_030_),
    .Q(\dpath.a_lt_b$in0[11] ),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hs__dfxtp_1 _552_ (.D(_031_),
    .Q(\dpath.a_lt_b$in0[12] ),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hs__dfxtp_1 _553_ (.D(_032_),
    .Q(\dpath.a_lt_b$in0[13] ),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _554_ (.D(_033_),
    .Q(\dpath.a_lt_b$in0[14] ),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hs__dfxtp_1 _555_ (.D(_034_),
    .Q(\dpath.a_lt_b$in0[15] ),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hs__tap_1 TAP_9 ();
 sky130_fd_sc_hs__tap_1 TAP_10 ();
 sky130_fd_sc_hs__tap_1 TAP_11 ();
 sky130_fd_sc_hs__tap_1 TAP_12 ();
 sky130_fd_sc_hs__tap_1 TAP_13 ();
 sky130_fd_sc_hs__tap_1 TAP_14 ();
 sky130_fd_sc_hs__tap_1 TAP_15 ();
 sky130_fd_sc_hs__tap_1 TAP_16 ();
 sky130_fd_sc_hs__tap_1 TAP_17 ();
 sky130_fd_sc_hs__tap_1 TAP_18 ();
 sky130_fd_sc_hs__tap_1 TAP_19 ();
 sky130_fd_sc_hs__tap_1 TAP_20 ();
 sky130_fd_sc_hs__tap_1 TAP_21 ();
 sky130_fd_sc_hs__tap_1 TAP_22 ();
 sky130_fd_sc_hs__tap_1 TAP_23 ();
 sky130_fd_sc_hs__tap_1 TAP_24 ();
 sky130_fd_sc_hs__tap_1 TAP_25 ();
 sky130_fd_sc_hs__tap_1 TAP_26 ();
 sky130_fd_sc_hs__tap_1 TAP_27 ();
 sky130_fd_sc_hs__tap_1 TAP_28 ();
 sky130_fd_sc_hs__tap_1 TAP_29 ();
 sky130_fd_sc_hs__tap_1 TAP_30 ();
 sky130_fd_sc_hs__tap_1 TAP_31 ();
 sky130_fd_sc_hs__tap_1 TAP_32 ();
 sky130_fd_sc_hs__tap_1 TAP_33 ();
 sky130_fd_sc_hs__tap_1 TAP_34 ();
 sky130_fd_sc_hs__tap_1 TAP_35 ();
 sky130_fd_sc_hs__tap_1 TAP_36 ();
 sky130_fd_sc_hs__tap_1 TAP_37 ();
 sky130_fd_sc_hs__tap_1 TAP_38 ();
 sky130_fd_sc_hs__tap_1 TAP_39 ();
 sky130_fd_sc_hs__tap_1 TAP_40 ();
 sky130_fd_sc_hs__tap_1 TAP_41 ();
 sky130_fd_sc_hs__tap_1 TAP_42 ();
 sky130_fd_sc_hs__tap_1 TAP_43 ();
 sky130_fd_sc_hs__tap_1 TAP_44 ();
 sky130_fd_sc_hs__tap_1 TAP_45 ();
 sky130_fd_sc_hs__tap_1 TAP_46 ();
 sky130_fd_sc_hs__tap_1 TAP_47 ();
 sky130_fd_sc_hs__tap_1 TAP_48 ();
 sky130_fd_sc_hs__tap_1 TAP_49 ();
 sky130_fd_sc_hs__tap_1 TAP_50 ();
 sky130_fd_sc_hs__tap_1 TAP_51 ();
 sky130_fd_sc_hs__tap_1 TAP_52 ();
 sky130_fd_sc_hs__tap_1 TAP_53 ();
 sky130_fd_sc_hs__tap_1 TAP_54 ();
 sky130_fd_sc_hs__tap_1 TAP_55 ();
 sky130_fd_sc_hs__tap_1 TAP_56 ();
 sky130_fd_sc_hs__tap_1 TAP_57 ();
 sky130_fd_sc_hs__tap_1 TAP_58 ();
 sky130_fd_sc_hs__tap_1 TAP_59 ();
 sky130_fd_sc_hs__tap_1 TAP_60 ();
 sky130_fd_sc_hs__tap_1 TAP_61 ();
 sky130_fd_sc_hs__tap_1 TAP_62 ();
 sky130_fd_sc_hs__tap_1 TAP_63 ();
 sky130_fd_sc_hs__tap_1 TAP_64 ();
 sky130_fd_sc_hs__tap_1 TAP_65 ();
 sky130_fd_sc_hs__tap_1 TAP_66 ();
 sky130_fd_sc_hs__tap_1 TAP_67 ();
 sky130_fd_sc_hs__tap_1 TAP_68 ();
 sky130_fd_sc_hs__tap_1 TAP_69 ();
 sky130_fd_sc_hs__tap_1 TAP_70 ();
 sky130_fd_sc_hs__tap_1 TAP_71 ();
 sky130_fd_sc_hs__tap_1 TAP_72 ();
 sky130_fd_sc_hs__tap_1 TAP_73 ();
 sky130_fd_sc_hs__tap_1 TAP_74 ();
 sky130_fd_sc_hs__tap_1 TAP_75 ();
 sky130_fd_sc_hs__tap_1 TAP_76 ();
 sky130_fd_sc_hs__tap_1 TAP_77 ();
 sky130_fd_sc_hs__tap_1 TAP_78 ();
 sky130_fd_sc_hs__tap_1 TAP_79 ();
 sky130_fd_sc_hs__tap_1 TAP_80 ();
 sky130_fd_sc_hs__tap_1 TAP_81 ();
 sky130_fd_sc_hs__tap_1 TAP_82 ();
 sky130_fd_sc_hs__tap_1 TAP_83 ();
 sky130_fd_sc_hs__tap_1 TAP_84 ();
 sky130_fd_sc_hs__tap_1 TAP_85 ();
 sky130_fd_sc_hs__tap_1 TAP_86 ();
 sky130_fd_sc_hs__tap_1 TAP_87 ();
 sky130_fd_sc_hs__tap_1 TAP_88 ();
 sky130_fd_sc_hs__tap_1 TAP_89 ();
 sky130_fd_sc_hs__tap_1 TAP_90 ();
 sky130_fd_sc_hs__tap_1 TAP_91 ();
 sky130_fd_sc_hs__tap_1 TAP_92 ();
 sky130_fd_sc_hs__tap_1 TAP_93 ();
 sky130_fd_sc_hs__tap_1 TAP_94 ();
 sky130_fd_sc_hs__tap_1 TAP_95 ();
 sky130_fd_sc_hs__tap_1 TAP_96 ();
 sky130_fd_sc_hs__tap_1 TAP_97 ();
 sky130_fd_sc_hs__tap_1 TAP_98 ();
 sky130_fd_sc_hs__tap_1 TAP_99 ();
 sky130_fd_sc_hs__tap_1 TAP_100 ();
 sky130_fd_sc_hs__tap_1 TAP_101 ();
 sky130_fd_sc_hs__tap_1 TAP_102 ();
 sky130_fd_sc_hs__tap_1 TAP_103 ();
 sky130_fd_sc_hs__tap_1 TAP_104 ();
 sky130_fd_sc_hs__tap_1 TAP_105 ();
 sky130_fd_sc_hs__tap_1 TAP_106 ();
 sky130_fd_sc_hs__tap_1 TAP_107 ();
 sky130_fd_sc_hs__tap_1 TAP_108 ();
 sky130_fd_sc_hs__tap_1 TAP_109 ();
 sky130_fd_sc_hs__tap_1 TAP_110 ();
 sky130_fd_sc_hs__tap_1 TAP_111 ();
 sky130_fd_sc_hs__tap_1 TAP_112 ();
 sky130_fd_sc_hs__tap_1 TAP_113 ();
 sky130_fd_sc_hs__tap_1 TAP_114 ();
 sky130_fd_sc_hs__tap_1 TAP_115 ();
 sky130_fd_sc_hs__tap_1 TAP_116 ();
 sky130_fd_sc_hs__tap_1 TAP_117 ();
 sky130_fd_sc_hs__tap_1 TAP_118 ();
 sky130_fd_sc_hs__tap_1 TAP_119 ();
 sky130_fd_sc_hs__tap_1 TAP_120 ();
 sky130_fd_sc_hs__tap_1 TAP_121 ();
 sky130_fd_sc_hs__tap_1 TAP_122 ();
 sky130_fd_sc_hs__tap_1 TAP_123 ();
 sky130_fd_sc_hs__tap_1 TAP_124 ();
 sky130_fd_sc_hs__tap_1 TAP_125 ();
 sky130_fd_sc_hs__tap_1 TAP_126 ();
 sky130_fd_sc_hs__tap_1 TAP_127 ();
 sky130_fd_sc_hs__tap_1 TAP_128 ();
 sky130_fd_sc_hs__tap_1 TAP_129 ();
 sky130_fd_sc_hs__tap_1 TAP_130 ();
 sky130_fd_sc_hs__tap_1 TAP_131 ();
 sky130_fd_sc_hs__tap_1 TAP_132 ();
 sky130_fd_sc_hs__tap_1 TAP_133 ();
 sky130_fd_sc_hs__tap_1 TAP_134 ();
 sky130_fd_sc_hs__tap_1 TAP_135 ();
 sky130_fd_sc_hs__tap_1 TAP_136 ();
 sky130_fd_sc_hs__tap_1 TAP_137 ();
 sky130_fd_sc_hs__tap_1 TAP_138 ();
 sky130_fd_sc_hs__tap_1 TAP_139 ();
 sky130_fd_sc_hs__tap_1 TAP_140 ();
 sky130_fd_sc_hs__tap_1 TAP_141 ();
 sky130_fd_sc_hs__tap_1 TAP_142 ();
 sky130_fd_sc_hs__tap_1 TAP_143 ();
 sky130_fd_sc_hs__tap_1 TAP_144 ();
 sky130_fd_sc_hs__tap_1 TAP_145 ();
 sky130_fd_sc_hs__tap_1 TAP_146 ();
 sky130_fd_sc_hs__tap_1 TAP_147 ();
 sky130_fd_sc_hs__tap_1 TAP_148 ();
 sky130_fd_sc_hs__tap_1 TAP_149 ();
 sky130_fd_sc_hs__tap_1 TAP_150 ();
 sky130_fd_sc_hs__tap_1 TAP_151 ();
 sky130_fd_sc_hs__tap_1 TAP_152 ();
 sky130_fd_sc_hs__tap_1 TAP_153 ();
 sky130_fd_sc_hs__tap_1 TAP_154 ();
 sky130_fd_sc_hs__tap_1 TAP_155 ();
 sky130_fd_sc_hs__tap_1 TAP_156 ();
 sky130_fd_sc_hs__tap_1 TAP_157 ();
 sky130_fd_sc_hs__tap_1 TAP_158 ();
 sky130_fd_sc_hs__tap_1 TAP_159 ();
 sky130_fd_sc_hs__tap_1 TAP_160 ();
 sky130_fd_sc_hs__tap_1 TAP_161 ();
 sky130_fd_sc_hs__tap_1 TAP_162 ();
 sky130_fd_sc_hs__tap_1 TAP_163 ();
 sky130_fd_sc_hs__tap_1 TAP_164 ();
 sky130_fd_sc_hs__tap_1 TAP_165 ();
 sky130_fd_sc_hs__tap_1 TAP_166 ();
 sky130_fd_sc_hs__tap_1 TAP_167 ();
 sky130_fd_sc_hs__tap_1 TAP_168 ();
 sky130_fd_sc_hs__tap_1 TAP_169 ();
 sky130_fd_sc_hs__tap_1 TAP_170 ();
 sky130_fd_sc_hs__tap_1 TAP_171 ();
 sky130_fd_sc_hs__tap_1 TAP_172 ();
 sky130_fd_sc_hs__tap_1 TAP_173 ();
 sky130_fd_sc_hs__tap_1 TAP_174 ();
 sky130_fd_sc_hs__tap_1 TAP_175 ();
 sky130_fd_sc_hs__tap_1 TAP_176 ();
 sky130_fd_sc_hs__tap_1 TAP_177 ();
 sky130_fd_sc_hs__tap_1 TAP_178 ();
 sky130_fd_sc_hs__tap_1 TAP_179 ();
 sky130_fd_sc_hs__tap_1 TAP_180 ();
 sky130_fd_sc_hs__tap_1 TAP_181 ();
 sky130_fd_sc_hs__tap_1 TAP_182 ();
 sky130_fd_sc_hs__tap_1 TAP_183 ();
 sky130_fd_sc_hs__tap_1 TAP_184 ();
 sky130_fd_sc_hs__tap_1 TAP_185 ();
 sky130_fd_sc_hs__tap_1 TAP_186 ();
 sky130_fd_sc_hs__tap_1 TAP_187 ();
 sky130_fd_sc_hs__tap_1 TAP_188 ();
 sky130_fd_sc_hs__tap_1 TAP_189 ();
 sky130_fd_sc_hs__tap_1 TAP_190 ();
 sky130_fd_sc_hs__tap_1 TAP_191 ();
 sky130_fd_sc_hs__tap_1 TAP_192 ();
 sky130_fd_sc_hs__tap_1 TAP_193 ();
 sky130_fd_sc_hs__tap_1 TAP_194 ();
 sky130_fd_sc_hs__tap_1 TAP_195 ();
 sky130_fd_sc_hs__tap_1 TAP_196 ();
 sky130_fd_sc_hs__tap_1 TAP_197 ();
 sky130_fd_sc_hs__tap_1 TAP_198 ();
 sky130_fd_sc_hs__tap_1 TAP_199 ();
 sky130_fd_sc_hs__tap_1 TAP_200 ();
 sky130_fd_sc_hs__tap_1 TAP_201 ();
 sky130_fd_sc_hs__tap_1 TAP_202 ();
 sky130_fd_sc_hs__tap_1 TAP_203 ();
 sky130_fd_sc_hs__tap_1 TAP_204 ();
 sky130_fd_sc_hs__tap_1 TAP_205 ();
 sky130_fd_sc_hs__tap_1 TAP_206 ();
 sky130_fd_sc_hs__tap_1 TAP_207 ();
 sky130_fd_sc_hs__tap_1 TAP_208 ();
 sky130_fd_sc_hs__tap_1 TAP_209 ();
 sky130_fd_sc_hs__tap_1 TAP_210 ();
 sky130_fd_sc_hs__tap_1 TAP_211 ();
 sky130_fd_sc_hs__tap_1 TAP_212 ();
 sky130_fd_sc_hs__tap_1 TAP_213 ();
 sky130_fd_sc_hs__tap_1 TAP_214 ();
 sky130_fd_sc_hs__tap_1 TAP_215 ();
 sky130_fd_sc_hs__tap_1 TAP_216 ();
 sky130_fd_sc_hs__tap_1 TAP_217 ();
 sky130_fd_sc_hs__tap_1 TAP_218 ();
 sky130_fd_sc_hs__tap_1 TAP_219 ();
 sky130_fd_sc_hs__tap_1 TAP_220 ();
 sky130_fd_sc_hs__tap_1 TAP_221 ();
 sky130_fd_sc_hs__tap_1 TAP_222 ();
 sky130_fd_sc_hs__tap_1 TAP_223 ();
 sky130_fd_sc_hs__tap_1 TAP_224 ();
 sky130_fd_sc_hs__tap_1 TAP_225 ();
 sky130_fd_sc_hs__tap_1 TAP_226 ();
 sky130_fd_sc_hs__tap_1 TAP_227 ();
 sky130_fd_sc_hs__tap_1 TAP_228 ();
 sky130_fd_sc_hs__tap_1 TAP_229 ();
 sky130_fd_sc_hs__tap_1 TAP_230 ();
 sky130_fd_sc_hs__tap_1 TAP_231 ();
 sky130_fd_sc_hs__tap_1 TAP_232 ();
 sky130_fd_sc_hs__tap_1 TAP_233 ();
 sky130_fd_sc_hs__tap_1 TAP_234 ();
 sky130_fd_sc_hs__tap_1 TAP_235 ();
 sky130_fd_sc_hs__tap_1 TAP_236 ();
 sky130_fd_sc_hs__tap_1 TAP_237 ();
 sky130_fd_sc_hs__tap_1 TAP_238 ();
 sky130_fd_sc_hs__tap_1 TAP_239 ();
 sky130_fd_sc_hs__tap_1 TAP_240 ();
 sky130_fd_sc_hs__tap_1 TAP_241 ();
 sky130_fd_sc_hs__tap_1 TAP_242 ();
 sky130_fd_sc_hs__tap_1 TAP_243 ();
 sky130_fd_sc_hs__tap_1 TAP_244 ();
 sky130_fd_sc_hs__tap_1 TAP_245 ();
 sky130_fd_sc_hs__tap_1 TAP_246 ();
 sky130_fd_sc_hs__tap_1 TAP_247 ();
 sky130_fd_sc_hs__tap_1 TAP_248 ();
 sky130_fd_sc_hs__tap_1 TAP_249 ();
 sky130_fd_sc_hs__tap_1 TAP_250 ();
 sky130_fd_sc_hs__tap_1 TAP_251 ();
 sky130_fd_sc_hs__tap_1 TAP_252 ();
 sky130_fd_sc_hs__tap_1 TAP_253 ();
 sky130_fd_sc_hs__tap_1 TAP_254 ();
 sky130_fd_sc_hs__tap_1 TAP_255 ();
 sky130_fd_sc_hs__tap_1 TAP_256 ();
 sky130_fd_sc_hs__tap_1 TAP_257 ();
 sky130_fd_sc_hs__tap_1 TAP_258 ();
 sky130_fd_sc_hs__tap_1 TAP_259 ();
 sky130_fd_sc_hs__tap_1 TAP_260 ();
 sky130_fd_sc_hs__tap_1 TAP_261 ();
 sky130_fd_sc_hs__tap_1 TAP_262 ();
 sky130_fd_sc_hs__tap_1 TAP_263 ();
 sky130_fd_sc_hs__tap_1 TAP_264 ();
 sky130_fd_sc_hs__tap_1 TAP_265 ();
 sky130_fd_sc_hs__tap_1 TAP_266 ();
 sky130_fd_sc_hs__tap_1 TAP_267 ();
 sky130_fd_sc_hs__tap_1 TAP_268 ();
 sky130_fd_sc_hs__tap_1 TAP_269 ();
 sky130_fd_sc_hs__tap_1 TAP_270 ();
 sky130_fd_sc_hs__tap_1 TAP_271 ();
 sky130_fd_sc_hs__tap_1 TAP_272 ();
 sky130_fd_sc_hs__tap_1 TAP_273 ();
 sky130_fd_sc_hs__tap_1 TAP_274 ();
 sky130_fd_sc_hs__tap_1 TAP_275 ();
 sky130_fd_sc_hs__tap_1 TAP_276 ();
 sky130_fd_sc_hs__tap_1 TAP_277 ();
 sky130_fd_sc_hs__tap_1 TAP_278 ();
 sky130_fd_sc_hs__tap_1 TAP_279 ();
 sky130_fd_sc_hs__tap_1 TAP_280 ();
 sky130_fd_sc_hs__tap_1 TAP_281 ();
 sky130_fd_sc_hs__tap_1 TAP_282 ();
 sky130_fd_sc_hs__tap_1 TAP_283 ();
 sky130_fd_sc_hs__tap_1 TAP_284 ();
 sky130_fd_sc_hs__tap_1 TAP_285 ();
 sky130_fd_sc_hs__tap_1 TAP_286 ();
 sky130_fd_sc_hs__tap_1 TAP_287 ();
 sky130_fd_sc_hs__tap_1 TAP_288 ();
 sky130_fd_sc_hs__tap_1 TAP_289 ();
 sky130_fd_sc_hs__tap_1 TAP_290 ();
 sky130_fd_sc_hs__tap_1 TAP_291 ();
 sky130_fd_sc_hs__tap_1 TAP_292 ();
 sky130_fd_sc_hs__tap_1 TAP_293 ();
 sky130_fd_sc_hs__tap_1 TAP_294 ();
 sky130_fd_sc_hs__tap_1 TAP_295 ();
 sky130_fd_sc_hs__tap_1 TAP_296 ();
 sky130_fd_sc_hs__tap_1 TAP_297 ();
 sky130_fd_sc_hs__tap_1 TAP_298 ();
 sky130_fd_sc_hs__tap_1 TAP_299 ();
 sky130_fd_sc_hs__tap_1 TAP_300 ();
 sky130_fd_sc_hs__tap_1 TAP_301 ();
 sky130_fd_sc_hs__tap_1 TAP_302 ();
 sky130_fd_sc_hs__tap_1 TAP_303 ();
 sky130_fd_sc_hs__tap_1 TAP_304 ();
 sky130_fd_sc_hs__tap_1 TAP_305 ();
 sky130_fd_sc_hs__tap_1 TAP_306 ();
 sky130_fd_sc_hs__tap_1 TAP_307 ();
 sky130_fd_sc_hs__tap_1 TAP_308 ();
 sky130_fd_sc_hs__tap_1 TAP_309 ();
 sky130_fd_sc_hs__tap_1 TAP_310 ();
 sky130_fd_sc_hs__tap_1 TAP_311 ();
 sky130_fd_sc_hs__tap_1 TAP_312 ();
 sky130_fd_sc_hs__tap_1 TAP_313 ();
 sky130_fd_sc_hs__tap_1 TAP_314 ();
 sky130_fd_sc_hs__tap_1 TAP_315 ();
 sky130_fd_sc_hs__tap_1 TAP_316 ();
 sky130_fd_sc_hs__tap_1 TAP_317 ();
 sky130_fd_sc_hs__tap_1 TAP_318 ();
 sky130_fd_sc_hs__tap_1 TAP_319 ();
 sky130_fd_sc_hs__tap_1 TAP_320 ();
 sky130_fd_sc_hs__tap_1 TAP_321 ();
 sky130_fd_sc_hs__tap_1 TAP_322 ();
 sky130_fd_sc_hs__tap_1 TAP_323 ();
 sky130_fd_sc_hs__tap_1 TAP_324 ();
 sky130_fd_sc_hs__tap_1 TAP_325 ();
 sky130_fd_sc_hs__tap_1 TAP_326 ();
 sky130_fd_sc_hs__tap_1 TAP_327 ();
 sky130_fd_sc_hs__tap_1 TAP_328 ();
 sky130_fd_sc_hs__tap_1 TAP_329 ();
 sky130_fd_sc_hs__tap_1 TAP_330 ();
 sky130_fd_sc_hs__tap_1 TAP_331 ();
 sky130_fd_sc_hs__tap_1 TAP_332 ();
 sky130_fd_sc_hs__tap_1 TAP_333 ();
 sky130_fd_sc_hs__tap_1 TAP_334 ();
 sky130_fd_sc_hs__tap_1 TAP_335 ();
 sky130_fd_sc_hs__tap_1 TAP_336 ();
 sky130_fd_sc_hs__tap_1 TAP_337 ();
 sky130_fd_sc_hs__tap_1 TAP_338 ();
 sky130_fd_sc_hs__tap_1 TAP_339 ();
 sky130_fd_sc_hs__tap_1 TAP_340 ();
 sky130_fd_sc_hs__tap_1 TAP_341 ();
 sky130_fd_sc_hs__tap_1 TAP_342 ();
 sky130_fd_sc_hs__tap_1 TAP_343 ();
 sky130_fd_sc_hs__tap_1 TAP_344 ();
 sky130_fd_sc_hs__tap_1 TAP_345 ();
 sky130_fd_sc_hs__tap_1 TAP_346 ();
 sky130_fd_sc_hs__tap_1 TAP_347 ();
 sky130_fd_sc_hs__tap_1 TAP_348 ();
 sky130_fd_sc_hs__tap_1 TAP_349 ();
 sky130_fd_sc_hs__tap_1 TAP_350 ();
 sky130_fd_sc_hs__tap_1 TAP_351 ();
 sky130_fd_sc_hs__tap_1 TAP_352 ();
 sky130_fd_sc_hs__tap_1 TAP_353 ();
 sky130_fd_sc_hs__tap_1 TAP_354 ();
 sky130_fd_sc_hs__tap_1 TAP_355 ();
 sky130_fd_sc_hs__tap_1 TAP_356 ();
 sky130_fd_sc_hs__tap_1 TAP_357 ();
 sky130_fd_sc_hs__tap_1 TAP_358 ();
 sky130_fd_sc_hs__tap_1 TAP_359 ();
 sky130_fd_sc_hs__tap_1 TAP_360 ();
 sky130_fd_sc_hs__tap_1 TAP_361 ();
 sky130_fd_sc_hs__tap_1 TAP_362 ();
 sky130_fd_sc_hs__tap_1 TAP_363 ();
 sky130_fd_sc_hs__tap_1 TAP_364 ();
 sky130_fd_sc_hs__tap_1 TAP_365 ();
 sky130_fd_sc_hs__tap_1 TAP_366 ();
 sky130_fd_sc_hs__tap_1 TAP_367 ();
 sky130_fd_sc_hs__tap_1 TAP_368 ();
 sky130_fd_sc_hs__tap_1 TAP_369 ();
 sky130_fd_sc_hs__tap_1 TAP_370 ();
 sky130_fd_sc_hs__tap_1 TAP_371 ();
 sky130_fd_sc_hs__tap_1 TAP_372 ();
 sky130_fd_sc_hs__tap_1 TAP_373 ();
 sky130_fd_sc_hs__tap_1 TAP_374 ();
 sky130_fd_sc_hs__tap_1 TAP_375 ();
 sky130_fd_sc_hs__tap_1 TAP_376 ();
 sky130_fd_sc_hs__tap_1 TAP_377 ();
 sky130_fd_sc_hs__tap_1 TAP_378 ();
 sky130_fd_sc_hs__tap_1 TAP_379 ();
 sky130_fd_sc_hs__tap_1 TAP_380 ();
 sky130_fd_sc_hs__tap_1 TAP_381 ();
 sky130_fd_sc_hs__tap_1 TAP_382 ();
 sky130_fd_sc_hs__tap_1 TAP_383 ();
 sky130_fd_sc_hs__tap_1 TAP_384 ();
 sky130_fd_sc_hs__tap_1 TAP_385 ();
 sky130_fd_sc_hs__tap_1 TAP_386 ();
 sky130_fd_sc_hs__tap_1 TAP_387 ();
 sky130_fd_sc_hs__tap_1 TAP_388 ();
 sky130_fd_sc_hs__tap_1 TAP_389 ();
 sky130_fd_sc_hs__tap_1 TAP_390 ();
 sky130_fd_sc_hs__tap_1 TAP_391 ();
 sky130_fd_sc_hs__tap_1 TAP_392 ();
 sky130_fd_sc_hs__tap_1 TAP_393 ();
 sky130_fd_sc_hs__tap_1 TAP_394 ();
 sky130_fd_sc_hs__tap_1 TAP_395 ();
 sky130_fd_sc_hs__tap_1 TAP_396 ();
 sky130_fd_sc_hs__tap_1 TAP_397 ();
 sky130_fd_sc_hs__tap_1 TAP_398 ();
 sky130_fd_sc_hs__tap_1 TAP_399 ();
 sky130_fd_sc_hs__tap_1 TAP_400 ();
 sky130_fd_sc_hs__tap_1 TAP_401 ();
 sky130_fd_sc_hs__tap_1 TAP_402 ();
 sky130_fd_sc_hs__tap_1 TAP_403 ();
 sky130_fd_sc_hs__tap_1 TAP_404 ();
 sky130_fd_sc_hs__tap_1 TAP_405 ();
 sky130_fd_sc_hs__tap_1 TAP_406 ();
 sky130_fd_sc_hs__tap_1 TAP_407 ();
 sky130_fd_sc_hs__tap_1 TAP_408 ();
 sky130_fd_sc_hs__tap_1 TAP_409 ();
 sky130_fd_sc_hs__tap_1 TAP_410 ();
 sky130_fd_sc_hs__tap_1 TAP_411 ();
 sky130_fd_sc_hs__tap_1 TAP_412 ();
 sky130_fd_sc_hs__tap_1 TAP_413 ();
 sky130_fd_sc_hs__tap_1 TAP_414 ();
 sky130_fd_sc_hs__tap_1 TAP_415 ();
 sky130_fd_sc_hs__tap_1 TAP_416 ();
 sky130_fd_sc_hs__tap_1 TAP_417 ();
 sky130_fd_sc_hs__tap_1 TAP_418 ();
 sky130_fd_sc_hs__tap_1 TAP_419 ();
 sky130_fd_sc_hs__tap_1 TAP_420 ();
 sky130_fd_sc_hs__tap_1 TAP_421 ();
 sky130_fd_sc_hs__tap_1 TAP_422 ();
 sky130_fd_sc_hs__tap_1 TAP_423 ();
 sky130_fd_sc_hs__tap_1 TAP_424 ();
 sky130_fd_sc_hs__tap_1 TAP_425 ();
 sky130_fd_sc_hs__tap_1 TAP_426 ();
 sky130_fd_sc_hs__tap_1 TAP_427 ();
 sky130_fd_sc_hs__tap_1 TAP_428 ();
 sky130_fd_sc_hs__tap_1 TAP_429 ();
 sky130_fd_sc_hs__tap_1 TAP_430 ();
 sky130_fd_sc_hs__tap_1 TAP_431 ();
 sky130_fd_sc_hs__tap_1 TAP_432 ();
 sky130_fd_sc_hs__tap_1 TAP_433 ();
 sky130_fd_sc_hs__tap_1 TAP_434 ();
 sky130_fd_sc_hs__tap_1 TAP_435 ();
 sky130_fd_sc_hs__tap_1 TAP_436 ();
 sky130_fd_sc_hs__tap_1 TAP_437 ();
 sky130_fd_sc_hs__tap_1 TAP_438 ();
 sky130_fd_sc_hs__tap_1 TAP_439 ();
 sky130_fd_sc_hs__tap_1 TAP_440 ();
 sky130_fd_sc_hs__tap_1 TAP_441 ();
 sky130_fd_sc_hs__tap_1 TAP_442 ();
 sky130_fd_sc_hs__tap_1 TAP_443 ();
 sky130_fd_sc_hs__tap_1 TAP_444 ();
 sky130_fd_sc_hs__tap_1 TAP_445 ();
 sky130_fd_sc_hs__tap_1 TAP_446 ();
 sky130_fd_sc_hs__tap_1 TAP_447 ();
 sky130_fd_sc_hs__tap_1 TAP_448 ();
 sky130_fd_sc_hs__tap_1 TAP_449 ();
 sky130_fd_sc_hs__tap_1 TAP_450 ();
 sky130_fd_sc_hs__tap_1 TAP_451 ();
 sky130_fd_sc_hs__tap_1 TAP_452 ();
 sky130_fd_sc_hs__tap_1 TAP_453 ();
 sky130_fd_sc_hs__tap_1 TAP_454 ();
 sky130_fd_sc_hs__tap_1 TAP_455 ();
 sky130_fd_sc_hs__tap_1 TAP_456 ();
 sky130_fd_sc_hs__tap_1 TAP_457 ();
 sky130_fd_sc_hs__tap_1 TAP_458 ();
 sky130_fd_sc_hs__tap_1 TAP_459 ();
 sky130_fd_sc_hs__tap_1 TAP_460 ();
 sky130_fd_sc_hs__tap_1 TAP_461 ();
 sky130_fd_sc_hs__tap_1 TAP_462 ();
 sky130_fd_sc_hs__tap_1 TAP_463 ();
 sky130_fd_sc_hs__tap_1 TAP_464 ();
 sky130_fd_sc_hs__tap_1 TAP_465 ();
 sky130_fd_sc_hs__tap_1 TAP_466 ();
 sky130_fd_sc_hs__tap_1 TAP_467 ();
 sky130_fd_sc_hs__tap_1 TAP_468 ();
 sky130_fd_sc_hs__tap_1 TAP_469 ();
 sky130_fd_sc_hs__tap_1 TAP_470 ();
 sky130_fd_sc_hs__tap_1 TAP_471 ();
 sky130_fd_sc_hs__tap_1 TAP_472 ();
 sky130_fd_sc_hs__tap_1 TAP_473 ();
 sky130_fd_sc_hs__tap_1 TAP_474 ();
 sky130_fd_sc_hs__tap_1 TAP_475 ();
 sky130_fd_sc_hs__tap_1 TAP_476 ();
 sky130_fd_sc_hs__tap_1 TAP_477 ();
 sky130_fd_sc_hs__tap_1 TAP_478 ();
 sky130_fd_sc_hs__tap_1 TAP_479 ();
 sky130_fd_sc_hs__tap_1 TAP_480 ();
 sky130_fd_sc_hs__tap_1 TAP_481 ();
 sky130_fd_sc_hs__tap_1 TAP_482 ();
 sky130_fd_sc_hs__tap_1 TAP_483 ();
 sky130_fd_sc_hs__tap_1 TAP_484 ();
 sky130_fd_sc_hs__tap_1 TAP_485 ();
 sky130_fd_sc_hs__tap_1 TAP_486 ();
 sky130_fd_sc_hs__tap_1 TAP_487 ();
 sky130_fd_sc_hs__tap_1 TAP_488 ();
 sky130_fd_sc_hs__tap_1 TAP_489 ();
 sky130_fd_sc_hs__tap_1 TAP_490 ();
 sky130_fd_sc_hs__tap_1 TAP_491 ();
 sky130_fd_sc_hs__tap_1 TAP_492 ();
 sky130_fd_sc_hs__tap_1 TAP_493 ();
 sky130_fd_sc_hs__tap_1 TAP_494 ();
 sky130_fd_sc_hs__tap_1 TAP_495 ();
 sky130_fd_sc_hs__tap_1 TAP_496 ();
 sky130_fd_sc_hs__tap_1 TAP_497 ();
 sky130_fd_sc_hs__tap_1 TAP_498 ();
 sky130_fd_sc_hs__tap_1 TAP_499 ();
 sky130_fd_sc_hs__tap_1 TAP_500 ();
 sky130_fd_sc_hs__tap_1 TAP_501 ();
 sky130_fd_sc_hs__tap_1 TAP_502 ();
 sky130_fd_sc_hs__tap_1 TAP_503 ();
 sky130_fd_sc_hs__tap_1 TAP_504 ();
 sky130_fd_sc_hs__tap_1 TAP_505 ();
 sky130_fd_sc_hs__tap_1 TAP_506 ();
 sky130_fd_sc_hs__tap_1 TAP_507 ();
 sky130_fd_sc_hs__tap_1 TAP_508 ();
 sky130_fd_sc_hs__tap_1 TAP_509 ();
 sky130_fd_sc_hs__tap_1 TAP_510 ();
 sky130_fd_sc_hs__tap_1 TAP_511 ();
 sky130_fd_sc_hs__tap_1 TAP_512 ();
 sky130_fd_sc_hs__tap_1 TAP_513 ();
 sky130_fd_sc_hs__tap_1 TAP_514 ();
 sky130_fd_sc_hs__tap_1 TAP_515 ();
 sky130_fd_sc_hs__tap_1 TAP_516 ();
 sky130_fd_sc_hs__tap_1 TAP_517 ();
 sky130_fd_sc_hs__tap_1 TAP_518 ();
 sky130_fd_sc_hs__tap_1 TAP_519 ();
 sky130_fd_sc_hs__tap_1 TAP_520 ();
 sky130_fd_sc_hs__tap_1 TAP_521 ();
 sky130_fd_sc_hs__tap_1 TAP_522 ();
 sky130_fd_sc_hs__tap_1 TAP_523 ();
 sky130_fd_sc_hs__tap_1 TAP_524 ();
 sky130_fd_sc_hs__tap_1 TAP_525 ();
 sky130_fd_sc_hs__tap_1 TAP_526 ();
 sky130_fd_sc_hs__tap_1 TAP_527 ();
 sky130_fd_sc_hs__tap_1 TAP_528 ();
 sky130_fd_sc_hs__tap_1 TAP_529 ();
 sky130_fd_sc_hs__tap_1 TAP_530 ();
 sky130_fd_sc_hs__tap_1 TAP_531 ();
 sky130_fd_sc_hs__tap_1 TAP_532 ();
 sky130_fd_sc_hs__tap_1 TAP_533 ();
 sky130_fd_sc_hs__tap_1 TAP_534 ();
 sky130_fd_sc_hs__tap_1 TAP_535 ();
 sky130_fd_sc_hs__tap_1 TAP_536 ();
 sky130_fd_sc_hs__tap_1 TAP_537 ();
 sky130_fd_sc_hs__tap_1 TAP_538 ();
 sky130_fd_sc_hs__tap_1 TAP_539 ();
 sky130_fd_sc_hs__tap_1 TAP_540 ();
 sky130_fd_sc_hs__tap_1 TAP_541 ();
 sky130_fd_sc_hs__tap_1 TAP_542 ();
 sky130_fd_sc_hs__tap_1 TAP_543 ();
 sky130_fd_sc_hs__tap_1 TAP_544 ();
 sky130_fd_sc_hs__tap_1 TAP_545 ();
 sky130_fd_sc_hs__tap_1 TAP_546 ();
 sky130_fd_sc_hs__tap_1 TAP_547 ();
 sky130_fd_sc_hs__tap_1 TAP_548 ();
 sky130_fd_sc_hs__tap_1 TAP_549 ();
 sky130_fd_sc_hs__tap_1 TAP_550 ();
 sky130_fd_sc_hs__tap_1 TAP_551 ();
 sky130_fd_sc_hs__tap_1 TAP_552 ();
 sky130_fd_sc_hs__tap_1 TAP_553 ();
 sky130_fd_sc_hs__tap_1 TAP_554 ();
 sky130_fd_sc_hs__tap_1 TAP_555 ();
 sky130_fd_sc_hs__tap_1 TAP_556 ();
 sky130_fd_sc_hs__tap_1 TAP_557 ();
 sky130_fd_sc_hs__tap_1 TAP_558 ();
 sky130_fd_sc_hs__tap_1 TAP_559 ();
 sky130_fd_sc_hs__tap_1 TAP_560 ();
 sky130_fd_sc_hs__tap_1 TAP_561 ();
 sky130_fd_sc_hs__tap_1 TAP_562 ();
 sky130_fd_sc_hs__tap_1 TAP_563 ();
 sky130_fd_sc_hs__tap_1 TAP_564 ();
 sky130_fd_sc_hs__tap_1 TAP_565 ();
 sky130_fd_sc_hs__tap_1 TAP_566 ();
 sky130_fd_sc_hs__tap_1 TAP_567 ();
 sky130_fd_sc_hs__tap_1 TAP_568 ();
 sky130_fd_sc_hs__tap_1 TAP_569 ();
 sky130_fd_sc_hs__tap_1 TAP_570 ();
 sky130_fd_sc_hs__tap_1 TAP_571 ();
 sky130_fd_sc_hs__tap_1 TAP_572 ();
 sky130_fd_sc_hs__tap_1 TAP_573 ();
 sky130_fd_sc_hs__tap_1 TAP_574 ();
 sky130_fd_sc_hs__tap_1 TAP_575 ();
 sky130_fd_sc_hs__tap_1 TAP_576 ();
 sky130_fd_sc_hs__tap_1 TAP_577 ();
 sky130_fd_sc_hs__tap_1 TAP_578 ();
 sky130_fd_sc_hs__tap_1 TAP_579 ();
 sky130_fd_sc_hs__tap_1 TAP_580 ();
 sky130_fd_sc_hs__tap_1 TAP_581 ();
 sky130_fd_sc_hs__tap_1 TAP_582 ();
 sky130_fd_sc_hs__tap_1 TAP_583 ();
 sky130_fd_sc_hs__tap_1 TAP_584 ();
 sky130_fd_sc_hs__tap_1 TAP_585 ();
 sky130_fd_sc_hs__tap_1 TAP_586 ();
 sky130_fd_sc_hs__tap_1 TAP_587 ();
 sky130_fd_sc_hs__tap_1 TAP_588 ();
 sky130_fd_sc_hs__tap_1 TAP_589 ();
 sky130_fd_sc_hs__tap_1 TAP_590 ();
 sky130_fd_sc_hs__tap_1 TAP_591 ();
 sky130_fd_sc_hs__tap_1 TAP_592 ();
 sky130_fd_sc_hs__tap_1 TAP_593 ();
 sky130_fd_sc_hs__tap_1 TAP_594 ();
 sky130_fd_sc_hs__tap_1 TAP_595 ();
 sky130_fd_sc_hs__tap_1 TAP_596 ();
 sky130_fd_sc_hs__tap_1 TAP_597 ();
 sky130_fd_sc_hs__tap_1 TAP_598 ();
 sky130_fd_sc_hs__tap_1 TAP_599 ();
 sky130_fd_sc_hs__tap_1 TAP_600 ();
 sky130_fd_sc_hs__tap_1 TAP_601 ();
 sky130_fd_sc_hs__tap_1 TAP_602 ();
 sky130_fd_sc_hs__tap_1 TAP_603 ();
 sky130_fd_sc_hs__tap_1 TAP_604 ();
 sky130_fd_sc_hs__tap_1 TAP_605 ();
 sky130_fd_sc_hs__tap_1 TAP_606 ();
 sky130_fd_sc_hs__tap_1 TAP_607 ();
 sky130_fd_sc_hs__tap_1 TAP_608 ();
 sky130_fd_sc_hs__tap_1 TAP_609 ();
 sky130_fd_sc_hs__tap_1 TAP_610 ();
 sky130_fd_sc_hs__tap_1 TAP_611 ();
 sky130_fd_sc_hs__tap_1 TAP_612 ();
 sky130_fd_sc_hs__tap_1 TAP_613 ();
 sky130_fd_sc_hs__tap_1 TAP_614 ();
 sky130_fd_sc_hs__tap_1 TAP_615 ();
 sky130_fd_sc_hs__tap_1 TAP_616 ();
 sky130_fd_sc_hs__tap_1 TAP_617 ();
 sky130_fd_sc_hs__tap_1 TAP_618 ();
 sky130_fd_sc_hs__tap_1 TAP_619 ();
 sky130_fd_sc_hs__tap_1 TAP_620 ();
 sky130_fd_sc_hs__tap_1 TAP_621 ();
 sky130_fd_sc_hs__tap_1 TAP_622 ();
 sky130_fd_sc_hs__tap_1 TAP_623 ();
 sky130_fd_sc_hs__tap_1 TAP_624 ();
 sky130_fd_sc_hs__tap_1 TAP_625 ();
 sky130_fd_sc_hs__tap_1 TAP_626 ();
 sky130_fd_sc_hs__tap_1 TAP_627 ();
 sky130_fd_sc_hs__tap_1 TAP_628 ();
 sky130_fd_sc_hs__tap_1 TAP_629 ();
 sky130_fd_sc_hs__tap_1 TAP_630 ();
 sky130_fd_sc_hs__tap_1 TAP_631 ();
 sky130_fd_sc_hs__tap_1 TAP_632 ();
 sky130_fd_sc_hs__tap_1 TAP_633 ();
 sky130_fd_sc_hs__tap_1 TAP_634 ();
 sky130_fd_sc_hs__tap_1 TAP_635 ();
 sky130_fd_sc_hs__tap_1 TAP_636 ();
 sky130_fd_sc_hs__tap_1 TAP_637 ();
 sky130_fd_sc_hs__tap_1 TAP_638 ();
 sky130_fd_sc_hs__tap_1 TAP_639 ();
 sky130_fd_sc_hs__tap_1 TAP_640 ();
 sky130_fd_sc_hs__tap_1 TAP_641 ();
 sky130_fd_sc_hs__tap_1 TAP_642 ();
 sky130_fd_sc_hs__tap_1 TAP_643 ();
 sky130_fd_sc_hs__tap_1 TAP_644 ();
 sky130_fd_sc_hs__tap_1 TAP_645 ();
 sky130_fd_sc_hs__tap_1 TAP_646 ();
 sky130_fd_sc_hs__tap_1 TAP_647 ();
 sky130_fd_sc_hs__tap_1 TAP_648 ();
 sky130_fd_sc_hs__tap_1 TAP_649 ();
 sky130_fd_sc_hs__tap_1 TAP_650 ();
 sky130_fd_sc_hs__tap_1 TAP_651 ();
 sky130_fd_sc_hs__tap_1 TAP_652 ();
 sky130_fd_sc_hs__tap_1 TAP_653 ();
 sky130_fd_sc_hs__tap_1 TAP_654 ();
 sky130_fd_sc_hs__tap_1 TAP_655 ();
 sky130_fd_sc_hs__tap_1 TAP_656 ();
 sky130_fd_sc_hs__tap_1 TAP_657 ();
 sky130_fd_sc_hs__tap_1 TAP_658 ();
 sky130_fd_sc_hs__tap_1 TAP_659 ();
 sky130_fd_sc_hs__tap_1 TAP_660 ();
 sky130_fd_sc_hs__tap_1 TAP_661 ();
 sky130_fd_sc_hs__tap_1 TAP_662 ();
 sky130_fd_sc_hs__tap_1 TAP_663 ();
 sky130_fd_sc_hs__tap_1 TAP_664 ();
 sky130_fd_sc_hs__tap_1 TAP_665 ();
 sky130_fd_sc_hs__tap_1 TAP_666 ();
 sky130_fd_sc_hs__tap_1 TAP_667 ();
 sky130_fd_sc_hs__tap_1 TAP_668 ();
 sky130_fd_sc_hs__tap_1 TAP_669 ();
 sky130_fd_sc_hs__tap_1 TAP_670 ();
 sky130_fd_sc_hs__tap_1 TAP_671 ();
 sky130_fd_sc_hs__tap_1 TAP_672 ();
 sky130_fd_sc_hs__tap_1 TAP_673 ();
 sky130_fd_sc_hs__tap_1 TAP_674 ();
 sky130_fd_sc_hs__tap_1 TAP_675 ();
 sky130_fd_sc_hs__tap_1 TAP_676 ();
 sky130_fd_sc_hs__tap_1 TAP_677 ();
 sky130_fd_sc_hs__tap_1 TAP_678 ();
 sky130_fd_sc_hs__tap_1 TAP_679 ();
 sky130_fd_sc_hs__tap_1 TAP_680 ();
 sky130_fd_sc_hs__tap_1 TAP_681 ();
 sky130_fd_sc_hs__tap_1 TAP_682 ();
 sky130_fd_sc_hs__tap_1 TAP_683 ();
 sky130_fd_sc_hs__tap_1 TAP_684 ();
 sky130_fd_sc_hs__tap_1 TAP_685 ();
 sky130_fd_sc_hs__tap_1 TAP_686 ();
 sky130_fd_sc_hs__tap_1 TAP_687 ();
 sky130_fd_sc_hs__tap_1 TAP_688 ();
 sky130_fd_sc_hs__tap_1 TAP_689 ();
 sky130_fd_sc_hs__tap_1 TAP_690 ();
 sky130_fd_sc_hs__tap_1 TAP_691 ();
 sky130_fd_sc_hs__tap_1 TAP_692 ();
 sky130_fd_sc_hs__tap_1 TAP_693 ();
 sky130_fd_sc_hs__tap_1 TAP_694 ();
 sky130_fd_sc_hs__tap_1 TAP_695 ();
 sky130_fd_sc_hs__tap_1 TAP_696 ();
 sky130_fd_sc_hs__tap_1 TAP_697 ();
 sky130_fd_sc_hs__tap_1 TAP_698 ();
 sky130_fd_sc_hs__tap_1 TAP_699 ();
 sky130_fd_sc_hs__tap_1 TAP_700 ();
 sky130_fd_sc_hs__tap_1 TAP_701 ();
 sky130_fd_sc_hs__tap_1 TAP_702 ();
 sky130_fd_sc_hs__tap_1 TAP_703 ();
 sky130_fd_sc_hs__tap_1 TAP_704 ();
 sky130_fd_sc_hs__tap_1 TAP_705 ();
 sky130_fd_sc_hs__tap_1 TAP_706 ();
 sky130_fd_sc_hs__tap_1 TAP_707 ();
 sky130_fd_sc_hs__tap_1 TAP_708 ();
 sky130_fd_sc_hs__tap_1 TAP_709 ();
 sky130_fd_sc_hs__tap_1 TAP_710 ();
 sky130_fd_sc_hs__tap_1 TAP_711 ();
 sky130_fd_sc_hs__tap_1 TAP_712 ();
 sky130_fd_sc_hs__tap_1 TAP_713 ();
 sky130_fd_sc_hs__tap_1 TAP_714 ();
 sky130_fd_sc_hs__tap_1 TAP_715 ();
 sky130_fd_sc_hs__tap_1 TAP_716 ();
 sky130_fd_sc_hs__tap_1 TAP_717 ();
 sky130_fd_sc_hs__tap_1 TAP_718 ();
 sky130_fd_sc_hs__tap_1 TAP_719 ();
 sky130_fd_sc_hs__tap_1 TAP_720 ();
 sky130_fd_sc_hs__tap_1 TAP_721 ();
 sky130_fd_sc_hs__tap_1 TAP_722 ();
 sky130_fd_sc_hs__tap_1 TAP_723 ();
 sky130_fd_sc_hs__tap_1 TAP_724 ();
 sky130_fd_sc_hs__tap_1 TAP_725 ();
 sky130_fd_sc_hs__tap_1 TAP_726 ();
 sky130_fd_sc_hs__tap_1 TAP_727 ();
 sky130_fd_sc_hs__tap_1 TAP_728 ();
 sky130_fd_sc_hs__tap_1 TAP_729 ();
 sky130_fd_sc_hs__tap_1 TAP_730 ();
 sky130_fd_sc_hs__tap_1 TAP_731 ();
 sky130_fd_sc_hs__tap_1 TAP_732 ();
 sky130_fd_sc_hs__tap_1 TAP_733 ();
 sky130_fd_sc_hs__tap_1 TAP_734 ();
 sky130_fd_sc_hs__tap_1 TAP_735 ();
 sky130_fd_sc_hs__tap_1 TAP_736 ();
 sky130_fd_sc_hs__tap_1 TAP_737 ();
 sky130_fd_sc_hs__tap_1 TAP_738 ();
 sky130_fd_sc_hs__tap_1 TAP_739 ();
 sky130_fd_sc_hs__tap_1 TAP_740 ();
 sky130_fd_sc_hs__tap_1 TAP_741 ();
 sky130_fd_sc_hs__tap_1 TAP_742 ();
 sky130_fd_sc_hs__tap_1 TAP_743 ();
 sky130_fd_sc_hs__tap_1 TAP_744 ();
 sky130_fd_sc_hs__tap_1 TAP_745 ();
 sky130_fd_sc_hs__tap_1 TAP_746 ();
 sky130_fd_sc_hs__tap_1 TAP_747 ();
 sky130_fd_sc_hs__tap_1 TAP_748 ();
 sky130_fd_sc_hs__tap_1 TAP_749 ();
 sky130_fd_sc_hs__tap_1 TAP_750 ();
 sky130_fd_sc_hs__tap_1 TAP_751 ();
 sky130_fd_sc_hs__tap_1 TAP_752 ();
 sky130_fd_sc_hs__tap_1 TAP_753 ();
 sky130_fd_sc_hs__tap_1 TAP_754 ();
 sky130_fd_sc_hs__tap_1 TAP_755 ();
 sky130_fd_sc_hs__tap_1 TAP_756 ();
 sky130_fd_sc_hs__tap_1 TAP_757 ();
 sky130_fd_sc_hs__tap_1 TAP_758 ();
 sky130_fd_sc_hs__tap_1 TAP_759 ();
 sky130_fd_sc_hs__tap_1 TAP_760 ();
 sky130_fd_sc_hs__tap_1 TAP_761 ();
 sky130_fd_sc_hs__tap_1 TAP_762 ();
 sky130_fd_sc_hs__tap_1 TAP_763 ();
 sky130_fd_sc_hs__tap_1 TAP_764 ();
 sky130_fd_sc_hs__tap_1 TAP_765 ();
 sky130_fd_sc_hs__tap_1 TAP_766 ();
 sky130_fd_sc_hs__tap_1 TAP_767 ();
 sky130_fd_sc_hs__tap_1 TAP_768 ();
 sky130_fd_sc_hs__tap_1 TAP_769 ();
 sky130_fd_sc_hs__tap_1 TAP_770 ();
 sky130_fd_sc_hs__tap_1 TAP_771 ();
 sky130_fd_sc_hs__tap_1 TAP_772 ();
 sky130_fd_sc_hs__tap_1 TAP_773 ();
 sky130_fd_sc_hs__tap_1 TAP_774 ();
 sky130_fd_sc_hs__tap_1 TAP_775 ();
 sky130_fd_sc_hs__tap_1 TAP_776 ();
 sky130_fd_sc_hs__tap_1 TAP_777 ();
 sky130_fd_sc_hs__tap_1 TAP_778 ();
 sky130_fd_sc_hs__tap_1 TAP_779 ();
 sky130_fd_sc_hs__tap_1 TAP_780 ();
 sky130_fd_sc_hs__tap_1 TAP_781 ();
 sky130_fd_sc_hs__tap_1 TAP_782 ();
 sky130_fd_sc_hs__tap_1 TAP_783 ();
 sky130_fd_sc_hs__tap_1 TAP_784 ();
 sky130_fd_sc_hs__tap_1 TAP_785 ();
 sky130_fd_sc_hs__tap_1 TAP_786 ();
 sky130_fd_sc_hs__tap_1 TAP_787 ();
 sky130_fd_sc_hs__tap_1 TAP_788 ();
 sky130_fd_sc_hs__tap_1 TAP_789 ();
 sky130_fd_sc_hs__tap_1 TAP_790 ();
 sky130_fd_sc_hs__tap_1 TAP_791 ();
 sky130_fd_sc_hs__tap_1 TAP_792 ();
 sky130_fd_sc_hs__tap_1 TAP_793 ();
 sky130_fd_sc_hs__tap_1 TAP_794 ();
 sky130_fd_sc_hs__tap_1 TAP_795 ();
 sky130_fd_sc_hs__tap_1 TAP_796 ();
 sky130_fd_sc_hs__tap_1 TAP_797 ();
 sky130_fd_sc_hs__tap_1 TAP_798 ();
 sky130_fd_sc_hs__tap_1 TAP_799 ();
 sky130_fd_sc_hs__tap_1 TAP_800 ();
 sky130_fd_sc_hs__tap_1 TAP_801 ();
 sky130_fd_sc_hs__tap_1 TAP_802 ();
 sky130_fd_sc_hs__tap_1 TAP_803 ();
 sky130_fd_sc_hs__tap_1 TAP_804 ();
 sky130_fd_sc_hs__tap_1 TAP_805 ();
 sky130_fd_sc_hs__tap_1 TAP_806 ();
 sky130_fd_sc_hs__tap_1 TAP_807 ();
 sky130_fd_sc_hs__tap_1 TAP_808 ();
 sky130_fd_sc_hs__tap_1 TAP_809 ();
 sky130_fd_sc_hs__tap_1 TAP_810 ();
 sky130_fd_sc_hs__tap_1 TAP_811 ();
 sky130_fd_sc_hs__tap_1 TAP_812 ();
 sky130_fd_sc_hs__tap_1 TAP_813 ();
 sky130_fd_sc_hs__tap_1 TAP_814 ();
 sky130_fd_sc_hs__tap_1 TAP_815 ();
 sky130_fd_sc_hs__tap_1 TAP_816 ();
 sky130_fd_sc_hs__tap_1 TAP_817 ();
 sky130_fd_sc_hs__tap_1 TAP_818 ();
 sky130_fd_sc_hs__tap_1 TAP_819 ();
 sky130_fd_sc_hs__tap_1 TAP_820 ();
 sky130_fd_sc_hs__tap_1 TAP_821 ();
 sky130_fd_sc_hs__tap_1 TAP_822 ();
 sky130_fd_sc_hs__tap_1 TAP_823 ();
 sky130_fd_sc_hs__tap_1 TAP_824 ();
 sky130_fd_sc_hs__tap_1 TAP_825 ();
 sky130_fd_sc_hs__tap_1 TAP_826 ();
 sky130_fd_sc_hs__tap_1 TAP_827 ();
 sky130_fd_sc_hs__tap_1 TAP_828 ();
 sky130_fd_sc_hs__tap_1 TAP_829 ();
 sky130_fd_sc_hs__tap_1 TAP_830 ();
 sky130_fd_sc_hs__tap_1 TAP_831 ();
 sky130_fd_sc_hs__tap_1 TAP_832 ();
 sky130_fd_sc_hs__tap_1 TAP_833 ();
 sky130_fd_sc_hs__tap_1 TAP_834 ();
 sky130_fd_sc_hs__tap_1 TAP_835 ();
 sky130_fd_sc_hs__tap_1 TAP_836 ();
 sky130_fd_sc_hs__tap_1 TAP_837 ();
 sky130_fd_sc_hs__tap_1 TAP_838 ();
 sky130_fd_sc_hs__tap_1 TAP_839 ();
 sky130_fd_sc_hs__tap_1 TAP_840 ();
 sky130_fd_sc_hs__tap_1 TAP_841 ();
 sky130_fd_sc_hs__tap_1 TAP_842 ();
 sky130_fd_sc_hs__tap_1 TAP_843 ();
 sky130_fd_sc_hs__tap_1 TAP_844 ();
 sky130_fd_sc_hs__tap_1 TAP_845 ();
 sky130_fd_sc_hs__tap_1 TAP_846 ();
 sky130_fd_sc_hs__tap_1 TAP_847 ();
 sky130_fd_sc_hs__tap_1 TAP_848 ();
 sky130_fd_sc_hs__tap_1 TAP_849 ();
 sky130_fd_sc_hs__clkbuf_4 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hs__clkbuf_4 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hs__clkbuf_4 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hs__clkbuf_4 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hs__clkbuf_4 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer1 (.A(\dpath.a_lt_b$in1[3] ),
    .X(net1));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer2 (.A(_039_),
    .X(net2));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer3 (.A(\dpath.a_lt_b$in1[2] ),
    .X(net3));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer4 (.A(_075_),
    .X(net4));
 sky130_fd_sc_hs__buf_2 rebuffer5 (.A(_098_),
    .X(net5));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer6 (.A(\dpath.a_lt_b$in1[7] ),
    .X(net6));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer7 (.A(_051_),
    .X(net7));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer8 (.A(_056_),
    .X(net8));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer9 (.A(\dpath.a_lt_b$in1[5] ),
    .X(net9));
 sky130_fd_sc_hs__clkbuf_2 rebuffer10 (.A(_112_),
    .X(net10));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer11 (.A(_042_),
    .X(net11));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer12 (.A(_123_),
    .X(net12));
 sky130_fd_sc_hs__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_0_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_46 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_75 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_104 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_133 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_162 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_191 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_220 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_249 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_278 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_307 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_336 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_365 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_394 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_423 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_452 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_481 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_510 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_539 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_0_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_1_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_1_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_1_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_1_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_1_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_1_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_1_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_1_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_1_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_1_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_1_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_2_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_2_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_2_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_2_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_2_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_2_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_2_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_2_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_2_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_2_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_2_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_2_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_2_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_3_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_3_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_3_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_3_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_3_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_3_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_3_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_3_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_3_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_3_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_3_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_4_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_4_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_4_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_4_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_4_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_4_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_4_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_4_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_4_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_4_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_4_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_4_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_4_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_5_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_5_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_5_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_5_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_5_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_5_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_5_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_5_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_5_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_5_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_5_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_6_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_6_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_6_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_6_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_6_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_6_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_6_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_6_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_6_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_6_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_6_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_6_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_6_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_7_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_7_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_7_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_7_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_7_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_7_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_7_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_7_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_7_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_7_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_7_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_8_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_8_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_8_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_8_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_8_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_8_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_8_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_8_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_8_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_8_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_8_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_8_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_8_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_8_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_9_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_9_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_9_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_9_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_9_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_9_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_9_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_9_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_9_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_9_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_9_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_10_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_10_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_10_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_10_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_10_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_10_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_10_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_10_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_10_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_10_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_10_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_10_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_10_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_10_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_11_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_11_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_11_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_11_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_11_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_11_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_11_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_11_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_11_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_11_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_11_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_12_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_12_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_12_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_12_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_12_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_12_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_12_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_12_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_12_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_12_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_12_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_12_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_12_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_12_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_13_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_13_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_13_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_13_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_13_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_13_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_13_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_13_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_13_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_13_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_13_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_14_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_14_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_14_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_14_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_14_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_14_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_14_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_14_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_14_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_14_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_14_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_14_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_14_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_15_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_15_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_15_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_15_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_15_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_291 ();
 sky130_fd_sc_hs__fill_1 FILLER_15_299 ();
 sky130_fd_sc_hs__fill_4 FILLER_15_303 ();
 sky130_fd_sc_hs__fill_2 FILLER_15_307 ();
 sky130_fd_sc_hs__fill_1 FILLER_15_309 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_336 ();
 sky130_fd_sc_hs__fill_4 FILLER_15_344 ();
 sky130_fd_sc_hs__fill_4 FILLER_15_349 ();
 sky130_fd_sc_hs__fill_2 FILLER_15_353 ();
 sky130_fd_sc_hs__fill_1 FILLER_15_355 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_362 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_370 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_394 ();
 sky130_fd_sc_hs__fill_4 FILLER_15_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_15_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_15_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_15_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_15_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_16_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_16_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_16_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_16_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_16_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_278 ();
 sky130_fd_sc_hs__fill_2 FILLER_16_286 ();
 sky130_fd_sc_hs__fill_1 FILLER_16_288 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_307 ();
 sky130_fd_sc_hs__fill_4 FILLER_16_315 ();
 sky130_fd_sc_hs__fill_4 FILLER_16_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_329 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_337 ();
 sky130_fd_sc_hs__fill_2 FILLER_16_345 ();
 sky130_fd_sc_hs__fill_1 FILLER_16_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_366 ();
 sky130_fd_sc_hs__fill_2 FILLER_16_374 ();
 sky130_fd_sc_hs__fill_1 FILLER_16_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_16_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_16_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_16_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_16_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_16_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_16_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_17_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_17_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_17_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_17_231 ();
 sky130_fd_sc_hs__fill_4 FILLER_17_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_242 ();
 sky130_fd_sc_hs__fill_4 FILLER_17_250 ();
 sky130_fd_sc_hs__fill_2 FILLER_17_254 ();
 sky130_fd_sc_hs__fill_4 FILLER_17_264 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_17_289 ();
 sky130_fd_sc_hs__fill_4 FILLER_17_291 ();
 sky130_fd_sc_hs__fill_2 FILLER_17_295 ();
 sky130_fd_sc_hs__fill_4 FILLER_17_316 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_17_347 ();
 sky130_fd_sc_hs__fill_4 FILLER_17_349 ();
 sky130_fd_sc_hs__fill_2 FILLER_17_353 ();
 sky130_fd_sc_hs__fill_1 FILLER_17_355 ();
 sky130_fd_sc_hs__fill_4 FILLER_17_359 ();
 sky130_fd_sc_hs__fill_4 FILLER_17_366 ();
 sky130_fd_sc_hs__fill_1 FILLER_17_370 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_17_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_431 ();
 sky130_fd_sc_hs__fill_4 FILLER_17_439 ();
 sky130_fd_sc_hs__fill_2 FILLER_17_443 ();
 sky130_fd_sc_hs__fill_1 FILLER_17_445 ();
 sky130_fd_sc_hs__fill_4 FILLER_17_449 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_456 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_17_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_17_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_17_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_18_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_18_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_18_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_18_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_18_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_220 ();
 sky130_fd_sc_hs__fill_1 FILLER_18_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_232 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_240 ();
 sky130_fd_sc_hs__fill_4 FILLER_18_248 ();
 sky130_fd_sc_hs__fill_2 FILLER_18_252 ();
 sky130_fd_sc_hs__fill_4 FILLER_18_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_262 ();
 sky130_fd_sc_hs__fill_1 FILLER_18_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_274 ();
 sky130_fd_sc_hs__fill_2 FILLER_18_282 ();
 sky130_fd_sc_hs__fill_4 FILLER_18_289 ();
 sky130_fd_sc_hs__fill_4 FILLER_18_297 ();
 sky130_fd_sc_hs__fill_2 FILLER_18_301 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_306 ();
 sky130_fd_sc_hs__fill_4 FILLER_18_314 ();
 sky130_fd_sc_hs__fill_1 FILLER_18_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_334 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_342 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_350 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_358 ();
 sky130_fd_sc_hs__fill_4 FILLER_18_366 ();
 sky130_fd_sc_hs__fill_4 FILLER_18_373 ();
 sky130_fd_sc_hs__fill_4 FILLER_18_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_385 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_393 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_401 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_409 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_417 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_425 ();
 sky130_fd_sc_hs__fill_2 FILLER_18_433 ();
 sky130_fd_sc_hs__fill_4 FILLER_18_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_443 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_457 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_481 ();
 sky130_fd_sc_hs__fill_4 FILLER_18_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_18_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_18_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_18_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_18_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_19_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_19_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_19_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_199 ();
 sky130_fd_sc_hs__fill_4 FILLER_19_207 ();
 sky130_fd_sc_hs__fill_2 FILLER_19_211 ();
 sky130_fd_sc_hs__fill_1 FILLER_19_213 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_221 ();
 sky130_fd_sc_hs__fill_2 FILLER_19_229 ();
 sky130_fd_sc_hs__fill_1 FILLER_19_231 ();
 sky130_fd_sc_hs__fill_4 FILLER_19_233 ();
 sky130_fd_sc_hs__fill_1 FILLER_19_237 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_243 ();
 sky130_fd_sc_hs__fill_4 FILLER_19_251 ();
 sky130_fd_sc_hs__fill_1 FILLER_19_255 ();
 sky130_fd_sc_hs__fill_4 FILLER_19_259 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_266 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_274 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_282 ();
 sky130_fd_sc_hs__fill_4 FILLER_19_291 ();
 sky130_fd_sc_hs__fill_1 FILLER_19_295 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_19_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_349 ();
 sky130_fd_sc_hs__fill_4 FILLER_19_357 ();
 sky130_fd_sc_hs__fill_2 FILLER_19_361 ();
 sky130_fd_sc_hs__fill_4 FILLER_19_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_391 ();
 sky130_fd_sc_hs__fill_4 FILLER_19_399 ();
 sky130_fd_sc_hs__fill_2 FILLER_19_403 ();
 sky130_fd_sc_hs__fill_1 FILLER_19_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_415 ();
 sky130_fd_sc_hs__fill_1 FILLER_19_423 ();
 sky130_fd_sc_hs__fill_4 FILLER_19_427 ();
 sky130_fd_sc_hs__fill_4 FILLER_19_436 ();
 sky130_fd_sc_hs__fill_4 FILLER_19_457 ();
 sky130_fd_sc_hs__fill_2 FILLER_19_461 ();
 sky130_fd_sc_hs__fill_1 FILLER_19_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_19_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_19_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_19_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_20_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_20_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_20_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_20_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_204 ();
 sky130_fd_sc_hs__fill_4 FILLER_20_212 ();
 sky130_fd_sc_hs__fill_2 FILLER_20_216 ();
 sky130_fd_sc_hs__fill_1 FILLER_20_218 ();
 sky130_fd_sc_hs__fill_4 FILLER_20_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_20_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_262 ();
 sky130_fd_sc_hs__fill_4 FILLER_20_270 ();
 sky130_fd_sc_hs__fill_2 FILLER_20_274 ();
 sky130_fd_sc_hs__fill_1 FILLER_20_276 ();
 sky130_fd_sc_hs__fill_4 FILLER_20_281 ();
 sky130_fd_sc_hs__fill_2 FILLER_20_285 ();
 sky130_fd_sc_hs__fill_1 FILLER_20_287 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_293 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_301 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_309 ();
 sky130_fd_sc_hs__fill_2 FILLER_20_317 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_360 ();
 sky130_fd_sc_hs__fill_2 FILLER_20_368 ();
 sky130_fd_sc_hs__fill_4 FILLER_20_373 ();
 sky130_fd_sc_hs__fill_4 FILLER_20_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_387 ();
 sky130_fd_sc_hs__fill_4 FILLER_20_395 ();
 sky130_fd_sc_hs__fill_1 FILLER_20_399 ();
 sky130_fd_sc_hs__fill_4 FILLER_20_419 ();
 sky130_fd_sc_hs__fill_4 FILLER_20_428 ();
 sky130_fd_sc_hs__fill_2 FILLER_20_432 ();
 sky130_fd_sc_hs__fill_1 FILLER_20_434 ();
 sky130_fd_sc_hs__fill_4 FILLER_20_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_457 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_481 ();
 sky130_fd_sc_hs__fill_4 FILLER_20_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_20_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_20_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_20_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_20_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_21_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_21_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_21_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_215 ();
 sky130_fd_sc_hs__fill_2 FILLER_21_223 ();
 sky130_fd_sc_hs__fill_4 FILLER_21_228 ();
 sky130_fd_sc_hs__fill_4 FILLER_21_233 ();
 sky130_fd_sc_hs__fill_2 FILLER_21_237 ();
 sky130_fd_sc_hs__fill_4 FILLER_21_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_21_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_299 ();
 sky130_fd_sc_hs__fill_4 FILLER_21_307 ();
 sky130_fd_sc_hs__fill_1 FILLER_21_311 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_317 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_325 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_333 ();
 sky130_fd_sc_hs__fill_4 FILLER_21_341 ();
 sky130_fd_sc_hs__fill_2 FILLER_21_345 ();
 sky130_fd_sc_hs__fill_1 FILLER_21_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_349 ();
 sky130_fd_sc_hs__fill_4 FILLER_21_357 ();
 sky130_fd_sc_hs__fill_4 FILLER_21_364 ();
 sky130_fd_sc_hs__fill_4 FILLER_21_385 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_393 ();
 sky130_fd_sc_hs__fill_4 FILLER_21_401 ();
 sky130_fd_sc_hs__fill_1 FILLER_21_405 ();
 sky130_fd_sc_hs__fill_4 FILLER_21_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_419 ();
 sky130_fd_sc_hs__fill_2 FILLER_21_427 ();
 sky130_fd_sc_hs__fill_1 FILLER_21_429 ();
 sky130_fd_sc_hs__fill_4 FILLER_21_435 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_452 ();
 sky130_fd_sc_hs__fill_4 FILLER_21_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_21_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_21_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_21_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_22_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_22_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_22_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_22_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_212 ();
 sky130_fd_sc_hs__fill_2 FILLER_22_220 ();
 sky130_fd_sc_hs__fill_4 FILLER_22_240 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_247 ();
 sky130_fd_sc_hs__fill_4 FILLER_22_255 ();
 sky130_fd_sc_hs__fill_2 FILLER_22_259 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_302 ();
 sky130_fd_sc_hs__fill_4 FILLER_22_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_320 ();
 sky130_fd_sc_hs__fill_4 FILLER_22_328 ();
 sky130_fd_sc_hs__fill_2 FILLER_22_332 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_337 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_345 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_353 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_361 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_369 ();
 sky130_fd_sc_hs__fill_4 FILLER_22_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_387 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_395 ();
 sky130_fd_sc_hs__fill_2 FILLER_22_403 ();
 sky130_fd_sc_hs__fill_1 FILLER_22_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_409 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_417 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_425 ();
 sky130_fd_sc_hs__fill_2 FILLER_22_433 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_436 ();
 sky130_fd_sc_hs__fill_4 FILLER_22_444 ();
 sky130_fd_sc_hs__fill_2 FILLER_22_448 ();
 sky130_fd_sc_hs__fill_1 FILLER_22_450 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_457 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_481 ();
 sky130_fd_sc_hs__fill_4 FILLER_22_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_22_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_22_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_22_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_22_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_23_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_23_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_23_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_207 ();
 sky130_fd_sc_hs__fill_2 FILLER_23_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_23_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_23_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_315 ();
 sky130_fd_sc_hs__fill_4 FILLER_23_323 ();
 sky130_fd_sc_hs__fill_1 FILLER_23_327 ();
 sky130_fd_sc_hs__fill_4 FILLER_23_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_340 ();
 sky130_fd_sc_hs__fill_4 FILLER_23_349 ();
 sky130_fd_sc_hs__fill_4 FILLER_23_356 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_363 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_371 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_379 ();
 sky130_fd_sc_hs__fill_2 FILLER_23_387 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_398 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_23_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_23_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_23_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_23_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_24_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_24_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_24_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_24_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_24_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_212 ();
 sky130_fd_sc_hs__fill_4 FILLER_24_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_229 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_237 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_245 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_253 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_24_318 ();
 sky130_fd_sc_hs__fill_4 FILLER_24_320 ();
 sky130_fd_sc_hs__fill_4 FILLER_24_338 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_355 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_363 ();
 sky130_fd_sc_hs__fill_4 FILLER_24_371 ();
 sky130_fd_sc_hs__fill_2 FILLER_24_375 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_24_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_24_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_24_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_24_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_24_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_24_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_25_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_25_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_25_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_25_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_265 ();
 sky130_fd_sc_hs__fill_4 FILLER_25_273 ();
 sky130_fd_sc_hs__fill_2 FILLER_25_277 ();
 sky130_fd_sc_hs__fill_4 FILLER_25_285 ();
 sky130_fd_sc_hs__fill_1 FILLER_25_289 ();
 sky130_fd_sc_hs__fill_4 FILLER_25_291 ();
 sky130_fd_sc_hs__fill_2 FILLER_25_295 ();
 sky130_fd_sc_hs__fill_1 FILLER_25_297 ();
 sky130_fd_sc_hs__fill_4 FILLER_25_315 ();
 sky130_fd_sc_hs__fill_4 FILLER_25_325 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_332 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_340 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_25_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_25_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_25_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_25_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_25_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_26_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_26_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_26_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_26_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_26_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_26_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_294 ();
 sky130_fd_sc_hs__fill_4 FILLER_26_302 ();
 sky130_fd_sc_hs__fill_4 FILLER_26_312 ();
 sky130_fd_sc_hs__fill_2 FILLER_26_316 ();
 sky130_fd_sc_hs__fill_1 FILLER_26_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_320 ();
 sky130_fd_sc_hs__fill_2 FILLER_26_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_365 ();
 sky130_fd_sc_hs__fill_4 FILLER_26_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_26_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_26_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_26_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_26_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_26_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_26_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_27_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_27_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_27_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_27_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_27_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_307 ();
 sky130_fd_sc_hs__fill_4 FILLER_27_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_322 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_330 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_338 ();
 sky130_fd_sc_hs__fill_2 FILLER_27_346 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_27_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_415 ();
 sky130_fd_sc_hs__fill_4 FILLER_27_423 ();
 sky130_fd_sc_hs__fill_1 FILLER_27_427 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_27_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_27_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_27_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_27_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_8 ();
 sky130_fd_sc_hs__fill_4 FILLER_28_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_28_25 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_28_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_28_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_28_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_204 ();
 sky130_fd_sc_hs__fill_2 FILLER_28_212 ();
 sky130_fd_sc_hs__fill_4 FILLER_28_219 ();
 sky130_fd_sc_hs__fill_1 FILLER_28_223 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_230 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_238 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_246 ();
 sky130_fd_sc_hs__fill_4 FILLER_28_254 ();
 sky130_fd_sc_hs__fill_2 FILLER_28_258 ();
 sky130_fd_sc_hs__fill_1 FILLER_28_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_28_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_28_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_418 ();
 sky130_fd_sc_hs__fill_1 FILLER_28_426 ();
 sky130_fd_sc_hs__fill_4 FILLER_28_431 ();
 sky130_fd_sc_hs__fill_4 FILLER_28_436 ();
 sky130_fd_sc_hs__fill_4 FILLER_28_445 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_28_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_28_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_28_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_28_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_28_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_29_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_29_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_29_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_191 ();
 sky130_fd_sc_hs__fill_2 FILLER_29_199 ();
 sky130_fd_sc_hs__fill_1 FILLER_29_201 ();
 sky130_fd_sc_hs__fill_4 FILLER_29_221 ();
 sky130_fd_sc_hs__fill_4 FILLER_29_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_257 ();
 sky130_fd_sc_hs__fill_4 FILLER_29_271 ();
 sky130_fd_sc_hs__fill_2 FILLER_29_275 ();
 sky130_fd_sc_hs__fill_1 FILLER_29_277 ();
 sky130_fd_sc_hs__fill_4 FILLER_29_284 ();
 sky130_fd_sc_hs__fill_2 FILLER_29_288 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_315 ();
 sky130_fd_sc_hs__fill_4 FILLER_29_323 ();
 sky130_fd_sc_hs__fill_2 FILLER_29_327 ();
 sky130_fd_sc_hs__fill_1 FILLER_29_329 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_335 ();
 sky130_fd_sc_hs__fill_4 FILLER_29_343 ();
 sky130_fd_sc_hs__fill_1 FILLER_29_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_365 ();
 sky130_fd_sc_hs__fill_1 FILLER_29_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_377 ();
 sky130_fd_sc_hs__fill_4 FILLER_29_385 ();
 sky130_fd_sc_hs__fill_1 FILLER_29_389 ();
 sky130_fd_sc_hs__fill_4 FILLER_29_393 ();
 sky130_fd_sc_hs__fill_4 FILLER_29_401 ();
 sky130_fd_sc_hs__fill_1 FILLER_29_405 ();
 sky130_fd_sc_hs__fill_4 FILLER_29_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_414 ();
 sky130_fd_sc_hs__fill_1 FILLER_29_422 ();
 sky130_fd_sc_hs__fill_4 FILLER_29_426 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_29_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_29_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_29_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_29_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_30_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_30_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_30_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_30_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_178 ();
 sky130_fd_sc_hs__fill_4 FILLER_30_186 ();
 sky130_fd_sc_hs__fill_2 FILLER_30_190 ();
 sky130_fd_sc_hs__fill_1 FILLER_30_192 ();
 sky130_fd_sc_hs__fill_4 FILLER_30_199 ();
 sky130_fd_sc_hs__fill_4 FILLER_30_204 ();
 sky130_fd_sc_hs__fill_2 FILLER_30_208 ();
 sky130_fd_sc_hs__fill_1 FILLER_30_210 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_229 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_237 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_245 ();
 sky130_fd_sc_hs__fill_1 FILLER_30_253 ();
 sky130_fd_sc_hs__fill_4 FILLER_30_257 ();
 sky130_fd_sc_hs__fill_4 FILLER_30_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_284 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_292 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_300 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_308 ();
 sky130_fd_sc_hs__fill_2 FILLER_30_316 ();
 sky130_fd_sc_hs__fill_1 FILLER_30_318 ();
 sky130_fd_sc_hs__fill_4 FILLER_30_320 ();
 sky130_fd_sc_hs__fill_1 FILLER_30_324 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_338 ();
 sky130_fd_sc_hs__fill_4 FILLER_30_346 ();
 sky130_fd_sc_hs__fill_1 FILLER_30_350 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_30_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_378 ();
 sky130_fd_sc_hs__fill_4 FILLER_30_390 ();
 sky130_fd_sc_hs__fill_4 FILLER_30_412 ();
 sky130_fd_sc_hs__fill_2 FILLER_30_416 ();
 sky130_fd_sc_hs__fill_4 FILLER_30_422 ();
 sky130_fd_sc_hs__fill_4 FILLER_30_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_444 ();
 sky130_fd_sc_hs__fill_1 FILLER_30_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_472 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_480 ();
 sky130_fd_sc_hs__fill_4 FILLER_30_488 ();
 sky130_fd_sc_hs__fill_1 FILLER_30_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_30_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_30_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_30_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_30_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_31_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_31_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_31_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_191 ();
 sky130_fd_sc_hs__fill_2 FILLER_31_199 ();
 sky130_fd_sc_hs__fill_4 FILLER_31_219 ();
 sky130_fd_sc_hs__fill_4 FILLER_31_226 ();
 sky130_fd_sc_hs__fill_2 FILLER_31_230 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_257 ();
 sky130_fd_sc_hs__fill_2 FILLER_31_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_272 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_280 ();
 sky130_fd_sc_hs__fill_2 FILLER_31_288 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_323 ();
 sky130_fd_sc_hs__fill_1 FILLER_31_331 ();
 sky130_fd_sc_hs__fill_4 FILLER_31_337 ();
 sky130_fd_sc_hs__fill_4 FILLER_31_344 ();
 sky130_fd_sc_hs__fill_4 FILLER_31_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_366 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_374 ();
 sky130_fd_sc_hs__fill_4 FILLER_31_382 ();
 sky130_fd_sc_hs__fill_1 FILLER_31_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_396 ();
 sky130_fd_sc_hs__fill_2 FILLER_31_404 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_407 ();
 sky130_fd_sc_hs__fill_4 FILLER_31_415 ();
 sky130_fd_sc_hs__fill_2 FILLER_31_419 ();
 sky130_fd_sc_hs__fill_1 FILLER_31_421 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_425 ();
 sky130_fd_sc_hs__fill_2 FILLER_31_433 ();
 sky130_fd_sc_hs__fill_1 FILLER_31_435 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_441 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_449 ();
 sky130_fd_sc_hs__fill_4 FILLER_31_457 ();
 sky130_fd_sc_hs__fill_2 FILLER_31_461 ();
 sky130_fd_sc_hs__fill_1 FILLER_31_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_31_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_31_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_31_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_32_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_32_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_32_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_32_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_32_202 ();
 sky130_fd_sc_hs__fill_4 FILLER_32_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_214 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_222 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_230 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_238 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_246 ();
 sky130_fd_sc_hs__fill_4 FILLER_32_254 ();
 sky130_fd_sc_hs__fill_2 FILLER_32_258 ();
 sky130_fd_sc_hs__fill_1 FILLER_32_260 ();
 sky130_fd_sc_hs__fill_4 FILLER_32_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_284 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_292 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_300 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_308 ();
 sky130_fd_sc_hs__fill_2 FILLER_32_316 ();
 sky130_fd_sc_hs__fill_1 FILLER_32_318 ();
 sky130_fd_sc_hs__fill_4 FILLER_32_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_337 ();
 sky130_fd_sc_hs__fill_2 FILLER_32_345 ();
 sky130_fd_sc_hs__fill_1 FILLER_32_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_351 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_359 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_367 ();
 sky130_fd_sc_hs__fill_2 FILLER_32_375 ();
 sky130_fd_sc_hs__fill_4 FILLER_32_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_399 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_423 ();
 sky130_fd_sc_hs__fill_4 FILLER_32_431 ();
 sky130_fd_sc_hs__fill_4 FILLER_32_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_445 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_453 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_461 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_469 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_477 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_485 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_32_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_32_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_32_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_32_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_33_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_33_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_33_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_199 ();
 sky130_fd_sc_hs__fill_2 FILLER_33_207 ();
 sky130_fd_sc_hs__fill_1 FILLER_33_209 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_221 ();
 sky130_fd_sc_hs__fill_2 FILLER_33_229 ();
 sky130_fd_sc_hs__fill_1 FILLER_33_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_268 ();
 sky130_fd_sc_hs__fill_4 FILLER_33_276 ();
 sky130_fd_sc_hs__fill_4 FILLER_33_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_315 ();
 sky130_fd_sc_hs__fill_4 FILLER_33_323 ();
 sky130_fd_sc_hs__fill_2 FILLER_33_327 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_334 ();
 sky130_fd_sc_hs__fill_4 FILLER_33_342 ();
 sky130_fd_sc_hs__fill_2 FILLER_33_346 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_33_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_415 ();
 sky130_fd_sc_hs__fill_4 FILLER_33_423 ();
 sky130_fd_sc_hs__fill_2 FILLER_33_427 ();
 sky130_fd_sc_hs__fill_1 FILLER_33_429 ();
 sky130_fd_sc_hs__fill_4 FILLER_33_443 ();
 sky130_fd_sc_hs__fill_2 FILLER_33_447 ();
 sky130_fd_sc_hs__fill_1 FILLER_33_449 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_33_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_33_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_33_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_33_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_34_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_34_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_34_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_34_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_34_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_34_260 ();
 sky130_fd_sc_hs__fill_4 FILLER_34_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_281 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_297 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_305 ();
 sky130_fd_sc_hs__fill_4 FILLER_34_313 ();
 sky130_fd_sc_hs__fill_2 FILLER_34_317 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_320 ();
 sky130_fd_sc_hs__fill_2 FILLER_34_328 ();
 sky130_fd_sc_hs__fill_1 FILLER_34_330 ();
 sky130_fd_sc_hs__fill_4 FILLER_34_339 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_346 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_354 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_362 ();
 sky130_fd_sc_hs__fill_4 FILLER_34_370 ();
 sky130_fd_sc_hs__fill_2 FILLER_34_374 ();
 sky130_fd_sc_hs__fill_1 FILLER_34_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_34_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_34_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_34_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_34_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_34_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_34_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_35_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_35_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_35_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_35_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_233 ();
 sky130_fd_sc_hs__fill_4 FILLER_35_241 ();
 sky130_fd_sc_hs__fill_2 FILLER_35_245 ();
 sky130_fd_sc_hs__fill_4 FILLER_35_266 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_277 ();
 sky130_fd_sc_hs__fill_4 FILLER_35_285 ();
 sky130_fd_sc_hs__fill_1 FILLER_35_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_35_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_35_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_439 ();
 sky130_fd_sc_hs__fill_2 FILLER_35_447 ();
 sky130_fd_sc_hs__fill_4 FILLER_35_452 ();
 sky130_fd_sc_hs__fill_4 FILLER_35_459 ();
 sky130_fd_sc_hs__fill_1 FILLER_35_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_35_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_35_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_35_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_36_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_36_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_36_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_36_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_36_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_36_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_262 ();
 sky130_fd_sc_hs__fill_1 FILLER_36_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_279 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_287 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_295 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_303 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_311 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_320 ();
 sky130_fd_sc_hs__fill_1 FILLER_36_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_343 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_351 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_359 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_367 ();
 sky130_fd_sc_hs__fill_2 FILLER_36_375 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_36_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_436 ();
 sky130_fd_sc_hs__fill_4 FILLER_36_450 ();
 sky130_fd_sc_hs__fill_2 FILLER_36_454 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_462 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_470 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_478 ();
 sky130_fd_sc_hs__fill_4 FILLER_36_486 ();
 sky130_fd_sc_hs__fill_2 FILLER_36_490 ();
 sky130_fd_sc_hs__fill_1 FILLER_36_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_36_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_36_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_36_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_36_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_37_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_37_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_37_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_191 ();
 sky130_fd_sc_hs__fill_2 FILLER_37_199 ();
 sky130_fd_sc_hs__fill_1 FILLER_37_201 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_221 ();
 sky130_fd_sc_hs__fill_2 FILLER_37_229 ();
 sky130_fd_sc_hs__fill_1 FILLER_37_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_241 ();
 sky130_fd_sc_hs__fill_2 FILLER_37_249 ();
 sky130_fd_sc_hs__fill_4 FILLER_37_269 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_278 ();
 sky130_fd_sc_hs__fill_4 FILLER_37_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_307 ();
 sky130_fd_sc_hs__fill_2 FILLER_37_315 ();
 sky130_fd_sc_hs__fill_1 FILLER_37_317 ();
 sky130_fd_sc_hs__fill_4 FILLER_37_321 ();
 sky130_fd_sc_hs__fill_4 FILLER_37_328 ();
 sky130_fd_sc_hs__fill_2 FILLER_37_332 ();
 sky130_fd_sc_hs__fill_1 FILLER_37_334 ();
 sky130_fd_sc_hs__fill_4 FILLER_37_344 ();
 sky130_fd_sc_hs__fill_4 FILLER_37_349 ();
 sky130_fd_sc_hs__fill_2 FILLER_37_353 ();
 sky130_fd_sc_hs__fill_1 FILLER_37_355 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_368 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_384 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_392 ();
 sky130_fd_sc_hs__fill_4 FILLER_37_400 ();
 sky130_fd_sc_hs__fill_2 FILLER_37_404 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_423 ();
 sky130_fd_sc_hs__fill_1 FILLER_37_431 ();
 sky130_fd_sc_hs__fill_4 FILLER_37_438 ();
 sky130_fd_sc_hs__fill_4 FILLER_37_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_37_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_37_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_37_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_38_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_38_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_38_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_38_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_38_202 ();
 sky130_fd_sc_hs__fill_4 FILLER_38_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_38_260 ();
 sky130_fd_sc_hs__fill_4 FILLER_38_262 ();
 sky130_fd_sc_hs__fill_4 FILLER_38_275 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_287 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_295 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_303 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_311 ();
 sky130_fd_sc_hs__fill_4 FILLER_38_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_343 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_351 ();
 sky130_fd_sc_hs__fill_4 FILLER_38_359 ();
 sky130_fd_sc_hs__fill_2 FILLER_38_363 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_38_376 ();
 sky130_fd_sc_hs__fill_4 FILLER_38_378 ();
 sky130_fd_sc_hs__fill_4 FILLER_38_385 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_392 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_400 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_408 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_416 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_424 ();
 sky130_fd_sc_hs__fill_2 FILLER_38_432 ();
 sky130_fd_sc_hs__fill_1 FILLER_38_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_436 ();
 sky130_fd_sc_hs__fill_2 FILLER_38_444 ();
 sky130_fd_sc_hs__fill_4 FILLER_38_465 ();
 sky130_fd_sc_hs__fill_4 FILLER_38_487 ();
 sky130_fd_sc_hs__fill_2 FILLER_38_491 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_38_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_38_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_38_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_38_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_39_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_39_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_39_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_183 ();
 sky130_fd_sc_hs__fill_2 FILLER_39_191 ();
 sky130_fd_sc_hs__fill_4 FILLER_39_196 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_219 ();
 sky130_fd_sc_hs__fill_4 FILLER_39_227 ();
 sky130_fd_sc_hs__fill_1 FILLER_39_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_233 ();
 sky130_fd_sc_hs__fill_4 FILLER_39_241 ();
 sky130_fd_sc_hs__fill_2 FILLER_39_245 ();
 sky130_fd_sc_hs__fill_1 FILLER_39_247 ();
 sky130_fd_sc_hs__fill_4 FILLER_39_253 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_275 ();
 sky130_fd_sc_hs__fill_4 FILLER_39_283 ();
 sky130_fd_sc_hs__fill_2 FILLER_39_287 ();
 sky130_fd_sc_hs__fill_1 FILLER_39_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_299 ();
 sky130_fd_sc_hs__fill_1 FILLER_39_307 ();
 sky130_fd_sc_hs__fill_4 FILLER_39_314 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_337 ();
 sky130_fd_sc_hs__fill_2 FILLER_39_345 ();
 sky130_fd_sc_hs__fill_1 FILLER_39_347 ();
 sky130_fd_sc_hs__fill_4 FILLER_39_349 ();
 sky130_fd_sc_hs__fill_4 FILLER_39_361 ();
 sky130_fd_sc_hs__fill_2 FILLER_39_365 ();
 sky130_fd_sc_hs__fill_4 FILLER_39_370 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_392 ();
 sky130_fd_sc_hs__fill_4 FILLER_39_400 ();
 sky130_fd_sc_hs__fill_2 FILLER_39_404 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_423 ();
 sky130_fd_sc_hs__fill_4 FILLER_39_431 ();
 sky130_fd_sc_hs__fill_4 FILLER_39_438 ();
 sky130_fd_sc_hs__fill_4 FILLER_39_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_39_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_39_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_39_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_40_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_40_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_40_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_40_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_186 ();
 sky130_fd_sc_hs__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hs__fill_4 FILLER_40_199 ();
 sky130_fd_sc_hs__fill_4 FILLER_40_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_223 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_239 ();
 sky130_fd_sc_hs__fill_2 FILLER_40_247 ();
 sky130_fd_sc_hs__fill_4 FILLER_40_257 ();
 sky130_fd_sc_hs__fill_4 FILLER_40_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_271 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_279 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_287 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_295 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_303 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_311 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_328 ();
 sky130_fd_sc_hs__fill_1 FILLER_40_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_356 ();
 sky130_fd_sc_hs__fill_4 FILLER_40_364 ();
 sky130_fd_sc_hs__fill_2 FILLER_40_368 ();
 sky130_fd_sc_hs__fill_4 FILLER_40_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_378 ();
 sky130_fd_sc_hs__fill_1 FILLER_40_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_413 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_421 ();
 sky130_fd_sc_hs__fill_4 FILLER_40_429 ();
 sky130_fd_sc_hs__fill_2 FILLER_40_433 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_436 ();
 sky130_fd_sc_hs__fill_1 FILLER_40_444 ();
 sky130_fd_sc_hs__fill_4 FILLER_40_450 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_457 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_481 ();
 sky130_fd_sc_hs__fill_4 FILLER_40_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_40_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_40_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_40_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_40_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_41_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_41_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_41_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_175 ();
 sky130_fd_sc_hs__fill_4 FILLER_41_183 ();
 sky130_fd_sc_hs__fill_2 FILLER_41_187 ();
 sky130_fd_sc_hs__fill_1 FILLER_41_189 ();
 sky130_fd_sc_hs__fill_4 FILLER_41_193 ();
 sky130_fd_sc_hs__fill_4 FILLER_41_217 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_224 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_271 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_279 ();
 sky130_fd_sc_hs__fill_2 FILLER_41_287 ();
 sky130_fd_sc_hs__fill_1 FILLER_41_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_307 ();
 sky130_fd_sc_hs__fill_4 FILLER_41_315 ();
 sky130_fd_sc_hs__fill_4 FILLER_41_322 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_335 ();
 sky130_fd_sc_hs__fill_4 FILLER_41_343 ();
 sky130_fd_sc_hs__fill_1 FILLER_41_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_357 ();
 sky130_fd_sc_hs__fill_4 FILLER_41_365 ();
 sky130_fd_sc_hs__fill_4 FILLER_41_387 ();
 sky130_fd_sc_hs__fill_2 FILLER_41_391 ();
 sky130_fd_sc_hs__fill_1 FILLER_41_393 ();
 sky130_fd_sc_hs__fill_4 FILLER_41_400 ();
 sky130_fd_sc_hs__fill_2 FILLER_41_404 ();
 sky130_fd_sc_hs__fill_4 FILLER_41_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_414 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_422 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_430 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_438 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_446 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_454 ();
 sky130_fd_sc_hs__fill_2 FILLER_41_462 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_41_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_41_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_41_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_42_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_42_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_42_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_42_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_170 ();
 sky130_fd_sc_hs__fill_2 FILLER_42_178 ();
 sky130_fd_sc_hs__fill_1 FILLER_42_180 ();
 sky130_fd_sc_hs__fill_4 FILLER_42_199 ();
 sky130_fd_sc_hs__fill_4 FILLER_42_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_213 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_221 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_229 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_237 ();
 sky130_fd_sc_hs__fill_4 FILLER_42_245 ();
 sky130_fd_sc_hs__fill_2 FILLER_42_249 ();
 sky130_fd_sc_hs__fill_1 FILLER_42_251 ();
 sky130_fd_sc_hs__fill_4 FILLER_42_257 ();
 sky130_fd_sc_hs__fill_4 FILLER_42_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_283 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_307 ();
 sky130_fd_sc_hs__fill_4 FILLER_42_315 ();
 sky130_fd_sc_hs__fill_4 FILLER_42_320 ();
 sky130_fd_sc_hs__fill_2 FILLER_42_324 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_339 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_355 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_363 ();
 sky130_fd_sc_hs__fill_4 FILLER_42_371 ();
 sky130_fd_sc_hs__fill_2 FILLER_42_375 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_378 ();
 sky130_fd_sc_hs__fill_2 FILLER_42_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_413 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_421 ();
 sky130_fd_sc_hs__fill_4 FILLER_42_429 ();
 sky130_fd_sc_hs__fill_2 FILLER_42_433 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_42_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_42_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_42_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_42_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_42_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_43_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_43_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_43_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_183 ();
 sky130_fd_sc_hs__fill_4 FILLER_43_197 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_220 ();
 sky130_fd_sc_hs__fill_4 FILLER_43_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_257 ();
 sky130_fd_sc_hs__fill_1 FILLER_43_265 ();
 sky130_fd_sc_hs__fill_4 FILLER_43_271 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_280 ();
 sky130_fd_sc_hs__fill_2 FILLER_43_288 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_43_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_381 ();
 sky130_fd_sc_hs__fill_4 FILLER_43_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_396 ();
 sky130_fd_sc_hs__fill_2 FILLER_43_404 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_43_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_43_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_43_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_43_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_44_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_44_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_44_86 ();
 sky130_fd_sc_hs__fill_4 FILLER_44_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_95 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_103 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_111 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_119 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_127 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_135 ();
 sky130_fd_sc_hs__fill_2 FILLER_44_143 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_178 ();
 sky130_fd_sc_hs__fill_4 FILLER_44_186 ();
 sky130_fd_sc_hs__fill_2 FILLER_44_190 ();
 sky130_fd_sc_hs__fill_1 FILLER_44_192 ();
 sky130_fd_sc_hs__fill_4 FILLER_44_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_244 ();
 sky130_fd_sc_hs__fill_2 FILLER_44_252 ();
 sky130_fd_sc_hs__fill_4 FILLER_44_257 ();
 sky130_fd_sc_hs__fill_4 FILLER_44_262 ();
 sky130_fd_sc_hs__fill_1 FILLER_44_266 ();
 sky130_fd_sc_hs__fill_4 FILLER_44_275 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_285 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_293 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_301 ();
 sky130_fd_sc_hs__fill_4 FILLER_44_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_44_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_44_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_44_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_44_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_44_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_44_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_44_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_45_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_45_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_45_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_45_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_257 ();
 sky130_fd_sc_hs__fill_1 FILLER_45_265 ();
 sky130_fd_sc_hs__fill_4 FILLER_45_269 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_276 ();
 sky130_fd_sc_hs__fill_4 FILLER_45_284 ();
 sky130_fd_sc_hs__fill_2 FILLER_45_288 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_323 ();
 sky130_fd_sc_hs__fill_4 FILLER_45_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_338 ();
 sky130_fd_sc_hs__fill_2 FILLER_45_346 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_45_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_440 ();
 sky130_fd_sc_hs__fill_2 FILLER_45_448 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_453 ();
 sky130_fd_sc_hs__fill_2 FILLER_45_461 ();
 sky130_fd_sc_hs__fill_1 FILLER_45_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_45_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_45_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_45_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_46_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_46_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_46_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_46_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_46_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_46_260 ();
 sky130_fd_sc_hs__fill_4 FILLER_46_262 ();
 sky130_fd_sc_hs__fill_2 FILLER_46_266 ();
 sky130_fd_sc_hs__fill_1 FILLER_46_268 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_275 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_283 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_307 ();
 sky130_fd_sc_hs__fill_4 FILLER_46_315 ();
 sky130_fd_sc_hs__fill_4 FILLER_46_320 ();
 sky130_fd_sc_hs__fill_4 FILLER_46_327 ();
 sky130_fd_sc_hs__fill_2 FILLER_46_331 ();
 sky130_fd_sc_hs__fill_4 FILLER_46_342 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_365 ();
 sky130_fd_sc_hs__fill_4 FILLER_46_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_378 ();
 sky130_fd_sc_hs__fill_4 FILLER_46_386 ();
 sky130_fd_sc_hs__fill_1 FILLER_46_390 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_396 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_404 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_412 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_420 ();
 sky130_fd_sc_hs__fill_4 FILLER_46_428 ();
 sky130_fd_sc_hs__fill_2 FILLER_46_432 ();
 sky130_fd_sc_hs__fill_1 FILLER_46_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_46_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_46_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_46_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_46_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_46_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_47_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_47_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_47_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_47_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_249 ();
 sky130_fd_sc_hs__fill_2 FILLER_47_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_277 ();
 sky130_fd_sc_hs__fill_4 FILLER_47_285 ();
 sky130_fd_sc_hs__fill_1 FILLER_47_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_299 ();
 sky130_fd_sc_hs__fill_4 FILLER_47_307 ();
 sky130_fd_sc_hs__fill_2 FILLER_47_311 ();
 sky130_fd_sc_hs__fill_4 FILLER_47_330 ();
 sky130_fd_sc_hs__fill_2 FILLER_47_334 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_47_347 ();
 sky130_fd_sc_hs__fill_4 FILLER_47_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_365 ();
 sky130_fd_sc_hs__fill_4 FILLER_47_373 ();
 sky130_fd_sc_hs__fill_2 FILLER_47_377 ();
 sky130_fd_sc_hs__fill_1 FILLER_47_379 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_47_405 ();
 sky130_fd_sc_hs__fill_4 FILLER_47_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_414 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_422 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_430 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_438 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_446 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_454 ();
 sky130_fd_sc_hs__fill_2 FILLER_47_462 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_47_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_47_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_47_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_48_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_48_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_48_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_48_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_48_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_48_260 ();
 sky130_fd_sc_hs__fill_4 FILLER_48_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_284 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_292 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_300 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_308 ();
 sky130_fd_sc_hs__fill_2 FILLER_48_316 ();
 sky130_fd_sc_hs__fill_1 FILLER_48_318 ();
 sky130_fd_sc_hs__fill_4 FILLER_48_320 ();
 sky130_fd_sc_hs__fill_4 FILLER_48_330 ();
 sky130_fd_sc_hs__fill_4 FILLER_48_337 ();
 sky130_fd_sc_hs__fill_2 FILLER_48_341 ();
 sky130_fd_sc_hs__fill_1 FILLER_48_343 ();
 sky130_fd_sc_hs__fill_4 FILLER_48_362 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_369 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_402 ();
 sky130_fd_sc_hs__fill_4 FILLER_48_430 ();
 sky130_fd_sc_hs__fill_1 FILLER_48_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_48_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_48_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_48_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_48_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_48_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_49_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_49_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_49_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_49_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_257 ();
 sky130_fd_sc_hs__fill_4 FILLER_49_265 ();
 sky130_fd_sc_hs__fill_4 FILLER_49_274 ();
 sky130_fd_sc_hs__fill_2 FILLER_49_278 ();
 sky130_fd_sc_hs__fill_4 FILLER_49_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_307 ();
 sky130_fd_sc_hs__fill_4 FILLER_49_315 ();
 sky130_fd_sc_hs__fill_2 FILLER_49_319 ();
 sky130_fd_sc_hs__fill_1 FILLER_49_321 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_325 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_333 ();
 sky130_fd_sc_hs__fill_4 FILLER_49_341 ();
 sky130_fd_sc_hs__fill_2 FILLER_49_345 ();
 sky130_fd_sc_hs__fill_1 FILLER_49_347 ();
 sky130_fd_sc_hs__fill_4 FILLER_49_349 ();
 sky130_fd_sc_hs__fill_2 FILLER_49_353 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_359 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_367 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_375 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_383 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_391 ();
 sky130_fd_sc_hs__fill_4 FILLER_49_399 ();
 sky130_fd_sc_hs__fill_2 FILLER_49_403 ();
 sky130_fd_sc_hs__fill_1 FILLER_49_405 ();
 sky130_fd_sc_hs__fill_4 FILLER_49_407 ();
 sky130_fd_sc_hs__fill_4 FILLER_49_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_428 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_452 ();
 sky130_fd_sc_hs__fill_4 FILLER_49_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_49_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_49_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_49_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_50_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_50_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_50_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_50_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_50_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_218 ();
 sky130_fd_sc_hs__fill_4 FILLER_50_226 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_50_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_270 ();
 sky130_fd_sc_hs__fill_4 FILLER_50_278 ();
 sky130_fd_sc_hs__fill_2 FILLER_50_282 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_290 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_298 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_306 ();
 sky130_fd_sc_hs__fill_4 FILLER_50_314 ();
 sky130_fd_sc_hs__fill_1 FILLER_50_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_50_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_394 ();
 sky130_fd_sc_hs__fill_4 FILLER_50_402 ();
 sky130_fd_sc_hs__fill_1 FILLER_50_406 ();
 sky130_fd_sc_hs__fill_4 FILLER_50_410 ();
 sky130_fd_sc_hs__fill_4 FILLER_50_431 ();
 sky130_fd_sc_hs__fill_4 FILLER_50_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_445 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_453 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_461 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_469 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_477 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_485 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_50_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_50_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_50_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_50_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_33 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_41 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_49 ();
 sky130_fd_sc_hs__fill_1 FILLER_51_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_51_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_51_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_199 ();
 sky130_fd_sc_hs__fill_2 FILLER_51_207 ();
 sky130_fd_sc_hs__fill_1 FILLER_51_209 ();
 sky130_fd_sc_hs__fill_4 FILLER_51_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_51_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_51_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_349 ();
 sky130_fd_sc_hs__fill_4 FILLER_51_357 ();
 sky130_fd_sc_hs__fill_2 FILLER_51_361 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_370 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_394 ();
 sky130_fd_sc_hs__fill_4 FILLER_51_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_426 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_442 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_450 ();
 sky130_fd_sc_hs__fill_4 FILLER_51_458 ();
 sky130_fd_sc_hs__fill_2 FILLER_51_462 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_51_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_51_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_51_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_52_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_52_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_52_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_52_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_52_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_204 ();
 sky130_fd_sc_hs__fill_4 FILLER_52_232 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_239 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_247 ();
 sky130_fd_sc_hs__fill_4 FILLER_52_255 ();
 sky130_fd_sc_hs__fill_2 FILLER_52_259 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_52_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_360 ();
 sky130_fd_sc_hs__fill_2 FILLER_52_368 ();
 sky130_fd_sc_hs__fill_4 FILLER_52_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_394 ();
 sky130_fd_sc_hs__fill_2 FILLER_52_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_407 ();
 sky130_fd_sc_hs__fill_2 FILLER_52_415 ();
 sky130_fd_sc_hs__fill_1 FILLER_52_417 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_422 ();
 sky130_fd_sc_hs__fill_4 FILLER_52_430 ();
 sky130_fd_sc_hs__fill_1 FILLER_52_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_52_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_52_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_52_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_52_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_52_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_53_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_53_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_53_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_199 ();
 sky130_fd_sc_hs__fill_4 FILLER_53_207 ();
 sky130_fd_sc_hs__fill_4 FILLER_53_216 ();
 sky130_fd_sc_hs__fill_4 FILLER_53_226 ();
 sky130_fd_sc_hs__fill_2 FILLER_53_230 ();
 sky130_fd_sc_hs__fill_4 FILLER_53_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_256 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_264 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_272 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_280 ();
 sky130_fd_sc_hs__fill_2 FILLER_53_288 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_53_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_389 ();
 sky130_fd_sc_hs__fill_4 FILLER_53_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_53_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_53_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_53_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_53_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_54_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_54_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_54_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_54_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_54_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_54_231 ();
 sky130_fd_sc_hs__fill_4 FILLER_54_235 ();
 sky130_fd_sc_hs__fill_4 FILLER_54_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_307 ();
 sky130_fd_sc_hs__fill_4 FILLER_54_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_54_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_422 ();
 sky130_fd_sc_hs__fill_4 FILLER_54_430 ();
 sky130_fd_sc_hs__fill_1 FILLER_54_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_54_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_54_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_54_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_54_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_54_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_55_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_55_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_55_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_55_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_265 ();
 sky130_fd_sc_hs__fill_2 FILLER_55_273 ();
 sky130_fd_sc_hs__fill_1 FILLER_55_275 ();
 sky130_fd_sc_hs__fill_4 FILLER_55_279 ();
 sky130_fd_sc_hs__fill_4 FILLER_55_286 ();
 sky130_fd_sc_hs__fill_4 FILLER_55_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_312 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_336 ();
 sky130_fd_sc_hs__fill_4 FILLER_55_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_55_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_55_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_55_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_55_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_55_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_56_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_56_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_56_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_56_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_56_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_56_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_262 ();
 sky130_fd_sc_hs__fill_4 FILLER_56_270 ();
 sky130_fd_sc_hs__fill_2 FILLER_56_274 ();
 sky130_fd_sc_hs__fill_4 FILLER_56_281 ();
 sky130_fd_sc_hs__fill_4 FILLER_56_293 ();
 sky130_fd_sc_hs__fill_4 FILLER_56_302 ();
 sky130_fd_sc_hs__fill_4 FILLER_56_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_352 ();
 sky130_fd_sc_hs__fill_4 FILLER_56_360 ();
 sky130_fd_sc_hs__fill_2 FILLER_56_364 ();
 sky130_fd_sc_hs__fill_4 FILLER_56_372 ();
 sky130_fd_sc_hs__fill_1 FILLER_56_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_56_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_56_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_56_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_56_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_56_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_56_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_57_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_57_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_57_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_57_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_265 ();
 sky130_fd_sc_hs__fill_4 FILLER_57_273 ();
 sky130_fd_sc_hs__fill_4 FILLER_57_286 ();
 sky130_fd_sc_hs__fill_4 FILLER_57_291 ();
 sky130_fd_sc_hs__fill_1 FILLER_57_295 ();
 sky130_fd_sc_hs__fill_4 FILLER_57_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_321 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_329 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_337 ();
 sky130_fd_sc_hs__fill_2 FILLER_57_345 ();
 sky130_fd_sc_hs__fill_1 FILLER_57_347 ();
 sky130_fd_sc_hs__fill_4 FILLER_57_349 ();
 sky130_fd_sc_hs__fill_2 FILLER_57_353 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_373 ();
 sky130_fd_sc_hs__fill_1 FILLER_57_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_57_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_415 ();
 sky130_fd_sc_hs__fill_2 FILLER_57_423 ();
 sky130_fd_sc_hs__fill_1 FILLER_57_425 ();
 sky130_fd_sc_hs__fill_4 FILLER_57_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_454 ();
 sky130_fd_sc_hs__fill_2 FILLER_57_462 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_57_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_57_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_57_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_58_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_58_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_58_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_58_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_58_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_58_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_270 ();
 sky130_fd_sc_hs__fill_2 FILLER_58_278 ();
 sky130_fd_sc_hs__fill_4 FILLER_58_285 ();
 sky130_fd_sc_hs__fill_4 FILLER_58_294 ();
 sky130_fd_sc_hs__fill_4 FILLER_58_303 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_58_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_328 ();
 sky130_fd_sc_hs__fill_4 FILLER_58_336 ();
 sky130_fd_sc_hs__fill_2 FILLER_58_340 ();
 sky130_fd_sc_hs__fill_1 FILLER_58_342 ();
 sky130_fd_sc_hs__fill_4 FILLER_58_362 ();
 sky130_fd_sc_hs__fill_4 FILLER_58_371 ();
 sky130_fd_sc_hs__fill_2 FILLER_58_375 ();
 sky130_fd_sc_hs__fill_4 FILLER_58_378 ();
 sky130_fd_sc_hs__fill_2 FILLER_58_382 ();
 sky130_fd_sc_hs__fill_4 FILLER_58_392 ();
 sky130_fd_sc_hs__fill_1 FILLER_58_396 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_413 ();
 sky130_fd_sc_hs__fill_4 FILLER_58_421 ();
 sky130_fd_sc_hs__fill_4 FILLER_58_431 ();
 sky130_fd_sc_hs__fill_4 FILLER_58_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_445 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_453 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_461 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_469 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_477 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_485 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_58_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_58_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_58_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_58_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_59_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_59_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_59_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_199 ();
 sky130_fd_sc_hs__fill_4 FILLER_59_207 ();
 sky130_fd_sc_hs__fill_1 FILLER_59_211 ();
 sky130_fd_sc_hs__fill_4 FILLER_59_218 ();
 sky130_fd_sc_hs__fill_4 FILLER_59_227 ();
 sky130_fd_sc_hs__fill_1 FILLER_59_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_233 ();
 sky130_fd_sc_hs__fill_2 FILLER_59_241 ();
 sky130_fd_sc_hs__fill_1 FILLER_59_243 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_249 ();
 sky130_fd_sc_hs__fill_4 FILLER_59_257 ();
 sky130_fd_sc_hs__fill_2 FILLER_59_261 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_268 ();
 sky130_fd_sc_hs__fill_2 FILLER_59_276 ();
 sky130_fd_sc_hs__fill_1 FILLER_59_278 ();
 sky130_fd_sc_hs__fill_4 FILLER_59_284 ();
 sky130_fd_sc_hs__fill_2 FILLER_59_288 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_291 ();
 sky130_fd_sc_hs__fill_2 FILLER_59_299 ();
 sky130_fd_sc_hs__fill_1 FILLER_59_301 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_310 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_326 ();
 sky130_fd_sc_hs__fill_4 FILLER_59_334 ();
 sky130_fd_sc_hs__fill_4 FILLER_59_344 ();
 sky130_fd_sc_hs__fill_4 FILLER_59_349 ();
 sky130_fd_sc_hs__fill_4 FILLER_59_371 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_59_405 ();
 sky130_fd_sc_hs__fill_4 FILLER_59_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_429 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_443 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_451 ();
 sky130_fd_sc_hs__fill_4 FILLER_59_459 ();
 sky130_fd_sc_hs__fill_1 FILLER_59_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_59_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_59_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_59_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_60_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_60_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_60_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_60_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_60_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_204 ();
 sky130_fd_sc_hs__fill_2 FILLER_60_212 ();
 sky130_fd_sc_hs__fill_4 FILLER_60_232 ();
 sky130_fd_sc_hs__fill_4 FILLER_60_239 ();
 sky130_fd_sc_hs__fill_2 FILLER_60_243 ();
 sky130_fd_sc_hs__fill_1 FILLER_60_245 ();
 sky130_fd_sc_hs__fill_4 FILLER_60_254 ();
 sky130_fd_sc_hs__fill_2 FILLER_60_258 ();
 sky130_fd_sc_hs__fill_1 FILLER_60_260 ();
 sky130_fd_sc_hs__fill_4 FILLER_60_262 ();
 sky130_fd_sc_hs__fill_2 FILLER_60_266 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_275 ();
 sky130_fd_sc_hs__fill_2 FILLER_60_283 ();
 sky130_fd_sc_hs__fill_1 FILLER_60_285 ();
 sky130_fd_sc_hs__fill_4 FILLER_60_291 ();
 sky130_fd_sc_hs__fill_2 FILLER_60_295 ();
 sky130_fd_sc_hs__fill_4 FILLER_60_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_328 ();
 sky130_fd_sc_hs__fill_4 FILLER_60_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_60_343 ();
 sky130_fd_sc_hs__fill_4 FILLER_60_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_369 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_410 ();
 sky130_fd_sc_hs__fill_1 FILLER_60_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_424 ();
 sky130_fd_sc_hs__fill_2 FILLER_60_432 ();
 sky130_fd_sc_hs__fill_1 FILLER_60_434 ();
 sky130_fd_sc_hs__fill_4 FILLER_60_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_443 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_451 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_459 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_467 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_475 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_483 ();
 sky130_fd_sc_hs__fill_2 FILLER_60_491 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_60_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_60_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_60_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_60_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_61_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_61_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_61_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_199 ();
 sky130_fd_sc_hs__fill_4 FILLER_61_207 ();
 sky130_fd_sc_hs__fill_4 FILLER_61_228 ();
 sky130_fd_sc_hs__fill_4 FILLER_61_233 ();
 sky130_fd_sc_hs__fill_1 FILLER_61_237 ();
 sky130_fd_sc_hs__fill_4 FILLER_61_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_248 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_256 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_264 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_272 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_280 ();
 sky130_fd_sc_hs__fill_2 FILLER_61_288 ();
 sky130_fd_sc_hs__fill_4 FILLER_61_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_298 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_306 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_314 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_322 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_330 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_338 ();
 sky130_fd_sc_hs__fill_2 FILLER_61_346 ();
 sky130_fd_sc_hs__fill_4 FILLER_61_349 ();
 sky130_fd_sc_hs__fill_2 FILLER_61_353 ();
 sky130_fd_sc_hs__fill_1 FILLER_61_355 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_359 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_367 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_375 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_383 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_391 ();
 sky130_fd_sc_hs__fill_4 FILLER_61_399 ();
 sky130_fd_sc_hs__fill_2 FILLER_61_403 ();
 sky130_fd_sc_hs__fill_1 FILLER_61_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_61_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_61_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_61_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_61_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_62_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_62_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_62_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_62_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_62_202 ();
 sky130_fd_sc_hs__fill_4 FILLER_62_204 ();
 sky130_fd_sc_hs__fill_2 FILLER_62_208 ();
 sky130_fd_sc_hs__fill_4 FILLER_62_216 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_226 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_234 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_242 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_250 ();
 sky130_fd_sc_hs__fill_2 FILLER_62_258 ();
 sky130_fd_sc_hs__fill_1 FILLER_62_260 ();
 sky130_fd_sc_hs__fill_4 FILLER_62_262 ();
 sky130_fd_sc_hs__fill_2 FILLER_62_266 ();
 sky130_fd_sc_hs__fill_1 FILLER_62_268 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_287 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_295 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_303 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_311 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_62_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_62_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_62_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_62_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_62_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_62_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_62_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_63_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_63_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_63_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_63_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_63_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_63_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_63_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_63_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_63_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_63_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_63_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_64_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_64_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_64_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_64_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_64_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_64_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_64_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_64_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_64_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_64_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_64_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_64_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_64_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_64_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_65_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_65_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_65_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_65_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_65_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_65_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_65_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_65_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_65_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_65_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_65_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_66_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_66_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_66_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_66_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_66_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_66_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_66_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_66_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_66_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_66_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_66_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_66_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_66_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_66_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_67_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_67_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_67_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_67_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_67_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_67_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_67_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_67_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_67_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_67_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_67_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_68_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_68_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_68_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_68_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_68_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_68_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_68_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_68_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_68_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_68_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_68_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_68_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_68_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_68_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_69_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_69_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_69_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_69_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_69_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_69_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_69_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_69_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_69_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_69_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_69_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_70_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_70_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_70_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_70_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_70_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_70_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_70_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_70_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_70_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_70_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_70_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_70_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_70_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_70_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_71_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_71_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_71_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_71_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_71_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_71_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_71_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_71_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_71_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_71_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_71_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_72_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_72_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_72_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_72_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_72_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_72_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_72_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_72_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_72_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_72_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_72_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_72_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_72_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_72_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_73_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_73_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_73_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_73_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_73_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_73_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_73_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_73_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_73_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_73_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_73_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_74_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_74_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_74_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_74_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_74_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_74_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_74_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_74_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_74_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_74_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_74_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_74_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_74_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_74_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_75_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_75_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_75_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_75_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_75_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_75_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_75_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_75_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_75_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_75_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_75_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_76_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_76_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_76_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_76_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_76_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_76_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_76_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_76_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_76_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_76_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_76_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_76_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_76_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_76_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_77_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_77_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_77_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_77_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_77_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_77_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_77_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_77_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_77_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_77_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_77_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_78_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_78_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_78_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_78_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_78_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_78_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_78_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_78_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_78_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_78_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_78_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_78_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_78_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_78_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_79_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_79_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_79_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_79_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_79_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_79_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_79_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_79_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_79_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_79_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_79_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_80_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_80_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_80_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_80_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_80_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_80_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_80_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_80_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_80_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_80_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_526 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_534 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_542 ();
 sky130_fd_sc_hs__fill_1 FILLER_80_550 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_80_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_80_580 ();
 sky130_fd_sc_hs__fill_1 FILLER_80_582 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_81_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_81_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_81_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_81_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_81_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_81_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_81_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_81_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_81_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_555 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_563 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_571 ();
 sky130_fd_sc_hs__fill_1 FILLER_81_579 ();
 sky130_fd_sc_hs__fill_2 FILLER_81_581 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_82_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_82_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_46 ();
 sky130_fd_sc_hs__fill_4 FILLER_82_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_75 ();
 sky130_fd_sc_hs__fill_4 FILLER_82_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_104 ();
 sky130_fd_sc_hs__fill_4 FILLER_82_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_133 ();
 sky130_fd_sc_hs__fill_4 FILLER_82_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_162 ();
 sky130_fd_sc_hs__fill_4 FILLER_82_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_191 ();
 sky130_fd_sc_hs__fill_4 FILLER_82_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_220 ();
 sky130_fd_sc_hs__fill_4 FILLER_82_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_249 ();
 sky130_fd_sc_hs__fill_4 FILLER_82_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_278 ();
 sky130_fd_sc_hs__fill_4 FILLER_82_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_307 ();
 sky130_fd_sc_hs__fill_4 FILLER_82_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_336 ();
 sky130_fd_sc_hs__fill_4 FILLER_82_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_365 ();
 sky130_fd_sc_hs__fill_4 FILLER_82_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_394 ();
 sky130_fd_sc_hs__fill_4 FILLER_82_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_423 ();
 sky130_fd_sc_hs__fill_4 FILLER_82_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_452 ();
 sky130_fd_sc_hs__fill_4 FILLER_82_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_481 ();
 sky130_fd_sc_hs__fill_4 FILLER_82_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_510 ();
 sky130_fd_sc_hs__fill_4 FILLER_82_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_539 ();
 sky130_fd_sc_hs__fill_4 FILLER_82_547 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_552 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_560 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_568 ();
 sky130_fd_sc_hs__fill_4 FILLER_82_576 ();
 sky130_fd_sc_hs__fill_2 FILLER_82_581 ();
endmodule
