VERSION 5.8 ;

SITE IOSite
  CLASS       PAD ;
  SYMMETRY    X Y R90 ;
  SIZE        0.010 BY 80.000 ;
END IOSite

SITE CornerSite
  CLASS       PAD ;
  SYMMETRY    X Y R90 ;
  SIZE        80.000 BY 80.000 ;
END CornerSite

MACRO PPAD_LONG
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN PPAD_LONG 0 0 ;
  SIZE 55 BY 80 ;
  SYMMETRY X Y R90 ;
  SITE IOSite ;
  PIN VDD
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.755 75.635 4.445 80 ;
        RECT 6.355 75.635 7.045 80 ;
        RECT 8.955 75.635 9.645 80 ;
        RECT 11.555 75.635 12.245 80 ;
        RECT 14.155 75.635 14.845 80 ;
        RECT 16.755 75.635 17.445 80 ;
        RECT 19.355 75.635 20.045 80 ;
        RECT 21.955 75.635 22.645 80 ;
        RECT 24.555 75.635 25.245 80 ;
        RECT 27.155 75.635 27.845 80 ;
        RECT 29.755 75.635 30.445 80 ;
        RECT 32.355 75.635 33.045 80 ;
        RECT 34.955 75.635 35.645 80 ;
        RECT 37.555 75.635 38.245 80 ;
        RECT 40.155 75.635 40.845 80 ;
        RECT 42.755 75.635 43.445 80 ;
        RECT 45.355 75.635 46.045 80 ;
        RECT 47.955 75.635 48.645 80 ;
        RECT 3.28 77.9 50.735 80 ;
        RECT 50.555 75.635 51.245 78.86 ;
      LAYER metal2 ;
        RECT 3.755 75.635 4.445 80 ;
        RECT 6.355 75.635 7.045 80 ;
        RECT 8.955 75.635 9.645 80 ;
        RECT 11.555 75.635 12.245 80 ;
        RECT 14.155 75.635 14.845 80 ;
        RECT 16.755 75.635 17.445 80 ;
        RECT 19.355 75.635 20.045 80 ;
        RECT 21.955 75.635 22.645 80 ;
        RECT 24.555 75.635 25.245 80 ;
        RECT 27.155 75.635 27.845 80 ;
        RECT 29.755 75.635 30.445 80 ;
        RECT 32.355 75.635 33.045 80 ;
        RECT 34.955 75.635 35.645 80 ;
        RECT 37.555 75.635 38.245 80 ;
        RECT 40.155 75.635 40.845 80 ;
        RECT 42.755 75.635 43.445 80 ;
        RECT 45.355 75.635 46.045 80 ;
        RECT 47.955 75.635 48.645 80 ;
        RECT 3.28 77.9 50.735 80 ;
        RECT 50.555 75.635 51.245 78.86 ;
      LAYER metal3 ;
        RECT 3.755 75.635 4.445 80 ;
        RECT 6.355 75.635 7.045 80 ;
        RECT 8.955 75.635 9.645 80 ;
        RECT 11.555 75.635 12.245 80 ;
        RECT 14.155 75.635 14.845 80 ;
        RECT 16.755 75.635 17.445 80 ;
        RECT 19.355 75.635 20.045 80 ;
        RECT 21.955 75.635 22.645 80 ;
        RECT 24.555 75.635 25.245 80 ;
        RECT 27.155 75.635 27.845 80 ;
        RECT 29.755 75.635 30.445 80 ;
        RECT 32.355 75.635 33.045 80 ;
        RECT 34.955 75.635 35.645 80 ;
        RECT 37.555 75.635 38.245 80 ;
        RECT 40.155 75.635 40.845 80 ;
        RECT 42.755 75.635 43.445 80 ;
        RECT 45.355 75.635 46.045 80 ;
        RECT 47.955 75.635 48.645 80 ;
        RECT 3.28 77.9 50.735 80 ;
        RECT 50.555 75.635 51.245 78.86 ;
      LAYER metal4 ;
        RECT 3.755 75.635 4.445 80 ;
        RECT 6.355 75.635 7.045 80 ;
        RECT 8.955 75.635 9.645 80 ;
        RECT 11.555 75.635 12.245 80 ;
        RECT 14.155 75.635 14.845 80 ;
        RECT 16.755 75.635 17.445 80 ;
        RECT 19.355 75.635 20.045 80 ;
        RECT 21.955 75.635 22.645 80 ;
        RECT 24.555 75.635 25.245 80 ;
        RECT 27.155 75.635 27.845 80 ;
        RECT 29.755 75.635 30.445 80 ;
        RECT 32.355 75.635 33.045 80 ;
        RECT 34.955 75.635 35.645 80 ;
        RECT 37.555 75.635 38.245 80 ;
        RECT 40.155 75.635 40.845 80 ;
        RECT 42.755 75.635 43.445 80 ;
        RECT 45.355 75.635 46.045 80 ;
        RECT 47.955 75.635 48.645 80 ;
        RECT 3.28 77.9 50.735 80 ;
        RECT 50.555 75.635 51.245 78.86 ;
    END
  END VDD
END PPAD_LONG

MACRO PPAD_SHORT
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN PPAD_SHORT 0 0 ;
  SIZE 55 BY 80 ;
  SYMMETRY X Y R90 ;
  SITE IOSite ;
  PIN VDD
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.755 75.635 4.445 80 ;
        RECT 6.355 75.635 7.045 80 ;
        RECT 8.955 75.635 9.645 80 ;
        RECT 11.555 75.635 12.245 80 ;
        RECT 14.155 75.635 14.845 80 ;
        RECT 16.755 75.635 17.445 80 ;
        RECT 19.355 75.635 20.045 80 ;
        RECT 21.955 75.635 22.645 80 ;
        RECT 24.555 75.635 25.245 80 ;
        RECT 27.155 75.635 27.845 80 ;
        RECT 29.755 75.635 30.445 80 ;
        RECT 32.355 75.635 33.045 80 ;
        RECT 34.955 75.635 35.645 80 ;
        RECT 37.555 75.635 38.245 80 ;
        RECT 40.155 75.635 40.845 80 ;
        RECT 42.755 75.635 43.445 80 ;
        RECT 45.355 75.635 46.045 80 ;
        RECT 47.955 75.635 48.645 80 ;
        RECT 50.555 75.635 51.245 78.86 ;
      LAYER metal2 ;
        RECT 3.755 75.635 4.445 80 ;
        RECT 6.355 75.635 7.045 80 ;
        RECT 8.955 75.635 9.645 80 ;
        RECT 11.555 75.635 12.245 80 ;
        RECT 14.155 75.635 14.845 80 ;
        RECT 16.755 75.635 17.445 80 ;
        RECT 19.355 75.635 20.045 80 ;
        RECT 21.955 75.635 22.645 80 ;
        RECT 24.555 75.635 25.245 80 ;
        RECT 27.155 75.635 27.845 80 ;
        RECT 29.755 75.635 30.445 80 ;
        RECT 32.355 75.635 33.045 80 ;
        RECT 34.955 75.635 35.645 80 ;
        RECT 37.555 75.635 38.245 80 ;
        RECT 40.155 75.635 40.845 80 ;
        RECT 42.755 75.635 43.445 80 ;
        RECT 45.355 75.635 46.045 80 ;
        RECT 47.955 75.635 48.645 80 ;
        RECT 50.555 75.635 51.245 78.86 ;
      LAYER metal3 ;
        RECT 3.755 75.635 4.445 80 ;
        RECT 6.355 75.635 7.045 80 ;
        RECT 8.955 75.635 9.645 80 ;
        RECT 11.555 75.635 12.245 80 ;
        RECT 14.155 75.635 14.845 80 ;
        RECT 16.755 75.635 17.445 80 ;
        RECT 19.355 75.635 20.045 80 ;
        RECT 21.955 75.635 22.645 80 ;
        RECT 24.555 75.635 25.245 80 ;
        RECT 27.155 75.635 27.845 80 ;
        RECT 29.755 75.635 30.445 80 ;
        RECT 32.355 75.635 33.045 80 ;
        RECT 34.955 75.635 35.645 80 ;
        RECT 37.555 75.635 38.245 80 ;
        RECT 40.155 75.635 40.845 80 ;
        RECT 42.755 75.635 43.445 80 ;
        RECT 45.355 75.635 46.045 80 ;
        RECT 47.955 75.635 48.645 80 ;
        RECT 50.555 75.635 51.245 78.86 ;
      LAYER metal4 ;
        RECT 3.755 75.635 4.445 80 ;
        RECT 6.355 75.635 7.045 80 ;
        RECT 8.955 75.635 9.645 80 ;
        RECT 11.555 75.635 12.245 80 ;
        RECT 14.155 75.635 14.845 80 ;
        RECT 16.755 75.635 17.445 80 ;
        RECT 19.355 75.635 20.045 80 ;
        RECT 21.955 75.635 22.645 80 ;
        RECT 24.555 75.635 25.245 80 ;
        RECT 27.155 75.635 27.845 80 ;
        RECT 29.755 75.635 30.445 80 ;
        RECT 32.355 75.635 33.045 80 ;
        RECT 34.955 75.635 35.645 80 ;
        RECT 37.555 75.635 38.245 80 ;
        RECT 40.155 75.635 40.845 80 ;
        RECT 42.755 75.635 43.445 80 ;
        RECT 45.355 75.635 46.045 80 ;
        RECT 47.955 75.635 48.645 80 ;
        RECT 50.555 75.635 51.245 78.86 ;
    END
  END VDD
END PPAD_SHORT

MACRO GPAD_LONG
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN GPAD_LONG 0 0 ;
  SIZE 55 BY 80 ;
  SYMMETRY X Y R90 ;
  SITE IOSite ;
  PIN VSS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.755 75.635 4.445 80 ;
        RECT 6.355 75.635 7.045 80 ;
        RECT 8.955 75.635 9.645 80 ;
        RECT 11.555 75.635 12.245 80 ;
        RECT 14.155 75.635 14.845 80 ;
        RECT 16.755 75.635 17.445 80 ;
        RECT 19.355 75.635 20.045 80 ;
        RECT 21.955 75.635 22.645 80 ;
        RECT 24.555 75.635 25.245 80 ;
        RECT 27.155 75.635 27.845 80 ;
        RECT 29.755 75.635 30.445 80 ;
        RECT 32.355 75.635 33.045 80 ;
        RECT 34.955 75.635 35.645 80 ;
        RECT 37.555 75.635 38.245 80 ;
        RECT 40.155 75.635 40.845 80 ;
        RECT 42.755 75.635 43.445 80 ;
        RECT 45.355 75.635 46.045 80 ;
        RECT 47.955 75.635 48.645 80 ;
        RECT 3.28 77.9 50.735 80 ;
        RECT 50.555 75.635 51.245 78.86 ;
      LAYER metal2 ;
        RECT 3.755 75.635 4.445 80 ;
        RECT 6.355 75.635 7.045 80 ;
        RECT 8.955 75.635 9.645 80 ;
        RECT 11.555 75.635 12.245 80 ;
        RECT 14.155 75.635 14.845 80 ;
        RECT 16.755 75.635 17.445 80 ;
        RECT 19.355 75.635 20.045 80 ;
        RECT 21.955 75.635 22.645 80 ;
        RECT 24.555 75.635 25.245 80 ;
        RECT 27.155 75.635 27.845 80 ;
        RECT 29.755 75.635 30.445 80 ;
        RECT 32.355 75.635 33.045 80 ;
        RECT 34.955 75.635 35.645 80 ;
        RECT 37.555 75.635 38.245 80 ;
        RECT 40.155 75.635 40.845 80 ;
        RECT 42.755 75.635 43.445 80 ;
        RECT 45.355 75.635 46.045 80 ;
        RECT 47.955 75.635 48.645 80 ;
        RECT 3.28 77.9 50.735 80 ;
        RECT 50.555 75.635 51.245 78.86 ;
      LAYER metal3 ;
        RECT 3.755 75.635 4.445 80 ;
        RECT 6.355 75.635 7.045 80 ;
        RECT 8.955 75.635 9.645 80 ;
        RECT 11.555 75.635 12.245 80 ;
        RECT 14.155 75.635 14.845 80 ;
        RECT 16.755 75.635 17.445 80 ;
        RECT 19.355 75.635 20.045 80 ;
        RECT 21.955 75.635 22.645 80 ;
        RECT 24.555 75.635 25.245 80 ;
        RECT 27.155 75.635 27.845 80 ;
        RECT 29.755 75.635 30.445 80 ;
        RECT 32.355 75.635 33.045 80 ;
        RECT 34.955 75.635 35.645 80 ;
        RECT 37.555 75.635 38.245 80 ;
        RECT 40.155 75.635 40.845 80 ;
        RECT 42.755 75.635 43.445 80 ;
        RECT 45.355 75.635 46.045 80 ;
        RECT 47.955 75.635 48.645 80 ;
        RECT 3.28 77.9 50.735 80 ;
        RECT 50.555 75.635 51.245 78.86 ;
      LAYER metal4 ;
        RECT 3.755 75.635 4.445 80 ;
        RECT 6.355 75.635 7.045 80 ;
        RECT 8.955 75.635 9.645 80 ;
        RECT 11.555 75.635 12.245 80 ;
        RECT 14.155 75.635 14.845 80 ;
        RECT 16.755 75.635 17.445 80 ;
        RECT 19.355 75.635 20.045 80 ;
        RECT 21.955 75.635 22.645 80 ;
        RECT 24.555 75.635 25.245 80 ;
        RECT 27.155 75.635 27.845 80 ;
        RECT 29.755 75.635 30.445 80 ;
        RECT 32.355 75.635 33.045 80 ;
        RECT 34.955 75.635 35.645 80 ;
        RECT 37.555 75.635 38.245 80 ;
        RECT 40.155 75.635 40.845 80 ;
        RECT 42.755 75.635 43.445 80 ;
        RECT 45.355 75.635 46.045 80 ;
        RECT 47.955 75.635 48.645 80 ;
        RECT 3.28 77.9 50.735 80 ;
        RECT 50.555 75.635 51.245 78.86 ;
    END
  END VSS
END GPAD_LONG

MACRO GPAD_SHORT
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN GPAD_SHORT 0 0 ;
  SIZE 55 BY 80 ;
  SYMMETRY X Y R90 ;
  SITE IOSite ;
  PIN VSS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.755 75.635 4.445 80 ;
        RECT 6.355 75.635 7.045 80 ;
        RECT 8.955 75.635 9.645 80 ;
        RECT 11.555 75.635 12.245 80 ;
        RECT 14.155 75.635 14.845 80 ;
        RECT 16.755 75.635 17.445 80 ;
        RECT 19.355 75.635 20.045 80 ;
        RECT 21.955 75.635 22.645 80 ;
        RECT 24.555 75.635 25.245 80 ;
        RECT 27.155 75.635 27.845 80 ;
        RECT 29.755 75.635 30.445 80 ;
        RECT 32.355 75.635 33.045 80 ;
        RECT 34.955 75.635 35.645 80 ;
        RECT 37.555 75.635 38.245 80 ;
        RECT 40.155 75.635 40.845 80 ;
        RECT 42.755 75.635 43.445 80 ;
        RECT 45.355 75.635 46.045 80 ;
        RECT 47.955 75.635 48.645 80 ;
        RECT 50.555 75.635 51.245 78.86 ;
      LAYER metal2 ;
        RECT 3.755 75.635 4.445 80 ;
        RECT 6.355 75.635 7.045 80 ;
        RECT 8.955 75.635 9.645 80 ;
        RECT 11.555 75.635 12.245 80 ;
        RECT 14.155 75.635 14.845 80 ;
        RECT 16.755 75.635 17.445 80 ;
        RECT 19.355 75.635 20.045 80 ;
        RECT 21.955 75.635 22.645 80 ;
        RECT 24.555 75.635 25.245 80 ;
        RECT 27.155 75.635 27.845 80 ;
        RECT 29.755 75.635 30.445 80 ;
        RECT 32.355 75.635 33.045 80 ;
        RECT 34.955 75.635 35.645 80 ;
        RECT 37.555 75.635 38.245 80 ;
        RECT 40.155 75.635 40.845 80 ;
        RECT 42.755 75.635 43.445 80 ;
        RECT 45.355 75.635 46.045 80 ;
        RECT 47.955 75.635 48.645 80 ;
        RECT 50.555 75.635 51.245 78.86 ;
      LAYER metal3 ;
        RECT 3.755 75.635 4.445 80 ;
        RECT 6.355 75.635 7.045 80 ;
        RECT 8.955 75.635 9.645 80 ;
        RECT 11.555 75.635 12.245 80 ;
        RECT 14.155 75.635 14.845 80 ;
        RECT 16.755 75.635 17.445 80 ;
        RECT 19.355 75.635 20.045 80 ;
        RECT 21.955 75.635 22.645 80 ;
        RECT 24.555 75.635 25.245 80 ;
        RECT 27.155 75.635 27.845 80 ;
        RECT 29.755 75.635 30.445 80 ;
        RECT 32.355 75.635 33.045 80 ;
        RECT 34.955 75.635 35.645 80 ;
        RECT 37.555 75.635 38.245 80 ;
        RECT 40.155 75.635 40.845 80 ;
        RECT 42.755 75.635 43.445 80 ;
        RECT 45.355 75.635 46.045 80 ;
        RECT 47.955 75.635 48.645 80 ;
        RECT 50.555 75.635 51.245 78.86 ;
      LAYER metal4 ;
        RECT 3.755 75.635 4.445 80 ;
        RECT 6.355 75.635 7.045 80 ;
        RECT 8.955 75.635 9.645 80 ;
        RECT 11.555 75.635 12.245 80 ;
        RECT 14.155 75.635 14.845 80 ;
        RECT 16.755 75.635 17.445 80 ;
        RECT 19.355 75.635 20.045 80 ;
        RECT 21.955 75.635 22.645 80 ;
        RECT 24.555 75.635 25.245 80 ;
        RECT 27.155 75.635 27.845 80 ;
        RECT 29.755 75.635 30.445 80 ;
        RECT 32.355 75.635 33.045 80 ;
        RECT 34.955 75.635 35.645 80 ;
        RECT 37.555 75.635 38.245 80 ;
        RECT 40.155 75.635 40.845 80 ;
        RECT 42.755 75.635 43.445 80 ;
        RECT 45.355 75.635 46.045 80 ;
        RECT 47.955 75.635 48.645 80 ;
        RECT 50.555 75.635 51.245 78.86 ;
    END
  END VSS
END GPAD_SHORT

END LIBRARY
