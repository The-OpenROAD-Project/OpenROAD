# macro with bus bit (intentionally reverse order of liberty)

VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MACRO bus16
 SIZE 50 BY 20 ;
 PIN in[0] DIRECTION INPUT ; END in[0]
 PIN in[1] DIRECTION INPUT ; END in[1]
 PIN in[2] DIRECTION INPUT ; END in[2]
 PIN in[3] DIRECTION INPUT ; END in[3]
 PIN in[4] DIRECTION INPUT ; END in[4]
 PIN in[5] DIRECTION INPUT ; END in[5]
 PIN in[6] DIRECTION INPUT ; END in[6]
 PIN in[7] DIRECTION INPUT ; END in[7]
 PIN in[8] DIRECTION INPUT ; END in[8]
 PIN in[9] DIRECTION INPUT ; END in[9]
 PIN in[10] DIRECTION INPUT ; END in[10]
 PIN in[11] DIRECTION INPUT ; END in[11]
 PIN in[12] DIRECTION INPUT ; END in[12]
 PIN in[13] DIRECTION INPUT ; END in[13]
 PIN in[14] DIRECTION INPUT ; END in[14]
 PIN in[15] DIRECTION INPUT ; END in[15]
 PIN out[0] DIRECTION OUTPUT ; END out[0]
 PIN out[1] DIRECTION OUTPUT ; END out[1]
 PIN out[2] DIRECTION OUTPUT ; END out[2]
 PIN out[3] DIRECTION OUTPUT ; END out[3]
 PIN out[4] DIRECTION OUTPUT ; END out[4]
 PIN out[5] DIRECTION OUTPUT ; END out[5]
 PIN out[6] DIRECTION OUTPUT ; END out[6]
 PIN out[7] DIRECTION OUTPUT ; END out[7]
 PIN out[8] DIRECTION OUTPUT ; END out[8]
 PIN out[9] DIRECTION OUTPUT ; END out[9]
 PIN out[10] DIRECTION OUTPUT ; END out[10]
 PIN out[11] DIRECTION OUTPUT ; END out[11]
 PIN out[12] DIRECTION OUTPUT ; END out[12]
 PIN out[13] DIRECTION OUTPUT ; END out[13]
 PIN out[14] DIRECTION OUTPUT ; END out[14]
 PIN out[15] DIRECTION OUTPUT ; END out[15]
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END bus16

END LIBRARY
