module test_no_sinks (clk);
 input clk;

 DFF_X1 ff1 .CK(clk);
endmodule
