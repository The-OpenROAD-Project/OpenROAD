VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  LAYER contactResistance REAL ;
END PROPERTYDEFINITIONS

UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MANUFACTURINGGRID 0.0025 ;
LAYER poly
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE NWELL ;" ;
END poly

LAYER contact
  TYPE CUT ;
  SPACING 0.075 ;
  PROPERTY contactResistance 10.5 ;
END contact

LAYER metal1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.19 ;
  WIDTH 0.065 ;
  SPACING 0.065 ;
  RESISTANCE RPERSQ 0.38 ;
  PROPERTY LEF58_SPACING "SPACING 1.3 ENDOFLINE 1.5 WITHIN 1.9 SAMEMASK EXCEPTEXACTWIDTH 0.5 0.3 PARALLELEDGE 0.2 WITHIN 9.1 PRL 81 MINLENGTH -0.1 TWOEDGES" ;
  PROPERTY LEF58_MINSTEP "MINSTEP 0.6 MAXEDGES 1 MINADJACENTLENGTH 1.0 CONVEXCORNER ;
                          MINSTEP 0.6 MINADJACENTLENGTH 1.0 0.15 ;
                          MINSTEP 0.6 MINBETWEENLENGTH 0.13 EXCEPTSAMECORNERS ;
                          MINSTEP 0.6 NOBETWEENEOL 0.5 ; " ;
  PROPERTY LEF58_CORNERSPACING
    "CORNERSPACING CONVEXCORNER EXCEPTEOL 0.090
      WIDTH 0.000 SPACING 0.110 ;" ;
  PROPERTY LEF58_SPACINGTABLE
    "SPACINGTABLE
      PARALLELRUNLENGTH WRONGDIRECTION
      EXCEPTEOL 0.090
                                                  0.00      0.07
         WIDTH 0.0                                0.05      0.05
         WIDTH 0.1   EXCEPTWITHIN 0.0 0.05        0.05      0.08 ;" ;
  PROPERTY LEF58_RIGHTWAYONGRIDONLY "RIGHTWAYONGRIDONLY CHECKMASK; " ;
  PROPERTY LEF58_RECTONLY "RECTONLY EXCEPTNONCOREPINS ; " ;
  PROPERTY LEF58_TYPE "TYPE MIMCAP ;" ;
  PROPERTY LEF58_EOLKEEPOUT "
    EOLKEEPOUT 0.2 EXTENSION 0.03 0.05 0.1 
    EXCEPTWITHIN -0.01 0.05
    CLASS EOL_WIDE ; 
  " ;
  PROPERTY LEF58_EOLEXTENSIONSPACING
    "EOLEXTENSIONSPACING 0.1 PARALLELONLY ENDOFLINE 0.11 EXTENSION 0.14 ;" ;
  PROPERTY LEF58_WIDTHTABLE
    "WIDTHTABLE 0.1 0.2 0.3 0.4 0.5 ORTHOGONAL ; " ;
  PROPERTY LEF58_MINIMUMCUT
    "MINIMUMCUT 2 WIDTH 0.09 WITHIN 0.05 FROMABOVE AREA 2.0 ; " ;
END metal1

LAYER via1
  TYPE CUT ;
  SPACING 0.075 ;
  PROPERTY contactResistance 5.69 ;
  PROPERTY LEF58_CUTCLASS 
  "CUTCLASS VA WIDTH 0.15 ; 
   CUTCLASS cls1 WIDTH 0.15 ; 
   CUTCLASS cls2 WIDTH 0.15 ; 
   CUTCLASS cls3 WIDTH 0.15 ; 
   CUTCLASS cls4 WIDTH 0.15 ; 
  " ;
  PROPERTY LEF58_SPACING
  "SPACING 0.12 MAXXY ;
   SPACING 0.3 SAMEMETAL LAYER metal1 STACK ;" ;
  PROPERTY LEF58_ENCLOSURE
    "ENCLOSURE CUTCLASS cls1 ABOVE 0.05 0.05
        WIDTH 0.2 INCLUDEABUTTED ; " ;
  PROPERTY LEF58_SPACINGTABLE
  "SPACINGTABLE ORTHOGONAL 
    WITHIN 0.2 SPACING 0.15
    WITHIN 0.3 SPACING 0.25 ;
  SPACINGTABLE DEFAULT 0.12 
    SAMEMASK
    SAMENET
    LAYER metal1 NOSTACK 
      PRLFORALIGNEDCUT cls1 TO cls2 cls3 TO cls4 
    PRL 0.14 MAXXY cls1 TO cls2 0.3
    CUTCLASS   cls1 SIDE  cls1 END   cls2
    cls3        0.1 0.2    0.3 -    0.4 0.5 
    cls4        0.6 -      0.7 -    0.8 0.9 ; " ;
  PROPERTY LEF58_ARRAYSPACING
  "ARRAYSPACING CUTCLASS VA PARALLELOVERLAP WIDTH 1.0 CUTSPACING 0.10
    ARRAYCUTS 3 SPACING 0.30 ; " ;
END via1

LAYER metal2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.19 ;
  WIDTH 0.07 ;
  SPACING 0.075 ;
  RESISTANCE RPERSQ 0.25 ;
END metal2

LAYER via2
  TYPE CUT ;
  SPACING 0.085 ;
  PROPERTY contactResistance 11.39 ;
END via2

LAYER metal3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.19 ;
  WIDTH 0.07 ;
  SPACING 0.07 ;
  RESISTANCE RPERSQ 0.25 ;
END metal3

LAYER via3
  TYPE CUT ;
  SPACING 0.085 ;
  PROPERTY contactResistance 16.73 ;
END via3

LAYER metal4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.285 ;
  WIDTH 0.14 ;
  SPACING 0.14 ;
  RESISTANCE RPERSQ 0.25 ;
END metal4

LAYER via4
  TYPE CUT ;
  SPACING 0.16 ;
  PROPERTY contactResistance 21.44 ;
END via4

LAYER metal5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.285 ;
  WIDTH 0.14 ;
  SPACING 0.14 ;
  RESISTANCE RPERSQ 0.25 ;
END metal5

LAYER via5
  TYPE CUT ;
  SPACING 0.16 ;
  PROPERTY contactResistance 24.08 ;
END via5

LAYER metal6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.285 ;
  WIDTH 0.14 ;
  SPACING 0.14 ;
  RESISTANCE RPERSQ 0.25 ;
END metal6

LAYER via6
  TYPE CUT ;
  SPACING 0.16 ;
  PROPERTY contactResistance 11.39 ;
END via6

LAYER metal7
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.855 ;
  WIDTH 0.4 ;
  SPACING 0.4 ;
  RESISTANCE RPERSQ 0.25 ;
END metal7

LAYER via7
  TYPE CUT ;
  SPACING 0.44 ;
  PROPERTY contactResistance 5.69 ;
END via7

LAYER metal8
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.855 ;
  WIDTH 0.4 ;
  SPACING 0.4 ;
  RESISTANCE RPERSQ 0.25 ;
END metal8

LAYER via8
  TYPE CUT ;
  SPACING 0.44 ;
  PROPERTY contactResistance 16.73 ;
END via8

LAYER metal9
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 1.71 ;
  WIDTH 0.8 ;
  SPACING 0.8 ;
  RESISTANCE RPERSQ 0.21 ;
END metal9

LAYER via9
  TYPE CUT ;
  SPACING 0.88 ;
  PROPERTY contactResistance 21.44 ;
END via9

LAYER metal10
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 1.71 ;
  WIDTH 0.8 ;
  SPACING 0.8 ;
  RESISTANCE RPERSQ 0.21 ;
END metal10

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA M2_M1_via DEFAULT
  LAYER metal1 ;
    RECT -0.0675 -0.0325 0.0675 0.0325 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
  LAYER metal2 ;
    RECT -0.035 -0.0675 0.035 0.0675 ;
END M2_M1_via

VIA M3_M2_via DEFAULT
  LAYER metal2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END M3_M2_via

VIA M4_M3_via DEFAULT
  LAYER metal3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END M4_M3_via

VIA M5_M4_via DEFAULT
  LAYER metal4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END M5_M4_via

VIA M6_M5_via DEFAULT
  LAYER metal5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END M6_M5_via

VIA M7_M6_via DEFAULT
  LAYER metal6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
END M7_M6_via

VIA M8_M7_via DEFAULT
  LAYER metal7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER via7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER metal8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
END M8_M7_via

VIA M9_M8_via DEFAULT
  LAYER metal8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER via8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER metal9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
END M9_M8_via

VIA M10_M9_via DEFAULT
  LAYER metal9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER via9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER metal10 ;
    RECT -0.4 -0.4 0.4 0.4 ;
END M10_M9_via

VIA M2_M1_viaB DEFAULT
  LAYER metal1 ;
    RECT -0.0675 -0.0325 0.0675 0.0325 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
  LAYER metal2 ;
    RECT -0.0675 -0.035 0.0675 0.035 ;
END M2_M1_viaB

VIA M2_M1_viaC DEFAULT
  LAYER metal1 ;
    RECT -0.0325 -0.0675 0.0325 0.0675 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
  LAYER metal2 ;
    RECT -0.035 -0.0675 0.035 0.0675 ;
END M2_M1_viaC

VIA M3_M2_viaB DEFAULT
  LAYER metal2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal3 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END M3_M2_viaB

VIA M3_M2_viaC DEFAULT
  LAYER metal2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END M3_M2_viaC

VIA M4_M3_viaB DEFAULT
  LAYER metal3 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END M4_M3_viaB

VIARULE M2_M1 GENERATE
  LAYER metal1 ;
    ENCLOSURE 0 0.035 ;
  LAYER metal2 ;
    ENCLOSURE 0 0.035 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
    SPACING 0.14 BY 0.14 ;
END M2_M1

VIARULE M3_M2 GENERATE
  LAYER metal2 ;
    ENCLOSURE 0 0.035 ;
  LAYER metal3 ;
    ENCLOSURE 0 0.035 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.155 BY 0.155 ;
END M3_M2

VIARULE M4_M3 GENERATE
  LAYER metal3 ;
    ENCLOSURE 0 0.035 ;
  LAYER metal4 ;
    ENCLOSURE 0 0 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.155 BY 0.155 ;
END M4_M3

VIARULE M5_M4 GENERATE
  LAYER metal4 ;
    ENCLOSURE 0 0 ;
  LAYER metal5 ;
    ENCLOSURE 0 0 ;
  LAYER via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END M5_M4

VIARULE M6_M5 GENERATE
  LAYER metal5 ;
    ENCLOSURE 0 0 ;
  LAYER metal6 ;
    ENCLOSURE 0 0 ;
  LAYER via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END M6_M5

VIARULE M7_M6 GENERATE
  LAYER metal6 ;
    ENCLOSURE 0 0 ;
  LAYER metal7 ;
    ENCLOSURE 0.13 0.13 ;
  LAYER via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END M7_M6

VIARULE M8_M7 GENERATE
  LAYER metal7 ;
    ENCLOSURE 0 0 ;
  LAYER metal8 ;
    ENCLOSURE 0 0 ;
  LAYER via7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.84 BY 0.84 ;
END M8_M7

VIARULE M9_M8 GENERATE
  LAYER metal8 ;
    ENCLOSURE 0 0 ;
  LAYER metal9 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER via8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.84 BY 0.84 ;
END M9_M8

VIARULE M10_M9 GENERATE
  LAYER metal9 ;
    ENCLOSURE 0 0 ;
  LAYER metal10 ;
    ENCLOSURE 0 0 ;
  LAYER via9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
    SPACING 1.68 BY 1.68 ;
END M10_M9

VIARULE M1_POLY GENERATE
  LAYER poly ;
    ENCLOSURE 0 0 ;
  LAYER metal1 ;
    ENCLOSURE 0 0.035 ;
  LAYER contact ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
    SPACING 0.14 BY 0.14 ;
END M1_POLY

SPACING
  SAMENET metal1 metal1 0.065 ;
  SAMENET metal2 metal2 0.07 ;
  SAMENET metal6 metal6 0.14 ;
  SAMENET metal5 metal5 0.14 ;
  SAMENET metal4 metal4 0.14 ;
  SAMENET metal3 metal3 0.07 ;
  SAMENET metal7 metal7 0.4 ;
  SAMENET metal8 metal8 0.4 ;
  SAMENET metal9 metal9 0.8 ;
  SAMENET metal10 metal10 0.8 ;
END SPACING

SITE CoreSite
  CLASS CORE ;
  SIZE 0.38 BY 2.47 ;
END CoreSite

MACRO AND2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X1 0 0 ;
  SIZE 1.14 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.1475 1.2275 0.2825 1.3625 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.3475 1.2275 0.4825 1.3625 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.9175 0.87 0.9825 2.1075 ;
    END
  END Y
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.7075 -0.065 0.7725 1.11 ;
        RECT 0 -0.065 1.14 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.1425 1.5575 0.2075 2.535 ;
        RECT 0.6225 1.5575 0.6875 2.535 ;
        RECT 0 2.405 1.14 2.535 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.1425 0.59 0.2075 1.145 ;
      RECT 0.1425 1.08 0.6425 1.145 ;
      RECT 0.5775 1.08 0.6425 1.4925 ;
      RECT 0.4375 1.4275 0.7775 1.4925 ;
      RECT 0.4375 1.4275 0.5025 2.1075 ;
  END
END AND2X1

MACRO AND2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X2 0 0 ;
  SIZE 0.95 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.1475 0.8475 0.2225 0.9825 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.4175 0.9175 0.6025 1.0525 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.7275 0.1725 0.7925 2.235 ;
        RECT 0.7275 1.1075 0.8025 2.235 ;
    END
  END Y
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.4425 -0.065 0.5075 0.7225 ;
        RECT 0 -0.065 0.95 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.0675 1.265 0.1325 2.535 ;
        RECT 0.4425 1.265 0.5075 2.535 ;
        RECT 0 2.405 0.95 2.535 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.0325 0.2075 0.1675 0.6925 ;
      RECT 0.0325 0.6275 0.3525 0.6925 ;
      RECT 0.2875 0.7875 0.5975 0.8525 ;
      RECT 0.2875 0.6275 0.3525 1.78 ;
      RECT 0.2175 1.295 0.3525 1.78 ;
  END
END AND2X2

MACRO AOI21X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21X1 0 0 ;
  SIZE 0.95 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.1575 0.8475 0.2825 0.9825 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.3475 0.7275 0.4475 0.8625 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.6675 0.8475 0.7925 0.9825 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.5125 0.1475 0.5775 0.9825 ;
        RECT 0.5375 0.9175 0.6025 1.15 ;
        RECT 0.5375 1.085 0.7675 1.15 ;
        RECT 0.7025 1.085 0.7675 2.235 ;
    END
  END Y
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.1375 -0.065 0.2025 0.7025 ;
        RECT 0.7525 -0.065 0.8175 0.6725 ;
        RECT 0 -0.065 0.95 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.3225 1.345 0.3875 2.535 ;
        RECT 0 2.405 0.95 2.535 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.1375 1.215 0.5775 1.28 ;
      RECT 0.1375 1.215 0.2025 2.235 ;
      RECT 0.5125 1.215 0.5775 2.235 ;
  END
END AOI21X1

MACRO AOI22X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22X1 0 0 ;
  SIZE 1.14 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.8575 0.7675 0.9825 0.9825 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.6675 0.7675 0.7925 0.9825 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.0325 0.7675 0.2225 0.9825 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.4775 0.7675 0.6025 0.9825 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.3475 0.13 0.4125 2.0675 ;
        RECT 0.3475 0.13 0.6 0.195 ;
        RECT 0.535 0.13 0.6 0.7025 ;
    END
  END Y
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.16 -0.065 0.225 0.7025 ;
        RECT 0.915 -0.065 0.98 0.7025 ;
        RECT 0 -0.065 1.14 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.725 1.1775 0.79 2.535 ;
        RECT 0 2.405 1.14 2.535 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.535 1.0475 0.98 1.1125 ;
      RECT 0.915 1.0475 0.98 2.0675 ;
      RECT 0.16 1.0475 0.225 2.1975 ;
      RECT 0.535 1.0475 0.6 2.1975 ;
      RECT 0.16 2.1325 0.6 2.1975 ;
  END
END AOI22X1

MACRO BUFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX2 0 0 ;
  SIZE 0.76 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.53 0.8975 0.645 1.0325 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.0325 0.13 0.0975 2.235 ;
        RECT 0.0325 0.13 0.225 0.7025 ;
        RECT 0.0325 0.7675 0.225 2.235 ;
    END
  END Y
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.345 -0.065 0.41 0.7025 ;
        RECT 0 -0.065 0.76 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.345 1.2275 0.41 2.535 ;
        RECT 0 2.405 0.76 2.535 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.53 0.13 0.705 0.8325 ;
      RECT 0.29 0.7675 0.705 0.8325 ;
      RECT 0.29 0.7675 0.465 0.9025 ;
      RECT 0.29 0.7675 0.355 1.1625 ;
      RECT 0.29 1.0975 0.705 1.1625 ;
      RECT 0.53 1.0975 0.705 1.815 ;
  END
END BUFX2

MACRO BUFX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX4 0 0 ;
  SIZE 1.14 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.85 1.0825 0.99 1.2175 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.215 0.4875 0.28 1.3325 ;
        RECT 0.215 0.4875 0.41 0.5525 ;
        RECT 0.215 1.2675 0.46 1.3325 ;
        RECT 0.345 0.4875 0.41 1.0425 ;
        RECT 0.215 1.1075 0.4125 1.1725 ;
        RECT 0.395 1.2675 0.46 2.2425 ;
    END
  END Y
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.0575 -0.065 0.1225 1.0375 ;
        RECT 0.585 -0.065 0.65 0.9275 ;
        RECT 1.03 -0.065 1.095 0.9275 ;
        RECT 0 -0.065 1.14 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.0475 1.1025 0.1125 2.535 ;
        RECT 0.585 1.2675 0.65 2.535 ;
        RECT 1.03 1.2825 1.095 2.535 ;
        RECT 0 2.405 1.14 2.535 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.715 0.3225 0.91 0.3875 ;
      RECT 0.845 0.3225 0.91 1.0175 ;
      RECT 0.4775 1.0675 0.78 1.1325 ;
      RECT 0.4775 1.0675 0.5425 1.2025 ;
      RECT 0.715 0.3225 0.78 1.3475 ;
      RECT 0.715 1.2825 0.91 1.3475 ;
      RECT 0.845 1.2825 0.91 1.6975 ;
  END
END BUFX4

MACRO CLKBUF1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUF1 0 0 ;
  SIZE 2.09 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.665 0.9175 1.7425 1.0525 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.1575 0.9175 0.24 0.9825 ;
        RECT 0.175 0.6575 0.24 1.28 ;
        RECT 0.175 1.215 0.37 1.28 ;
        RECT 0.305 0.1675 0.37 0.7225 ;
        RECT 0.175 0.6575 0.37 0.7225 ;
        RECT 0.305 1.215 0.37 2.235 ;
    END
  END Y
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.045 -0.065 0.11 0.7225 ;
        RECT 0.565 -0.065 0.63 0.7225 ;
        RECT 1.045 -0.065 1.11 0.7225 ;
        RECT 1.53 -0.065 1.595 0.7225 ;
        RECT 1.905 -0.065 1.97 0.7225 ;
        RECT 0 -0.065 2.09 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.12 1.345 0.185 2.535 ;
        RECT 0.54 1.345 0.605 2.535 ;
        RECT 1.045 1.345 1.11 2.535 ;
        RECT 1.525 1.345 1.59 2.535 ;
        RECT 1.905 1.345 1.97 2.535 ;
        RECT 0 2.405 2.09 2.535 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.435 0.7475 0.5 0.8825 ;
      RECT 0.75 0.1725 0.815 0.8825 ;
      RECT 0.435 0.8175 0.815 0.8825 ;
      RECT 0.62 0.8175 0.685 1.28 ;
      RECT 0.62 1.215 0.885 1.28 ;
      RECT 0.75 1.215 0.885 2.2 ;
      RECT 1.305 0.2075 1.44 0.6925 ;
      RECT 1.175 0.6275 1.44 0.6925 ;
      RECT 0.77 0.9475 1.24 1.0125 ;
      RECT 1.175 0.6275 1.24 1.325 ;
      RECT 1.175 1.26 1.4 1.325 ;
      RECT 1.335 1.26 1.4 2.235 ;
      RECT 1.4 0.7825 1.465 0.9175 ;
      RECT 1.535 0.7875 1.78 0.8525 ;
      RECT 1.715 0.1725 1.78 0.8525 ;
      RECT 1.4 0.8525 1.6 0.9175 ;
      RECT 1.535 0.7875 1.6 1.28 ;
      RECT 1.535 1.215 1.815 1.28 ;
      RECT 1.68 1.215 1.815 2.2 ;
  END
END CLKBUF1

MACRO CLKBUF2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUF2 0 0 ;
  SIZE 2.85 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.1575 0.9175 0.35 1.0525 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.48 0.1725 2.545 0.7275 ;
        RECT 2.48 0.6625 2.675 0.7275 ;
        RECT 2.55 1.215 2.615 2.235 ;
        RECT 2.61 0.6625 2.675 0.9825 ;
        RECT 2.61 0.9175 2.745 0.9825 ;
        RECT 2.68 0.9175 2.745 1.28 ;
        RECT 2.55 1.215 2.745 1.28 ;
    END
  END Y
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.045 -0.065 0.11 0.7225 ;
        RECT 0.42 -0.065 0.485 0.7225 ;
        RECT 0.8 -0.065 0.865 0.7225 ;
        RECT 1.305 -0.065 1.37 0.7225 ;
        RECT 1.785 -0.065 1.85 0.7225 ;
        RECT 2.29 -0.065 2.355 0.7225 ;
        RECT 2.74 -0.065 2.805 0.7225 ;
        RECT 0 -0.065 2.85 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.045 1.345 0.11 2.535 ;
        RECT 0.42 1.345 0.485 2.535 ;
        RECT 0.8 1.345 0.865 2.535 ;
        RECT 1.305 1.345 1.37 2.535 ;
        RECT 1.785 1.345 1.85 2.535 ;
        RECT 2.29 1.345 2.355 2.535 ;
        RECT 2.735 1.345 2.8 2.535 ;
        RECT 0 2.405 2.85 2.535 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.235 0.1725 0.3 0.8525 ;
      RECT 0.235 0.7875 0.48 0.8525 ;
      RECT 0.415 0.9525 0.61 1.0175 ;
      RECT 0.545 0.9525 0.61 1.0875 ;
      RECT 0.415 0.7875 0.48 1.28 ;
      RECT 0.2 1.215 0.48 1.28 ;
      RECT 0.2 1.215 0.335 2.2 ;
      RECT 0.615 0.1725 0.68 0.8875 ;
      RECT 1.045 0.7525 1.11 0.8875 ;
      RECT 0.615 0.8225 1.11 0.8875 ;
      RECT 0.775 0.8225 0.84 1.28 ;
      RECT 0.575 1.215 0.84 1.28 ;
      RECT 0.575 1.215 0.71 2.2 ;
      RECT 0.975 0.2025 1.11 0.6875 ;
      RECT 0.975 0.6225 1.24 0.6875 ;
      RECT 1.175 0.9525 1.645 1.0175 ;
      RECT 1.175 0.6225 1.24 1.36 ;
      RECT 0.975 1.295 1.24 1.36 ;
      RECT 0.975 1.295 1.11 2.2 ;
      RECT 1.6 0.1725 1.665 0.8875 ;
      RECT 2.03 0.7525 2.095 0.8875 ;
      RECT 1.6 0.8225 2.095 0.8875 ;
      RECT 1.73 0.8225 1.795 1.28 ;
      RECT 1.53 1.215 1.795 1.28 ;
      RECT 1.53 1.215 1.665 2.2 ;
      RECT 1.96 0.2025 2.095 0.6875 ;
      RECT 1.96 0.6225 2.225 0.6875 ;
      RECT 2.16 0.7925 2.485 0.8575 ;
      RECT 2.42 0.7925 2.485 0.9275 ;
      RECT 2.16 0.6225 2.225 1.36 ;
      RECT 1.96 1.295 2.225 1.36 ;
      RECT 1.96 1.295 2.095 2.2 ;
  END
END CLKBUF2

MACRO CLKBUF3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUF3 0 0 ;
  SIZE 3.61 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.1575 0.9175 0.35 1.0525 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.24 0.1725 3.305 0.7275 ;
        RECT 3.24 0.6625 3.435 0.7275 ;
        RECT 3.31 1.215 3.375 2.235 ;
        RECT 3.37 0.6625 3.435 0.9825 ;
        RECT 3.37 0.9175 3.505 0.9825 ;
        RECT 3.44 0.9175 3.505 1.28 ;
        RECT 3.31 1.215 3.505 1.28 ;
    END
  END Y
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.045 -0.065 0.11 0.7225 ;
        RECT 0.42 -0.065 0.485 0.7225 ;
        RECT 0.8 -0.065 0.865 0.7225 ;
        RECT 1.305 -0.065 1.37 0.7225 ;
        RECT 1.68 -0.065 1.745 0.7225 ;
        RECT 2.06 -0.065 2.125 0.7225 ;
        RECT 2.545 -0.065 2.61 0.7225 ;
        RECT 3.05 -0.065 3.115 0.7225 ;
        RECT 3.5 -0.065 3.565 0.7225 ;
        RECT 0 -0.065 3.61 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.045 1.345 0.11 2.535 ;
        RECT 0.42 1.345 0.485 2.535 ;
        RECT 0.8 1.345 0.865 2.535 ;
        RECT 1.305 1.345 1.37 2.535 ;
        RECT 1.68 1.345 1.745 2.535 ;
        RECT 2.06 1.345 2.125 2.535 ;
        RECT 2.545 1.345 2.61 2.535 ;
        RECT 3.05 1.345 3.115 2.535 ;
        RECT 3.495 1.345 3.56 2.535 ;
        RECT 0 2.405 3.61 2.535 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.235 0.1725 0.3 0.8525 ;
      RECT 0.235 0.7875 0.48 0.8525 ;
      RECT 0.415 0.9525 0.61 1.0175 ;
      RECT 0.545 0.9525 0.61 1.0875 ;
      RECT 0.415 0.7875 0.48 1.28 ;
      RECT 0.2 1.215 0.48 1.28 ;
      RECT 0.2 1.215 0.335 2.2 ;
      RECT 0.615 0.1725 0.68 0.8875 ;
      RECT 1.045 0.7525 1.11 0.8875 ;
      RECT 0.615 0.8225 1.11 0.8875 ;
      RECT 0.775 0.8225 0.84 1.28 ;
      RECT 0.575 1.215 0.84 1.28 ;
      RECT 0.575 1.215 0.71 2.2 ;
      RECT 0.975 0.2025 1.11 0.6875 ;
      RECT 0.975 0.6225 1.24 0.6875 ;
      RECT 1.175 0.9175 1.5 0.9825 ;
      RECT 1.435 0.9175 1.5 1.0525 ;
      RECT 1.175 0.6225 1.24 1.36 ;
      RECT 0.975 1.295 1.24 1.36 ;
      RECT 0.975 1.295 1.11 2.2 ;
      RECT 1.495 0.1725 1.56 0.8525 ;
      RECT 1.495 0.7875 1.72 0.8525 ;
      RECT 1.655 0.9175 1.92 0.9825 ;
      RECT 1.655 0.7875 1.72 1.28 ;
      RECT 1.455 1.215 1.72 1.28 ;
      RECT 1.455 1.215 1.59 2.2 ;
      RECT 1.875 0.1725 1.94 0.8525 ;
      RECT 1.875 0.7875 2.1 0.8525 ;
      RECT 2.035 0.9525 2.405 1.0175 ;
      RECT 2.035 0.7875 2.1 1.28 ;
      RECT 1.835 1.215 2.1 1.28 ;
      RECT 1.835 1.215 1.97 2.2 ;
      RECT 2.36 0.1725 2.425 0.8875 ;
      RECT 2.79 0.7525 2.855 0.8875 ;
      RECT 2.36 0.8225 2.855 0.8875 ;
      RECT 2.49 0.8225 2.555 1.28 ;
      RECT 2.29 1.215 2.555 1.28 ;
      RECT 2.29 1.215 2.425 2.2 ;
      RECT 2.72 0.2025 2.855 0.6875 ;
      RECT 2.72 0.6225 2.985 0.6875 ;
      RECT 2.92 0.7925 3.245 0.8575 ;
      RECT 3.18 0.7925 3.245 0.9275 ;
      RECT 2.92 0.6225 2.985 1.36 ;
      RECT 2.72 1.295 2.985 1.36 ;
      RECT 2.72 1.295 2.855 2.2 ;
  END
END CLKBUF3

MACRO DFFNEGX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNEGX1 0 0 ;
  SIZE 2.85 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER metal1 ;
        RECT 2.0575 2.0575 2.255 2.1925 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.6225 1.0375 2.7 1.1725 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.065 0.2175 0.13 2.2375 ;
        RECT 0.065 0.9175 0.2225 0.9825 ;
        RECT 0.065 1.625 0.525 1.69 ;
    END
  END Q
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2875 -0.065 0.3525 0.8475 ;
        RECT 0.815 -0.065 0.88 0.4675 ;
        RECT 1.34 -0.065 1.405 0.8125 ;
        RECT 1.955 -0.065 2.02 0.5475 ;
        RECT 2.74 -0.065 2.805 0.9375 ;
        RECT 0 -0.065 2.85 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.25 1.9075 0.315 2.535 ;
        RECT 1.34 2.0475 1.405 2.535 ;
        RECT 1.875 1.3875 1.94 2.535 ;
        RECT 2.74 1.3875 2.805 2.535 ;
        RECT 0 2.405 2.85 2.535 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.38 1.755 0.515 1.96 ;
      RECT 0.38 1.755 0.445 2.13 ;
      RECT 0.38 2.065 0.515 2.13 ;
      RECT 0.405 1.365 0.67 1.43 ;
      RECT 0.605 1.365 0.67 2.115 ;
      RECT 0.58 1.84 0.67 2.115 ;
      RECT 0.63 0.2275 0.695 0.5025 ;
      RECT 0.43 0.4375 0.695 0.5025 ;
      RECT 0.43 0.4375 0.565 0.8875 ;
      RECT 0.67 0.6825 0.805 0.8875 ;
      RECT 0.67 0.6825 0.735 1.0175 ;
      RECT 0.34 0.9525 0.735 1.0175 ;
      RECT 0.34 0.9525 0.405 1.1475 ;
      RECT 0.25 1.0825 0.405 1.1475 ;
      RECT 0.25 1.0825 0.315 1.56 ;
      RECT 0.25 1.495 0.515 1.56 ;
      RECT 0.735 1.3575 1.275 1.8425 ;
      RECT 1.21 1.3575 1.275 2.26 ;
      RECT 0.38 2.195 1.275 2.26 ;
      RECT 0.38 2.195 1.145 2.33 ;
      RECT 1.655 0.8725 1.79 0.9375 ;
      RECT 1.69 1.0125 2.03 1.0775 ;
      RECT 1.165 1.2125 1.405 1.2775 ;
      RECT 1.34 1.2125 1.405 1.9775 ;
      RECT 1.69 0.8725 1.755 1.9775 ;
      RECT 1.34 1.9125 1.755 1.9775 ;
      RECT 1.525 0.7425 2.285 0.8075 ;
      RECT 0.87 0.5425 1.005 0.9525 ;
      RECT 0.87 0.8875 1.59 0.9525 ;
      RECT 2.22 0.7425 2.285 1.1175 ;
      RECT 2.22 1.0525 2.355 1.1175 ;
      RECT 0.605 1.0825 1.59 1.1475 ;
      RECT 0.605 1.0825 0.67 1.2975 ;
      RECT 1.525 0.3975 1.59 1.8475 ;
      RECT 1.895 1.2525 2.425 1.3175 ;
      RECT 2.36 1.2525 2.425 1.9375 ;
      RECT 1.795 0.5225 1.86 0.6775 ;
      RECT 1.795 0.6125 2.425 0.6775 ;
      RECT 2.36 0.6125 2.425 0.8775 ;
    LAYER metal2 ;
      RECT 0.41 1.46 0.48 1.995 ;
      RECT 0.345 2.065 0.515 2.135 ;
      RECT 0.345 2.065 0.415 2.295 ;
      RECT 0.345 2.225 1.18 2.295 ;
    LAYER via1 ;
      RECT 0.38 2.23 0.445 2.295 ;
      RECT 0.415 2.065 0.48 2.13 ;
      RECT 0.415 1.895 0.48 1.96 ;
      RECT 0.415 1.755 0.48 1.82 ;
      RECT 0.415 1.495 0.48 1.56 ;
      RECT 0.52 2.23 0.585 2.295 ;
      RECT 0.66 2.23 0.725 2.295 ;
      RECT 0.8 2.23 0.865 2.295 ;
      RECT 0.94 2.23 1.005 2.295 ;
      RECT 1.08 2.23 1.145 2.295 ;
  END
END DFFNEGX1

MACRO DFFPOSX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFPOSX1 0 0 ;
  SIZE 2.66 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER metal2 ;
        RECT 1.4675 1.4275 1.5375 1.9975 ;
        RECT 1.4675 1.4275 1.5525 1.7025 ;
      LAYER metal1 ;
        RECT 0.5075 0.9275 0.5725 1.1925 ;
        RECT 0.4375 1.1275 0.5725 1.1925 ;
        RECT 0.5075 0.9275 0.9825 0.9925 ;
        RECT 0.7875 0.9275 0.9825 1.2075 ;
        RECT 1.2125 1.015 1.3475 1.2075 ;
        RECT 0.7875 1.1425 1.3475 1.2075 ;
        RECT 1.2825 1.015 1.3475 1.5275 ;
        RECT 1.2825 1.4625 1.5875 1.5275 ;
        RECT 1.4525 1.4625 1.5875 1.6675 ;
        RECT 1.4675 1.8625 1.5325 2.1875 ;
        RECT 2.2225 1.1175 2.3725 1.1825 ;
        RECT 2.3075 1.1175 2.3725 2.1875 ;
        RECT 1.4675 2.1225 2.3725 2.1875 ;
      LAYER via1 ;
        RECT 1.4675 1.8975 1.5325 1.9625 ;
        RECT 1.4875 1.6025 1.5525 1.6675 ;
        RECT 1.4875 1.4625 1.5525 1.5275 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.4375 1.0375 2.515 1.1725 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.0525 0.2175 0.1175 2.2375 ;
        RECT 0.0525 0.9175 0.2225 0.9825 ;
        RECT 0.0525 1.6475 0.4475 1.7125 ;
    END
  END Q
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2875 -0.065 0.3525 0.9875 ;
        RECT 0.7725 -0.065 0.8375 0.4675 ;
        RECT 1.1375 -0.065 1.2025 0.7925 ;
        RECT 1.7075 -0.065 1.8425 0.235 ;
        RECT 2.5275 -0.065 2.5925 0.845 ;
        RECT 0 -0.065 2.66 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2375 1.9075 0.3025 2.535 ;
        RECT 1.1375 1.7225 1.2025 2.535 ;
        RECT 1.7025 2.2525 1.8375 2.535 ;
        RECT 2.5275 1.2675 2.5925 2.535 ;
        RECT 0 2.405 2.66 2.535 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.3675 1.7775 0.4325 2.1275 ;
      RECT 0.3225 1.3875 0.5875 1.4525 ;
      RECT 0.5225 1.3875 0.5875 2.1375 ;
      RECT 0.4975 1.8625 0.5875 2.1375 ;
      RECT 0.5875 0.2275 0.6525 0.5025 ;
      RECT 0.4575 0.4375 0.6525 0.5025 ;
      RECT 0.4575 0.4375 0.5225 0.7625 ;
      RECT 0.1925 1.0575 0.3575 1.1925 ;
      RECT 0.6425 1.0575 0.7075 1.3225 ;
      RECT 0.1925 1.2575 0.7075 1.3225 ;
      RECT 0.1925 1.0575 0.2575 1.5825 ;
      RECT 0.1925 1.5175 0.4575 1.5825 ;
      RECT 0.6475 0.5875 0.7125 0.8625 ;
      RECT 0.6525 1.4425 0.9125 1.8575 ;
      RECT 0.8475 1.4425 0.9125 2.2675 ;
      RECT 0.3675 2.2025 0.9125 2.2675 ;
      RECT 1.0825 0.885 1.5425 0.95 ;
      RECT 1.4775 0.95 1.8175 1.015 ;
      RECT 1.0825 0.885 1.1475 1.0775 ;
      RECT 1.4775 0.685 1.5425 1.3975 ;
      RECT 1.5475 0.465 2.2125 0.53 ;
      RECT 2.1475 0.465 2.2125 0.845 ;
      RECT 2.1525 1.3825 2.2425 1.7975 ;
      RECT 1.5975 1.9225 1.6625 2.0575 ;
      RECT 2.1775 1.3825 2.2425 2.0575 ;
      RECT 1.5975 1.9925 2.2425 2.0575 ;
      RECT 1.3225 0.335 2.3425 0.4 ;
      RECT 1.3225 0.335 1.3875 0.7925 ;
      RECT 2.2775 0.335 2.3425 0.975 ;
      RECT 1.9775 0.91 2.3425 0.975 ;
      RECT 0.9775 1.5925 1.3875 1.6575 ;
      RECT 1.3225 1.7325 2.0425 1.7975 ;
      RECT 1.9775 0.91 2.0425 1.9275 ;
      RECT 1.9775 1.8625 2.1125 1.9275 ;
      RECT 0.9775 1.5925 1.0425 2.0725 ;
      RECT 1.3225 1.5925 1.3875 2.1475 ;
    LAYER metal2 ;
      RECT 0.3575 1.4825 0.4275 1.9125 ;
      RECT 0.3575 1.7775 0.4325 1.9125 ;
      RECT 0.6425 0.5875 0.7125 1.1925 ;
      RECT 0.3675 1.9925 0.4375 2.2675 ;
      RECT 0.3675 2.1975 0.7825 2.2675 ;
    LAYER via1 ;
      RECT 0.3575 1.5175 0.4225 1.5825 ;
      RECT 0.3675 2.0275 0.4325 2.0925 ;
      RECT 0.3675 1.8125 0.4325 1.8775 ;
      RECT 0.4025 2.2025 0.4675 2.2675 ;
      RECT 0.5425 2.2025 0.6075 2.2675 ;
      RECT 0.6425 1.0925 0.7075 1.1575 ;
      RECT 0.6475 0.7625 0.7125 0.8275 ;
      RECT 0.6475 0.6225 0.7125 0.6875 ;
      RECT 0.6825 2.2025 0.7475 2.2675 ;
      RECT 1.4675 1.8975 1.5325 1.9625 ;
      RECT 1.4875 1.6025 1.5525 1.6675 ;
      RECT 1.4875 1.4625 1.5525 1.5275 ;
  END
END DFFPOSX1

MACRO DFFSR
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSR 0 0 ;
  SIZE 4.18 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER metal1 ;
        RECT 0.3475 1.015 0.4125 1.1725 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.5375 0.7275 0.6025 1.075 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.94 0.3925 4.005 0.6025 ;
        RECT 3.9575 0.5375 4.0225 1.8425 ;
        RECT 3.9225 1.2875 4.0225 1.8425 ;
        RECT 4.07 0.1825 4.135 0.4575 ;
        RECT 3.94 0.3925 4.135 0.4575 ;
    END
  END Q
  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.3625 1.815 1.4275 1.95 ;
        RECT 1.3625 1.885 3.5225 1.95 ;
        RECT 3.3875 1.885 3.5225 2.1225 ;
    END
  END R
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.4375 0.9175 2.5725 1.055 ;
        RECT 2.4375 0.945 2.8975 1.01 ;
    END
  END S
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.4075 -0.065 0.4725 0.9 ;
        RECT 0.6675 -0.065 0.7325 0.51 ;
        RECT 1.7075 -0.065 1.7725 0.51 ;
        RECT 3.2475 -0.065 3.3125 0.405 ;
        RECT 3.81 -0.065 3.875 0.4225 ;
        RECT 0 -0.065 4.18 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.4025 1.58 0.4675 2.535 ;
        RECT 1.2025 1.7675 1.2675 2.535 ;
        RECT 1.5175 2.015 1.5825 2.535 ;
        RECT 2.0375 2.015 2.1025 2.535 ;
        RECT 2.6175 2.1425 2.6825 2.535 ;
        RECT 3.2575 2.015 3.3225 2.535 ;
        RECT 3.7375 1.2875 3.8025 2.535 ;
        RECT 0 2.405 4.18 2.535 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.6675 0.64 0.7325 1.3725 ;
      RECT 0.7925 1.5675 0.9275 2.1925 ;
      RECT 0.8625 1.5675 0.9275 2.3225 ;
      RECT 1.0175 1.7675 1.0825 2.3225 ;
      RECT 0.8625 2.2575 1.0825 2.3225 ;
      RECT 0.9275 0.27 1.1525 0.335 ;
      RECT 1.0875 0.27 1.1525 0.405 ;
      RECT 0.9275 0.27 0.9925 0.545 ;
      RECT 0.7975 0.48 0.9925 0.545 ;
      RECT 0.7975 0.48 0.8625 1.3725 ;
      RECT 0.7975 0.7475 0.9325 1.3725 ;
      RECT 0.2175 0.66 0.2875 0.935 ;
      RECT 1.1675 0.835 1.2325 1.115 ;
      RECT 1.1275 1.05 1.2625 1.115 ;
      RECT 1.1275 1.05 1.1925 1.5025 ;
      RECT 0.2175 1.4375 1.1925 1.5025 ;
      RECT 0.2175 0.66 0.2825 1.71 ;
      RECT 1.2975 0.835 1.4325 0.9 ;
      RECT 1.2575 1.27 1.7875 1.335 ;
      RECT 1.3275 0.835 1.3925 1.455 ;
      RECT 1.2575 1.18 1.3925 1.455 ;
      RECT 1.7225 1.27 1.7875 1.685 ;
      RECT 0.9975 0.705 1.8275 0.77 ;
      RECT 0.9975 0.66 1.1025 0.935 ;
      RECT 1.7625 0.705 1.8275 1.075 ;
      RECT 0.9975 0.66 1.0625 1.31 ;
      RECT 1.6025 0.94 1.6675 1.205 ;
      RECT 2.3075 0.375 2.3725 1.205 ;
      RECT 1.6025 1.14 2.3725 1.205 ;
      RECT 2.2425 1.14 2.3075 1.82 ;
      RECT 1.6225 1.755 2.3075 1.82 ;
      RECT 2.4925 1.12 2.5575 1.815 ;
      RECT 0.8125 0.13 1.5125 0.195 ;
      RECT 2.1775 0.1675 2.7025 0.2325 ;
      RECT 1.4475 0.13 1.5125 0.64 ;
      RECT 1.1675 0.505 1.5125 0.64 ;
      RECT 2.1775 0.1675 2.2425 0.64 ;
      RECT 1.1675 0.575 2.2425 0.64 ;
      RECT 2.4925 0.1675 2.5575 0.8525 ;
      RECT 2.8375 0.73 3.0275 0.795 ;
      RECT 2.9625 0.73 3.0275 1.6625 ;
      RECT 2.8275 1.3175 3.0275 1.6625 ;
      RECT 3.4975 0.165 3.6625 0.23 ;
      RECT 3.4975 0.165 3.5625 0.585 ;
      RECT 2.6825 0.52 3.5625 0.585 ;
      RECT 2.6825 0.52 2.7475 0.795 ;
      RECT 2.6225 1.3175 2.6875 1.7925 ;
      RECT 3.6075 1.0875 3.6725 1.7925 ;
      RECT 2.6225 1.7275 3.6725 1.7925 ;
      RECT 3.6275 0.53 3.7325 0.805 ;
      RECT 3.6275 0.53 3.6925 0.935 ;
      RECT 3.1325 0.87 3.8925 0.935 ;
      RECT 3.4775 0.87 3.5425 1.5625 ;
    LAYER metal2 ;
      RECT 0.8275 0.7125 0.8975 2.2275 ;
      RECT 1.1675 0.505 1.5125 0.64 ;
      RECT 1.1675 0.505 1.2375 0.97 ;
      RECT 2.4875 0.2975 2.5575 1.815 ;
    LAYER via1 ;
      RECT 0.8275 2.1275 0.8925 2.1925 ;
      RECT 0.8275 1.9875 0.8925 2.0525 ;
      RECT 0.8275 1.8475 0.8925 1.9125 ;
      RECT 0.8275 1.7075 0.8925 1.7725 ;
      RECT 0.8275 1.5675 0.8925 1.6325 ;
      RECT 0.8325 1.3075 0.8975 1.3725 ;
      RECT 0.8325 1.1675 0.8975 1.2325 ;
      RECT 0.8325 1.0275 0.8975 1.0925 ;
      RECT 0.8325 0.8875 0.8975 0.9525 ;
      RECT 0.8325 0.7475 0.8975 0.8125 ;
      RECT 1.1675 0.87 1.2325 0.935 ;
      RECT 1.1675 0.54 1.2325 0.605 ;
      RECT 1.3075 0.54 1.3725 0.605 ;
      RECT 1.4475 0.54 1.5125 0.605 ;
      RECT 2.4925 1.715 2.5575 1.78 ;
      RECT 2.4925 1.575 2.5575 1.64 ;
      RECT 2.4925 1.435 2.5575 1.5 ;
      RECT 2.4925 1.295 2.5575 1.36 ;
      RECT 2.4925 1.155 2.5575 1.22 ;
      RECT 2.4925 0.7525 2.5575 0.8175 ;
      RECT 2.4925 0.6125 2.5575 0.6775 ;
      RECT 2.4925 0.4725 2.5575 0.5375 ;
      RECT 2.4925 0.3325 2.5575 0.3975 ;
  END
END DFFSR

MACRO FAX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FAX1 0 0 ;
  SIZE 3.61 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.255 1.1075 0.955 1.1725 ;
        RECT 0.89 0.8275 0.955 1.4325 ;
        RECT 0.89 0.8275 2.205 0.8925 ;
        RECT 2.14 0.8275 2.205 0.9725 ;
        RECT 3.075 0.9225 3.14 1.4325 ;
        RECT 0.89 1.3675 3.14 1.4325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.3475 0.1575 0.47 0.2925 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.02 0.9575 1.085 1.1425 ;
        RECT 1.02 0.9575 1.755 1.0225 ;
        RECT 1.69 0.9575 1.755 1.2925 ;
        RECT 2.775 0.8975 2.84 1.2925 ;
        RECT 1.69 1.2275 2.84 1.2925 ;
        RECT 2.775 0.8975 2.8825 1.0325 ;
    END
  END C
  PIN YC
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 1.41 0.1025 1.48 1.3275 ;
      LAYER metal1 ;
        RECT 1.38 0.1375 1.515 0.7625 ;
        RECT 1.38 1.0875 1.5525 1.3025 ;
      LAYER via1 ;
        RECT 1.415 1.2275 1.48 1.2925 ;
        RECT 1.415 1.0875 1.48 1.1525 ;
        RECT 1.415 0.6975 1.48 0.7625 ;
        RECT 1.415 0.5575 1.48 0.6225 ;
        RECT 1.415 0.4175 1.48 0.4825 ;
        RECT 1.415 0.2775 1.48 0.3425 ;
        RECT 1.415 0.1375 1.48 0.2025 ;
    END
  END YC
  PIN YS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.3875 1.1075 3.565 1.1725 ;
        RECT 3.5 0.5575 3.565 1.865 ;
    END
  END YS
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.05 -0.065 0.115 0.9975 ;
        RECT 0.535 -0.065 0.6 0.5775 ;
        RECT 1.71 -0.065 1.775 0.6875 ;
        RECT 2.085 -0.065 2.15 0.5475 ;
        RECT 3.205 -0.065 3.27 0.6875 ;
        RECT 0 -0.065 3.61 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.05 1.3475 0.115 2.535 ;
        RECT 0.53 2.1875 0.595 2.535 ;
        RECT 1.71 1.6075 1.775 2.535 ;
        RECT 2.185 1.7075 2.25 2.535 ;
        RECT 3.205 1.0675 3.27 2.535 ;
        RECT 0 2.405 3.61 2.535 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.915 0.2625 1.065 0.3275 ;
      RECT 0.915 0.2625 0.98 0.5775 ;
      RECT 0.345 2.0475 1.165 2.1125 ;
      RECT 0.345 1.2625 0.41 2.2375 ;
      RECT 1.1 1.6275 1.165 2.3225 ;
      RECT 1.1 0.4425 1.165 0.7175 ;
      RECT 0.345 0.6525 1.165 0.7175 ;
      RECT 0.345 0.4425 0.41 0.9975 ;
      RECT 0.88 1.4975 1.34 1.5625 ;
      RECT 1.275 1.4975 1.34 1.7225 ;
      RECT 0.88 1.4975 1.015 1.9825 ;
      RECT 1.865 1.4975 2.435 1.5625 ;
      RECT 1.865 1.4975 2 1.9825 ;
      RECT 2.37 1.4975 2.435 2.0525 ;
      RECT 1.9 0.2725 1.965 0.6875 ;
      RECT 1.9 0.6225 2.485 0.6875 ;
      RECT 2.42 0.2725 2.485 0.8275 ;
      RECT 2.615 0.7675 3.29 0.8325 ;
      RECT 3.225 0.7675 3.29 0.9625 ;
      RECT 3.225 0.8975 3.36 0.9625 ;
      RECT 2.615 0.2775 2.68 1.1625 ;
      RECT 2.575 1.0975 2.71 1.1625 ;
    LAYER via1 ;
      RECT 1.415 1.2275 1.48 1.2925 ;
      RECT 1.415 1.0875 1.48 1.1525 ;
      RECT 1.415 0.6975 1.48 0.7625 ;
      RECT 1.415 0.5575 1.48 0.6225 ;
      RECT 1.415 0.4175 1.48 0.4825 ;
      RECT 1.415 0.2775 1.48 0.3425 ;
      RECT 1.415 0.1375 1.48 0.2025 ;
  END
END FAX1

MACRO FILL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL 0 0 ;
  SIZE 0.38 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.065 0.38 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 2.405 0.38 2.535 ;
    END
  END vdd
END FILL

MACRO HAX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HAX1 0 0 ;
  SIZE 2.09 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.1075 0.8725 1.1725 1.0075 ;
        RECT 1.1075 0.9425 1.6575 1.0075 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.9125 0.8475 0.9825 0.9825 ;
        RECT 0.9175 0.8475 0.9825 1.1375 ;
        RECT 0.9175 1.0725 1.3075 1.1375 ;
    END
  END B
  PIN YC
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.8675 0.9175 2.0425 0.9825 ;
        RECT 1.9775 0.4775 2.0425 1.8175 ;
    END
  END YC
  PIN YS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.0775 0.5375 0.1525 0.8125 ;
        RECT 0.0875 0.5375 0.1525 1.8175 ;
        RECT 0.0875 0.9175 0.2225 0.9825 ;
    END
  END YS
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2625 -0.065 0.3275 0.7775 ;
        RECT 1.6825 -0.065 1.7475 0.7475 ;
        RECT 0 -0.065 2.09 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2725 1.2675 0.3375 2.535 ;
        RECT 1.1525 1.3475 1.2175 2.535 ;
        RECT 1.6375 1.2675 1.7025 2.535 ;
        RECT 0 2.405 2.09 2.535 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.7125 0.2925 0.8475 0.9375 ;
      RECT 0.3925 0.8725 0.8475 0.9375 ;
      RECT 0.3925 0.8725 0.4575 1.2025 ;
      RECT 0.3175 1.0675 0.4575 1.2025 ;
      RECT 0.3175 1.1375 0.6225 1.2025 ;
      RECT 0.5575 1.1375 0.6225 1.8175 ;
      RECT 0.5625 0.1625 1.2175 0.2275 ;
      RECT 0.5625 0.1625 0.6275 0.8075 ;
      RECT 1.1525 0.1625 1.2175 0.8075 ;
      RECT 1.3075 0.1975 1.3725 0.8775 ;
      RECT 1.3075 0.8125 1.8025 0.8775 ;
      RECT 0.5775 1.0075 0.8425 1.0725 ;
      RECT 0.7775 1.0075 0.8425 1.2675 ;
      RECT 1.4475 1.1375 1.8025 1.2025 ;
      RECT 1.7375 0.8125 1.8025 1.2025 ;
      RECT 0.7775 1.2025 1.5125 1.2675 ;
      RECT 1.4475 1.1375 1.5125 1.8175 ;
  END
END HAX1

MACRO INVX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX1 0 0 ;
  SIZE 0.57 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.1575 0.4875 0.2575 0.6225 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.3475 0.2175 0.4125 1.815 ;
        RECT 0.3125 0.2175 0.4475 0.4225 ;
    END
  END Y
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.1625 -0.065 0.2275 0.4225 ;
        RECT 0 -0.065 0.57 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.1625 1.265 0.2275 2.535 ;
        RECT 0 2.405 0.57 2.535 ;
    END
  END vdd
END INVX1

MACRO INVX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX2 0 0 ;
  SIZE 0.57 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.145 0.8475 0.28 0.9825 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.345 0.1825 0.41 2.235 ;
        RECT 0.345 1.26 0.4125 2.235 ;
        RECT 0.31 0.1825 0.445 0.6675 ;
    END
  END Y
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.16 -0.065 0.225 0.7025 ;
        RECT 0 -0.065 0.57 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.16 1.26 0.225 2.535 ;
        RECT 0 2.405 0.57 2.535 ;
    END
  END vdd
END INVX2

MACRO INVX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX4 0 0 ;
  SIZE 0.76 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.51 0.9175 0.645 1.0525 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.335 0.2975 0.4 1.28 ;
        RECT 0.335 0.9175 0.4125 0.9825 ;
        RECT 0.335 0.2975 0.53 0.3625 ;
        RECT 0.335 1.215 0.53 1.28 ;
        RECT 0.465 0.2975 0.53 0.8525 ;
        RECT 0.465 1.215 0.53 2.235 ;
    END
  END Y
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.205 -0.065 0.27 0.8475 ;
        RECT 0.65 -0.065 0.715 0.8475 ;
        RECT 0 -0.065 0.76 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.275 1.345 0.34 2.535 ;
        RECT 0.65 1.345 0.715 2.535 ;
        RECT 0 2.405 0.76 2.535 ;
    END
  END vdd
END INVX4

MACRO INVX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX8 0 0 ;
  SIZE 1.33 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.3475 1.0425 0.6625 1.1725 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2175 0.18 0.2825 1.3625 ;
        RECT 0.2175 0.18 0.5725 0.245 ;
        RECT 0.5075 0.18 0.5725 0.975 ;
        RECT 0.4775 1.2975 0.6125 2.2025 ;
        RECT 0.2175 1.2975 0.9875 1.3625 ;
        RECT 0.8875 0.18 0.9525 0.975 ;
        RECT 0.5075 0.91 0.9525 0.975 ;
        RECT 0.8525 1.295 0.9875 2.2 ;
    END
  END Y
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.0875 -0.065 0.1525 0.8425 ;
        RECT 0.6975 -0.065 0.7625 0.845 ;
        RECT 0 -0.065 1.33 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.0875 1.26 0.1525 2.535 ;
        RECT 0.6975 1.4275 0.7625 2.535 ;
        RECT 1.0775 1.26 1.1425 2.535 ;
        RECT 0 2.405 1.33 2.535 ;
    END
  END vdd
END INVX8

MACRO LATCH
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LATCH 0 0 ;
  SIZE 1.71 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER metal1 ;
        RECT 0.7025 0.7275 0.7675 1.0675 ;
        RECT 0.3275 1.0025 0.7675 1.0675 ;
        RECT 0.7025 0.7275 0.8375 0.9375 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.4875 0.7275 0.6225 0.9375 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.3325 0.8625 1.3975 0.9975 ;
        RECT 1.3325 0.9175 1.6375 0.9825 ;
        RECT 1.5725 0.2775 1.6375 2.2375 ;
    END
  END Q
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.3075 -0.065 0.3725 0.8275 ;
        RECT 1.2775 -0.065 1.3425 0.7975 ;
        RECT 0 -0.065 1.71 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.3075 1.3475 0.3725 2.535 ;
        RECT 1.3875 1.3475 1.4525 2.535 ;
        RECT 0 2.405 1.71 2.535 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.0325 0.13 0.1875 0.195 ;
      RECT 0.1225 1.1575 0.7875 1.2225 ;
      RECT 0.1225 0.13 0.1875 2.2375 ;
      RECT 0.9025 0.5575 0.9675 0.8325 ;
      RECT 0.9025 0.7675 1.0975 0.8325 ;
      RECT 1.0325 1.0625 1.4325 1.1275 ;
      RECT 1.0325 0.7675 1.0975 1.3625 ;
      RECT 0.8125 1.2975 1.0975 1.3625 ;
      RECT 0.8125 1.2975 0.9475 1.7825 ;
  END
END LATCH

MACRO MUX2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX2X1 0 0 ;
  SIZE 1.52 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.5375 0.5375 0.6525 0.6025 ;
        RECT 0.5875 0.5375 0.6525 0.92 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.1825 0.8475 1.3625 0.9825 ;
    END
  END B
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.3475 0.915 0.4925 1.05 ;
        RECT 0.7175 0.13 0.7825 1.05 ;
        RECT 0.3475 0.985 0.7825 1.05 ;
        RECT 0.7175 0.84 0.8525 0.905 ;
        RECT 0.7175 0.13 1.1125 0.195 ;
        RECT 1.0475 0.13 1.1125 1.25 ;
    END
  END S
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.8475 0.26 0.9825 0.745 ;
        RECT 0.9175 0.26 0.9825 2.29 ;
        RECT 0.8925 1.315 0.9825 2.29 ;
    END
  END Y
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.3725 -0.065 0.4375 0.745 ;
        RECT 1.2575 -0.065 1.3225 0.775 ;
        RECT 0 -0.065 1.52 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.3725 1.26 0.4375 2.535 ;
        RECT 1.2875 1.34 1.3525 2.535 ;
        RECT 0 2.405 1.52 2.535 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.1875 1.115 0.8475 1.18 ;
      RECT 0.7825 1.115 0.8475 1.25 ;
      RECT 0.1875 0.505 0.2525 1.81 ;
  END
END MUX2X1

MACRO NAND2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X1 0 0 ;
  SIZE 0.76 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.045 0.7725 0.235 0.9825 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.43 0.7775 0.6025 0.9825 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.3 0.1575 0.365 1.78 ;
        RECT 0.285 1.0475 0.42 1.78 ;
        RECT 0.3 0.1575 0.6 0.2225 ;
        RECT 0.535 0.1575 0.6 0.7125 ;
    END
  END Y
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.16 -0.065 0.225 0.7075 ;
        RECT 0 -0.065 0.76 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.135 1.0475 0.2 2.535 ;
        RECT 0.51 1.0475 0.575 2.535 ;
        RECT 0 2.405 0.76 2.535 ;
    END
  END vdd
END NAND2X1

MACRO NAND3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3X1 0 0 ;
  SIZE 0.95 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.0325 0.9075 0.2225 1.0975 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2925 0.13 0.4675 1.0975 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.5325 0.13 0.6575 1.0975 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.3475 1.1625 0.4125 1.8425 ;
        RECT 0.3475 1.1625 0.7925 1.2275 ;
        RECT 0.7275 0.13 0.7925 1.8425 ;
    END
  END Y
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.1625 -0.065 0.2275 0.8425 ;
        RECT 0 -0.065 0.95 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.1625 1.1625 0.2275 2.535 ;
        RECT 0.5375 1.2925 0.6025 2.535 ;
        RECT 0 2.405 0.95 2.535 ;
    END
  END vdd
END NAND3X1

MACRO NOR2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X1 0 0 ;
  SIZE 0.76 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.1575 0.4875 0.2825 0.6225 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.4775 0.4875 0.6025 0.6225 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.3475 0.2175 0.4125 0.7925 ;
        RECT 0.31 0.2175 0.445 0.4225 ;
        RECT 0.3475 0.7275 0.6 0.7925 ;
        RECT 0.535 0.7275 0.6 1.7025 ;
    END
  END Y
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.16 -0.065 0.225 0.4225 ;
        RECT 0.535 -0.065 0.6 0.4225 ;
        RECT 0 -0.065 0.76 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.16 0.7275 0.225 2.535 ;
        RECT 0 2.405 0.76 2.535 ;
    END
  END vdd
END NOR2X1

MACRO NOR3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3X1 0 0 ;
  SIZE 0.95 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.07 0.525 0.2225 0.6025 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.3475 0.6225 0.465 0.7925 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.5375 0.6225 0.66 0.7925 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.35 0.1875 0.415 0.5575 ;
        RECT 0.35 0.4925 0.79 0.5575 ;
        RECT 0.725 0.1875 0.79 2.3225 ;
        RECT 0.725 0.7875 0.7925 2.3225 ;
    END
  END Y
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.16 -0.065 0.225 0.4275 ;
        RECT 0.535 -0.065 0.6 0.4275 ;
        RECT 0 -0.065 0.95 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.16 0.7875 0.225 2.535 ;
        RECT 0 2.405 0.95 2.535 ;
    END
  END vdd
END NOR3X1

MACRO OAI21X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21X1 0 0 ;
  SIZE 0.95 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.1575 1.0375 0.2675 1.1725 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.3475 1.0375 0.4275 1.1725 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.6675 1.0675 0.7925 1.2025 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.5375 0.9375 0.6025 1.7825 ;
        RECT 0.4675 1.2975 0.6025 1.7825 ;
        RECT 0.6875 0.1925 0.7525 1.0025 ;
        RECT 0.5375 0.9375 0.7525 1.0025 ;
    END
  END Y
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.3075 -0.065 0.3725 0.7425 ;
        RECT 0 -0.065 0.95 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.1225 1.3475 0.1875 2.535 ;
        RECT 0.6875 1.2675 0.7525 2.535 ;
        RECT 0 2.405 0.95 2.535 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.1225 0.1925 0.1875 0.8725 ;
      RECT 0.4975 0.1925 0.5625 0.8725 ;
      RECT 0.1225 0.8075 0.5625 0.8725 ;
  END
END OAI21X1

MACRO OAI22X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22X1 0 0 ;
  SIZE 1.14 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.8575 1.0475 0.9825 1.1825 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.6675 1.0475 0.7925 1.1825 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.1575 0.9175 0.2825 1.0525 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.4775 1.0475 0.6025 1.1825 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.3475 0.3025 0.4125 1.325 ;
        RECT 0.3475 1.26 0.6025 1.325 ;
        RECT 0.5375 1.26 0.6025 2.235 ;
    END
  END Y
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.7275 -0.065 0.7925 0.8525 ;
        RECT 0 -0.065 1.14 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.1625 1.345 0.2275 2.535 ;
        RECT 0.9175 1.345 0.9825 2.535 ;
        RECT 0 2.405 1.14 2.535 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.1625 0.1725 0.6025 0.2375 ;
      RECT 0.1625 0.1725 0.2275 0.8525 ;
      RECT 0.5375 0.1725 0.6025 0.9825 ;
      RECT 0.9175 0.3025 0.9825 0.9825 ;
      RECT 0.5375 0.9175 0.9825 0.9825 ;
  END
END OAI22X1

MACRO OR2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X1 0 0 ;
  SIZE 1.14 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.3475 0.9175 0.4125 1.0525 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.5075 0.9175 0.6025 1.0525 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.8725 0.5175 0.9375 1.815 ;
        RECT 0.8725 1.1075 0.9825 1.815 ;
        RECT 0.8725 0.5175 1.0075 0.7225 ;
    END
  END Y
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2375 -0.065 0.3025 0.7225 ;
        RECT 0.6125 -0.065 0.6775 0.7225 ;
        RECT 0 -0.065 1.14 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.5925 1.345 0.6575 2.535 ;
        RECT 0 2.405 1.14 2.535 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.4225 0.4825 0.4875 0.8525 ;
      RECT 0.2175 0.7875 0.7325 0.8525 ;
      RECT 0.6675 0.7875 0.7325 1.0525 ;
      RECT 0.2175 0.7875 0.2825 2.235 ;
  END
END OR2X1

MACRO OR2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X2 0 0 ;
  SIZE 0.95 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.0325 0.7375 0.2225 0.9825 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2875 0.8975 0.5 1.0125 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.7275 0.13 0.7925 2.235 ;
        RECT 0.7275 0.13 0.895 0.7025 ;
        RECT 0.7275 0.7675 0.895 2.235 ;
    END
  END Y
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.16 -0.065 0.225 0.6725 ;
        RECT 0.535 -0.065 0.6 0.6725 ;
        RECT 0 -0.065 0.95 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.535 1.2275 0.6 2.535 ;
        RECT 0 2.405 0.95 2.535 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.345 0.13 0.41 0.8325 ;
      RECT 0.345 0.7675 0.655 0.8325 ;
      RECT 0.59 0.7675 0.655 1.1625 ;
      RECT 0.16 1.0975 0.655 1.1625 ;
      RECT 0.16 1.0975 0.225 2.235 ;
  END
END OR2X2

MACRO TBUFX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX1 0 0 ;
  SIZE 0.95 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.4875 0.9175 0.6025 1.0525 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.3475 0.7875 0.4125 1.0525 ;
        RECT 0.3475 0.7875 0.7425 0.8525 ;
    END
  END EN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.7775 0.1675 0.8725 0.7225 ;
        RECT 0.8075 0.1675 0.8725 2.24 ;
        RECT 0.7275 1.265 0.8725 2.24 ;
    END
  END Y
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.3975 -0.065 0.4625 0.6925 ;
        RECT 0 -0.065 0.95 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.3975 1.265 0.4625 2.535 ;
        RECT 0 2.405 0.95 2.535 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.6725 0.935 0.7375 1.2 ;
      RECT 0.2125 1.135 0.7375 1.2 ;
      RECT 0.2125 0.4475 0.2775 1.815 ;
  END
END TBUFX1

MACRO TBUFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX2 0 0 ;
  SIZE 1.33 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.4675 0.1675 0.5325 0.9825 ;
        RECT 0.3975 0.9175 0.5325 0.9825 ;
        RECT 0.4675 0.1675 0.9825 0.2325 ;
        RECT 0.9175 0.1675 0.9825 1.0525 ;
        RECT 0.9175 0.9175 1.0625 1.0525 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.1375 0.1525 0.2725 0.2225 ;
    END
  END EN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.7275 0.2975 0.7925 2.255 ;
    END
  END Y
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.3375 -0.065 0.4025 0.8525 ;
        RECT 1.1025 -0.065 1.1675 0.8525 ;
        RECT 0 -0.065 1.33 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.3375 1.345 0.4025 2.535 ;
        RECT 1.1025 1.345 1.1675 2.535 ;
        RECT 0 2.405 1.33 2.535 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.1175 0.3375 0.2525 0.8225 ;
      RECT 0.1525 1.12 0.6625 1.185 ;
      RECT 0.5975 1.12 0.6625 1.255 ;
      RECT 0.1525 0.3375 0.2175 2.235 ;
  END
END TBUFX2

MACRO XNOR2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2X1 0 0 ;
  SIZE 1.71 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.1075 0.7275 1.2875 0.9575 ;
        RECT 0.8575 0.8925 1.2875 0.9575 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.3475 1.1075 0.5325 1.1725 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.7275 0.2725 0.7925 1.9575 ;
        RECT 0.7275 0.2725 0.8225 0.8275 ;
        RECT 0.7275 1.2625 0.8225 1.9575 ;
    END
  END Y
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.3225 -0.065 0.3875 0.8275 ;
        RECT 1.1325 -0.065 1.1975 0.5475 ;
        RECT 0 -0.065 1.71 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.3775 2.1875 0.4425 2.535 ;
        RECT 1.1925 1.3475 1.2575 2.535 ;
        RECT 0 2.405 1.71 2.535 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.1375 0.2775 0.2025 0.9575 ;
      RECT 0.1375 0.8925 0.6625 0.9575 ;
      RECT 0.9975 1.1575 1.1325 1.2225 ;
      RECT 0.5975 0.8925 0.6625 2.0875 ;
      RECT 0.9975 1.1575 1.0625 2.0875 ;
      RECT 0.1925 2.0225 1.0625 2.0875 ;
      RECT 0.1925 1.2625 0.2575 2.2375 ;
      RECT 1.4275 0.13 1.5825 0.195 ;
      RECT 0.8675 1.0275 1.4925 1.0925 ;
      RECT 0.8675 1.0275 0.9325 1.1725 ;
      RECT 1.4275 0.13 1.4925 2.2375 ;
  END
END XNOR2X1

MACRO XOR2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2X1 0 0 ;
  SIZE 1.71 BY 2.47 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.5975 0.1675 0.6625 1.0125 ;
        RECT 0.5975 0.1675 0.9325 0.2325 ;
        RECT 0.8675 0.1675 0.9325 1.2225 ;
        RECT 0.8675 1.1575 1.0025 1.2225 ;
        RECT 0.8675 1.0275 1.3475 1.0925 ;
        RECT 1.2825 1.0275 1.3475 1.3625 ;
        RECT 1.2825 1.1575 1.4175 1.3625 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2575 0.9175 0.4125 1.1125 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.7275 0.2975 0.7925 1.5625 ;
        RECT 0.7275 1.2875 0.8475 1.5625 ;
    END
  END Y
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2925 -0.065 0.3575 0.8525 ;
        RECT 1.1025 -0.065 1.1675 0.7125 ;
        RECT 0 -0.065 1.71 0.065 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.2375 1.7675 0.3025 2.535 ;
        RECT 1.1975 1.4875 1.2625 2.535 ;
        RECT 0 2.405 1.71 2.535 ;
    END
  END vdd
  OBS
    LAYER metal1 ;
      RECT 0.0525 0.13 0.1875 0.195 ;
      RECT 1.0675 1.1575 1.2025 1.2225 ;
      RECT 1.0675 1.1575 1.1325 1.6925 ;
      RECT 0.0525 1.6275 1.1325 1.6925 ;
      RECT 0.0525 0.13 0.1175 2.2375 ;
      RECT 1.5225 0.3375 1.6575 0.8225 ;
      RECT 1.5225 0.3375 1.5875 0.9625 ;
      RECT 1.1225 0.8975 1.6225 0.9625 ;
      RECT 1.5575 0.8975 1.6225 2.2375 ;
  END
END XOR2X1

END LIBRARY
