VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO BUMP
  CLASS COVER BUMP ;
  ORIGIN 0 0 ;
  FOREIGN BUMP 0 0 ;
  SIZE 29 BY 29 ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT -5 -5 5 5 ;
    END
  END PAD
END BUMP