VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  LAYER LEF58_TYPE STRING ;
  LAYER LEF58_ENCLOSURE STRING ;
  LAYER LEF58_VOLTAGESPACING STRING ;
  LAYER LEF58_SPACING STRING ;
  LAYER LEF58_WIDTH STRING ;
  LAYER LEF58_ARRAYSPACING STRING ;
END PROPERTYDEFINITIONS

UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.005 ;
USEMINSPACING OBS OFF ;

LAYER M1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.770 0.770 ;
  WIDTH 0.395 ;
  OFFSET 0.385 0.000 ;
  AREA 0.230 ;
  SPACING 0.340 ;
  SPACING 0.340 LENGTHTHRESHOLD 1.880 RANGE 0.565 18.800 ;
  SPACING 0.415 RANGE 0.565 18.800 USELENGTHTHRESHOLD ;
  SPACING 1.130 RANGE 18.800 18800.000 ;
  SPACING 0.340 RANGE 0.000 18.800 INFLUENCE 0.340 ;
  SPACING 1.130 RANGE 18.800 18800.000 INFLUENCE 0.340 ;
  MINIMUMCUT 2 WIDTH 0.300 FROMABOVE ;
  MINWIDTH 0.300 ;
  MINENCLOSEDAREA 0.375 ;
END M1

LAYER V1
  TYPE CUT ;
  SPACING 0.415 ;
  WIDTH 0.355 ;
  ENCLOSURE BELOW 0.095 0.020 ;
  ENCLOSURE ABOVE 0.095 0.010 ;
END V1

LAYER M2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.770 0.770 ;
  WIDTH 0.375 ;
  OFFSET 0.385 0.000 ;
  AREA 0.270 ;
  SPACING 0.395 ;
  SPACING 0.395 LENGTHTHRESHOLD 1.880 RANGE 0.735 18.800 ;
  SPACING 0.450 RANGE 0.735 18.800 USELENGTHTHRESHOLD ;
  SPACING 1.130 RANGE 18.800 18800.000 ;
  SPACING 0.395 RANGE 0.000 18.800 INFLUENCE 0.395 ;
  SPACING 1.130 RANGE 18.800 18800.000 INFLUENCE 0.395 ;
  MINIMUMCUT 2 WIDTH 0.300 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 0.375 FROMABOVE ;
  MINENCLOSEDAREA 0.500 ;
END M2

LAYER V2
  TYPE CUT ;
  SPACING 0.415 ;
  WIDTH 0.355 ;
  ENCLOSURE BELOW 0.095 0.010 ;
  ENCLOSURE ABOVE 0.095 0.010 ;
END V2

LAYER M3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.770 0.770 ;
  WIDTH 0.375 ;
  OFFSET 0.385 0.000 ;
  AREA 0.270 ;
  SPACING 0.395 ;
  SPACING 0.395 LENGTHTHRESHOLD 1.880 RANGE 0.735 18.800 ;
  SPACING 0.450 RANGE 0.735 18.800 USELENGTHTHRESHOLD ;
  SPACING 1.130 RANGE 18.800 18800.000 ;
  SPACING 0.395 RANGE 0.000 18.800 INFLUENCE 0.395 ;
  SPACING 1.130 RANGE 18.800 18800.000 INFLUENCE 0.395 ;
  MINIMUMCUT 2 WIDTH 0.375 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 0.375 FROMABOVE ;
  MINIMUMCUT 3 WIDTH 3.950 FROMABOVE ;
  MINENCLOSEDAREA 0.500 ;
END M3

LAYER V3
  TYPE CUT ;
  SPACING 0.525 ;
  WIDTH 0.525 ;
  ENCLOSURE BELOW 0.245 0.190 ;
  ENCLOSURE ABOVE 1.270 1.270 WIDTH 3.760 ;
  ENCLOSURE ABOVE 2.115 2.115 WIDTH 7.520 ;
  ENCLOSURE ABOVE 3.150 3.150 WIDTH 13.160 ;
  ENCLOSURE ABOVE 4.090 4.090 WIDTH 52.640 ;
  ENCLOSURE ABOVE 0.675 1.130 ;
END V3

LAYER M4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 3.855 3.855 ;
  WIDTH 1.880 ;
  OFFSET 0.385 0.000 ;
  AREA 5.395 ;
  SPACING 1.880 ;
  SPACING 3.760 RANGE 13.160 26.320 ;
  SPACING 7.520 RANGE 26.320 52.640 ;
  SPACING 15.040 RANGE 52.640 105.280 ;
  SPACING 20.680 RANGE 105.280 161.680 ;
  SPACING 26.320 RANGE 161.680 18800.000 ;
  MINIMUMCUT 2 WIDTH 0.375 FROMBELOW ;
  MINIMUMCUT 3 WIDTH 3.950 FROMBELOW ;
  MINSTEP 0.470 MAXEDGES 0.000 ;
END M4

VIA M2_M1_VH_via DEFAULT
  LAYER M2 ;
    RECT -0.190 -0.275 0.190 0.275 ;
  LAYER M1 ;
    RECT -0.275 -0.195 0.275 0.195 ;
  LAYER V1 ;
    RECT -0.180 -0.180 0.180 0.180 ;
  RESISTANCE 2.630 ;
END M2_M1_VH_via

VIA M3_M2_HV_via DEFAULT
  LAYER M3 ;
    RECT -0.275 -0.190 0.275 0.190 ;
  LAYER M2 ;
    RECT -0.190 -0.275 0.190 0.275 ;
  LAYER V2 ;
    RECT -0.180 -0.180 0.180 0.180 ;
  RESISTANCE 2.630 ;
END M3_M2_HV_via

VIA M4_M3_CUT1
  LAYER V3 ;
    RECT -0.790 -0.265 -0.265 0.265 ;
  LAYER M4 ;
    RECT -1.920 -0.940 1.920 0.940 ;
  LAYER M3 ;
   RECT -1.035 -0.450 1.035 0.450 ;
  RESISTANCE 1.130 ;
END M4_M3_CUT1

SITE CORE
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.770 BY 9.250 ;
END CORE

MACRO CELL
  CLASS BLOCK ;
  ORIGIN 0.000 0.000 ;
  FOREIGN CELL 0.000 0.000 ;
  SIZE 788.230 BY 910.880 ;
  SYMMETRY X Y R90 ;
  PIN erase
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000 294.990 1.880 296.120 ;
      LAYER M2 ;
        RECT 0.000 294.990 1.880 296.120 ;
    END
  END erase
  PIN GND_0
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M3 ;
        RECT 92.610 903.380 111.410 910.880 ;
      LAYER M4 ;
        RECT 97.310 903.380 106.710 910.880 ;
    END
  END GND_0
  PIN VDD_0
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M3 ;
        RECT 780.710 394.840 788.230 413.640 ;
      LAYER M4 ;
        RECT 780.710 399.540 788.230 408.940 ;
    END
  END VDD_0
  OBS
    LAYER M1 ;
      RECT 0.000 0.000 788.230 910.880 ;
    LAYER M2 ;
      RECT 0.000 0.000 788.230 910.880 ;
    LAYER M3 ;
      RECT 0.000 0.000 788.230 910.880 ;
    LAYER M4 ;
      RECT 0.000 0.000 788.230 910.880 ;
    LAYER V1 ;
      RECT 0.000 0.000 788.230 910.880 ;
    LAYER V2 ;
      RECT 0.000 0.000 788.230 910.880 ;
    LAYER V3 ;
      RECT 0.000 0.000 788.230 910.880 ;
 END

END CELL

END LIBRARY
