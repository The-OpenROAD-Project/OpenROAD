VERSION 5.6 ;
#  NOWIREEXTENSIONATPIN ON ;
#  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
  DIVIDERCHAR "/" ;

#UNITS
#  DATABASE MICRONS 200 ;
#END UNITS

#LAYER via2
#  TYPE CUT ;
#END via2

#LAYER via
#  TYPE CUT ;
#END via

#LAYER nwell
#  TYPE MASTERSLICE ;
#END nwell

#LAYER via3
#  TYPE CUT ;
#END via3

#LAYER pwell
#  TYPE MASTERSLICE ;
#END pwell

#LAYER via4
#  TYPE CUT ;
#END via4

#LAYER mcon
#  TYPE CUT ;
#END mcon

#LAYER met6
#  TYPE ROUTING ;
#  WIDTH 0.030000 ;
#  SPACING 0.040000 ;
#  DIRECTION HORIZONTAL ;
#END met6

#LAYER met1
#  TYPE ROUTING ;
#  WIDTH 0.140000 ;
#  SPACING 0.140000 ;
#  DIRECTION HORIZONTAL ;
#END met1

#LAYER met3
#  TYPE ROUTING ;
#  WIDTH 0.300000 ;
#  SPACING 0.300000 ;
#  DIRECTION HORIZONTAL ;
#END met3

#LAYER met2
#  TYPE ROUTING ;
#  WIDTH 0.140000 ;
#  SPACING 0.140000 ;
#  DIRECTION HORIZONTAL ;
#END met2

#LAYER met4
#  TYPE ROUTING ;
#  WIDTH 0.300000 ;
#  SPACING 0.300000 ;
#  DIRECTION HORIZONTAL ;
#END met4

#LAYER met5
#  TYPE ROUTING ;
#  WIDTH 1.600000 ;
#  SPACING 1.600000 ;
#  DIRECTION HORIZONTAL ;
#END met5

#LAYER li1
#  TYPE ROUTING ;
#  WIDTH 0.170000 ;
#  SPACING 0.170000 ;
#  DIRECTION HORIZONTAL ;
#END li1

MACRO PT_UNIT_CELL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN PT_UNIT_CELL 0 0 ;
  SIZE 1.440 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN CTRL
#    ANTENNAGATEAREA 0.375000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.260 2.085 0.840 2.355 ;
    END
  END CTRL
  PIN VREG
 #   ANTENNAGATEAREA 0.375000 ;
 #   ANTENNADIFFAREA 0.213750 ;
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.940 2.655 1.345 3.480 ;
        RECT 1.025 1.715 1.345 2.655 ;
        RECT 0.500 1.380 1.345 1.715 ;
    END
  END VREG
  PIN vgnd
  #  ANTENNADIFFAREA 0.427500 ;
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.255 0.625 1.210 ;
        RECT 0.830 0.255 1.350 1.210 ;
      LAYER mcon ;
        RECT 0.280 0.310 0.450 0.480 ;
        RECT 1.060 0.310 1.230 0.480 ;
      LAYER met1 ;
        RECT 0.000 0.255 1.440 0.625 ;
    END
  END vgnd
  PIN vpb
#    ANTENNADIFFAREA 0.244800 ;
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      #LAYER nwell ;
      #  RECT -0.330 1.885 1.770 4.490 ;
      LAYER li1 ;
        RECT 0.000 3.985 1.440 4.155 ;
      LAYER mcon ;
        RECT 0.155 3.985 0.325 4.155 ;
        RECT 0.635 3.985 0.805 4.155 ;
        RECT 1.115 3.985 1.285 4.155 ;
      LAYER met1 ;
        RECT 0.000 3.955 1.440 4.185 ;
    END
  END vpb
  PIN vnb
#    ANTENNADIFFAREA 0.244800 ;
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      #LAYER pwell ;
      #  RECT 0.090 0.215 1.420 1.415 ;
      #  RECT -0.130 -0.215 1.570 0.215 ;
      LAYER li1 ;
        RECT 0.000 -0.085 1.440 0.085 ;
      LAYER mcon ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.115 1.440 0.115 ;
    END
  END vnb
  PIN vpwr
#    ANTENNADIFFAREA 0.213750 ;
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.090 2.655 0.680 3.730 ;
      LAYER mcon ;
        RECT 0.120 3.500 0.290 3.670 ;
        RECT 0.480 3.500 0.650 3.670 ;
      LAYER met1 ;
        RECT 0.000 3.445 1.440 3.815 ;
    END
  END vpwr
END PT_UNIT_CELL
END LIBRARY

