VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 2000 ;
END UNITS

MACRO BLOCK1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SIZE 50 BY 50 ;
  PIN A
    DIRECTION INPUT ;
  END A
  PIN Z
    DIRECTION OUTPUT ;
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
  END VSS
END BLOCK1
