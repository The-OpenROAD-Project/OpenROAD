../../../test/pad.lef