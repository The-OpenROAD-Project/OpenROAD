# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_io__overlay_vdda_hvc
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 200 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 1.270000 56.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 53.125000 75.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 1.270000 51.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 48.365000 75.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 8.885000 1.270000 13.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 8.885000 75.000000 13.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 8.985000 1.270000 13.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 8.985000 75.000000 13.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2.035000 1.270000 7.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 2.035000 75.000000 7.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 2.135000 1.270000 7.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 2.135000 75.000000 7.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.495000 14.940000 24.395000 18.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390000 14.940000 74.290000 18.380000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 14.935000 24.370000 18.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.415000 14.935000 75.000000 18.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 15.035000 0.965000 18.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 15.035000 75.000000 18.285000 ;
    END
    PORT
      LAYER via3 ;
        RECT  0.585000 15.020000  0.785000 15.220000 ;
        RECT  0.585000 15.460000  0.785000 15.660000 ;
        RECT  0.585000 15.900000  0.785000 16.100000 ;
        RECT  0.585000 16.340000  0.785000 16.540000 ;
        RECT  0.585000 16.780000  0.785000 16.980000 ;
        RECT  0.585000 17.220000  0.785000 17.420000 ;
        RECT  0.585000 17.660000  0.785000 17.860000 ;
        RECT  0.585000 18.100000  0.785000 18.300000 ;
        RECT  0.995000 15.020000  1.195000 15.220000 ;
        RECT  0.995000 15.460000  1.195000 15.660000 ;
        RECT  0.995000 15.900000  1.195000 16.100000 ;
        RECT  0.995000 16.340000  1.195000 16.540000 ;
        RECT  0.995000 16.780000  1.195000 16.980000 ;
        RECT  0.995000 17.220000  1.195000 17.420000 ;
        RECT  0.995000 17.660000  1.195000 17.860000 ;
        RECT  0.995000 18.100000  1.195000 18.300000 ;
        RECT  1.405000 15.020000  1.605000 15.220000 ;
        RECT  1.405000 15.460000  1.605000 15.660000 ;
        RECT  1.405000 15.900000  1.605000 16.100000 ;
        RECT  1.405000 16.340000  1.605000 16.540000 ;
        RECT  1.405000 16.780000  1.605000 16.980000 ;
        RECT  1.405000 17.220000  1.605000 17.420000 ;
        RECT  1.405000 17.660000  1.605000 17.860000 ;
        RECT  1.405000 18.100000  1.605000 18.300000 ;
        RECT  1.815000 15.020000  2.015000 15.220000 ;
        RECT  1.815000 15.460000  2.015000 15.660000 ;
        RECT  1.815000 15.900000  2.015000 16.100000 ;
        RECT  1.815000 16.340000  2.015000 16.540000 ;
        RECT  1.815000 16.780000  2.015000 16.980000 ;
        RECT  1.815000 17.220000  2.015000 17.420000 ;
        RECT  1.815000 17.660000  2.015000 17.860000 ;
        RECT  1.815000 18.100000  2.015000 18.300000 ;
        RECT  2.225000 15.020000  2.425000 15.220000 ;
        RECT  2.225000 15.460000  2.425000 15.660000 ;
        RECT  2.225000 15.900000  2.425000 16.100000 ;
        RECT  2.225000 16.340000  2.425000 16.540000 ;
        RECT  2.225000 16.780000  2.425000 16.980000 ;
        RECT  2.225000 17.220000  2.425000 17.420000 ;
        RECT  2.225000 17.660000  2.425000 17.860000 ;
        RECT  2.225000 18.100000  2.425000 18.300000 ;
        RECT  2.635000 15.020000  2.835000 15.220000 ;
        RECT  2.635000 15.460000  2.835000 15.660000 ;
        RECT  2.635000 15.900000  2.835000 16.100000 ;
        RECT  2.635000 16.340000  2.835000 16.540000 ;
        RECT  2.635000 16.780000  2.835000 16.980000 ;
        RECT  2.635000 17.220000  2.835000 17.420000 ;
        RECT  2.635000 17.660000  2.835000 17.860000 ;
        RECT  2.635000 18.100000  2.835000 18.300000 ;
        RECT  3.045000 15.020000  3.245000 15.220000 ;
        RECT  3.045000 15.460000  3.245000 15.660000 ;
        RECT  3.045000 15.900000  3.245000 16.100000 ;
        RECT  3.045000 16.340000  3.245000 16.540000 ;
        RECT  3.045000 16.780000  3.245000 16.980000 ;
        RECT  3.045000 17.220000  3.245000 17.420000 ;
        RECT  3.045000 17.660000  3.245000 17.860000 ;
        RECT  3.045000 18.100000  3.245000 18.300000 ;
        RECT  3.450000 15.020000  3.650000 15.220000 ;
        RECT  3.450000 15.460000  3.650000 15.660000 ;
        RECT  3.450000 15.900000  3.650000 16.100000 ;
        RECT  3.450000 16.340000  3.650000 16.540000 ;
        RECT  3.450000 16.780000  3.650000 16.980000 ;
        RECT  3.450000 17.220000  3.650000 17.420000 ;
        RECT  3.450000 17.660000  3.650000 17.860000 ;
        RECT  3.450000 18.100000  3.650000 18.300000 ;
        RECT  3.855000 15.020000  4.055000 15.220000 ;
        RECT  3.855000 15.460000  4.055000 15.660000 ;
        RECT  3.855000 15.900000  4.055000 16.100000 ;
        RECT  3.855000 16.340000  4.055000 16.540000 ;
        RECT  3.855000 16.780000  4.055000 16.980000 ;
        RECT  3.855000 17.220000  4.055000 17.420000 ;
        RECT  3.855000 17.660000  4.055000 17.860000 ;
        RECT  3.855000 18.100000  4.055000 18.300000 ;
        RECT  4.260000 15.020000  4.460000 15.220000 ;
        RECT  4.260000 15.460000  4.460000 15.660000 ;
        RECT  4.260000 15.900000  4.460000 16.100000 ;
        RECT  4.260000 16.340000  4.460000 16.540000 ;
        RECT  4.260000 16.780000  4.460000 16.980000 ;
        RECT  4.260000 17.220000  4.460000 17.420000 ;
        RECT  4.260000 17.660000  4.460000 17.860000 ;
        RECT  4.260000 18.100000  4.460000 18.300000 ;
        RECT  4.665000 15.020000  4.865000 15.220000 ;
        RECT  4.665000 15.460000  4.865000 15.660000 ;
        RECT  4.665000 15.900000  4.865000 16.100000 ;
        RECT  4.665000 16.340000  4.865000 16.540000 ;
        RECT  4.665000 16.780000  4.865000 16.980000 ;
        RECT  4.665000 17.220000  4.865000 17.420000 ;
        RECT  4.665000 17.660000  4.865000 17.860000 ;
        RECT  4.665000 18.100000  4.865000 18.300000 ;
        RECT  5.070000 15.020000  5.270000 15.220000 ;
        RECT  5.070000 15.460000  5.270000 15.660000 ;
        RECT  5.070000 15.900000  5.270000 16.100000 ;
        RECT  5.070000 16.340000  5.270000 16.540000 ;
        RECT  5.070000 16.780000  5.270000 16.980000 ;
        RECT  5.070000 17.220000  5.270000 17.420000 ;
        RECT  5.070000 17.660000  5.270000 17.860000 ;
        RECT  5.070000 18.100000  5.270000 18.300000 ;
        RECT  5.475000 15.020000  5.675000 15.220000 ;
        RECT  5.475000 15.460000  5.675000 15.660000 ;
        RECT  5.475000 15.900000  5.675000 16.100000 ;
        RECT  5.475000 16.340000  5.675000 16.540000 ;
        RECT  5.475000 16.780000  5.675000 16.980000 ;
        RECT  5.475000 17.220000  5.675000 17.420000 ;
        RECT  5.475000 17.660000  5.675000 17.860000 ;
        RECT  5.475000 18.100000  5.675000 18.300000 ;
        RECT  5.880000 15.020000  6.080000 15.220000 ;
        RECT  5.880000 15.460000  6.080000 15.660000 ;
        RECT  5.880000 15.900000  6.080000 16.100000 ;
        RECT  5.880000 16.340000  6.080000 16.540000 ;
        RECT  5.880000 16.780000  6.080000 16.980000 ;
        RECT  5.880000 17.220000  6.080000 17.420000 ;
        RECT  5.880000 17.660000  6.080000 17.860000 ;
        RECT  5.880000 18.100000  6.080000 18.300000 ;
        RECT  6.285000 15.020000  6.485000 15.220000 ;
        RECT  6.285000 15.460000  6.485000 15.660000 ;
        RECT  6.285000 15.900000  6.485000 16.100000 ;
        RECT  6.285000 16.340000  6.485000 16.540000 ;
        RECT  6.285000 16.780000  6.485000 16.980000 ;
        RECT  6.285000 17.220000  6.485000 17.420000 ;
        RECT  6.285000 17.660000  6.485000 17.860000 ;
        RECT  6.285000 18.100000  6.485000 18.300000 ;
        RECT  6.690000 15.020000  6.890000 15.220000 ;
        RECT  6.690000 15.460000  6.890000 15.660000 ;
        RECT  6.690000 15.900000  6.890000 16.100000 ;
        RECT  6.690000 16.340000  6.890000 16.540000 ;
        RECT  6.690000 16.780000  6.890000 16.980000 ;
        RECT  6.690000 17.220000  6.890000 17.420000 ;
        RECT  6.690000 17.660000  6.890000 17.860000 ;
        RECT  6.690000 18.100000  6.890000 18.300000 ;
        RECT  7.095000 15.020000  7.295000 15.220000 ;
        RECT  7.095000 15.460000  7.295000 15.660000 ;
        RECT  7.095000 15.900000  7.295000 16.100000 ;
        RECT  7.095000 16.340000  7.295000 16.540000 ;
        RECT  7.095000 16.780000  7.295000 16.980000 ;
        RECT  7.095000 17.220000  7.295000 17.420000 ;
        RECT  7.095000 17.660000  7.295000 17.860000 ;
        RECT  7.095000 18.100000  7.295000 18.300000 ;
        RECT  7.500000 15.020000  7.700000 15.220000 ;
        RECT  7.500000 15.460000  7.700000 15.660000 ;
        RECT  7.500000 15.900000  7.700000 16.100000 ;
        RECT  7.500000 16.340000  7.700000 16.540000 ;
        RECT  7.500000 16.780000  7.700000 16.980000 ;
        RECT  7.500000 17.220000  7.700000 17.420000 ;
        RECT  7.500000 17.660000  7.700000 17.860000 ;
        RECT  7.500000 18.100000  7.700000 18.300000 ;
        RECT  7.905000 15.020000  8.105000 15.220000 ;
        RECT  7.905000 15.460000  8.105000 15.660000 ;
        RECT  7.905000 15.900000  8.105000 16.100000 ;
        RECT  7.905000 16.340000  8.105000 16.540000 ;
        RECT  7.905000 16.780000  8.105000 16.980000 ;
        RECT  7.905000 17.220000  8.105000 17.420000 ;
        RECT  7.905000 17.660000  8.105000 17.860000 ;
        RECT  7.905000 18.100000  8.105000 18.300000 ;
        RECT  8.310000 15.020000  8.510000 15.220000 ;
        RECT  8.310000 15.460000  8.510000 15.660000 ;
        RECT  8.310000 15.900000  8.510000 16.100000 ;
        RECT  8.310000 16.340000  8.510000 16.540000 ;
        RECT  8.310000 16.780000  8.510000 16.980000 ;
        RECT  8.310000 17.220000  8.510000 17.420000 ;
        RECT  8.310000 17.660000  8.510000 17.860000 ;
        RECT  8.310000 18.100000  8.510000 18.300000 ;
        RECT  8.715000 15.020000  8.915000 15.220000 ;
        RECT  8.715000 15.460000  8.915000 15.660000 ;
        RECT  8.715000 15.900000  8.915000 16.100000 ;
        RECT  8.715000 16.340000  8.915000 16.540000 ;
        RECT  8.715000 16.780000  8.915000 16.980000 ;
        RECT  8.715000 17.220000  8.915000 17.420000 ;
        RECT  8.715000 17.660000  8.915000 17.860000 ;
        RECT  8.715000 18.100000  8.915000 18.300000 ;
        RECT  9.120000 15.020000  9.320000 15.220000 ;
        RECT  9.120000 15.460000  9.320000 15.660000 ;
        RECT  9.120000 15.900000  9.320000 16.100000 ;
        RECT  9.120000 16.340000  9.320000 16.540000 ;
        RECT  9.120000 16.780000  9.320000 16.980000 ;
        RECT  9.120000 17.220000  9.320000 17.420000 ;
        RECT  9.120000 17.660000  9.320000 17.860000 ;
        RECT  9.120000 18.100000  9.320000 18.300000 ;
        RECT  9.525000 15.020000  9.725000 15.220000 ;
        RECT  9.525000 15.460000  9.725000 15.660000 ;
        RECT  9.525000 15.900000  9.725000 16.100000 ;
        RECT  9.525000 16.340000  9.725000 16.540000 ;
        RECT  9.525000 16.780000  9.725000 16.980000 ;
        RECT  9.525000 17.220000  9.725000 17.420000 ;
        RECT  9.525000 17.660000  9.725000 17.860000 ;
        RECT  9.525000 18.100000  9.725000 18.300000 ;
        RECT  9.930000 15.020000 10.130000 15.220000 ;
        RECT  9.930000 15.460000 10.130000 15.660000 ;
        RECT  9.930000 15.900000 10.130000 16.100000 ;
        RECT  9.930000 16.340000 10.130000 16.540000 ;
        RECT  9.930000 16.780000 10.130000 16.980000 ;
        RECT  9.930000 17.220000 10.130000 17.420000 ;
        RECT  9.930000 17.660000 10.130000 17.860000 ;
        RECT  9.930000 18.100000 10.130000 18.300000 ;
        RECT 10.335000 15.020000 10.535000 15.220000 ;
        RECT 10.335000 15.460000 10.535000 15.660000 ;
        RECT 10.335000 15.900000 10.535000 16.100000 ;
        RECT 10.335000 16.340000 10.535000 16.540000 ;
        RECT 10.335000 16.780000 10.535000 16.980000 ;
        RECT 10.335000 17.220000 10.535000 17.420000 ;
        RECT 10.335000 17.660000 10.535000 17.860000 ;
        RECT 10.335000 18.100000 10.535000 18.300000 ;
        RECT 10.740000 15.020000 10.940000 15.220000 ;
        RECT 10.740000 15.460000 10.940000 15.660000 ;
        RECT 10.740000 15.900000 10.940000 16.100000 ;
        RECT 10.740000 16.340000 10.940000 16.540000 ;
        RECT 10.740000 16.780000 10.940000 16.980000 ;
        RECT 10.740000 17.220000 10.940000 17.420000 ;
        RECT 10.740000 17.660000 10.940000 17.860000 ;
        RECT 10.740000 18.100000 10.940000 18.300000 ;
        RECT 11.145000 15.020000 11.345000 15.220000 ;
        RECT 11.145000 15.460000 11.345000 15.660000 ;
        RECT 11.145000 15.900000 11.345000 16.100000 ;
        RECT 11.145000 16.340000 11.345000 16.540000 ;
        RECT 11.145000 16.780000 11.345000 16.980000 ;
        RECT 11.145000 17.220000 11.345000 17.420000 ;
        RECT 11.145000 17.660000 11.345000 17.860000 ;
        RECT 11.145000 18.100000 11.345000 18.300000 ;
        RECT 11.550000 15.020000 11.750000 15.220000 ;
        RECT 11.550000 15.460000 11.750000 15.660000 ;
        RECT 11.550000 15.900000 11.750000 16.100000 ;
        RECT 11.550000 16.340000 11.750000 16.540000 ;
        RECT 11.550000 16.780000 11.750000 16.980000 ;
        RECT 11.550000 17.220000 11.750000 17.420000 ;
        RECT 11.550000 17.660000 11.750000 17.860000 ;
        RECT 11.550000 18.100000 11.750000 18.300000 ;
        RECT 11.955000 15.020000 12.155000 15.220000 ;
        RECT 11.955000 15.460000 12.155000 15.660000 ;
        RECT 11.955000 15.900000 12.155000 16.100000 ;
        RECT 11.955000 16.340000 12.155000 16.540000 ;
        RECT 11.955000 16.780000 12.155000 16.980000 ;
        RECT 11.955000 17.220000 12.155000 17.420000 ;
        RECT 11.955000 17.660000 12.155000 17.860000 ;
        RECT 11.955000 18.100000 12.155000 18.300000 ;
        RECT 12.360000 15.020000 12.560000 15.220000 ;
        RECT 12.360000 15.460000 12.560000 15.660000 ;
        RECT 12.360000 15.900000 12.560000 16.100000 ;
        RECT 12.360000 16.340000 12.560000 16.540000 ;
        RECT 12.360000 16.780000 12.560000 16.980000 ;
        RECT 12.360000 17.220000 12.560000 17.420000 ;
        RECT 12.360000 17.660000 12.560000 17.860000 ;
        RECT 12.360000 18.100000 12.560000 18.300000 ;
        RECT 12.765000 15.020000 12.965000 15.220000 ;
        RECT 12.765000 15.460000 12.965000 15.660000 ;
        RECT 12.765000 15.900000 12.965000 16.100000 ;
        RECT 12.765000 16.340000 12.965000 16.540000 ;
        RECT 12.765000 16.780000 12.965000 16.980000 ;
        RECT 12.765000 17.220000 12.965000 17.420000 ;
        RECT 12.765000 17.660000 12.965000 17.860000 ;
        RECT 12.765000 18.100000 12.965000 18.300000 ;
        RECT 13.170000 15.020000 13.370000 15.220000 ;
        RECT 13.170000 15.460000 13.370000 15.660000 ;
        RECT 13.170000 15.900000 13.370000 16.100000 ;
        RECT 13.170000 16.340000 13.370000 16.540000 ;
        RECT 13.170000 16.780000 13.370000 16.980000 ;
        RECT 13.170000 17.220000 13.370000 17.420000 ;
        RECT 13.170000 17.660000 13.370000 17.860000 ;
        RECT 13.170000 18.100000 13.370000 18.300000 ;
        RECT 13.575000 15.020000 13.775000 15.220000 ;
        RECT 13.575000 15.460000 13.775000 15.660000 ;
        RECT 13.575000 15.900000 13.775000 16.100000 ;
        RECT 13.575000 16.340000 13.775000 16.540000 ;
        RECT 13.575000 16.780000 13.775000 16.980000 ;
        RECT 13.575000 17.220000 13.775000 17.420000 ;
        RECT 13.575000 17.660000 13.775000 17.860000 ;
        RECT 13.575000 18.100000 13.775000 18.300000 ;
        RECT 13.980000 15.020000 14.180000 15.220000 ;
        RECT 13.980000 15.460000 14.180000 15.660000 ;
        RECT 13.980000 15.900000 14.180000 16.100000 ;
        RECT 13.980000 16.340000 14.180000 16.540000 ;
        RECT 13.980000 16.780000 14.180000 16.980000 ;
        RECT 13.980000 17.220000 14.180000 17.420000 ;
        RECT 13.980000 17.660000 14.180000 17.860000 ;
        RECT 13.980000 18.100000 14.180000 18.300000 ;
        RECT 14.385000 15.020000 14.585000 15.220000 ;
        RECT 14.385000 15.460000 14.585000 15.660000 ;
        RECT 14.385000 15.900000 14.585000 16.100000 ;
        RECT 14.385000 16.340000 14.585000 16.540000 ;
        RECT 14.385000 16.780000 14.585000 16.980000 ;
        RECT 14.385000 17.220000 14.585000 17.420000 ;
        RECT 14.385000 17.660000 14.585000 17.860000 ;
        RECT 14.385000 18.100000 14.585000 18.300000 ;
        RECT 14.790000 15.020000 14.990000 15.220000 ;
        RECT 14.790000 15.460000 14.990000 15.660000 ;
        RECT 14.790000 15.900000 14.990000 16.100000 ;
        RECT 14.790000 16.340000 14.990000 16.540000 ;
        RECT 14.790000 16.780000 14.990000 16.980000 ;
        RECT 14.790000 17.220000 14.990000 17.420000 ;
        RECT 14.790000 17.660000 14.990000 17.860000 ;
        RECT 14.790000 18.100000 14.990000 18.300000 ;
        RECT 15.195000 15.020000 15.395000 15.220000 ;
        RECT 15.195000 15.460000 15.395000 15.660000 ;
        RECT 15.195000 15.900000 15.395000 16.100000 ;
        RECT 15.195000 16.340000 15.395000 16.540000 ;
        RECT 15.195000 16.780000 15.395000 16.980000 ;
        RECT 15.195000 17.220000 15.395000 17.420000 ;
        RECT 15.195000 17.660000 15.395000 17.860000 ;
        RECT 15.195000 18.100000 15.395000 18.300000 ;
        RECT 15.600000 15.020000 15.800000 15.220000 ;
        RECT 15.600000 15.460000 15.800000 15.660000 ;
        RECT 15.600000 15.900000 15.800000 16.100000 ;
        RECT 15.600000 16.340000 15.800000 16.540000 ;
        RECT 15.600000 16.780000 15.800000 16.980000 ;
        RECT 15.600000 17.220000 15.800000 17.420000 ;
        RECT 15.600000 17.660000 15.800000 17.860000 ;
        RECT 15.600000 18.100000 15.800000 18.300000 ;
        RECT 16.005000 15.020000 16.205000 15.220000 ;
        RECT 16.005000 15.460000 16.205000 15.660000 ;
        RECT 16.005000 15.900000 16.205000 16.100000 ;
        RECT 16.005000 16.340000 16.205000 16.540000 ;
        RECT 16.005000 16.780000 16.205000 16.980000 ;
        RECT 16.005000 17.220000 16.205000 17.420000 ;
        RECT 16.005000 17.660000 16.205000 17.860000 ;
        RECT 16.005000 18.100000 16.205000 18.300000 ;
        RECT 16.410000 15.020000 16.610000 15.220000 ;
        RECT 16.410000 15.460000 16.610000 15.660000 ;
        RECT 16.410000 15.900000 16.610000 16.100000 ;
        RECT 16.410000 16.340000 16.610000 16.540000 ;
        RECT 16.410000 16.780000 16.610000 16.980000 ;
        RECT 16.410000 17.220000 16.610000 17.420000 ;
        RECT 16.410000 17.660000 16.610000 17.860000 ;
        RECT 16.410000 18.100000 16.610000 18.300000 ;
        RECT 16.815000 15.020000 17.015000 15.220000 ;
        RECT 16.815000 15.460000 17.015000 15.660000 ;
        RECT 16.815000 15.900000 17.015000 16.100000 ;
        RECT 16.815000 16.340000 17.015000 16.540000 ;
        RECT 16.815000 16.780000 17.015000 16.980000 ;
        RECT 16.815000 17.220000 17.015000 17.420000 ;
        RECT 16.815000 17.660000 17.015000 17.860000 ;
        RECT 16.815000 18.100000 17.015000 18.300000 ;
        RECT 17.220000 15.020000 17.420000 15.220000 ;
        RECT 17.220000 15.460000 17.420000 15.660000 ;
        RECT 17.220000 15.900000 17.420000 16.100000 ;
        RECT 17.220000 16.340000 17.420000 16.540000 ;
        RECT 17.220000 16.780000 17.420000 16.980000 ;
        RECT 17.220000 17.220000 17.420000 17.420000 ;
        RECT 17.220000 17.660000 17.420000 17.860000 ;
        RECT 17.220000 18.100000 17.420000 18.300000 ;
        RECT 17.625000 15.020000 17.825000 15.220000 ;
        RECT 17.625000 15.460000 17.825000 15.660000 ;
        RECT 17.625000 15.900000 17.825000 16.100000 ;
        RECT 17.625000 16.340000 17.825000 16.540000 ;
        RECT 17.625000 16.780000 17.825000 16.980000 ;
        RECT 17.625000 17.220000 17.825000 17.420000 ;
        RECT 17.625000 17.660000 17.825000 17.860000 ;
        RECT 17.625000 18.100000 17.825000 18.300000 ;
        RECT 18.030000 15.020000 18.230000 15.220000 ;
        RECT 18.030000 15.460000 18.230000 15.660000 ;
        RECT 18.030000 15.900000 18.230000 16.100000 ;
        RECT 18.030000 16.340000 18.230000 16.540000 ;
        RECT 18.030000 16.780000 18.230000 16.980000 ;
        RECT 18.030000 17.220000 18.230000 17.420000 ;
        RECT 18.030000 17.660000 18.230000 17.860000 ;
        RECT 18.030000 18.100000 18.230000 18.300000 ;
        RECT 18.435000 15.020000 18.635000 15.220000 ;
        RECT 18.435000 15.460000 18.635000 15.660000 ;
        RECT 18.435000 15.900000 18.635000 16.100000 ;
        RECT 18.435000 16.340000 18.635000 16.540000 ;
        RECT 18.435000 16.780000 18.635000 16.980000 ;
        RECT 18.435000 17.220000 18.635000 17.420000 ;
        RECT 18.435000 17.660000 18.635000 17.860000 ;
        RECT 18.435000 18.100000 18.635000 18.300000 ;
        RECT 18.840000 15.020000 19.040000 15.220000 ;
        RECT 18.840000 15.460000 19.040000 15.660000 ;
        RECT 18.840000 15.900000 19.040000 16.100000 ;
        RECT 18.840000 16.340000 19.040000 16.540000 ;
        RECT 18.840000 16.780000 19.040000 16.980000 ;
        RECT 18.840000 17.220000 19.040000 17.420000 ;
        RECT 18.840000 17.660000 19.040000 17.860000 ;
        RECT 18.840000 18.100000 19.040000 18.300000 ;
        RECT 19.245000 15.020000 19.445000 15.220000 ;
        RECT 19.245000 15.460000 19.445000 15.660000 ;
        RECT 19.245000 15.900000 19.445000 16.100000 ;
        RECT 19.245000 16.340000 19.445000 16.540000 ;
        RECT 19.245000 16.780000 19.445000 16.980000 ;
        RECT 19.245000 17.220000 19.445000 17.420000 ;
        RECT 19.245000 17.660000 19.445000 17.860000 ;
        RECT 19.245000 18.100000 19.445000 18.300000 ;
        RECT 19.650000 15.020000 19.850000 15.220000 ;
        RECT 19.650000 15.460000 19.850000 15.660000 ;
        RECT 19.650000 15.900000 19.850000 16.100000 ;
        RECT 19.650000 16.340000 19.850000 16.540000 ;
        RECT 19.650000 16.780000 19.850000 16.980000 ;
        RECT 19.650000 17.220000 19.850000 17.420000 ;
        RECT 19.650000 17.660000 19.850000 17.860000 ;
        RECT 19.650000 18.100000 19.850000 18.300000 ;
        RECT 20.055000 15.020000 20.255000 15.220000 ;
        RECT 20.055000 15.460000 20.255000 15.660000 ;
        RECT 20.055000 15.900000 20.255000 16.100000 ;
        RECT 20.055000 16.340000 20.255000 16.540000 ;
        RECT 20.055000 16.780000 20.255000 16.980000 ;
        RECT 20.055000 17.220000 20.255000 17.420000 ;
        RECT 20.055000 17.660000 20.255000 17.860000 ;
        RECT 20.055000 18.100000 20.255000 18.300000 ;
        RECT 20.460000 15.020000 20.660000 15.220000 ;
        RECT 20.460000 15.460000 20.660000 15.660000 ;
        RECT 20.460000 15.900000 20.660000 16.100000 ;
        RECT 20.460000 16.340000 20.660000 16.540000 ;
        RECT 20.460000 16.780000 20.660000 16.980000 ;
        RECT 20.460000 17.220000 20.660000 17.420000 ;
        RECT 20.460000 17.660000 20.660000 17.860000 ;
        RECT 20.460000 18.100000 20.660000 18.300000 ;
        RECT 20.865000 15.020000 21.065000 15.220000 ;
        RECT 20.865000 15.460000 21.065000 15.660000 ;
        RECT 20.865000 15.900000 21.065000 16.100000 ;
        RECT 20.865000 16.340000 21.065000 16.540000 ;
        RECT 20.865000 16.780000 21.065000 16.980000 ;
        RECT 20.865000 17.220000 21.065000 17.420000 ;
        RECT 20.865000 17.660000 21.065000 17.860000 ;
        RECT 20.865000 18.100000 21.065000 18.300000 ;
        RECT 21.270000 15.020000 21.470000 15.220000 ;
        RECT 21.270000 15.460000 21.470000 15.660000 ;
        RECT 21.270000 15.900000 21.470000 16.100000 ;
        RECT 21.270000 16.340000 21.470000 16.540000 ;
        RECT 21.270000 16.780000 21.470000 16.980000 ;
        RECT 21.270000 17.220000 21.470000 17.420000 ;
        RECT 21.270000 17.660000 21.470000 17.860000 ;
        RECT 21.270000 18.100000 21.470000 18.300000 ;
        RECT 21.675000 15.020000 21.875000 15.220000 ;
        RECT 21.675000 15.460000 21.875000 15.660000 ;
        RECT 21.675000 15.900000 21.875000 16.100000 ;
        RECT 21.675000 16.340000 21.875000 16.540000 ;
        RECT 21.675000 16.780000 21.875000 16.980000 ;
        RECT 21.675000 17.220000 21.875000 17.420000 ;
        RECT 21.675000 17.660000 21.875000 17.860000 ;
        RECT 21.675000 18.100000 21.875000 18.300000 ;
        RECT 22.080000 15.020000 22.280000 15.220000 ;
        RECT 22.080000 15.460000 22.280000 15.660000 ;
        RECT 22.080000 15.900000 22.280000 16.100000 ;
        RECT 22.080000 16.340000 22.280000 16.540000 ;
        RECT 22.080000 16.780000 22.280000 16.980000 ;
        RECT 22.080000 17.220000 22.280000 17.420000 ;
        RECT 22.080000 17.660000 22.280000 17.860000 ;
        RECT 22.080000 18.100000 22.280000 18.300000 ;
        RECT 22.485000 15.020000 22.685000 15.220000 ;
        RECT 22.485000 15.460000 22.685000 15.660000 ;
        RECT 22.485000 15.900000 22.685000 16.100000 ;
        RECT 22.485000 16.340000 22.685000 16.540000 ;
        RECT 22.485000 16.780000 22.685000 16.980000 ;
        RECT 22.485000 17.220000 22.685000 17.420000 ;
        RECT 22.485000 17.660000 22.685000 17.860000 ;
        RECT 22.485000 18.100000 22.685000 18.300000 ;
        RECT 22.890000 15.020000 23.090000 15.220000 ;
        RECT 22.890000 15.460000 23.090000 15.660000 ;
        RECT 22.890000 15.900000 23.090000 16.100000 ;
        RECT 22.890000 16.340000 23.090000 16.540000 ;
        RECT 22.890000 16.780000 23.090000 16.980000 ;
        RECT 22.890000 17.220000 23.090000 17.420000 ;
        RECT 22.890000 17.660000 23.090000 17.860000 ;
        RECT 22.890000 18.100000 23.090000 18.300000 ;
        RECT 23.295000 15.020000 23.495000 15.220000 ;
        RECT 23.295000 15.460000 23.495000 15.660000 ;
        RECT 23.295000 15.900000 23.495000 16.100000 ;
        RECT 23.295000 16.340000 23.495000 16.540000 ;
        RECT 23.295000 16.780000 23.495000 16.980000 ;
        RECT 23.295000 17.220000 23.495000 17.420000 ;
        RECT 23.295000 17.660000 23.495000 17.860000 ;
        RECT 23.295000 18.100000 23.495000 18.300000 ;
        RECT 23.700000 15.020000 23.900000 15.220000 ;
        RECT 23.700000 15.460000 23.900000 15.660000 ;
        RECT 23.700000 15.900000 23.900000 16.100000 ;
        RECT 23.700000 16.340000 23.900000 16.540000 ;
        RECT 23.700000 16.780000 23.900000 16.980000 ;
        RECT 23.700000 17.220000 23.900000 17.420000 ;
        RECT 23.700000 17.660000 23.900000 17.860000 ;
        RECT 23.700000 18.100000 23.900000 18.300000 ;
        RECT 24.105000 15.020000 24.305000 15.220000 ;
        RECT 24.105000 15.460000 24.305000 15.660000 ;
        RECT 24.105000 15.900000 24.305000 16.100000 ;
        RECT 24.105000 16.340000 24.305000 16.540000 ;
        RECT 24.105000 16.780000 24.305000 16.980000 ;
        RECT 24.105000 17.220000 24.305000 17.420000 ;
        RECT 24.105000 17.660000 24.305000 17.860000 ;
        RECT 24.105000 18.100000 24.305000 18.300000 ;
        RECT 50.480000 15.020000 50.680000 15.220000 ;
        RECT 50.480000 15.460000 50.680000 15.660000 ;
        RECT 50.480000 15.900000 50.680000 16.100000 ;
        RECT 50.480000 16.340000 50.680000 16.540000 ;
        RECT 50.480000 16.780000 50.680000 16.980000 ;
        RECT 50.480000 17.220000 50.680000 17.420000 ;
        RECT 50.480000 17.660000 50.680000 17.860000 ;
        RECT 50.480000 18.100000 50.680000 18.300000 ;
        RECT 50.890000 15.020000 51.090000 15.220000 ;
        RECT 50.890000 15.460000 51.090000 15.660000 ;
        RECT 50.890000 15.900000 51.090000 16.100000 ;
        RECT 50.890000 16.340000 51.090000 16.540000 ;
        RECT 50.890000 16.780000 51.090000 16.980000 ;
        RECT 50.890000 17.220000 51.090000 17.420000 ;
        RECT 50.890000 17.660000 51.090000 17.860000 ;
        RECT 50.890000 18.100000 51.090000 18.300000 ;
        RECT 51.300000 15.020000 51.500000 15.220000 ;
        RECT 51.300000 15.460000 51.500000 15.660000 ;
        RECT 51.300000 15.900000 51.500000 16.100000 ;
        RECT 51.300000 16.340000 51.500000 16.540000 ;
        RECT 51.300000 16.780000 51.500000 16.980000 ;
        RECT 51.300000 17.220000 51.500000 17.420000 ;
        RECT 51.300000 17.660000 51.500000 17.860000 ;
        RECT 51.300000 18.100000 51.500000 18.300000 ;
        RECT 51.710000 15.020000 51.910000 15.220000 ;
        RECT 51.710000 15.460000 51.910000 15.660000 ;
        RECT 51.710000 15.900000 51.910000 16.100000 ;
        RECT 51.710000 16.340000 51.910000 16.540000 ;
        RECT 51.710000 16.780000 51.910000 16.980000 ;
        RECT 51.710000 17.220000 51.910000 17.420000 ;
        RECT 51.710000 17.660000 51.910000 17.860000 ;
        RECT 51.710000 18.100000 51.910000 18.300000 ;
        RECT 52.120000 15.020000 52.320000 15.220000 ;
        RECT 52.120000 15.460000 52.320000 15.660000 ;
        RECT 52.120000 15.900000 52.320000 16.100000 ;
        RECT 52.120000 16.340000 52.320000 16.540000 ;
        RECT 52.120000 16.780000 52.320000 16.980000 ;
        RECT 52.120000 17.220000 52.320000 17.420000 ;
        RECT 52.120000 17.660000 52.320000 17.860000 ;
        RECT 52.120000 18.100000 52.320000 18.300000 ;
        RECT 52.530000 15.020000 52.730000 15.220000 ;
        RECT 52.530000 15.460000 52.730000 15.660000 ;
        RECT 52.530000 15.900000 52.730000 16.100000 ;
        RECT 52.530000 16.340000 52.730000 16.540000 ;
        RECT 52.530000 16.780000 52.730000 16.980000 ;
        RECT 52.530000 17.220000 52.730000 17.420000 ;
        RECT 52.530000 17.660000 52.730000 17.860000 ;
        RECT 52.530000 18.100000 52.730000 18.300000 ;
        RECT 52.940000 15.020000 53.140000 15.220000 ;
        RECT 52.940000 15.460000 53.140000 15.660000 ;
        RECT 52.940000 15.900000 53.140000 16.100000 ;
        RECT 52.940000 16.340000 53.140000 16.540000 ;
        RECT 52.940000 16.780000 53.140000 16.980000 ;
        RECT 52.940000 17.220000 53.140000 17.420000 ;
        RECT 52.940000 17.660000 53.140000 17.860000 ;
        RECT 52.940000 18.100000 53.140000 18.300000 ;
        RECT 53.345000 15.020000 53.545000 15.220000 ;
        RECT 53.345000 15.460000 53.545000 15.660000 ;
        RECT 53.345000 15.900000 53.545000 16.100000 ;
        RECT 53.345000 16.340000 53.545000 16.540000 ;
        RECT 53.345000 16.780000 53.545000 16.980000 ;
        RECT 53.345000 17.220000 53.545000 17.420000 ;
        RECT 53.345000 17.660000 53.545000 17.860000 ;
        RECT 53.345000 18.100000 53.545000 18.300000 ;
        RECT 53.750000 15.020000 53.950000 15.220000 ;
        RECT 53.750000 15.460000 53.950000 15.660000 ;
        RECT 53.750000 15.900000 53.950000 16.100000 ;
        RECT 53.750000 16.340000 53.950000 16.540000 ;
        RECT 53.750000 16.780000 53.950000 16.980000 ;
        RECT 53.750000 17.220000 53.950000 17.420000 ;
        RECT 53.750000 17.660000 53.950000 17.860000 ;
        RECT 53.750000 18.100000 53.950000 18.300000 ;
        RECT 54.155000 15.020000 54.355000 15.220000 ;
        RECT 54.155000 15.460000 54.355000 15.660000 ;
        RECT 54.155000 15.900000 54.355000 16.100000 ;
        RECT 54.155000 16.340000 54.355000 16.540000 ;
        RECT 54.155000 16.780000 54.355000 16.980000 ;
        RECT 54.155000 17.220000 54.355000 17.420000 ;
        RECT 54.155000 17.660000 54.355000 17.860000 ;
        RECT 54.155000 18.100000 54.355000 18.300000 ;
        RECT 54.560000 15.020000 54.760000 15.220000 ;
        RECT 54.560000 15.460000 54.760000 15.660000 ;
        RECT 54.560000 15.900000 54.760000 16.100000 ;
        RECT 54.560000 16.340000 54.760000 16.540000 ;
        RECT 54.560000 16.780000 54.760000 16.980000 ;
        RECT 54.560000 17.220000 54.760000 17.420000 ;
        RECT 54.560000 17.660000 54.760000 17.860000 ;
        RECT 54.560000 18.100000 54.760000 18.300000 ;
        RECT 54.965000 15.020000 55.165000 15.220000 ;
        RECT 54.965000 15.460000 55.165000 15.660000 ;
        RECT 54.965000 15.900000 55.165000 16.100000 ;
        RECT 54.965000 16.340000 55.165000 16.540000 ;
        RECT 54.965000 16.780000 55.165000 16.980000 ;
        RECT 54.965000 17.220000 55.165000 17.420000 ;
        RECT 54.965000 17.660000 55.165000 17.860000 ;
        RECT 54.965000 18.100000 55.165000 18.300000 ;
        RECT 55.370000 15.020000 55.570000 15.220000 ;
        RECT 55.370000 15.460000 55.570000 15.660000 ;
        RECT 55.370000 15.900000 55.570000 16.100000 ;
        RECT 55.370000 16.340000 55.570000 16.540000 ;
        RECT 55.370000 16.780000 55.570000 16.980000 ;
        RECT 55.370000 17.220000 55.570000 17.420000 ;
        RECT 55.370000 17.660000 55.570000 17.860000 ;
        RECT 55.370000 18.100000 55.570000 18.300000 ;
        RECT 55.775000 15.020000 55.975000 15.220000 ;
        RECT 55.775000 15.460000 55.975000 15.660000 ;
        RECT 55.775000 15.900000 55.975000 16.100000 ;
        RECT 55.775000 16.340000 55.975000 16.540000 ;
        RECT 55.775000 16.780000 55.975000 16.980000 ;
        RECT 55.775000 17.220000 55.975000 17.420000 ;
        RECT 55.775000 17.660000 55.975000 17.860000 ;
        RECT 55.775000 18.100000 55.975000 18.300000 ;
        RECT 56.180000 15.020000 56.380000 15.220000 ;
        RECT 56.180000 15.460000 56.380000 15.660000 ;
        RECT 56.180000 15.900000 56.380000 16.100000 ;
        RECT 56.180000 16.340000 56.380000 16.540000 ;
        RECT 56.180000 16.780000 56.380000 16.980000 ;
        RECT 56.180000 17.220000 56.380000 17.420000 ;
        RECT 56.180000 17.660000 56.380000 17.860000 ;
        RECT 56.180000 18.100000 56.380000 18.300000 ;
        RECT 56.585000 15.020000 56.785000 15.220000 ;
        RECT 56.585000 15.460000 56.785000 15.660000 ;
        RECT 56.585000 15.900000 56.785000 16.100000 ;
        RECT 56.585000 16.340000 56.785000 16.540000 ;
        RECT 56.585000 16.780000 56.785000 16.980000 ;
        RECT 56.585000 17.220000 56.785000 17.420000 ;
        RECT 56.585000 17.660000 56.785000 17.860000 ;
        RECT 56.585000 18.100000 56.785000 18.300000 ;
        RECT 56.990000 15.020000 57.190000 15.220000 ;
        RECT 56.990000 15.460000 57.190000 15.660000 ;
        RECT 56.990000 15.900000 57.190000 16.100000 ;
        RECT 56.990000 16.340000 57.190000 16.540000 ;
        RECT 56.990000 16.780000 57.190000 16.980000 ;
        RECT 56.990000 17.220000 57.190000 17.420000 ;
        RECT 56.990000 17.660000 57.190000 17.860000 ;
        RECT 56.990000 18.100000 57.190000 18.300000 ;
        RECT 57.395000 15.020000 57.595000 15.220000 ;
        RECT 57.395000 15.460000 57.595000 15.660000 ;
        RECT 57.395000 15.900000 57.595000 16.100000 ;
        RECT 57.395000 16.340000 57.595000 16.540000 ;
        RECT 57.395000 16.780000 57.595000 16.980000 ;
        RECT 57.395000 17.220000 57.595000 17.420000 ;
        RECT 57.395000 17.660000 57.595000 17.860000 ;
        RECT 57.395000 18.100000 57.595000 18.300000 ;
        RECT 57.800000 15.020000 58.000000 15.220000 ;
        RECT 57.800000 15.460000 58.000000 15.660000 ;
        RECT 57.800000 15.900000 58.000000 16.100000 ;
        RECT 57.800000 16.340000 58.000000 16.540000 ;
        RECT 57.800000 16.780000 58.000000 16.980000 ;
        RECT 57.800000 17.220000 58.000000 17.420000 ;
        RECT 57.800000 17.660000 58.000000 17.860000 ;
        RECT 57.800000 18.100000 58.000000 18.300000 ;
        RECT 58.205000 15.020000 58.405000 15.220000 ;
        RECT 58.205000 15.460000 58.405000 15.660000 ;
        RECT 58.205000 15.900000 58.405000 16.100000 ;
        RECT 58.205000 16.340000 58.405000 16.540000 ;
        RECT 58.205000 16.780000 58.405000 16.980000 ;
        RECT 58.205000 17.220000 58.405000 17.420000 ;
        RECT 58.205000 17.660000 58.405000 17.860000 ;
        RECT 58.205000 18.100000 58.405000 18.300000 ;
        RECT 58.610000 15.020000 58.810000 15.220000 ;
        RECT 58.610000 15.460000 58.810000 15.660000 ;
        RECT 58.610000 15.900000 58.810000 16.100000 ;
        RECT 58.610000 16.340000 58.810000 16.540000 ;
        RECT 58.610000 16.780000 58.810000 16.980000 ;
        RECT 58.610000 17.220000 58.810000 17.420000 ;
        RECT 58.610000 17.660000 58.810000 17.860000 ;
        RECT 58.610000 18.100000 58.810000 18.300000 ;
        RECT 59.015000 15.020000 59.215000 15.220000 ;
        RECT 59.015000 15.460000 59.215000 15.660000 ;
        RECT 59.015000 15.900000 59.215000 16.100000 ;
        RECT 59.015000 16.340000 59.215000 16.540000 ;
        RECT 59.015000 16.780000 59.215000 16.980000 ;
        RECT 59.015000 17.220000 59.215000 17.420000 ;
        RECT 59.015000 17.660000 59.215000 17.860000 ;
        RECT 59.015000 18.100000 59.215000 18.300000 ;
        RECT 59.420000 15.020000 59.620000 15.220000 ;
        RECT 59.420000 15.460000 59.620000 15.660000 ;
        RECT 59.420000 15.900000 59.620000 16.100000 ;
        RECT 59.420000 16.340000 59.620000 16.540000 ;
        RECT 59.420000 16.780000 59.620000 16.980000 ;
        RECT 59.420000 17.220000 59.620000 17.420000 ;
        RECT 59.420000 17.660000 59.620000 17.860000 ;
        RECT 59.420000 18.100000 59.620000 18.300000 ;
        RECT 59.825000 15.020000 60.025000 15.220000 ;
        RECT 59.825000 15.460000 60.025000 15.660000 ;
        RECT 59.825000 15.900000 60.025000 16.100000 ;
        RECT 59.825000 16.340000 60.025000 16.540000 ;
        RECT 59.825000 16.780000 60.025000 16.980000 ;
        RECT 59.825000 17.220000 60.025000 17.420000 ;
        RECT 59.825000 17.660000 60.025000 17.860000 ;
        RECT 59.825000 18.100000 60.025000 18.300000 ;
        RECT 60.230000 15.020000 60.430000 15.220000 ;
        RECT 60.230000 15.460000 60.430000 15.660000 ;
        RECT 60.230000 15.900000 60.430000 16.100000 ;
        RECT 60.230000 16.340000 60.430000 16.540000 ;
        RECT 60.230000 16.780000 60.430000 16.980000 ;
        RECT 60.230000 17.220000 60.430000 17.420000 ;
        RECT 60.230000 17.660000 60.430000 17.860000 ;
        RECT 60.230000 18.100000 60.430000 18.300000 ;
        RECT 60.635000 15.020000 60.835000 15.220000 ;
        RECT 60.635000 15.460000 60.835000 15.660000 ;
        RECT 60.635000 15.900000 60.835000 16.100000 ;
        RECT 60.635000 16.340000 60.835000 16.540000 ;
        RECT 60.635000 16.780000 60.835000 16.980000 ;
        RECT 60.635000 17.220000 60.835000 17.420000 ;
        RECT 60.635000 17.660000 60.835000 17.860000 ;
        RECT 60.635000 18.100000 60.835000 18.300000 ;
        RECT 61.040000 15.020000 61.240000 15.220000 ;
        RECT 61.040000 15.460000 61.240000 15.660000 ;
        RECT 61.040000 15.900000 61.240000 16.100000 ;
        RECT 61.040000 16.340000 61.240000 16.540000 ;
        RECT 61.040000 16.780000 61.240000 16.980000 ;
        RECT 61.040000 17.220000 61.240000 17.420000 ;
        RECT 61.040000 17.660000 61.240000 17.860000 ;
        RECT 61.040000 18.100000 61.240000 18.300000 ;
        RECT 61.445000 15.020000 61.645000 15.220000 ;
        RECT 61.445000 15.460000 61.645000 15.660000 ;
        RECT 61.445000 15.900000 61.645000 16.100000 ;
        RECT 61.445000 16.340000 61.645000 16.540000 ;
        RECT 61.445000 16.780000 61.645000 16.980000 ;
        RECT 61.445000 17.220000 61.645000 17.420000 ;
        RECT 61.445000 17.660000 61.645000 17.860000 ;
        RECT 61.445000 18.100000 61.645000 18.300000 ;
        RECT 61.850000 15.020000 62.050000 15.220000 ;
        RECT 61.850000 15.460000 62.050000 15.660000 ;
        RECT 61.850000 15.900000 62.050000 16.100000 ;
        RECT 61.850000 16.340000 62.050000 16.540000 ;
        RECT 61.850000 16.780000 62.050000 16.980000 ;
        RECT 61.850000 17.220000 62.050000 17.420000 ;
        RECT 61.850000 17.660000 62.050000 17.860000 ;
        RECT 61.850000 18.100000 62.050000 18.300000 ;
        RECT 62.255000 15.020000 62.455000 15.220000 ;
        RECT 62.255000 15.460000 62.455000 15.660000 ;
        RECT 62.255000 15.900000 62.455000 16.100000 ;
        RECT 62.255000 16.340000 62.455000 16.540000 ;
        RECT 62.255000 16.780000 62.455000 16.980000 ;
        RECT 62.255000 17.220000 62.455000 17.420000 ;
        RECT 62.255000 17.660000 62.455000 17.860000 ;
        RECT 62.255000 18.100000 62.455000 18.300000 ;
        RECT 62.660000 15.020000 62.860000 15.220000 ;
        RECT 62.660000 15.460000 62.860000 15.660000 ;
        RECT 62.660000 15.900000 62.860000 16.100000 ;
        RECT 62.660000 16.340000 62.860000 16.540000 ;
        RECT 62.660000 16.780000 62.860000 16.980000 ;
        RECT 62.660000 17.220000 62.860000 17.420000 ;
        RECT 62.660000 17.660000 62.860000 17.860000 ;
        RECT 62.660000 18.100000 62.860000 18.300000 ;
        RECT 63.065000 15.020000 63.265000 15.220000 ;
        RECT 63.065000 15.460000 63.265000 15.660000 ;
        RECT 63.065000 15.900000 63.265000 16.100000 ;
        RECT 63.065000 16.340000 63.265000 16.540000 ;
        RECT 63.065000 16.780000 63.265000 16.980000 ;
        RECT 63.065000 17.220000 63.265000 17.420000 ;
        RECT 63.065000 17.660000 63.265000 17.860000 ;
        RECT 63.065000 18.100000 63.265000 18.300000 ;
        RECT 63.470000 15.020000 63.670000 15.220000 ;
        RECT 63.470000 15.460000 63.670000 15.660000 ;
        RECT 63.470000 15.900000 63.670000 16.100000 ;
        RECT 63.470000 16.340000 63.670000 16.540000 ;
        RECT 63.470000 16.780000 63.670000 16.980000 ;
        RECT 63.470000 17.220000 63.670000 17.420000 ;
        RECT 63.470000 17.660000 63.670000 17.860000 ;
        RECT 63.470000 18.100000 63.670000 18.300000 ;
        RECT 63.875000 15.020000 64.075000 15.220000 ;
        RECT 63.875000 15.460000 64.075000 15.660000 ;
        RECT 63.875000 15.900000 64.075000 16.100000 ;
        RECT 63.875000 16.340000 64.075000 16.540000 ;
        RECT 63.875000 16.780000 64.075000 16.980000 ;
        RECT 63.875000 17.220000 64.075000 17.420000 ;
        RECT 63.875000 17.660000 64.075000 17.860000 ;
        RECT 63.875000 18.100000 64.075000 18.300000 ;
        RECT 64.280000 15.020000 64.480000 15.220000 ;
        RECT 64.280000 15.460000 64.480000 15.660000 ;
        RECT 64.280000 15.900000 64.480000 16.100000 ;
        RECT 64.280000 16.340000 64.480000 16.540000 ;
        RECT 64.280000 16.780000 64.480000 16.980000 ;
        RECT 64.280000 17.220000 64.480000 17.420000 ;
        RECT 64.280000 17.660000 64.480000 17.860000 ;
        RECT 64.280000 18.100000 64.480000 18.300000 ;
        RECT 64.685000 15.020000 64.885000 15.220000 ;
        RECT 64.685000 15.460000 64.885000 15.660000 ;
        RECT 64.685000 15.900000 64.885000 16.100000 ;
        RECT 64.685000 16.340000 64.885000 16.540000 ;
        RECT 64.685000 16.780000 64.885000 16.980000 ;
        RECT 64.685000 17.220000 64.885000 17.420000 ;
        RECT 64.685000 17.660000 64.885000 17.860000 ;
        RECT 64.685000 18.100000 64.885000 18.300000 ;
        RECT 65.090000 15.020000 65.290000 15.220000 ;
        RECT 65.090000 15.460000 65.290000 15.660000 ;
        RECT 65.090000 15.900000 65.290000 16.100000 ;
        RECT 65.090000 16.340000 65.290000 16.540000 ;
        RECT 65.090000 16.780000 65.290000 16.980000 ;
        RECT 65.090000 17.220000 65.290000 17.420000 ;
        RECT 65.090000 17.660000 65.290000 17.860000 ;
        RECT 65.090000 18.100000 65.290000 18.300000 ;
        RECT 65.495000 15.020000 65.695000 15.220000 ;
        RECT 65.495000 15.460000 65.695000 15.660000 ;
        RECT 65.495000 15.900000 65.695000 16.100000 ;
        RECT 65.495000 16.340000 65.695000 16.540000 ;
        RECT 65.495000 16.780000 65.695000 16.980000 ;
        RECT 65.495000 17.220000 65.695000 17.420000 ;
        RECT 65.495000 17.660000 65.695000 17.860000 ;
        RECT 65.495000 18.100000 65.695000 18.300000 ;
        RECT 65.900000 15.020000 66.100000 15.220000 ;
        RECT 65.900000 15.460000 66.100000 15.660000 ;
        RECT 65.900000 15.900000 66.100000 16.100000 ;
        RECT 65.900000 16.340000 66.100000 16.540000 ;
        RECT 65.900000 16.780000 66.100000 16.980000 ;
        RECT 65.900000 17.220000 66.100000 17.420000 ;
        RECT 65.900000 17.660000 66.100000 17.860000 ;
        RECT 65.900000 18.100000 66.100000 18.300000 ;
        RECT 66.305000 15.020000 66.505000 15.220000 ;
        RECT 66.305000 15.460000 66.505000 15.660000 ;
        RECT 66.305000 15.900000 66.505000 16.100000 ;
        RECT 66.305000 16.340000 66.505000 16.540000 ;
        RECT 66.305000 16.780000 66.505000 16.980000 ;
        RECT 66.305000 17.220000 66.505000 17.420000 ;
        RECT 66.305000 17.660000 66.505000 17.860000 ;
        RECT 66.305000 18.100000 66.505000 18.300000 ;
        RECT 66.710000 15.020000 66.910000 15.220000 ;
        RECT 66.710000 15.460000 66.910000 15.660000 ;
        RECT 66.710000 15.900000 66.910000 16.100000 ;
        RECT 66.710000 16.340000 66.910000 16.540000 ;
        RECT 66.710000 16.780000 66.910000 16.980000 ;
        RECT 66.710000 17.220000 66.910000 17.420000 ;
        RECT 66.710000 17.660000 66.910000 17.860000 ;
        RECT 66.710000 18.100000 66.910000 18.300000 ;
        RECT 67.115000 15.020000 67.315000 15.220000 ;
        RECT 67.115000 15.460000 67.315000 15.660000 ;
        RECT 67.115000 15.900000 67.315000 16.100000 ;
        RECT 67.115000 16.340000 67.315000 16.540000 ;
        RECT 67.115000 16.780000 67.315000 16.980000 ;
        RECT 67.115000 17.220000 67.315000 17.420000 ;
        RECT 67.115000 17.660000 67.315000 17.860000 ;
        RECT 67.115000 18.100000 67.315000 18.300000 ;
        RECT 67.520000 15.020000 67.720000 15.220000 ;
        RECT 67.520000 15.460000 67.720000 15.660000 ;
        RECT 67.520000 15.900000 67.720000 16.100000 ;
        RECT 67.520000 16.340000 67.720000 16.540000 ;
        RECT 67.520000 16.780000 67.720000 16.980000 ;
        RECT 67.520000 17.220000 67.720000 17.420000 ;
        RECT 67.520000 17.660000 67.720000 17.860000 ;
        RECT 67.520000 18.100000 67.720000 18.300000 ;
        RECT 67.925000 15.020000 68.125000 15.220000 ;
        RECT 67.925000 15.460000 68.125000 15.660000 ;
        RECT 67.925000 15.900000 68.125000 16.100000 ;
        RECT 67.925000 16.340000 68.125000 16.540000 ;
        RECT 67.925000 16.780000 68.125000 16.980000 ;
        RECT 67.925000 17.220000 68.125000 17.420000 ;
        RECT 67.925000 17.660000 68.125000 17.860000 ;
        RECT 67.925000 18.100000 68.125000 18.300000 ;
        RECT 68.330000 15.020000 68.530000 15.220000 ;
        RECT 68.330000 15.460000 68.530000 15.660000 ;
        RECT 68.330000 15.900000 68.530000 16.100000 ;
        RECT 68.330000 16.340000 68.530000 16.540000 ;
        RECT 68.330000 16.780000 68.530000 16.980000 ;
        RECT 68.330000 17.220000 68.530000 17.420000 ;
        RECT 68.330000 17.660000 68.530000 17.860000 ;
        RECT 68.330000 18.100000 68.530000 18.300000 ;
        RECT 68.735000 15.020000 68.935000 15.220000 ;
        RECT 68.735000 15.460000 68.935000 15.660000 ;
        RECT 68.735000 15.900000 68.935000 16.100000 ;
        RECT 68.735000 16.340000 68.935000 16.540000 ;
        RECT 68.735000 16.780000 68.935000 16.980000 ;
        RECT 68.735000 17.220000 68.935000 17.420000 ;
        RECT 68.735000 17.660000 68.935000 17.860000 ;
        RECT 68.735000 18.100000 68.935000 18.300000 ;
        RECT 69.140000 15.020000 69.340000 15.220000 ;
        RECT 69.140000 15.460000 69.340000 15.660000 ;
        RECT 69.140000 15.900000 69.340000 16.100000 ;
        RECT 69.140000 16.340000 69.340000 16.540000 ;
        RECT 69.140000 16.780000 69.340000 16.980000 ;
        RECT 69.140000 17.220000 69.340000 17.420000 ;
        RECT 69.140000 17.660000 69.340000 17.860000 ;
        RECT 69.140000 18.100000 69.340000 18.300000 ;
        RECT 69.545000 15.020000 69.745000 15.220000 ;
        RECT 69.545000 15.460000 69.745000 15.660000 ;
        RECT 69.545000 15.900000 69.745000 16.100000 ;
        RECT 69.545000 16.340000 69.745000 16.540000 ;
        RECT 69.545000 16.780000 69.745000 16.980000 ;
        RECT 69.545000 17.220000 69.745000 17.420000 ;
        RECT 69.545000 17.660000 69.745000 17.860000 ;
        RECT 69.545000 18.100000 69.745000 18.300000 ;
        RECT 69.950000 15.020000 70.150000 15.220000 ;
        RECT 69.950000 15.460000 70.150000 15.660000 ;
        RECT 69.950000 15.900000 70.150000 16.100000 ;
        RECT 69.950000 16.340000 70.150000 16.540000 ;
        RECT 69.950000 16.780000 70.150000 16.980000 ;
        RECT 69.950000 17.220000 70.150000 17.420000 ;
        RECT 69.950000 17.660000 70.150000 17.860000 ;
        RECT 69.950000 18.100000 70.150000 18.300000 ;
        RECT 70.355000 15.020000 70.555000 15.220000 ;
        RECT 70.355000 15.460000 70.555000 15.660000 ;
        RECT 70.355000 15.900000 70.555000 16.100000 ;
        RECT 70.355000 16.340000 70.555000 16.540000 ;
        RECT 70.355000 16.780000 70.555000 16.980000 ;
        RECT 70.355000 17.220000 70.555000 17.420000 ;
        RECT 70.355000 17.660000 70.555000 17.860000 ;
        RECT 70.355000 18.100000 70.555000 18.300000 ;
        RECT 70.760000 15.020000 70.960000 15.220000 ;
        RECT 70.760000 15.460000 70.960000 15.660000 ;
        RECT 70.760000 15.900000 70.960000 16.100000 ;
        RECT 70.760000 16.340000 70.960000 16.540000 ;
        RECT 70.760000 16.780000 70.960000 16.980000 ;
        RECT 70.760000 17.220000 70.960000 17.420000 ;
        RECT 70.760000 17.660000 70.960000 17.860000 ;
        RECT 70.760000 18.100000 70.960000 18.300000 ;
        RECT 71.165000 15.020000 71.365000 15.220000 ;
        RECT 71.165000 15.460000 71.365000 15.660000 ;
        RECT 71.165000 15.900000 71.365000 16.100000 ;
        RECT 71.165000 16.340000 71.365000 16.540000 ;
        RECT 71.165000 16.780000 71.365000 16.980000 ;
        RECT 71.165000 17.220000 71.365000 17.420000 ;
        RECT 71.165000 17.660000 71.365000 17.860000 ;
        RECT 71.165000 18.100000 71.365000 18.300000 ;
        RECT 71.570000 15.020000 71.770000 15.220000 ;
        RECT 71.570000 15.460000 71.770000 15.660000 ;
        RECT 71.570000 15.900000 71.770000 16.100000 ;
        RECT 71.570000 16.340000 71.770000 16.540000 ;
        RECT 71.570000 16.780000 71.770000 16.980000 ;
        RECT 71.570000 17.220000 71.770000 17.420000 ;
        RECT 71.570000 17.660000 71.770000 17.860000 ;
        RECT 71.570000 18.100000 71.770000 18.300000 ;
        RECT 71.975000 15.020000 72.175000 15.220000 ;
        RECT 71.975000 15.460000 72.175000 15.660000 ;
        RECT 71.975000 15.900000 72.175000 16.100000 ;
        RECT 71.975000 16.340000 72.175000 16.540000 ;
        RECT 71.975000 16.780000 72.175000 16.980000 ;
        RECT 71.975000 17.220000 72.175000 17.420000 ;
        RECT 71.975000 17.660000 72.175000 17.860000 ;
        RECT 71.975000 18.100000 72.175000 18.300000 ;
        RECT 72.380000 15.020000 72.580000 15.220000 ;
        RECT 72.380000 15.460000 72.580000 15.660000 ;
        RECT 72.380000 15.900000 72.580000 16.100000 ;
        RECT 72.380000 16.340000 72.580000 16.540000 ;
        RECT 72.380000 16.780000 72.580000 16.980000 ;
        RECT 72.380000 17.220000 72.580000 17.420000 ;
        RECT 72.380000 17.660000 72.580000 17.860000 ;
        RECT 72.380000 18.100000 72.580000 18.300000 ;
        RECT 72.785000 15.020000 72.985000 15.220000 ;
        RECT 72.785000 15.460000 72.985000 15.660000 ;
        RECT 72.785000 15.900000 72.985000 16.100000 ;
        RECT 72.785000 16.340000 72.985000 16.540000 ;
        RECT 72.785000 16.780000 72.985000 16.980000 ;
        RECT 72.785000 17.220000 72.985000 17.420000 ;
        RECT 72.785000 17.660000 72.985000 17.860000 ;
        RECT 72.785000 18.100000 72.985000 18.300000 ;
        RECT 73.190000 15.020000 73.390000 15.220000 ;
        RECT 73.190000 15.460000 73.390000 15.660000 ;
        RECT 73.190000 15.900000 73.390000 16.100000 ;
        RECT 73.190000 16.340000 73.390000 16.540000 ;
        RECT 73.190000 16.780000 73.390000 16.980000 ;
        RECT 73.190000 17.220000 73.390000 17.420000 ;
        RECT 73.190000 17.660000 73.390000 17.860000 ;
        RECT 73.190000 18.100000 73.390000 18.300000 ;
        RECT 73.595000 15.020000 73.795000 15.220000 ;
        RECT 73.595000 15.460000 73.795000 15.660000 ;
        RECT 73.595000 15.900000 73.795000 16.100000 ;
        RECT 73.595000 16.340000 73.795000 16.540000 ;
        RECT 73.595000 16.780000 73.795000 16.980000 ;
        RECT 73.595000 17.220000 73.795000 17.420000 ;
        RECT 73.595000 17.660000 73.795000 17.860000 ;
        RECT 73.595000 18.100000 73.795000 18.300000 ;
        RECT 74.000000 15.020000 74.200000 15.220000 ;
        RECT 74.000000 15.460000 74.200000 15.660000 ;
        RECT 74.000000 15.900000 74.200000 16.100000 ;
        RECT 74.000000 16.340000 74.200000 16.540000 ;
        RECT 74.000000 16.780000 74.200000 16.980000 ;
        RECT 74.000000 17.220000 74.200000 17.420000 ;
        RECT 74.000000 17.660000 74.200000 17.860000 ;
        RECT 74.000000 18.100000 74.200000 18.300000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 19.785000 1.270000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 70.035000 1.270000 95.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 19.785000 75.000000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 70.035000 75.000000 95.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 19.885000 1.270000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 70.035000 1.270000 94.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 19.885000 75.000000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 70.035000 75.000000 94.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 64.085000 1.270000 68.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 64.085000 75.000000 68.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 64.185000 1.270000 68.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 64.185000 75.000000 68.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 36.735000 1.270000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 47.735000 1.270000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 51.645000 1.270000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 56.405000 1.270000 56.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 36.735000 75.000000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 47.735000 75.000000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.645000 75.000000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 56.405000 75.000000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 36.840000 1.270000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 47.735000 1.270000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 36.840000 75.000000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 47.735000 75.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 41.585000 1.270000 46.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 41.585000 75.000000 46.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 41.685000 1.270000 46.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 41.685000 75.000000 46.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 25.835000 1.270000 30.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 25.835000 75.000000 30.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 25.935000 1.270000 30.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 25.935000 75.000000 30.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 58.235000 1.270000 62.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 58.235000 75.000000 62.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 58.335000 1.270000 62.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 58.335000 75.000000 62.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 31.885000 1.270000 35.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 31.885000 75.000000 35.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 31.985000 1.270000 35.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 31.985000 75.000000 35.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met1 ;
      RECT 0.000000 0.000000 75.000000 200.000000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 75.000000 200.000000 ;
    LAYER met3 ;
      RECT  0.000000  0.000000 75.000000  14.540000 ;
      RECT  0.000000 18.780000 75.000000 200.000000 ;
      RECT 24.795000 14.540000 49.990000  18.780000 ;
      RECT 74.690000 14.540000 75.000000  18.780000 ;
    LAYER met4 ;
      RECT  0.000000   0.000000  1.670000   1.635000 ;
      RECT  0.000000   7.885000  1.670000   8.485000 ;
      RECT  0.000000  13.935000  1.670000  14.535000 ;
      RECT  0.000000  18.785000  1.670000  19.385000 ;
      RECT  0.000000  24.835000  1.670000  25.435000 ;
      RECT  0.000000  30.885000  1.670000  31.485000 ;
      RECT  0.000000  35.735000  1.670000  36.335000 ;
      RECT  0.000000  40.585000  1.670000  41.185000 ;
      RECT  0.000000  46.635000  1.670000  47.335000 ;
      RECT  0.000000  57.135000  1.670000  57.835000 ;
      RECT  0.000000  63.085000  1.670000  63.685000 ;
      RECT  0.000000  68.935000  1.670000  69.635000 ;
      RECT  0.000000  95.400000 75.000000 175.385000 ;
      RECT  1.670000   0.000000 73.330000  14.535000 ;
      RECT  1.670000  18.785000 73.330000  95.400000 ;
      RECT  1.670000 175.385000 73.330000 200.000000 ;
      RECT 24.770000  14.535000 50.015000  18.785000 ;
      RECT 73.330000   0.000000 75.000000   1.635000 ;
      RECT 73.330000   7.885000 75.000000   8.485000 ;
      RECT 73.330000  13.935000 75.000000  14.535000 ;
      RECT 73.330000  18.785000 75.000000  19.385000 ;
      RECT 73.330000  24.835000 75.000000  25.435000 ;
      RECT 73.330000  30.885000 75.000000  31.485000 ;
      RECT 73.330000  35.735000 75.000000  36.335000 ;
      RECT 73.330000  40.585000 75.000000  41.185000 ;
      RECT 73.330000  46.635000 75.000000  47.335000 ;
      RECT 73.330000  57.135000 75.000000  57.835000 ;
      RECT 73.330000  63.085000 75.000000  63.685000 ;
      RECT 73.330000  68.935000 75.000000  69.635000 ;
    LAYER met5 ;
      RECT 0.000000   0.000000 75.000000   1.335000 ;
      RECT 0.000000  95.785000 75.000000 174.985000 ;
      RECT 1.765000  14.235000 73.235000  19.085000 ;
      RECT 2.070000   1.335000 72.930000  14.235000 ;
      RECT 2.070000  19.085000 72.930000  95.785000 ;
      RECT 2.070000 174.985000 72.930000 200.000000 ;
  END
END sky130_fd_io__overlay_vdda_hvc
END LIBRARY
