VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO HEADER
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HEADER 0 0 ;
  SIZE 12.42 BY 2.72 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.045 0.71 9.81 0.88 ;
        RECT 8.605 0.71 8.775 1.34 ;
        RECT 7.045 0.71 7.215 1.34 ;
    END
  END VIN
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 11.585 0.265 11.875 0.81 ;
        RECT 0.545 0.265 0.835 0.81 ;
    END
  END VNB
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 -0.24 12.42 0.24 ;
      LAYER li1 ;
        RECT 0 -0.085 12.42 0.085 ;
        RECT 5.395 1.89 10.15 2.06 ;
        RECT 9.98 -0.085 10.15 2.06 ;
        RECT 5.395 1.51 5.565 2.06 ;
      LAYER mcon ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 12.42 2.96 ;
      LAYER li1 ;
        RECT 0 2.635 12.42 2.805 ;
        RECT 4.92 1.05 5.09 2.805 ;
        RECT 3.36 1.51 5.09 1.68 ;
        RECT 3.36 1.05 3.53 2.805 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 6.265 1.51 9.555 1.68 ;
      RECT 9.385 1.05 9.555 1.68 ;
      RECT 7.825 1.05 7.995 1.68 ;
      RECT 6.265 0.71 6.435 1.68 ;
      RECT 5.7 0.71 5.87 1.34 ;
      RECT 4.14 0.71 4.31 1.34 ;
      RECT 2.58 0.71 2.75 1.34 ;
      RECT 2.58 0.71 6.435 0.88 ;
      RECT 11.585 1.47 11.875 2.455 ;
      RECT 0.545 1.47 0.835 2.455 ;
  END
END HEADER

END LIBRARY
