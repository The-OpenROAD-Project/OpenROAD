module empty ();
endmodule
