module gcd (
	resp_val,
	resp_rdy,
	resp_msg,
	reset,
	req_val,
	req_rdy,
	req_msg,
	clk);
   output resp_val;
   input resp_rdy;
   output [15:0] resp_msg;
   input reset;
   input req_val;
   output req_rdy;
   input [31:0] req_msg;
   input clk;

   // Internal wires
   wire resp_val;
   wire resp_rdy;
   wire [15:0] resp_msg;
   wire reset;
   wire req_val;
   wire req_rdy;
   wire [31:0] req_msg;
   wire net9;
   wire net8;
   wire net7;
   wire net6;
   wire net53;
   wire net52;
   wire net51;
   wire net50;
   wire net5;
   wire net49;
   wire net48;
   wire net47;
   wire net46;
   wire net45;
   wire net44;
   wire net43;
   wire net42;
   wire net41;
   wire net40;
   wire net4;
   wire net39;
   wire net38;
   wire net37;
   wire net36;
   wire net35;
   wire net34;
   wire net33;
   wire net32;
   wire net31;
   wire net30;
   wire net3;
   wire net29;
   wire net28;
   wire net27;
   wire net26;
   wire net25;
   wire net24;
   wire net23;
   wire net22;
   wire net21;
   wire net20;
   wire net2;
   wire net19;
   wire net18;
   wire net17;
   wire net16;
   wire net15;
   wire net14;
   wire net13;
   wire net12;
   wire net11;
   wire net10;
   wire net1;
   wire \dpath.a_lt_b$in1\[9\] ;
   wire \dpath.a_lt_b$in1\[8\] ;
   wire \dpath.a_lt_b$in1\[7\] ;
   wire \dpath.a_lt_b$in1\[6\] ;
   wire \dpath.a_lt_b$in1\[5\] ;
   wire \dpath.a_lt_b$in1\[4\] ;
   wire \dpath.a_lt_b$in1\[3\] ;
   wire \dpath.a_lt_b$in1\[2\] ;
   wire \dpath.a_lt_b$in1\[1\] ;
   wire \dpath.a_lt_b$in1\[15\] ;
   wire \dpath.a_lt_b$in1\[14\] ;
   wire \dpath.a_lt_b$in1\[13\] ;
   wire \dpath.a_lt_b$in1\[12\] ;
   wire \dpath.a_lt_b$in1\[11\] ;
   wire \dpath.a_lt_b$in1\[10\] ;
   wire \dpath.a_lt_b$in1\[0\] ;
   wire \dpath.a_lt_b$in0\[9\] ;
   wire \dpath.a_lt_b$in0\[8\] ;
   wire \dpath.a_lt_b$in0\[7\] ;
   wire \dpath.a_lt_b$in0\[6\] ;
   wire \dpath.a_lt_b$in0\[5\] ;
   wire \dpath.a_lt_b$in0\[4\] ;
   wire \dpath.a_lt_b$in0\[3\] ;
   wire \dpath.a_lt_b$in0\[2\] ;
   wire \dpath.a_lt_b$in0\[1\] ;
   wire \dpath.a_lt_b$in0\[15\] ;
   wire \dpath.a_lt_b$in0\[14\] ;
   wire \dpath.a_lt_b$in0\[13\] ;
   wire \dpath.a_lt_b$in0\[12\] ;
   wire \dpath.a_lt_b$in0\[11\] ;
   wire \dpath.a_lt_b$in0\[10\] ;
   wire \dpath.a_lt_b$in0\[0\] ;
   wire \ctrl.state.out\[2\] ;
   wire \ctrl.state.out\[1\] ;
   wire clk;
   wire _437_;
   wire _436_;
   wire _435_;
   wire _434_;
   wire _433_;
   wire _432_;
   wire _431_;
   wire _430_;
   wire _429_;
   wire _428_;
   wire _427_;
   wire _426_;
   wire _425_;
   wire _424_;
   wire _423_;
   wire _422_;
   wire _421_;
   wire _420_;
   wire _419_;
   wire _418_;
   wire _417_;
   wire _416_;
   wire _415_;
   wire _414_;
   wire _413_;
   wire _412_;
   wire _411_;
   wire _410_;
   wire _409_;
   wire _408_;
   wire _407_;
   wire _406_;
   wire _405_;
   wire _404_;
   wire _403_;
   wire _402_;
   wire _401_;
   wire _400_;
   wire _399_;
   wire _398_;
   wire _397_;
   wire _396_;
   wire _395_;
   wire _394_;
   wire _393_;
   wire _392_;
   wire _391_;
   wire _390_;
   wire _389_;
   wire _388_;
   wire _387_;
   wire _386_;
   wire _385_;
   wire _384_;
   wire _383_;
   wire _382_;
   wire _381_;
   wire _380_;
   wire _379_;
   wire _378_;
   wire _377_;
   wire _376_;
   wire _375_;
   wire _374_;
   wire _373_;
   wire _372_;
   wire _371_;
   wire _370_;
   wire _369_;
   wire _368_;
   wire _367_;
   wire _366_;
   wire _365_;
   wire _364_;
   wire _363_;
   wire _362_;
   wire _361_;
   wire _360_;
   wire _359_;
   wire _358_;
   wire _357_;
   wire _356_;
   wire _355_;
   wire _354_;
   wire _353_;
   wire _352_;
   wire _351_;
   wire _350_;
   wire _349_;
   wire _348_;
   wire _347_;
   wire _346_;
   wire _345_;
   wire _344_;
   wire _343_;
   wire _342_;
   wire _341_;
   wire _340_;
   wire _339_;
   wire _338_;
   wire _337_;
   wire _336_;
   wire _335_;
   wire _334_;
   wire _333_;
   wire _332_;
   wire _331_;
   wire _330_;
   wire _329_;
   wire _328_;
   wire _327_;
   wire _326_;
   wire _325_;
   wire _324_;
   wire _323_;
   wire _322_;
   wire _321_;
   wire _320_;
   wire _319_;
   wire _318_;
   wire _317_;
   wire _316_;
   wire _315_;
   wire _314_;
   wire _313_;
   wire _312_;
   wire _311_;
   wire _310_;
   wire _309_;
   wire _308_;
   wire _307_;
   wire _306_;
   wire _305_;
   wire _304_;
   wire _303_;
   wire _302_;
   wire _301_;
   wire _300_;
   wire _299_;
   wire _298_;
   wire _297_;
   wire _296_;
   wire _295_;
   wire _294_;
   wire _293_;
   wire _292_;
   wire _291_;
   wire _290_;
   wire _289_;
   wire _288_;
   wire _287_;
   wire _286_;
   wire _285_;
   wire _284_;
   wire _283_;
   wire _282_;
   wire _281_;
   wire _280_;
   wire _279_;
   wire _278_;
   wire _277_;
   wire _276_;
   wire _275_;
   wire _274_;
   wire _273_;
   wire _272_;
   wire _271_;
   wire _270_;
   wire _269_;
   wire _268_;
   wire _267_;
   wire _266_;
   wire _265_;
   wire _264_;
   wire _263_;
   wire _262_;
   wire _261_;
   wire _260_;
   wire _259_;
   wire _258_;
   wire _257_;
   wire _256_;
   wire _255_;
   wire _254_;
   wire _253_;
   wire _252_;
   wire _251_;
   wire _250_;
   wire _249_;
   wire _248_;
   wire _247_;
   wire _246_;
   wire _245_;
   wire _244_;
   wire _243_;
   wire _242_;
   wire _241_;
   wire _240_;
   wire _239_;
   wire _238_;
   wire _237_;
   wire _236_;
   wire _235_;
   wire _234_;
   wire _233_;
   wire _232_;
   wire _231_;
   wire _230_;
   wire _229_;
   wire _228_;
   wire _227_;
   wire _226_;
   wire _225_;
   wire _224_;
   wire _223_;
   wire _222_;
   wire _221_;
   wire _220_;
   wire _219_;
   wire _218_;
   wire _217_;
   wire _216_;
   wire _215_;
   wire _214_;
   wire _213_;
   wire _212_;
   wire _211_;
   wire _210_;
   wire _209_;
   wire _208_;
   wire _207_;
   wire _206_;
   wire _205_;
   wire _204_;
   wire _203_;
   wire _202_;
   wire _201_;
   wire _200_;
   wire _199_;
   wire _198_;
   wire _197_;
   wire _196_;
   wire _195_;
   wire _194_;
   wire _193_;
   wire _192_;
   wire _191_;
   wire _190_;
   wire _189_;
   wire _188_;
   wire _187_;
   wire _186_;
   wire _185_;
   wire _184_;
   wire _183_;
   wire _182_;
   wire _181_;
   wire _180_;
   wire _179_;
   wire _178_;
   wire _177_;
   wire _176_;
   wire _175_;
   wire _174_;
   wire _173_;
   wire _172_;
   wire _171_;
   wire _170_;
   wire _169_;
   wire _168_;
   wire _167_;
   wire _166_;
   wire _165_;
   wire _164_;
   wire _163_;
   wire _162_;
   wire _161_;
   wire _160_;
   wire _159_;
   wire _158_;
   wire _157_;
   wire _156_;
   wire _155_;
   wire _154_;
   wire _153_;
   wire _152_;
   wire _151_;
   wire _150_;
   wire _149_;
   wire _148_;
   wire _147_;
   wire _146_;
   wire _145_;
   wire _144_;
   wire _143_;
   wire _142_;
   wire _141_;
   wire _140_;
   wire _139_;
   wire _138_;
   wire _137_;
   wire _136_;
   wire _135_;
   wire _134_;
   wire _133_;
   wire _132_;
   wire _131_;
   wire _130_;
   wire _129_;
   wire _128_;
   wire _127_;
   wire _126_;
   wire _125_;
   wire _124_;
   wire _123_;
   wire _122_;
   wire _121_;
   wire _120_;
   wire _119_;
   wire _118_;
   wire _117_;
   wire _116_;
   wire _115_;
   wire _114_;
   wire _113_;
   wire _112_;
   wire _111_;
   wire _110_;
   wire _109_;
   wire _108_;
   wire _107_;
   wire _106_;
   wire _105_;
   wire _104_;
   wire _103_;
   wire _102_;
   wire _101_;
   wire _100_;
   wire _099_;
   wire _098_;
   wire _097_;
   wire _096_;
   wire _095_;
   wire _094_;
   wire _093_;
   wire _092_;
   wire _091_;
   wire _090_;
   wire _089_;
   wire _088_;
   wire _087_;
   wire _086_;
   wire _085_;
   wire _084_;
   wire _083_;
   wire _082_;
   wire _081_;
   wire _080_;
   wire _079_;
   wire _078_;
   wire _077_;
   wire _076_;
   wire _075_;
   wire _074_;
   wire _073_;
   wire _072_;
   wire _071_;
   wire _070_;
   wire _069_;
   wire _068_;
   wire _067_;
   wire _066_;
   wire _065_;
   wire _064_;
   wire _063_;
   wire _062_;
   wire _061_;
   wire _060_;
   wire _059_;
   wire _058_;
   wire _057_;
   wire _056_;
   wire _055_;
   wire _054_;
   wire _053_;
   wire _052_;
   wire _051_;
   wire _050_;
   wire _049_;
   wire _048_;
   wire _047_;
   wire _046_;
   wire _045_;
   wire _044_;
   wire _043_;
   wire _042_;
   wire _041_;
   wire _040_;
   wire _039_;
   wire _038_;
   wire _037_;
   wire _036_;
   wire _035_;
   wire _034_;
   wire _033_;
   wire _032_;
   wire _031_;
   wire _030_;
   wire _029_;
   wire _028_;
   wire _027_;
   wire _026_;
   wire _025_;
   wire _024_;
   wire _023_;
   wire _022_;
   wire _021_;
   wire _020_;
   wire _019_;
   wire _018_;
   wire _017_;
   wire _016_;
   wire _015_;
   wire _014_;
   wire _013_;
   wire _012_;
   wire _011_;
   wire _010_;
   wire _009_;
   wire _008_;
   wire _007_;
   wire _006_;
   wire _005_;
   wire _004_;
   wire _003_;
   wire _002_;
   wire _001_;
   wire _000_;

   // Assignments 

   // Module instantiations
   BUF_X4 buffer9 (
	   .Z (net9),
	   .A (req_msg[23]) );
   BUF_X4 buffer8 (
	   .Z (net8),
	   .A (req_msg[24]) );
   BUF_X4 buffer7 (
	   .Z (net7),
	   .A (req_msg[25]) );
   BUF_X4 buffer6 (
	   .Z (net6),
	   .A (req_msg[26]) );
   BUF_X4 buffer53 (
	   .Z (resp_val),
	   .A (net53) );
   BUF_X4 buffer52 (
	   .Z (resp_msg[0]),
	   .A (net52) );
   BUF_X4 buffer51 (
	   .Z (resp_msg[1]),
	   .A (net51) );
   BUF_X4 buffer50 (
	   .Z (resp_msg[2]),
	   .A (net50) );
   BUF_X4 buffer5 (
	   .Z (net5),
	   .A (req_msg[27]) );
   BUF_X4 buffer49 (
	   .Z (resp_msg[3]),
	   .A (net49) );
   BUF_X4 buffer48 (
	   .Z (resp_msg[4]),
	   .A (net48) );
   BUF_X4 buffer47 (
	   .Z (resp_msg[5]),
	   .A (net47) );
   BUF_X4 buffer46 (
	   .Z (resp_msg[6]),
	   .A (net46) );
   BUF_X4 buffer45 (
	   .Z (resp_msg[7]),
	   .A (net45) );
   BUF_X4 buffer44 (
	   .Z (resp_msg[8]),
	   .A (net44) );
   BUF_X4 buffer43 (
	   .Z (resp_msg[9]),
	   .A (net43) );
   BUF_X4 buffer42 (
	   .Z (resp_msg[10]),
	   .A (net42) );
   BUF_X4 buffer41 (
	   .Z (resp_msg[11]),
	   .A (net41) );
   BUF_X4 buffer40 (
	   .Z (resp_msg[12]),
	   .A (net40) );
   BUF_X4 buffer4 (
	   .Z (net4),
	   .A (req_msg[28]) );
   BUF_X4 buffer39 (
	   .Z (resp_msg[13]),
	   .A (net39) );
   BUF_X4 buffer38 (
	   .Z (resp_msg[14]),
	   .A (net38) );
   BUF_X4 buffer37 (
	   .Z (resp_msg[15]),
	   .A (net37) );
   BUF_X4 buffer36 (
	   .Z (req_rdy),
	   .A (net36) );
   BUF_X4 buffer35 (
	   .Z (net35),
	   .A (resp_rdy) );
   BUF_X4 buffer34 (
	   .Z (net34),
	   .A (reset) );
   BUF_X4 buffer33 (
	   .Z (net33),
	   .A (req_val) );
   BUF_X4 buffer32 (
	   .Z (net32),
	   .A (req_msg[0]) );
   BUF_X4 buffer31 (
	   .Z (net31),
	   .A (req_msg[1]) );
   BUF_X4 buffer30 (
	   .Z (net30),
	   .A (req_msg[2]) );
   BUF_X4 buffer3 (
	   .Z (net3),
	   .A (req_msg[29]) );
   BUF_X4 buffer29 (
	   .Z (net29),
	   .A (req_msg[3]) );
   BUF_X4 buffer28 (
	   .Z (net28),
	   .A (req_msg[4]) );
   BUF_X4 buffer27 (
	   .Z (net27),
	   .A (req_msg[5]) );
   BUF_X4 buffer26 (
	   .Z (net26),
	   .A (req_msg[6]) );
   BUF_X4 buffer25 (
	   .Z (net25),
	   .A (req_msg[7]) );
   BUF_X4 buffer24 (
	   .Z (net24),
	   .A (req_msg[8]) );
   BUF_X4 buffer23 (
	   .Z (net23),
	   .A (req_msg[9]) );
   BUF_X4 buffer22 (
	   .Z (net22),
	   .A (req_msg[10]) );
   BUF_X4 buffer21 (
	   .Z (net21),
	   .A (req_msg[11]) );
   BUF_X4 buffer20 (
	   .Z (net20),
	   .A (req_msg[12]) );
   BUF_X4 buffer2 (
	   .Z (net2),
	   .A (req_msg[30]) );
   BUF_X4 buffer19 (
	   .Z (net19),
	   .A (req_msg[13]) );
   BUF_X4 buffer18 (
	   .Z (net18),
	   .A (req_msg[14]) );
   BUF_X4 buffer17 (
	   .Z (net17),
	   .A (req_msg[15]) );
   BUF_X4 buffer16 (
	   .Z (net16),
	   .A (req_msg[16]) );
   BUF_X4 buffer15 (
	   .Z (net15),
	   .A (req_msg[17]) );
   BUF_X4 buffer14 (
	   .Z (net14),
	   .A (req_msg[18]) );
   BUF_X4 buffer13 (
	   .Z (net13),
	   .A (req_msg[19]) );
   BUF_X4 buffer12 (
	   .Z (net12),
	   .A (req_msg[20]) );
   BUF_X4 buffer11 (
	   .Z (net11),
	   .A (req_msg[21]) );
   BUF_X4 buffer10 (
	   .Z (net10),
	   .A (req_msg[22]) );
   BUF_X4 buffer1 (
	   .Z (net1),
	   .A (req_msg[31]) );
   DFF_X1 _892_ (
	   .QN (_021_),
	   .Q (\dpath.a_lt_b$in1\[15\] ),
	   .D (_044_),
	   .CK (clk) );
   DFF_X1 _891_ (
	   .QN (_020_),
	   .Q (\dpath.a_lt_b$in1\[14\] ),
	   .D (_043_),
	   .CK (clk) );
   DFF_X1 _890_ (
	   .QN (_019_),
	   .Q (\dpath.a_lt_b$in1\[13\] ),
	   .D (_042_),
	   .CK (clk) );
   DFF_X1 _889_ (
	   .QN (_018_),
	   .Q (\dpath.a_lt_b$in1\[12\] ),
	   .D (_041_),
	   .CK (clk) );
   DFF_X1 _888_ (
	   .QN (_017_),
	   .Q (\dpath.a_lt_b$in1\[11\] ),
	   .D (_040_),
	   .CK (clk) );
   DFF_X1 _887_ (
	   .QN (_016_),
	   .Q (\dpath.a_lt_b$in1\[10\] ),
	   .D (_039_),
	   .CK (clk) );
   DFF_X1 _886_ (
	   .QN (_015_),
	   .Q (\dpath.a_lt_b$in1\[9\] ),
	   .D (_053_),
	   .CK (clk) );
   DFF_X1 _885_ (
	   .QN (_014_),
	   .Q (\dpath.a_lt_b$in1\[8\] ),
	   .D (_052_),
	   .CK (clk) );
   DFF_X1 _884_ (
	   .QN (_013_),
	   .Q (\dpath.a_lt_b$in1\[7\] ),
	   .D (_051_),
	   .CK (clk) );
   DFF_X1 _883_ (
	   .QN (_012_),
	   .Q (\dpath.a_lt_b$in1\[6\] ),
	   .D (_050_),
	   .CK (clk) );
   DFF_X1 _882_ (
	   .QN (_011_),
	   .Q (\dpath.a_lt_b$in1\[5\] ),
	   .D (_049_),
	   .CK (clk) );
   DFF_X1 _881_ (
	   .QN (_010_),
	   .Q (\dpath.a_lt_b$in1\[4\] ),
	   .D (_048_),
	   .CK (clk) );
   DFF_X1 _880_ (
	   .QN (_009_),
	   .Q (\dpath.a_lt_b$in1\[3\] ),
	   .D (_047_),
	   .CK (clk) );
   DFF_X1 _879_ (
	   .QN (_008_),
	   .Q (\dpath.a_lt_b$in1\[2\] ),
	   .D (_046_),
	   .CK (clk) );
   DFF_X1 _878_ (
	   .QN (_007_),
	   .Q (\dpath.a_lt_b$in1\[1\] ),
	   .D (_045_),
	   .CK (clk) );
   DFF_X1 _877_ (
	   .QN (_006_),
	   .Q (\dpath.a_lt_b$in1\[0\] ),
	   .D (_038_),
	   .CK (clk) );
   DFF_X1 _876_ (
	   .QN (_437_),
	   .Q (\dpath.a_lt_b$in0\[15\] ),
	   .D (_028_),
	   .CK (clk) );
   DFF_X1 _875_ (
	   .QN (_436_),
	   .Q (\dpath.a_lt_b$in0\[14\] ),
	   .D (_027_),
	   .CK (clk) );
   DFF_X1 _874_ (
	   .QN (_435_),
	   .Q (\dpath.a_lt_b$in0\[13\] ),
	   .D (_026_),
	   .CK (clk) );
   DFF_X1 _873_ (
	   .QN (_434_),
	   .Q (\dpath.a_lt_b$in0\[12\] ),
	   .D (_025_),
	   .CK (clk) );
   DFF_X1 _872_ (
	   .QN (_433_),
	   .Q (\dpath.a_lt_b$in0\[11\] ),
	   .D (_024_),
	   .CK (clk) );
   DFF_X1 _871_ (
	   .QN (_432_),
	   .Q (\dpath.a_lt_b$in0\[10\] ),
	   .D (_023_),
	   .CK (clk) );
   DFF_X1 _870_ (
	   .QN (_431_),
	   .Q (\dpath.a_lt_b$in0\[9\] ),
	   .D (_037_),
	   .CK (clk) );
   DFF_X1 _869_ (
	   .QN (_430_),
	   .Q (\dpath.a_lt_b$in0\[8\] ),
	   .D (_036_),
	   .CK (clk) );
   DFF_X1 _868_ (
	   .QN (_429_),
	   .Q (\dpath.a_lt_b$in0\[7\] ),
	   .D (_035_),
	   .CK (clk) );
   DFF_X1 _867_ (
	   .QN (_428_),
	   .Q (\dpath.a_lt_b$in0\[6\] ),
	   .D (_034_),
	   .CK (clk) );
   DFF_X1 _866_ (
	   .QN (_427_),
	   .Q (\dpath.a_lt_b$in0\[5\] ),
	   .D (_033_),
	   .CK (clk) );
   DFF_X1 _865_ (
	   .QN (_426_),
	   .Q (\dpath.a_lt_b$in0\[4\] ),
	   .D (_032_),
	   .CK (clk) );
   DFF_X1 _864_ (
	   .QN (_425_),
	   .Q (\dpath.a_lt_b$in0\[3\] ),
	   .D (_031_),
	   .CK (clk) );
   DFF_X1 _863_ (
	   .QN (_424_),
	   .Q (\dpath.a_lt_b$in0\[2\] ),
	   .D (_030_),
	   .CK (clk) );
   DFF_X1 _862_ (
	   .QN (_423_),
	   .Q (\dpath.a_lt_b$in0\[1\] ),
	   .D (_029_),
	   .CK (clk) );
   DFF_X1 _861_ (
	   .QN (_422_),
	   .Q (\dpath.a_lt_b$in0\[0\] ),
	   .D (_022_),
	   .CK (clk) );
   DFF_X1 _860_ (
	   .QN (_004_),
	   .Q (\ctrl.state.out\[2\] ),
	   .D (_002_),
	   .CK (clk) );
   DFF_X1 _859_ (
	   .QN (_003_),
	   .Q (\ctrl.state.out\[1\] ),
	   .D (_001_),
	   .CK (clk) );
   DFF_X1 _858_ (
	   .QN (_005_),
	   .Q (net36),
	   .D (_000_),
	   .CK (clk) );
   CLKBUF_X1 _857_ (
	   .Z (net37),
	   .A (_410_) );
   CLKBUF_X1 _856_ (
	   .Z (net38),
	   .A (_409_) );
   CLKBUF_X1 _855_ (
	   .Z (net39),
	   .A (_408_) );
   CLKBUF_X1 _854_ (
	   .Z (net40),
	   .A (_407_) );
   CLKBUF_X1 _853_ (
	   .Z (net41),
	   .A (_406_) );
   CLKBUF_X1 _852_ (
	   .Z (net42),
	   .A (_405_) );
   CLKBUF_X1 _851_ (
	   .Z (net43),
	   .A (_419_) );
   CLKBUF_X1 _850_ (
	   .Z (net44),
	   .A (_418_) );
   CLKBUF_X1 _849_ (
	   .Z (net45),
	   .A (_417_) );
   CLKBUF_X1 _848_ (
	   .Z (net46),
	   .A (_416_) );
   CLKBUF_X1 _847_ (
	   .Z (net47),
	   .A (_415_) );
   CLKBUF_X1 _846_ (
	   .Z (net48),
	   .A (_414_) );
   CLKBUF_X1 _845_ (
	   .Z (net49),
	   .A (_413_) );
   CLKBUF_X1 _844_ (
	   .Z (net50),
	   .A (_412_) );
   CLKBUF_X1 _843_ (
	   .Z (net51),
	   .A (_411_) );
   CLKBUF_X1 _842_ (
	   .Z (_044_),
	   .A (_098_) );
   CLKBUF_X1 _841_ (
	   .Z (_375_),
	   .A (net17) );
   CLKBUF_X1 _840_ (
	   .Z (_043_),
	   .A (_097_) );
   CLKBUF_X1 _839_ (
	   .Z (_374_),
	   .A (net18) );
   CLKBUF_X1 _838_ (
	   .Z (_042_),
	   .A (_096_) );
   CLKBUF_X1 _837_ (
	   .Z (_373_),
	   .A (net19) );
   CLKBUF_X1 _836_ (
	   .Z (_041_),
	   .A (_095_) );
   CLKBUF_X1 _835_ (
	   .Z (_372_),
	   .A (net20) );
   CLKBUF_X1 _834_ (
	   .Z (_040_),
	   .A (_094_) );
   CLKBUF_X1 _833_ (
	   .Z (_371_),
	   .A (net21) );
   CLKBUF_X1 _832_ (
	   .Z (_039_),
	   .A (_093_) );
   CLKBUF_X1 _831_ (
	   .Z (_370_),
	   .A (net22) );
   CLKBUF_X1 _830_ (
	   .Z (_053_),
	   .A (_107_) );
   CLKBUF_X1 _829_ (
	   .Z (_400_),
	   .A (net23) );
   CLKBUF_X1 _828_ (
	   .Z (_052_),
	   .A (_106_) );
   CLKBUF_X1 _827_ (
	   .Z (_399_),
	   .A (net24) );
   CLKBUF_X1 _826_ (
	   .Z (_051_),
	   .A (_105_) );
   CLKBUF_X1 _825_ (
	   .Z (_398_),
	   .A (net25) );
   CLKBUF_X1 _824_ (
	   .Z (_050_),
	   .A (_104_) );
   CLKBUF_X1 _823_ (
	   .Z (_397_),
	   .A (net26) );
   CLKBUF_X1 _822_ (
	   .Z (_049_),
	   .A (_103_) );
   CLKBUF_X1 _821_ (
	   .Z (_396_),
	   .A (net27) );
   CLKBUF_X1 _820_ (
	   .Z (_048_),
	   .A (_102_) );
   CLKBUF_X1 _819_ (
	   .Z (_395_),
	   .A (net28) );
   CLKBUF_X1 _818_ (
	   .Z (_047_),
	   .A (_101_) );
   CLKBUF_X1 _817_ (
	   .Z (_394_),
	   .A (net29) );
   CLKBUF_X1 _816_ (
	   .Z (_046_),
	   .A (_100_) );
   CLKBUF_X1 _815_ (
	   .Z (_391_),
	   .A (net30) );
   CLKBUF_X1 _814_ (
	   .Z (_045_),
	   .A (_099_) );
   CLKBUF_X1 _813_ (
	   .Z (_380_),
	   .A (net31) );
   CLKBUF_X1 _812_ (
	   .Z (_038_),
	   .A (_092_) );
   CLKBUF_X1 _811_ (
	   .Z (_369_),
	   .A (net32) );
   CLKBUF_X1 _810_ (
	   .Z (_028_),
	   .A (_082_) );
   CLKBUF_X1 _809_ (
	   .Z (_393_),
	   .A (net1) );
   CLKBUF_X1 _808_ (
	   .Z (_075_),
	   .A (_021_) );
   CLKBUF_X1 _807_ (
	   .Z (_027_),
	   .A (_081_) );
   CLKBUF_X1 _806_ (
	   .Z (_392_),
	   .A (net2) );
   CLKBUF_X1 _805_ (
	   .Z (_074_),
	   .A (_020_) );
   CLKBUF_X1 _804_ (
	   .Z (_026_),
	   .A (_080_) );
   CLKBUF_X1 _803_ (
	   .Z (_390_),
	   .A (net3) );
   CLKBUF_X1 _802_ (
	   .Z (_073_),
	   .A (_019_) );
   CLKBUF_X1 _801_ (
	   .Z (_025_),
	   .A (_079_) );
   CLKBUF_X1 _800_ (
	   .Z (_389_),
	   .A (net4) );
   CLKBUF_X1 _799_ (
	   .Z (_072_),
	   .A (_018_) );
   CLKBUF_X1 _798_ (
	   .Z (_024_),
	   .A (_078_) );
   CLKBUF_X1 _797_ (
	   .Z (_388_),
	   .A (net5) );
   CLKBUF_X1 _796_ (
	   .Z (_071_),
	   .A (_017_) );
   CLKBUF_X1 _795_ (
	   .Z (_023_),
	   .A (_077_) );
   CLKBUF_X1 _794_ (
	   .Z (_387_),
	   .A (net6) );
   CLKBUF_X1 _793_ (
	   .Z (_070_),
	   .A (_016_) );
   CLKBUF_X1 _792_ (
	   .Z (_037_),
	   .A (_091_) );
   CLKBUF_X1 _791_ (
	   .Z (_386_),
	   .A (net7) );
   CLKBUF_X1 _790_ (
	   .Z (_069_),
	   .A (_015_) );
   CLKBUF_X1 _789_ (
	   .Z (_036_),
	   .A (_090_) );
   CLKBUF_X1 _788_ (
	   .Z (_385_),
	   .A (net8) );
   CLKBUF_X1 _787_ (
	   .Z (_068_),
	   .A (_014_) );
   CLKBUF_X1 _786_ (
	   .Z (_035_),
	   .A (_089_) );
   CLKBUF_X1 _785_ (
	   .Z (_384_),
	   .A (net9) );
   CLKBUF_X1 _784_ (
	   .Z (_067_),
	   .A (_013_) );
   CLKBUF_X1 _783_ (
	   .Z (_034_),
	   .A (_088_) );
   CLKBUF_X1 _782_ (
	   .Z (_383_),
	   .A (net10) );
   CLKBUF_X1 _781_ (
	   .Z (_066_),
	   .A (_012_) );
   CLKBUF_X1 _780_ (
	   .Z (_033_),
	   .A (_087_) );
   CLKBUF_X1 _779_ (
	   .Z (_382_),
	   .A (net11) );
   CLKBUF_X1 _778_ (
	   .Z (_065_),
	   .A (_011_) );
   CLKBUF_X1 _777_ (
	   .Z (_032_),
	   .A (_086_) );
   CLKBUF_X1 _776_ (
	   .Z (_381_),
	   .A (net12) );
   CLKBUF_X1 _775_ (
	   .Z (_064_),
	   .A (_010_) );
   CLKBUF_X1 _774_ (
	   .Z (_031_),
	   .A (_085_) );
   CLKBUF_X1 _773_ (
	   .Z (_379_),
	   .A (net13) );
   CLKBUF_X1 _772_ (
	   .Z (_063_),
	   .A (_009_) );
   CLKBUF_X1 _771_ (
	   .Z (_030_),
	   .A (_084_) );
   CLKBUF_X1 _770_ (
	   .Z (_378_),
	   .A (net14) );
   CLKBUF_X1 _769_ (
	   .Z (_062_),
	   .A (_008_) );
   CLKBUF_X1 _768_ (
	   .Z (_029_),
	   .A (_083_) );
   CLKBUF_X1 _767_ (
	   .Z (_377_),
	   .A (net15) );
   CLKBUF_X1 _766_ (
	   .Z (_061_),
	   .A (_007_) );
   CLKBUF_X1 _765_ (
	   .Z (_022_),
	   .A (_076_) );
   CLKBUF_X1 _764_ (
	   .Z (_376_),
	   .A (net16) );
   CLKBUF_X1 _763_ (
	   .Z (_060_),
	   .A (_006_) );
   CLKBUF_X1 _762_ (
	   .Z (_000_),
	   .A (_054_) );
   CLKBUF_X1 _761_ (
	   .Z (_002_),
	   .A (_056_) );
   CLKBUF_X1 _760_ (
	   .Z (_402_),
	   .A (net33) );
   BUF_X2 _759_ (
	   .Z (_401_),
	   .A (net36) );
   CLKBUF_X1 _758_ (
	   .Z (_001_),
	   .A (_055_) );
   CLKBUF_X1 _757_ (
	   .Z (_057_),
	   .A (_003_) );
   CLKBUF_X1 _756_ (
	   .Z (_058_),
	   .A (_004_) );
   CLKBUF_X1 _755_ (
	   .Z (net52),
	   .A (_404_) );
   BUF_X1 _754_ (
	   .Z (_126_),
	   .A (\dpath.a_lt_b$in1\[0\] ) );
   CLKBUF_X1 _753_ (
	   .Z (_110_),
	   .A (\dpath.a_lt_b$in0\[0\] ) );
   BUF_X1 _752_ (
	   .Z (_133_),
	   .A (\dpath.a_lt_b$in1\[1\] ) );
   BUF_X1 _751_ (
	   .Z (_117_),
	   .A (\dpath.a_lt_b$in0\[1\] ) );
   CLKBUF_X1 _750_ (
	   .Z (_134_),
	   .A (\dpath.a_lt_b$in1\[2\] ) );
   CLKBUF_X1 _749_ (
	   .Z (_118_),
	   .A (\dpath.a_lt_b$in0\[2\] ) );
   CLKBUF_X1 _748_ (
	   .Z (_135_),
	   .A (\dpath.a_lt_b$in1\[3\] ) );
   BUF_X1 _747_ (
	   .Z (_119_),
	   .A (\dpath.a_lt_b$in0\[3\] ) );
   CLKBUF_X1 _746_ (
	   .Z (_136_),
	   .A (\dpath.a_lt_b$in1\[4\] ) );
   CLKBUF_X1 _745_ (
	   .Z (_120_),
	   .A (\dpath.a_lt_b$in0\[4\] ) );
   BUF_X1 _744_ (
	   .Z (_137_),
	   .A (\dpath.a_lt_b$in1\[5\] ) );
   CLKBUF_X1 _743_ (
	   .Z (_121_),
	   .A (\dpath.a_lt_b$in0\[5\] ) );
   BUF_X1 _742_ (
	   .Z (_138_),
	   .A (\dpath.a_lt_b$in1\[6\] ) );
   CLKBUF_X1 _741_ (
	   .Z (_122_),
	   .A (\dpath.a_lt_b$in0\[6\] ) );
   BUF_X1 _740_ (
	   .Z (_139_),
	   .A (\dpath.a_lt_b$in1\[7\] ) );
   BUF_X1 _739_ (
	   .Z (_123_),
	   .A (\dpath.a_lt_b$in0\[7\] ) );
   CLKBUF_X1 _738_ (
	   .Z (_140_),
	   .A (\dpath.a_lt_b$in1\[8\] ) );
   CLKBUF_X1 _737_ (
	   .Z (_124_),
	   .A (\dpath.a_lt_b$in0\[8\] ) );
   BUF_X1 _736_ (
	   .Z (_141_),
	   .A (\dpath.a_lt_b$in1\[9\] ) );
   CLKBUF_X1 _735_ (
	   .Z (_125_),
	   .A (\dpath.a_lt_b$in0\[9\] ) );
   BUF_X1 _734_ (
	   .Z (_127_),
	   .A (\dpath.a_lt_b$in1\[10\] ) );
   CLKBUF_X1 _733_ (
	   .Z (_111_),
	   .A (\dpath.a_lt_b$in0\[10\] ) );
   BUF_X1 _732_ (
	   .Z (_128_),
	   .A (\dpath.a_lt_b$in1\[11\] ) );
   CLKBUF_X1 _731_ (
	   .Z (_112_),
	   .A (\dpath.a_lt_b$in0\[11\] ) );
   BUF_X1 _730_ (
	   .Z (_129_),
	   .A (\dpath.a_lt_b$in1\[12\] ) );
   CLKBUF_X1 _729_ (
	   .Z (_113_),
	   .A (\dpath.a_lt_b$in0\[12\] ) );
   CLKBUF_X2 _728_ (
	   .Z (_130_),
	   .A (\dpath.a_lt_b$in1\[13\] ) );
   BUF_X1 _727_ (
	   .Z (_114_),
	   .A (\dpath.a_lt_b$in0\[13\] ) );
   BUF_X1 _726_ (
	   .Z (_131_),
	   .A (\dpath.a_lt_b$in1\[14\] ) );
   CLKBUF_X1 _725_ (
	   .Z (_115_),
	   .A (\dpath.a_lt_b$in0\[14\] ) );
   BUF_X1 _724_ (
	   .Z (_132_),
	   .A (\dpath.a_lt_b$in1\[15\] ) );
   CLKBUF_X1 _723_ (
	   .Z (_116_),
	   .A (\dpath.a_lt_b$in0\[15\] ) );
   CLKBUF_X1 _722_ (
	   .Z (_420_),
	   .A (net35) );
   CLKBUF_X1 _721_ (
	   .Z (net53),
	   .A (_421_) );
   BUF_X1 _720_ (
	   .Z (_059_),
	   .A (_005_) );
   CLKBUF_X1 _719_ (
	   .Z (_108_),
	   .A (\ctrl.state.out\[1\] ) );
   CLKBUF_X1 _718_ (
	   .Z (_109_),
	   .A (\ctrl.state.out\[2\] ) );
   CLKBUF_X1 _717_ (
	   .Z (_403_),
	   .A (net34) );
   MUX2_X1 _716_ (
	   .Z (_098_),
	   .S (_352_),
	   .B (_368_),
	   .A (_132_) );
   MUX2_X1 _715_ (
	   .Z (_368_),
	   .S (_401_),
	   .B (_375_),
	   .A (_116_) );
   MUX2_X1 _714_ (
	   .Z (_097_),
	   .S (_352_),
	   .B (_367_),
	   .A (_131_) );
   MUX2_X1 _713_ (
	   .Z (_367_),
	   .S (_401_),
	   .B (_374_),
	   .A (_115_) );
   MUX2_X1 _712_ (
	   .Z (_096_),
	   .S (_352_),
	   .B (_366_),
	   .A (_130_) );
   MUX2_X1 _711_ (
	   .Z (_366_),
	   .S (_401_),
	   .B (_373_),
	   .A (_114_) );
   MUX2_X1 _710_ (
	   .Z (_095_),
	   .S (_352_),
	   .B (_365_),
	   .A (_129_) );
   MUX2_X1 _709_ (
	   .Z (_365_),
	   .S (_401_),
	   .B (_372_),
	   .A (_113_) );
   MUX2_X1 _708_ (
	   .Z (_094_),
	   .S (_352_),
	   .B (_364_),
	   .A (_128_) );
   MUX2_X1 _707_ (
	   .Z (_364_),
	   .S (_401_),
	   .B (_371_),
	   .A (_112_) );
   MUX2_X1 _706_ (
	   .Z (_093_),
	   .S (_352_),
	   .B (_363_),
	   .A (_127_) );
   MUX2_X1 _705_ (
	   .Z (_363_),
	   .S (_401_),
	   .B (_370_),
	   .A (_111_) );
   MUX2_X1 _704_ (
	   .Z (_107_),
	   .S (_353_),
	   .B (_362_),
	   .A (_141_) );
   MUX2_X1 _703_ (
	   .Z (_362_),
	   .S (_401_),
	   .B (_400_),
	   .A (_125_) );
   MUX2_X1 _702_ (
	   .Z (_106_),
	   .S (_353_),
	   .B (_361_),
	   .A (_140_) );
   MUX2_X1 _701_ (
	   .Z (_361_),
	   .S (_401_),
	   .B (_399_),
	   .A (_124_) );
   MUX2_X1 _700_ (
	   .Z (_105_),
	   .S (_353_),
	   .B (_360_),
	   .A (_139_) );
   MUX2_X1 _699_ (
	   .Z (_360_),
	   .S (_160_),
	   .B (_398_),
	   .A (_123_) );
   MUX2_X1 _698_ (
	   .Z (_104_),
	   .S (_353_),
	   .B (_359_),
	   .A (_138_) );
   MUX2_X1 _697_ (
	   .Z (_359_),
	   .S (_160_),
	   .B (_397_),
	   .A (_122_) );
   MUX2_X1 _696_ (
	   .Z (_103_),
	   .S (_353_),
	   .B (_358_),
	   .A (_137_) );
   MUX2_X1 _695_ (
	   .Z (_358_),
	   .S (_160_),
	   .B (_396_),
	   .A (_121_) );
   MUX2_X1 _694_ (
	   .Z (_102_),
	   .S (_353_),
	   .B (_357_),
	   .A (_136_) );
   MUX2_X1 _693_ (
	   .Z (_357_),
	   .S (_160_),
	   .B (_395_),
	   .A (_120_) );
   MUX2_X1 _692_ (
	   .Z (_101_),
	   .S (_353_),
	   .B (_356_),
	   .A (_135_) );
   MUX2_X1 _691_ (
	   .Z (_356_),
	   .S (_160_),
	   .B (_394_),
	   .A (_119_) );
   MUX2_X1 _690_ (
	   .Z (_100_),
	   .S (_353_),
	   .B (_355_),
	   .A (_134_) );
   MUX2_X1 _689_ (
	   .Z (_355_),
	   .S (_160_),
	   .B (_391_),
	   .A (_118_) );
   MUX2_X1 _688_ (
	   .Z (_099_),
	   .S (_353_),
	   .B (_354_),
	   .A (_133_) );
   MUX2_X1 _687_ (
	   .Z (_354_),
	   .S (_160_),
	   .B (_380_),
	   .A (_117_) );
   MUX2_X1 _686_ (
	   .Z (_092_),
	   .S (_353_),
	   .B (_351_),
	   .A (_126_) );
   BUF_X2 _685_ (
	   .Z (_353_),
	   .A (_352_) );
   NAND2_X2 _684_ (
	   .ZN (_352_),
	   .A2 (_059_),
	   .A1 (_243_) );
   MUX2_X1 _683_ (
	   .Z (_351_),
	   .S (_160_),
	   .B (_369_),
	   .A (_110_) );
   OAI21_X1 _682_ (
	   .ZN (_082_),
	   .B2 (_249_),
	   .B1 (_167_),
	   .A (_350_) );
   OAI21_X1 _681_ (
	   .ZN (_350_),
	   .B2 (_349_),
	   .B1 (_347_),
	   .A (_249_) );
   OAI21_X1 _680_ (
	   .ZN (_349_),
	   .B2 (_075_),
	   .B1 (_245_),
	   .A (_348_) );
   OAI21_X1 _679_ (
	   .ZN (_348_),
	   .B2 (_159_),
	   .B1 (_165_),
	   .A (_393_) );
   AND2_X1 _678_ (
	   .ZN (_347_),
	   .A2 (_253_),
	   .A1 (_410_) );
   XNOR2_X1 _677_ (
	   .ZN (_410_),
	   .B (_207_),
	   .A (_346_) );
   NOR2_X1 _676_ (
	   .ZN (_346_),
	   .A2 (_345_),
	   .A1 (_341_) );
   NOR2_X1 _675_ (
	   .ZN (_345_),
	   .A2 (_131_),
	   .A1 (_227_) );
   MUX2_X1 _674_ (
	   .Z (_081_),
	   .S (_248_),
	   .B (_344_),
	   .A (_115_) );
   OAI211_X1 _673_ (
	   .ZN (_344_),
	   .C2 (_244_),
	   .C1 (_074_),
	   .B (_343_),
	   .A (_342_) );
   OAI21_X1 _672_ (
	   .ZN (_343_),
	   .B2 (_158_),
	   .B1 (_142_),
	   .A (_392_) );
   NAND2_X1 _671_ (
	   .ZN (_342_),
	   .A2 (_252_),
	   .A1 (_409_) );
   NOR2_X1 _670_ (
	   .ZN (_409_),
	   .A2 (_341_),
	   .A1 (_340_) );
   AOI21_X1 _669_ (
	   .ZN (_341_),
	   .B2 (_339_),
	   .B1 (_337_),
	   .A (_338_) );
   AND3_X1 _668_ (
	   .ZN (_340_),
	   .A3 (_339_),
	   .A2 (_338_),
	   .A1 (_337_) );
   AOI22_X1 _667_ (
	   .ZN (_339_),
	   .B2 (_073_),
	   .B1 (_114_),
	   .A2 (_332_),
	   .A1 (_209_) );
   INV_X1 _666_ (
	   .ZN (_338_),
	   .A (_206_) );
   OR3_X1 _665_ (
	   .ZN (_337_),
	   .A3 (_212_),
	   .A2 (_210_),
	   .A1 (_327_) );
   MUX2_X1 _664_ (
	   .Z (_080_),
	   .S (_248_),
	   .B (_336_),
	   .A (_114_) );
   OAI211_X1 _663_ (
	   .ZN (_336_),
	   .C2 (_244_),
	   .C1 (_073_),
	   .B (_335_),
	   .A (_334_) );
   OAI21_X1 _662_ (
	   .ZN (_335_),
	   .B2 (_158_),
	   .B1 (_142_),
	   .A (_390_) );
   NAND2_X1 _661_ (
	   .ZN (_334_),
	   .A2 (_252_),
	   .A1 (_408_) );
   XNOR2_X1 _660_ (
	   .ZN (_408_),
	   .B (_209_),
	   .A (_333_) );
   NOR2_X1 _659_ (
	   .ZN (_333_),
	   .A2 (_332_),
	   .A1 (_331_) );
   NOR2_X1 _658_ (
	   .ZN (_332_),
	   .A2 (_129_),
	   .A1 (_233_) );
   NOR2_X1 _657_ (
	   .ZN (_331_),
	   .A2 (_212_),
	   .A1 (_327_) );
   MUX2_X1 _656_ (
	   .Z (_079_),
	   .S (_248_),
	   .B (_330_),
	   .A (_113_) );
   OAI211_X1 _655_ (
	   .ZN (_330_),
	   .C2 (_072_),
	   .C1 (_244_),
	   .B (_329_),
	   .A (_328_) );
   OAI21_X1 _654_ (
	   .ZN (_329_),
	   .B2 (_158_),
	   .B1 (_142_),
	   .A (_389_) );
   NAND2_X1 _653_ (
	   .ZN (_328_),
	   .A2 (_252_),
	   .A1 (_407_) );
   XNOR2_X1 _652_ (
	   .ZN (_407_),
	   .B (_211_),
	   .A (_327_) );
   AND3_X1 _651_ (
	   .ZN (_327_),
	   .A3 (_326_),
	   .A2 (_325_),
	   .A1 (_324_) );
   AOI21_X1 _650_ (
	   .ZN (_326_),
	   .B2 (_318_),
	   .B1 (_201_),
	   .A (_222_) );
   NAND2_X1 _649_ (
	   .ZN (_325_),
	   .A2 (_202_),
	   .A1 (_311_) );
   INV_X1 _648_ (
	   .ZN (_324_),
	   .A (_323_) );
   AND2_X1 _647_ (
	   .ZN (_323_),
	   .A2 (_205_),
	   .A1 (_298_) );
   OAI21_X1 _646_ (
	   .ZN (_078_),
	   .B2 (_249_),
	   .B1 (_221_),
	   .A (_322_) );
   OAI21_X1 _645_ (
	   .ZN (_322_),
	   .B2 (_321_),
	   .B1 (_316_),
	   .A (_249_) );
   AND2_X1 _644_ (
	   .ZN (_321_),
	   .A2 (_253_),
	   .A1 (_406_) );
   XNOR2_X1 _643_ (
	   .ZN (_406_),
	   .B (_201_),
	   .A (_320_) );
   AND2_X1 _642_ (
	   .ZN (_320_),
	   .A2 (_319_),
	   .A1 (_317_) );
   INV_X1 _641_ (
	   .ZN (_319_),
	   .A (_318_) );
   NOR2_X1 _640_ (
	   .ZN (_318_),
	   .A2 (_127_),
	   .A1 (_223_) );
   OAI21_X1 _639_ (
	   .ZN (_317_),
	   .B2 (_311_),
	   .B1 (_302_),
	   .A (_200_) );
   OAI21_X1 _638_ (
	   .ZN (_316_),
	   .B2 (_071_),
	   .B1 (_245_),
	   .A (_315_) );
   OAI21_X1 _637_ (
	   .ZN (_315_),
	   .B2 (_159_),
	   .B1 (_165_),
	   .A (_388_) );
   MUX2_X1 _636_ (
	   .Z (_077_),
	   .S (_248_),
	   .B (_314_),
	   .A (_111_) );
   OAI211_X1 _635_ (
	   .ZN (_314_),
	   .C2 (_070_),
	   .C1 (_244_),
	   .B (_313_),
	   .A (_308_) );
   NAND2_X1 _634_ (
	   .ZN (_313_),
	   .A2 (_405_),
	   .A1 (_252_) );
   XNOR2_X1 _633_ (
	   .ZN (_405_),
	   .B (_200_),
	   .A (_312_) );
   NOR2_X1 _632_ (
	   .ZN (_312_),
	   .A2 (_311_),
	   .A1 (_302_) );
   INV_X1 _631_ (
	   .ZN (_311_),
	   .A (_310_) );
   AOI21_X1 _630_ (
	   .ZN (_310_),
	   .B2 (_304_),
	   .B1 (_203_),
	   .A (_309_) );
   NOR2_X1 _629_ (
	   .ZN (_309_),
	   .A2 (_141_),
	   .A1 (_218_) );
   OAI21_X1 _628_ (
	   .ZN (_308_),
	   .B2 (_158_),
	   .B1 (_142_),
	   .A (_387_) );
   MUX2_X1 _627_ (
	   .Z (_091_),
	   .S (_248_),
	   .B (_307_),
	   .A (_125_) );
   OAI211_X1 _626_ (
	   .ZN (_307_),
	   .C2 (_069_),
	   .C1 (_244_),
	   .B (_306_),
	   .A (_301_) );
   NAND2_X1 _625_ (
	   .ZN (_306_),
	   .A2 (_252_),
	   .A1 (_419_) );
   AOI211_X1 _624_ (
	   .ZN (_419_),
	   .C2 (_304_),
	   .C1 (_203_),
	   .B (_305_),
	   .A (_302_) );
   NOR3_X1 _623_ (
	   .ZN (_305_),
	   .A3 (_304_),
	   .A2 (_203_),
	   .A1 (_303_) );
   NOR2_X1 _622_ (
	   .ZN (_304_),
	   .A2 (_140_),
	   .A1 (_216_) );
   AND2_X1 _621_ (
	   .ZN (_303_),
	   .A2 (_204_),
	   .A1 (_298_) );
   AND3_X1 _620_ (
	   .ZN (_302_),
	   .A3 (_204_),
	   .A2 (_203_),
	   .A1 (_298_) );
   OAI21_X1 _619_ (
	   .ZN (_301_),
	   .B2 (_158_),
	   .B1 (_142_),
	   .A (_386_) );
   MUX2_X1 _618_ (
	   .Z (_090_),
	   .S (_248_),
	   .B (_300_),
	   .A (_124_) );
   OAI211_X1 _617_ (
	   .ZN (_300_),
	   .C2 (_068_),
	   .C1 (_244_),
	   .B (_299_),
	   .A (_294_) );
   NAND2_X1 _616_ (
	   .ZN (_299_),
	   .A2 (_418_),
	   .A1 (_253_) );
   XOR2_X1 _615_ (
	   .Z (_418_),
	   .B (_204_),
	   .A (_298_) );
   NAND2_X1 _614_ (
	   .ZN (_298_),
	   .A2 (_297_),
	   .A1 (_295_) );
   AOI221_X1 _613_ (
	   .ZN (_297_),
	   .C2 (_171_),
	   .C1 (_283_),
	   .B2 (_190_),
	   .B1 (_123_),
	   .A (_296_) );
   AND2_X1 _612_ (
	   .ZN (_296_),
	   .A2 (_289_),
	   .A1 (_169_) );
   NAND2_X1 _611_ (
	   .ZN (_295_),
	   .A2 (_237_),
	   .A1 (_272_) );
   OAI21_X1 _610_ (
	   .ZN (_294_),
	   .B2 (_158_),
	   .B1 (_142_),
	   .A (_385_) );
   MUX2_X1 _609_ (
	   .Z (_089_),
	   .S (_248_),
	   .B (_293_),
	   .A (_123_) );
   OAI211_X1 _608_ (
	   .ZN (_293_),
	   .C2 (_067_),
	   .C1 (_245_),
	   .B (_292_),
	   .A (_287_) );
   NAND2_X1 _607_ (
	   .ZN (_292_),
	   .A2 (_417_),
	   .A1 (_253_) );
   XNOR2_X1 _606_ (
	   .ZN (_417_),
	   .B (_169_),
	   .A (_291_) );
   NOR2_X1 _605_ (
	   .ZN (_291_),
	   .A2 (_289_),
	   .A1 (_290_) );
   NOR3_X1 _604_ (
	   .ZN (_290_),
	   .A3 (_289_),
	   .A2 (_288_),
	   .A1 (_284_) );
   NOR2_X1 _603_ (
	   .ZN (_289_),
	   .A2 (_138_),
	   .A1 (_193_) );
   AND2_X1 _602_ (
	   .ZN (_288_),
	   .A2 (_138_),
	   .A1 (_193_) );
   OAI21_X1 _601_ (
	   .ZN (_287_),
	   .B2 (_158_),
	   .B1 (_165_),
	   .A (_384_) );
   MUX2_X1 _600_ (
	   .Z (_088_),
	   .S (_248_),
	   .B (_286_),
	   .A (_122_) );
   OAI211_X1 _599_ (
	   .ZN (_286_),
	   .C2 (_066_),
	   .C1 (_245_),
	   .B (_285_),
	   .A (_281_) );
   NAND2_X1 _598_ (
	   .ZN (_285_),
	   .A2 (_416_),
	   .A1 (_253_) );
   XNOR2_X1 _597_ (
	   .ZN (_416_),
	   .B (_170_),
	   .A (_284_) );
   AOI21_X1 _596_ (
	   .ZN (_284_),
	   .B2 (_177_),
	   .B1 (_272_),
	   .A (_283_) );
   OAI21_X1 _595_ (
	   .ZN (_283_),
	   .B2 (_137_),
	   .B1 (_187_),
	   .A (_282_) );
   NAND2_X1 _594_ (
	   .ZN (_282_),
	   .A2 (_277_),
	   .A1 (_175_) );
   OAI21_X1 _593_ (
	   .ZN (_281_),
	   .B2 (_159_),
	   .B1 (_165_),
	   .A (_383_) );
   MUX2_X1 _592_ (
	   .Z (_087_),
	   .S (_249_),
	   .B (_280_),
	   .A (_121_) );
   OAI211_X1 _591_ (
	   .ZN (_280_),
	   .C2 (_065_),
	   .C1 (_245_),
	   .B (_279_),
	   .A (_275_) );
   NAND2_X1 _590_ (
	   .ZN (_279_),
	   .A2 (_415_),
	   .A1 (_253_) );
   AOI221_X4 _589_ (
	   .ZN (_415_),
	   .C2 (_272_),
	   .C1 (_177_),
	   .B2 (_277_),
	   .B1 (_175_),
	   .A (_278_) );
   NOR3_X1 _588_ (
	   .ZN (_278_),
	   .A3 (_277_),
	   .A2 (_175_),
	   .A1 (_276_) );
   NOR2_X1 _587_ (
	   .ZN (_277_),
	   .A2 (_136_),
	   .A1 (_185_) );
   AND2_X1 _586_ (
	   .ZN (_276_),
	   .A2 (_176_),
	   .A1 (_272_) );
   OAI21_X1 _585_ (
	   .ZN (_275_),
	   .B2 (_159_),
	   .B1 (_165_),
	   .A (_382_) );
   MUX2_X1 _584_ (
	   .Z (_086_),
	   .S (_249_),
	   .B (_274_),
	   .A (_120_) );
   OAI211_X1 _583_ (
	   .ZN (_274_),
	   .C2 (_064_),
	   .C1 (_245_),
	   .B (_273_),
	   .A (_268_) );
   NAND2_X1 _582_ (
	   .ZN (_273_),
	   .A2 (_414_),
	   .A1 (_253_) );
   XOR2_X1 _581_ (
	   .Z (_414_),
	   .B (_176_),
	   .A (_272_) );
   NAND2_X1 _580_ (
	   .ZN (_272_),
	   .A2 (_271_),
	   .A1 (_270_) );
   NAND2_X1 _579_ (
	   .ZN (_271_),
	   .A2 (_174_),
	   .A1 (_262_) );
   AOI21_X1 _578_ (
	   .ZN (_270_),
	   .B2 (_144_),
	   .B1 (_119_),
	   .A (_269_) );
   AND2_X1 _577_ (
	   .ZN (_269_),
	   .A2 (_264_),
	   .A1 (_172_) );
   OAI21_X1 _576_ (
	   .ZN (_268_),
	   .B2 (_159_),
	   .B1 (_165_),
	   .A (_381_) );
   MUX2_X1 _575_ (
	   .Z (_085_),
	   .S (_249_),
	   .B (_267_),
	   .A (_119_) );
   OAI211_X1 _574_ (
	   .ZN (_267_),
	   .C2 (_063_),
	   .C1 (_245_),
	   .B (_266_),
	   .A (_261_) );
   NAND2_X1 _573_ (
	   .ZN (_266_),
	   .A2 (_413_),
	   .A1 (_253_) );
   XNOR2_X1 _572_ (
	   .ZN (_413_),
	   .B (_172_),
	   .A (_265_) );
   NOR2_X1 _571_ (
	   .ZN (_265_),
	   .A2 (_264_),
	   .A1 (_263_) );
   AND2_X1 _570_ (
	   .ZN (_264_),
	   .A2 (_118_),
	   .A1 (_145_) );
   AND2_X1 _569_ (
	   .ZN (_263_),
	   .A2 (_173_),
	   .A1 (_262_) );
   INV_X1 _568_ (
	   .ZN (_262_),
	   .A (_258_) );
   OAI21_X1 _567_ (
	   .ZN (_261_),
	   .B2 (_159_),
	   .B1 (_165_),
	   .A (_379_) );
   MUX2_X1 _566_ (
	   .Z (_084_),
	   .S (_249_),
	   .B (_260_),
	   .A (_118_) );
   OAI211_X1 _565_ (
	   .ZN (_260_),
	   .C2 (_062_),
	   .C1 (_245_),
	   .B (_259_),
	   .A (_257_) );
   NAND2_X1 _564_ (
	   .ZN (_259_),
	   .A2 (_412_),
	   .A1 (_253_) );
   XNOR2_X1 _563_ (
	   .ZN (_412_),
	   .B (_173_),
	   .A (_258_) );
   AOI21_X1 _562_ (
	   .ZN (_258_),
	   .B2 (_254_),
	   .B1 (_239_),
	   .A (_180_) );
   OAI21_X1 _561_ (
	   .ZN (_257_),
	   .B2 (_159_),
	   .B1 (_165_),
	   .A (_378_) );
   MUX2_X1 _560_ (
	   .Z (_083_),
	   .S (_249_),
	   .B (_256_),
	   .A (_117_) );
   OAI211_X1 _559_ (
	   .ZN (_256_),
	   .C2 (_061_),
	   .C1 (_245_),
	   .B (_255_),
	   .A (_250_) );
   NAND2_X1 _558_ (
	   .ZN (_255_),
	   .A2 (_411_),
	   .A1 (_253_) );
   XOR2_X1 _557_ (
	   .Z (_411_),
	   .B (_254_),
	   .A (_239_) );
   NAND2_X1 _556_ (
	   .ZN (_254_),
	   .A2 (_126_),
	   .A1 (_182_) );
   CLKBUF_X2 _555_ (
	   .Z (_253_),
	   .A (_252_) );
   NOR2_X2 _554_ (
	   .ZN (_252_),
	   .A2 (_251_),
	   .A1 (_242_) );
   INV_X1 _553_ (
	   .ZN (_251_),
	   .A (_230_) );
   OAI21_X1 _552_ (
	   .ZN (_250_),
	   .B2 (_159_),
	   .B1 (_165_),
	   .A (_377_) );
   MUX2_X1 _551_ (
	   .Z (_076_),
	   .S (_249_),
	   .B (_246_),
	   .A (_110_) );
   BUF_X2 _550_ (
	   .Z (_249_),
	   .A (_248_) );
   BUF_X2 _549_ (
	   .Z (_248_),
	   .A (_247_) );
   OR2_X1 _548_ (
	   .ZN (_247_),
	   .A2 (_401_),
	   .A1 (_109_) );
   OAI211_X1 _547_ (
	   .ZN (_246_),
	   .C2 (_060_),
	   .C1 (_245_),
	   .B (_236_),
	   .A (_166_) );
   BUF_X2 _546_ (
	   .Z (_245_),
	   .A (_244_) );
   OR2_X2 _545_ (
	   .ZN (_244_),
	   .A2 (_158_),
	   .A1 (_243_) );
   NAND2_X1 _544_ (
	   .ZN (_243_),
	   .A2 (_109_),
	   .A1 (_242_) );
   AOI21_X1 _543_ (
	   .ZN (_242_),
	   .B2 (_235_),
	   .B1 (_229_),
	   .A (_241_) );
   NOR3_X1 _542_ (
	   .ZN (_241_),
	   .A3 (_240_),
	   .A2 (_404_),
	   .A1 (_238_) );
   INV_X1 _541_ (
	   .ZN (_240_),
	   .A (_239_) );
   XNOR2_X2 _540_ (
	   .ZN (_239_),
	   .B (_133_),
	   .A (_117_) );
   NAND4_X1 _539_ (
	   .ZN (_238_),
	   .A4 (_174_),
	   .A3 (_213_),
	   .A2 (_237_),
	   .A1 (_205_) );
   AND2_X1 _538_ (
	   .ZN (_237_),
	   .A2 (_177_),
	   .A1 (_171_) );
   NAND4_X1 _537_ (
	   .ZN (_236_),
	   .A4 (_235_),
	   .A3 (_230_),
	   .A2 (_404_),
	   .A1 (_229_) );
   OR3_X1 _536_ (
	   .ZN (_235_),
	   .A3 (_234_),
	   .A2 (_232_),
	   .A1 (_208_) );
   AOI22_X1 _535_ (
	   .ZN (_234_),
	   .B2 (_129_),
	   .B1 (_233_),
	   .A2 (_130_),
	   .A1 (_231_) );
   INV_X1 _534_ (
	   .ZN (_233_),
	   .A (_113_) );
   NOR2_X1 _533_ (
	   .ZN (_232_),
	   .A2 (_130_),
	   .A1 (_231_) );
   INV_X1 _532_ (
	   .ZN (_231_),
	   .A (_114_) );
   AND2_X1 _531_ (
	   .ZN (_230_),
	   .A2 (_059_),
	   .A1 (_109_) );
   AND4_X1 _530_ (
	   .ZN (_229_),
	   .A4 (_228_),
	   .A3 (_226_),
	   .A2 (_215_),
	   .A1 (_168_) );
   NAND3_X1 _529_ (
	   .ZN (_228_),
	   .A3 (_131_),
	   .A2 (_227_),
	   .A1 (_207_) );
   INV_X1 _528_ (
	   .ZN (_227_),
	   .A (_115_) );
   NAND2_X1 _527_ (
	   .ZN (_226_),
	   .A2 (_213_),
	   .A1 (_225_) );
   OAI21_X1 _526_ (
	   .ZN (_225_),
	   .B2 (_224_),
	   .B1 (_222_),
	   .A (_220_) );
   AOI22_X1 _525_ (
	   .ZN (_224_),
	   .B2 (_127_),
	   .B1 (_223_),
	   .A2 (_128_),
	   .A1 (_221_) );
   INV_X1 _524_ (
	   .ZN (_223_),
	   .A (_111_) );
   NOR2_X1 _523_ (
	   .ZN (_222_),
	   .A2 (_128_),
	   .A1 (_221_) );
   INV_X1 _522_ (
	   .ZN (_221_),
	   .A (_112_) );
   OAI21_X1 _521_ (
	   .ZN (_220_),
	   .B2 (_219_),
	   .B1 (_217_),
	   .A (_202_) );
   AND2_X1 _520_ (
	   .ZN (_219_),
	   .A2 (_141_),
	   .A1 (_218_) );
   INV_X1 _519_ (
	   .ZN (_218_),
	   .A (_125_) );
   AND3_X1 _518_ (
	   .ZN (_217_),
	   .A3 (_140_),
	   .A2 (_216_),
	   .A1 (_203_) );
   INV_X1 _517_ (
	   .ZN (_216_),
	   .A (_124_) );
   NAND2_X1 _516_ (
	   .ZN (_215_),
	   .A2 (_214_),
	   .A1 (_199_) );
   AND2_X1 _515_ (
	   .ZN (_214_),
	   .A2 (_213_),
	   .A1 (_205_) );
   NOR3_X1 _514_ (
	   .ZN (_213_),
	   .A3 (_212_),
	   .A2 (_210_),
	   .A1 (_208_) );
   INV_X1 _513_ (
	   .ZN (_212_),
	   .A (_211_) );
   XNOR2_X1 _512_ (
	   .ZN (_211_),
	   .B (_129_),
	   .A (_113_) );
   INV_X1 _511_ (
	   .ZN (_210_),
	   .A (_209_) );
   XNOR2_X2 _510_ (
	   .ZN (_209_),
	   .B (_130_),
	   .A (_114_) );
   NAND2_X1 _509_ (
	   .ZN (_208_),
	   .A2 (_207_),
	   .A1 (_206_) );
   XNOR2_X2 _508_ (
	   .ZN (_207_),
	   .B (_132_),
	   .A (_116_) );
   XNOR2_X1 _507_ (
	   .ZN (_206_),
	   .B (_131_),
	   .A (_115_) );
   AND3_X1 _506_ (
	   .ZN (_205_),
	   .A3 (_204_),
	   .A2 (_203_),
	   .A1 (_202_) );
   XNOR2_X1 _505_ (
	   .ZN (_204_),
	   .B (_140_),
	   .A (_124_) );
   XNOR2_X2 _504_ (
	   .ZN (_203_),
	   .B (_141_),
	   .A (_125_) );
   AND2_X1 _503_ (
	   .ZN (_202_),
	   .A2 (_201_),
	   .A1 (_200_) );
   XNOR2_X1 _502_ (
	   .ZN (_201_),
	   .B (_128_),
	   .A (_112_) );
   XNOR2_X1 _501_ (
	   .ZN (_200_),
	   .B (_127_),
	   .A (_111_) );
   NAND3_X1 _500_ (
	   .ZN (_199_),
	   .A3 (_198_),
	   .A2 (_195_),
	   .A1 (_184_) );
   OAI211_X1 _499_ (
	   .ZN (_198_),
	   .C2 (_197_),
	   .C1 (_196_),
	   .B (_177_),
	   .A (_171_) );
   AOI211_X1 _498_ (
	   .ZN (_197_),
	   .C2 (_144_),
	   .C1 (_119_),
	   .B (_145_),
	   .A (_118_) );
   NOR2_X1 _497_ (
	   .ZN (_196_),
	   .A2 (_119_),
	   .A1 (_144_) );
   AND3_X1 _496_ (
	   .ZN (_195_),
	   .A3 (_194_),
	   .A2 (_192_),
	   .A1 (_189_) );
   NAND3_X1 _495_ (
	   .ZN (_194_),
	   .A3 (_138_),
	   .A2 (_193_),
	   .A1 (_169_) );
   INV_X1 _494_ (
	   .ZN (_193_),
	   .A (_122_) );
   INV_X1 _493_ (
	   .ZN (_192_),
	   .A (_191_) );
   NOR2_X1 _492_ (
	   .ZN (_191_),
	   .A2 (_123_),
	   .A1 (_190_) );
   INV_X1 _491_ (
	   .ZN (_190_),
	   .A (_139_) );
   OAI21_X1 _490_ (
	   .ZN (_189_),
	   .B2 (_188_),
	   .B1 (_186_),
	   .A (_171_) );
   AND2_X1 _489_ (
	   .ZN (_188_),
	   .A2 (_137_),
	   .A1 (_187_) );
   INV_X1 _488_ (
	   .ZN (_187_),
	   .A (_121_) );
   AND3_X1 _487_ (
	   .ZN (_186_),
	   .A3 (_136_),
	   .A2 (_185_),
	   .A1 (_175_) );
   INV_X1 _486_ (
	   .ZN (_185_),
	   .A (_120_) );
   OR3_X1 _485_ (
	   .ZN (_184_),
	   .A3 (_183_),
	   .A2 (_180_),
	   .A1 (_178_) );
   NOR3_X1 _484_ (
	   .ZN (_183_),
	   .A3 (_126_),
	   .A2 (_182_),
	   .A1 (_181_) );
   INV_X1 _483_ (
	   .ZN (_182_),
	   .A (_110_) );
   NOR2_X1 _482_ (
	   .ZN (_181_),
	   .A2 (_117_),
	   .A1 (_179_) );
   AND2_X1 _481_ (
	   .ZN (_180_),
	   .A2 (_117_),
	   .A1 (_179_) );
   INV_X1 _480_ (
	   .ZN (_179_),
	   .A (_133_) );
   NAND3_X1 _479_ (
	   .ZN (_178_),
	   .A3 (_177_),
	   .A2 (_174_),
	   .A1 (_171_) );
   AND2_X1 _478_ (
	   .ZN (_177_),
	   .A2 (_176_),
	   .A1 (_175_) );
   XNOR2_X1 _477_ (
	   .ZN (_176_),
	   .B (_136_),
	   .A (_120_) );
   XNOR2_X2 _476_ (
	   .ZN (_175_),
	   .B (_137_),
	   .A (_121_) );
   AND2_X1 _475_ (
	   .ZN (_174_),
	   .A2 (_173_),
	   .A1 (_172_) );
   XNOR2_X1 _474_ (
	   .ZN (_173_),
	   .B (_134_),
	   .A (_118_) );
   XNOR2_X1 _473_ (
	   .ZN (_172_),
	   .B (_135_),
	   .A (_119_) );
   AND2_X1 _472_ (
	   .ZN (_171_),
	   .A2 (_170_),
	   .A1 (_169_) );
   XNOR2_X1 _471_ (
	   .ZN (_170_),
	   .B (_138_),
	   .A (_122_) );
   XNOR2_X2 _470_ (
	   .ZN (_169_),
	   .B (_139_),
	   .A (_123_) );
   NAND2_X1 _469_ (
	   .ZN (_168_),
	   .A2 (_132_),
	   .A1 (_167_) );
   INV_X1 _468_ (
	   .ZN (_167_),
	   .A (_116_) );
   OAI21_X1 _467_ (
	   .ZN (_166_),
	   .B2 (_159_),
	   .B1 (_165_),
	   .A (_376_) );
   BUF_X2 _466_ (
	   .Z (_165_),
	   .A (_142_) );
   OR3_X1 _465_ (
	   .ZN (_054_),
	   .A3 (_164_),
	   .A2 (_403_),
	   .A1 (_163_) );
   AOI211_X1 _464_ (
	   .ZN (_164_),
	   .C2 (_402_),
	   .C1 (_160_),
	   .B (_059_),
	   .A (_403_) );
   NOR2_X1 _463_ (
	   .ZN (_163_),
	   .A2 (_057_),
	   .A1 (_162_) );
   NAND3_X1 _462_ (
	   .ZN (_162_),
	   .A3 (_420_),
	   .A2 (_152_),
	   .A1 (_421_) );
   NAND2_X1 _461_ (
	   .ZN (_056_),
	   .A2 (_161_),
	   .A1 (_157_) );
   NAND4_X1 _460_ (
	   .ZN (_161_),
	   .A4 (_402_),
	   .A3 (_160_),
	   .A2 (_159_),
	   .A1 (_152_) );
   BUF_X2 _459_ (
	   .Z (_160_),
	   .A (_401_) );
   BUF_X2 _458_ (
	   .Z (_159_),
	   .A (_158_) );
   INV_X2 _457_ (
	   .ZN (_158_),
	   .A (_059_) );
   OAI211_X1 _456_ (
	   .ZN (_157_),
	   .C2 (_150_),
	   .C1 (_147_),
	   .B (_153_),
	   .A (_152_) );
   NAND2_X1 _455_ (
	   .ZN (_055_),
	   .A2 (_156_),
	   .A1 (_154_) );
   OR3_X1 _454_ (
	   .ZN (_156_),
	   .A3 (_057_),
	   .A2 (_403_),
	   .A1 (_155_) );
   AND2_X1 _453_ (
	   .ZN (_155_),
	   .A2 (_420_),
	   .A1 (_421_) );
   NAND3_X1 _452_ (
	   .ZN (_154_),
	   .A3 (_153_),
	   .A2 (_152_),
	   .A1 (_151_) );
   INV_X1 _451_ (
	   .ZN (_153_),
	   .A (_058_) );
   INV_X1 _450_ (
	   .ZN (_152_),
	   .A (_403_) );
   NOR2_X1 _449_ (
	   .ZN (_151_),
	   .A2 (_150_),
	   .A1 (_147_) );
   NAND2_X1 _448_ (
	   .ZN (_150_),
	   .A2 (_149_),
	   .A1 (_148_) );
   NOR4_X1 _447_ (
	   .ZN (_149_),
	   .A4 (_129_),
	   .A3 (_130_),
	   .A2 (_131_),
	   .A1 (_132_) );
   NOR4_X1 _446_ (
	   .ZN (_148_),
	   .A4 (_140_),
	   .A3 (_141_),
	   .A2 (_127_),
	   .A1 (_128_) );
   NAND4_X1 _445_ (
	   .ZN (_147_),
	   .A4 (_146_),
	   .A3 (_145_),
	   .A2 (_144_),
	   .A1 (_143_) );
   NOR2_X1 _444_ (
	   .ZN (_146_),
	   .A2 (_126_),
	   .A1 (_133_) );
   INV_X1 _443_ (
	   .ZN (_145_),
	   .A (_134_) );
   INV_X1 _442_ (
	   .ZN (_144_),
	   .A (_135_) );
   NOR4_X1 _441_ (
	   .ZN (_143_),
	   .A4 (_136_),
	   .A3 (_137_),
	   .A2 (_138_),
	   .A1 (_139_) );
   XOR2_X1 _440_ (
	   .Z (_404_),
	   .B (_126_),
	   .A (_110_) );
   AND3_X1 _439_ (
	   .ZN (_421_),
	   .A3 (_059_),
	   .A2 (_108_),
	   .A1 (_142_) );
   INV_X2 _438_ (
	   .ZN (_142_),
	   .A (_109_) );
endmodule

