// Used to silence warnings.
module TAPCELL_ASAP7_75t_R ();
  // silence eqy
  wire dummy_wire;
  assign dummy_wire = 1'b0;
endmodule
module FILLERxp5_ASAP7_75t_R;
  // silence eqy
  wire dummy_wire;
  assign dummy_wire = 1'b0;
endmodule
module FILLER_ASAP7_75t_R ();
  // silence eqy
  wire dummy_wire;
  assign dummy_wire = 1'b0;
endmodule
module DECAPx1_ASAP7_75t_R ();
  // silence eqy
  wire dummy_wire;
  assign dummy_wire = 1'b0;
endmodule
module DECAPx2_ASAP7_75t_R ();
  // silence eqy
  wire dummy_wire;
  assign dummy_wire = 1'b0;
endmodule
module DECAPx4_ASAP7_75t_R ();
  // silence eqy
  wire dummy_wire;
  assign dummy_wire = 1'b0;
endmodule
module DECAPx6_ASAP7_75t_R ();
  // silence eqy
  wire dummy_wire;
  assign dummy_wire = 1'b0;
endmodule
module DECAPx10_ASAP7_75t_R ();
  // silence eqy
  wire dummy_wire;
  assign dummy_wire = 1'b0;
endmodule
