VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 2000 ;
END UNITS

MACRO ENDCAP_X1_TOPEDGE
  PROPERTY LEF58_CLASS " CLASS ENDCAP TOPEDGE ; " ;
  ORIGIN 0 0 ;
  FOREIGN ENDCAP_X1_TOPEDGE 0 0 ;
  SIZE 0.19 BY 1.4 ;
  SYMMETRY X ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.19 1.485 ;
        RECT 0.06 0.975 0.13 1.315 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.19 0.085 ;
        RECT 0.06 0.085 0.13 0.425 ;
    END
  END VSS
END ENDCAP_X1_TOPEDGE
MACRO ENDCAP_X1_BOTTOMEDGE
  PROPERTY LEF58_CLASS " CLASS ENDCAP BOTTOMEDGE ; " ;
  ORIGIN 0 0 ;
  FOREIGN ENDCAP_X1_BOTTOMEDGE 0 0 ;
  SIZE 0.19 BY 1.4 ;
  SYMMETRY X ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.19 1.485 ;
        RECT 0.06 0.975 0.13 1.315 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.19 0.085 ;
        RECT 0.06 0.085 0.13 0.425 ;
    END
  END VSS
END ENDCAP_X1_BOTTOMEDGE

MACRO ENDCAP_X4_RIGHTTOPCORNER
  PROPERTY LEF58_CLASS " CLASS ENDCAP RIGHTTOPCORNER ; " ;
  ORIGIN 0 0 ;
  FOREIGN ENDCAP_X4 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.76 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.76 0.085 ;
    END
  END VSS
END ENDCAP_X4_RIGHTTOPCORNER

MACRO ENDCAP_X4_RIGHTBOTTOMCORNER
  PROPERTY LEF58_CLASS " CLASS ENDCAP RIGHTBOTTOMCORNER ; " ;
  ORIGIN 0 0 ;
  FOREIGN ENDCAP_X4 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.76 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.76 0.085 ;
    END
  END VSS
END ENDCAP_X4_RIGHTBOTTOMCORNER
MACRO ENDCAP_X4_LEFTBOTTOMCORNER
  PROPERTY LEF58_CLASS " CLASS ENDCAP LEFTBOTTOMCORNER ; " ;
  ORIGIN 0 0 ;
  FOREIGN ENDCAP_X4 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.76 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.76 0.085 ;
    END
  END VSS
END ENDCAP_X4_LEFTBOTTOMCORNER
MACRO ENDCAP_X4_RIGHTTOPCORNER
  PROPERTY LEF58_CLASS " CLASS ENDCAP RIGHTTOPCORNER ; " ;
  ORIGIN 0 0 ;
  FOREIGN ENDCAP_X4 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.76 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.76 0.085 ;
    END
  END VSS
END ENDCAP_X4_RIGHTTOPCORNER
MACRO ENDCAP_X4_LEFTTOPCORNER
  PROPERTY LEF58_CLASS " CLASS ENDCAP LEFTTOPCORNER ; " ;
  ORIGIN 0 0 ;
  FOREIGN ENDCAP_X4 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.76 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.76 0.085 ;
    END
  END VSS
END ENDCAP_X4_LEFTTOPCORNER

MACRO ENDCAP_X4_RIGHTBOTTOMEDGE
  PROPERTY LEF58_CLASS " CLASS ENDCAP RIGHTBOTTOMEDGE ; " ;
  ORIGIN 0 0 ;
  FOREIGN ENDCAP_X4 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.76 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.76 0.085 ;
    END
  END VSS
END ENDCAP_X4_RIGHTBOTTOMEDGE
MACRO ENDCAP_X4_LEFTBOTTOMEDGE
  PROPERTY LEF58_CLASS " CLASS ENDCAP LEFTBOTTOMEDGE ; " ;
  ORIGIN 0 0 ;
  FOREIGN ENDCAP_X4 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.76 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.76 0.085 ;
    END
  END VSS
END ENDCAP_X4_LEFTBOTTOMEDGE
MACRO ENDCAP_X4_RIGHTTOPEDGE
  PROPERTY LEF58_CLASS " CLASS ENDCAP RIGHTTOPEDGE ; " ;
  ORIGIN 0 0 ;
  FOREIGN ENDCAP_X4 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.76 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.76 0.085 ;
    END
  END VSS
END ENDCAP_X4_RIGHTTOPEDGE
MACRO ENDCAP_X4_LEFTTOPEDGE
  PROPERTY LEF58_CLASS " CLASS ENDCAP LEFTTOPEDGE ; " ;
  ORIGIN 0 0 ;
  FOREIGN ENDCAP_X4 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.76 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.76 0.085 ;
    END
  END VSS
END ENDCAP_X4_LEFTTOPEDGE

MACRO ENDCAP_X4_RIGHTEDGE
  PROPERTY LEF58_CLASS " CLASS ENDCAP RIGHTEDGE ; " ;
  ORIGIN 0 0 ;
  FOREIGN ENDCAP_X4 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.76 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.76 0.085 ;
    END
  END VSS
END ENDCAP_X4_RIGHTEDGE
MACRO ENDCAP_X4_LEFTEDGE
  PROPERTY LEF58_CLASS " CLASS ENDCAP LEFTEDGE ; " ;
  ORIGIN 0 0 ;
  FOREIGN ENDCAP_X4 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.76 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.76 0.085 ;
    END
  END VSS
END ENDCAP_X4_LEFTEDGE

END LIBRARY
#
# End of file
#
