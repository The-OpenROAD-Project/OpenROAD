VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO HM_100x400_4x4
  CLASS BLOCK ;
  FOREIGN HM_100x400_4x4 0 0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SIZE 100 BY 400 ;
  PIN I1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 0 200 1 201  ;
    END
  END I1
  PIN I2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 0 210 1 211  ;
    END
  END I2 
  PIN I3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 0 220 1 221  ;
    END
  END I3 
  PIN I4
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 0 230 1 231  ;
    END
  END I4 
  PIN O1 
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 99 200 100 201  ;
    END
  END O1 
  PIN O2 
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 99 210 100 211  ;
    END
  END O2 
  PIN O3 
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 99 220 100 221  ;
    END
  END O3 
  PIN O4 
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 99 230 100 231  ;
    END
  END O4
  OBS
      LAYER metal1 ;
        POLYGON 0.235 0.84 0.47 0.84 0.47 0.46 0.045 0.46 0.045 0.19 0.115 0.19 0.115 0.39 0.54 0.39 0.54 0.91 0.305 0.91 0.305 1.25 0.235 1.25  ;
  END
END HM_100x400_4x4 

MACRO HM_100x100_1x1
  CLASS BLOCK ;
  FOREIGN HM_100x100_1x1 0 0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SIZE 100 BY 100 ;
  PIN I1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 0 50 1 51  ;
    END
  END I1
  PIN O1 
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 99 50 100 51  ;
    END
  END O1 
  OBS
      LAYER metal1 ;
        POLYGON 0.235 0.84 0.47 0.84 0.47 0.46 0.045 0.46 0.045 0.19 0.115 0.19 0.115 0.39 0.54 0.39 0.54 0.91 0.305 0.91 0.305 1.25 0.235 1.25  ;
  END
END HM_100x100_1x1 

SITE SingleHeightSite
  SYMMETRY y ;
  CLASS core ;
  SIZE 0.19 BY 1.4 ;
END SingleHeightSite

SITE DoubleHeightSite
  SYMMETRY y ;
  CLASS core ;
  SIZE 0.19 BY 2.8 ;
END DoubleHeightSite


site TripleHeightSite
  SYMMETRY y ;
  CLASS core ;
  SIZE 0.19 BY 4.2 ;
END TripleHeightSite

MACRO MOCK_DOUBLE
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2_X1 0 0 ;
  SIZE 0.76 BY 2.8 ;
  SYMMETRY X Y ;
  SITE DoubleHeightSite ;
  PIN A1 
  END A1
  PIN A2 
  END A2
  PIN ZN 
  END ZN
  PIN VDD 
  END VDD
  PIN VSS 
  END VSS
END MOCK_DOUBLE

MACRO MOCK_TRIPLE
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2_X1 0 0 ;
  SIZE 0.76 BY 4.2 ;
  SYMMETRY X Y ;
  SITE TripleHeightSite ;
  PIN A1 
  END A1
  PIN A2 
  END A2
  PIN ZN 
  END ZN
  PIN VDD 
  END VDD
  PIN VSS 
  END VSS
END MOCK_TRIPLE

MACRO MOCK_SINGLE
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2_X1 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X Y ;
  SITE SingleHeightSite ;
  PIN A1 
  END A1
  PIN A2 
  END A2
  PIN ZN 
  END ZN
  PIN VDD 
  END VDD
  PIN VSS 
  END VSS
END MOCK_SINGLE
