VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 2000 ;
END UNITS

MANUFACTURINGGRID 0.0050 ;

SITE FreePDK45_38x28_10R_NP_162NW_34O_DoubleHeight
  SYMMETRY y ;
  CLASS core ;
  SIZE 0.19 BY 2.8 ;
END FreePDK45_38x28_10R_NP_162NW_34O_DoubleHeight
