VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram7_256x32
  FOREIGN fakeram7_256x32 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 4.180 BY 67.200 ;
  CLASS BLOCK ;
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.048 0.024 0.072 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.912 0.024 0.936 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.776 0.024 1.800 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.640 0.024 2.664 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.504 0.024 3.528 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.368 0.024 4.392 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.232 0.024 5.256 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.096 0.024 6.120 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.960 0.024 6.984 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.824 0.024 7.848 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.688 0.024 8.712 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.552 0.024 9.576 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.416 0.024 10.440 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.280 0.024 11.304 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.144 0.024 12.168 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.008 0.024 13.032 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.872 0.024 13.896 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.736 0.024 14.760 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 15.600 0.024 15.624 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.464 0.024 16.488 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 17.328 0.024 17.352 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.192 0.024 18.216 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.056 0.024 19.080 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.920 0.024 19.944 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.784 0.024 20.808 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.648 0.024 21.672 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.512 0.024 22.536 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.376 0.024 23.400 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 24.240 0.024 24.264 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 25.104 0.024 25.128 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 25.968 0.024 25.992 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 26.832 0.024 26.856 ;
    END
  END rd_out[31]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 27.408 0.024 27.432 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 28.272 0.024 28.296 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 29.136 0.024 29.160 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 30.000 0.024 30.024 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 30.864 0.024 30.888 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 31.728 0.024 31.752 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 32.592 0.024 32.616 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 33.456 0.024 33.480 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 34.320 0.024 34.344 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 35.184 0.024 35.208 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 36.048 0.024 36.072 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 36.912 0.024 36.936 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 37.776 0.024 37.800 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 38.640 0.024 38.664 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 39.504 0.024 39.528 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 40.368 0.024 40.392 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 41.232 0.024 41.256 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 42.096 0.024 42.120 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 42.960 0.024 42.984 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 43.824 0.024 43.848 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 44.688 0.024 44.712 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 45.552 0.024 45.576 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 46.416 0.024 46.440 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 47.280 0.024 47.304 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 48.144 0.024 48.168 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 49.008 0.024 49.032 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 49.872 0.024 49.896 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 50.736 0.024 50.760 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 51.600 0.024 51.624 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 52.464 0.024 52.488 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 53.328 0.024 53.352 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 54.192 0.024 54.216 ;
    END
  END wd_in[31]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 54.768 0.024 54.792 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 55.632 0.024 55.656 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 56.496 0.024 56.520 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 57.360 0.024 57.384 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 58.224 0.024 58.248 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 59.088 0.024 59.112 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 59.952 0.024 59.976 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 60.816 0.024 60.840 ;
    END
  END addr_in[7]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 61.392 0.024 61.416 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 62.256 0.024 62.280 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 63.120 0.024 63.144 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 0.048 0.000 4.132 0.096 ;
      RECT 0.048 0.768 4.132 0.864 ;
      RECT 0.048 1.536 4.132 1.632 ;
      RECT 0.048 2.304 4.132 2.400 ;
      RECT 0.048 3.072 4.132 3.168 ;
      RECT 0.048 3.840 4.132 3.936 ;
      RECT 0.048 4.608 4.132 4.704 ;
      RECT 0.048 5.376 4.132 5.472 ;
      RECT 0.048 6.144 4.132 6.240 ;
      RECT 0.048 6.912 4.132 7.008 ;
      RECT 0.048 7.680 4.132 7.776 ;
      RECT 0.048 8.448 4.132 8.544 ;
      RECT 0.048 9.216 4.132 9.312 ;
      RECT 0.048 9.984 4.132 10.080 ;
      RECT 0.048 10.752 4.132 10.848 ;
      RECT 0.048 11.520 4.132 11.616 ;
      RECT 0.048 12.288 4.132 12.384 ;
      RECT 0.048 13.056 4.132 13.152 ;
      RECT 0.048 13.824 4.132 13.920 ;
      RECT 0.048 14.592 4.132 14.688 ;
      RECT 0.048 15.360 4.132 15.456 ;
      RECT 0.048 16.128 4.132 16.224 ;
      RECT 0.048 16.896 4.132 16.992 ;
      RECT 0.048 17.664 4.132 17.760 ;
      RECT 0.048 18.432 4.132 18.528 ;
      RECT 0.048 19.200 4.132 19.296 ;
      RECT 0.048 19.968 4.132 20.064 ;
      RECT 0.048 20.736 4.132 20.832 ;
      RECT 0.048 21.504 4.132 21.600 ;
      RECT 0.048 22.272 4.132 22.368 ;
      RECT 0.048 23.040 4.132 23.136 ;
      RECT 0.048 23.808 4.132 23.904 ;
      RECT 0.048 24.576 4.132 24.672 ;
      RECT 0.048 25.344 4.132 25.440 ;
      RECT 0.048 26.112 4.132 26.208 ;
      RECT 0.048 26.880 4.132 26.976 ;
      RECT 0.048 27.648 4.132 27.744 ;
      RECT 0.048 28.416 4.132 28.512 ;
      RECT 0.048 29.184 4.132 29.280 ;
      RECT 0.048 29.952 4.132 30.048 ;
      RECT 0.048 30.720 4.132 30.816 ;
      RECT 0.048 31.488 4.132 31.584 ;
      RECT 0.048 32.256 4.132 32.352 ;
      RECT 0.048 33.024 4.132 33.120 ;
      RECT 0.048 33.792 4.132 33.888 ;
      RECT 0.048 34.560 4.132 34.656 ;
      RECT 0.048 35.328 4.132 35.424 ;
      RECT 0.048 36.096 4.132 36.192 ;
      RECT 0.048 36.864 4.132 36.960 ;
      RECT 0.048 37.632 4.132 37.728 ;
      RECT 0.048 38.400 4.132 38.496 ;
      RECT 0.048 39.168 4.132 39.264 ;
      RECT 0.048 39.936 4.132 40.032 ;
      RECT 0.048 40.704 4.132 40.800 ;
      RECT 0.048 41.472 4.132 41.568 ;
      RECT 0.048 42.240 4.132 42.336 ;
      RECT 0.048 43.008 4.132 43.104 ;
      RECT 0.048 43.776 4.132 43.872 ;
      RECT 0.048 44.544 4.132 44.640 ;
      RECT 0.048 45.312 4.132 45.408 ;
      RECT 0.048 46.080 4.132 46.176 ;
      RECT 0.048 46.848 4.132 46.944 ;
      RECT 0.048 47.616 4.132 47.712 ;
      RECT 0.048 48.384 4.132 48.480 ;
      RECT 0.048 49.152 4.132 49.248 ;
      RECT 0.048 49.920 4.132 50.016 ;
      RECT 0.048 50.688 4.132 50.784 ;
      RECT 0.048 51.456 4.132 51.552 ;
      RECT 0.048 52.224 4.132 52.320 ;
      RECT 0.048 52.992 4.132 53.088 ;
      RECT 0.048 53.760 4.132 53.856 ;
      RECT 0.048 54.528 4.132 54.624 ;
      RECT 0.048 55.296 4.132 55.392 ;
      RECT 0.048 56.064 4.132 56.160 ;
      RECT 0.048 56.832 4.132 56.928 ;
      RECT 0.048 57.600 4.132 57.696 ;
      RECT 0.048 58.368 4.132 58.464 ;
      RECT 0.048 59.136 4.132 59.232 ;
      RECT 0.048 59.904 4.132 60.000 ;
      RECT 0.048 60.672 4.132 60.768 ;
      RECT 0.048 61.440 4.132 61.536 ;
      RECT 0.048 62.208 4.132 62.304 ;
      RECT 0.048 62.976 4.132 63.072 ;
      RECT 0.048 63.744 4.132 63.840 ;
      RECT 0.048 64.512 4.132 64.608 ;
      RECT 0.048 65.280 4.132 65.376 ;
      RECT 0.048 66.048 4.132 66.144 ;
      RECT 0.048 66.816 4.132 66.912 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.048 0.384 4.132 0.480 ;
      RECT 0.048 1.152 4.132 1.248 ;
      RECT 0.048 1.920 4.132 2.016 ;
      RECT 0.048 2.688 4.132 2.784 ;
      RECT 0.048 3.456 4.132 3.552 ;
      RECT 0.048 4.224 4.132 4.320 ;
      RECT 0.048 4.992 4.132 5.088 ;
      RECT 0.048 5.760 4.132 5.856 ;
      RECT 0.048 6.528 4.132 6.624 ;
      RECT 0.048 7.296 4.132 7.392 ;
      RECT 0.048 8.064 4.132 8.160 ;
      RECT 0.048 8.832 4.132 8.928 ;
      RECT 0.048 9.600 4.132 9.696 ;
      RECT 0.048 10.368 4.132 10.464 ;
      RECT 0.048 11.136 4.132 11.232 ;
      RECT 0.048 11.904 4.132 12.000 ;
      RECT 0.048 12.672 4.132 12.768 ;
      RECT 0.048 13.440 4.132 13.536 ;
      RECT 0.048 14.208 4.132 14.304 ;
      RECT 0.048 14.976 4.132 15.072 ;
      RECT 0.048 15.744 4.132 15.840 ;
      RECT 0.048 16.512 4.132 16.608 ;
      RECT 0.048 17.280 4.132 17.376 ;
      RECT 0.048 18.048 4.132 18.144 ;
      RECT 0.048 18.816 4.132 18.912 ;
      RECT 0.048 19.584 4.132 19.680 ;
      RECT 0.048 20.352 4.132 20.448 ;
      RECT 0.048 21.120 4.132 21.216 ;
      RECT 0.048 21.888 4.132 21.984 ;
      RECT 0.048 22.656 4.132 22.752 ;
      RECT 0.048 23.424 4.132 23.520 ;
      RECT 0.048 24.192 4.132 24.288 ;
      RECT 0.048 24.960 4.132 25.056 ;
      RECT 0.048 25.728 4.132 25.824 ;
      RECT 0.048 26.496 4.132 26.592 ;
      RECT 0.048 27.264 4.132 27.360 ;
      RECT 0.048 28.032 4.132 28.128 ;
      RECT 0.048 28.800 4.132 28.896 ;
      RECT 0.048 29.568 4.132 29.664 ;
      RECT 0.048 30.336 4.132 30.432 ;
      RECT 0.048 31.104 4.132 31.200 ;
      RECT 0.048 31.872 4.132 31.968 ;
      RECT 0.048 32.640 4.132 32.736 ;
      RECT 0.048 33.408 4.132 33.504 ;
      RECT 0.048 34.176 4.132 34.272 ;
      RECT 0.048 34.944 4.132 35.040 ;
      RECT 0.048 35.712 4.132 35.808 ;
      RECT 0.048 36.480 4.132 36.576 ;
      RECT 0.048 37.248 4.132 37.344 ;
      RECT 0.048 38.016 4.132 38.112 ;
      RECT 0.048 38.784 4.132 38.880 ;
      RECT 0.048 39.552 4.132 39.648 ;
      RECT 0.048 40.320 4.132 40.416 ;
      RECT 0.048 41.088 4.132 41.184 ;
      RECT 0.048 41.856 4.132 41.952 ;
      RECT 0.048 42.624 4.132 42.720 ;
      RECT 0.048 43.392 4.132 43.488 ;
      RECT 0.048 44.160 4.132 44.256 ;
      RECT 0.048 44.928 4.132 45.024 ;
      RECT 0.048 45.696 4.132 45.792 ;
      RECT 0.048 46.464 4.132 46.560 ;
      RECT 0.048 47.232 4.132 47.328 ;
      RECT 0.048 48.000 4.132 48.096 ;
      RECT 0.048 48.768 4.132 48.864 ;
      RECT 0.048 49.536 4.132 49.632 ;
      RECT 0.048 50.304 4.132 50.400 ;
      RECT 0.048 51.072 4.132 51.168 ;
      RECT 0.048 51.840 4.132 51.936 ;
      RECT 0.048 52.608 4.132 52.704 ;
      RECT 0.048 53.376 4.132 53.472 ;
      RECT 0.048 54.144 4.132 54.240 ;
      RECT 0.048 54.912 4.132 55.008 ;
      RECT 0.048 55.680 4.132 55.776 ;
      RECT 0.048 56.448 4.132 56.544 ;
      RECT 0.048 57.216 4.132 57.312 ;
      RECT 0.048 57.984 4.132 58.080 ;
      RECT 0.048 58.752 4.132 58.848 ;
      RECT 0.048 59.520 4.132 59.616 ;
      RECT 0.048 60.288 4.132 60.384 ;
      RECT 0.048 61.056 4.132 61.152 ;
      RECT 0.048 61.824 4.132 61.920 ;
      RECT 0.048 62.592 4.132 62.688 ;
      RECT 0.048 63.360 4.132 63.456 ;
      RECT 0.048 64.128 4.132 64.224 ;
      RECT 0.048 64.896 4.132 64.992 ;
      RECT 0.048 65.664 4.132 65.760 ;
      RECT 0.048 66.432 4.132 66.528 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 4.180 67.200 ;
    LAYER M2 ;
    RECT 0 0 4.180 67.200 ;
    LAYER M3 ;
    RECT 0 0 4.180 67.200 ;
    LAYER M4 ;
    RECT 0.1 0 4.080 67.200 ;
    LAYER M5 ;
    RECT 0.048 0 4.132 67.200 ;
  END
END fakeram7_256x32

END LIBRARY
