module gcd (clk,
    req_rdy,
    req_val,
    reset,
    resp_rdy,
    resp_val,
    req_msg,
    resp_msg);
 input clk;
 output req_rdy;
 input req_val;
 input reset;
 input resp_rdy;
 output resp_val;
 input [31:0] req_msg;
 output [15:0] resp_msg;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire net2;
 wire net1;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire clknet_2_3__leaf_clk;
 wire _171_;
 wire _172_;
 wire clknet_2_2__leaf_clk;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire clknet_2_1__leaf_clk;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire clknet_2_0__leaf_clk;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire clknet_0_clk;
 wire _205_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire \ctrl.state.out[1] ;
 wire \ctrl.state.out[2] ;
 wire \dpath.a_lt_b$in0[0] ;
 wire \dpath.a_lt_b$in0[10] ;
 wire \dpath.a_lt_b$in0[11] ;
 wire \dpath.a_lt_b$in0[12] ;
 wire \dpath.a_lt_b$in0[13] ;
 wire \dpath.a_lt_b$in0[14] ;
 wire \dpath.a_lt_b$in0[15] ;
 wire \dpath.a_lt_b$in0[1] ;
 wire \dpath.a_lt_b$in0[2] ;
 wire \dpath.a_lt_b$in0[3] ;
 wire \dpath.a_lt_b$in0[4] ;
 wire \dpath.a_lt_b$in0[5] ;
 wire \dpath.a_lt_b$in0[6] ;
 wire \dpath.a_lt_b$in0[7] ;
 wire \dpath.a_lt_b$in0[8] ;
 wire \dpath.a_lt_b$in0[9] ;
 wire \dpath.a_lt_b$in1[0] ;
 wire \dpath.a_lt_b$in1[10] ;
 wire \dpath.a_lt_b$in1[11] ;
 wire \dpath.a_lt_b$in1[12] ;
 wire \dpath.a_lt_b$in1[13] ;
 wire \dpath.a_lt_b$in1[14] ;
 wire \dpath.a_lt_b$in1[15] ;
 wire \dpath.a_lt_b$in1[1] ;
 wire \dpath.a_lt_b$in1[2] ;
 wire \dpath.a_lt_b$in1[3] ;
 wire \dpath.a_lt_b$in1[4] ;
 wire \dpath.a_lt_b$in1[5] ;
 wire \dpath.a_lt_b$in1[6] ;
 wire \dpath.a_lt_b$in1[7] ;
 wire \dpath.a_lt_b$in1[8] ;
 wire \dpath.a_lt_b$in1[9] ;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;

 sky130_fd_sc_hs__nor2b_4 _252_ (.A(\dpath.a_lt_b$in0[0] ),
    .B_N(\dpath.a_lt_b$in1[0] ),
    .Y(_035_));
 sky130_fd_sc_hs__nor2b_2 _253_ (.A(\dpath.a_lt_b$in0[1] ),
    .B_N(\dpath.a_lt_b$in1[1] ),
    .Y(_036_));
 sky130_fd_sc_hs__inv_2 _254_ (.A(\dpath.a_lt_b$in1[1] ),
    .Y(_037_));
 sky130_fd_sc_hs__nand2_1 _255_ (.A(_037_),
    .B(\dpath.a_lt_b$in0[1] ),
    .Y(_038_));
 sky130_fd_sc_hs__o21ai_4 _256_ (.A1(_036_),
    .A2(_035_),
    .B1(_038_),
    .Y(_039_));
 sky130_fd_sc_hs__nand2b_1 _257_ (.A_N(\dpath.a_lt_b$in1[3] ),
    .B(\dpath.a_lt_b$in0[3] ),
    .Y(_040_));
 sky130_fd_sc_hs__nand2b_1 _258_ (.A_N(\dpath.a_lt_b$in0[3] ),
    .B(net18),
    .Y(_041_));
 sky130_fd_sc_hs__nand2_2 _259_ (.A(_041_),
    .B(_040_),
    .Y(_042_));
 sky130_fd_sc_hs__nand2b_2 _260_ (.A_N(\dpath.a_lt_b$in1[2] ),
    .B(\dpath.a_lt_b$in0[2] ),
    .Y(_043_));
 sky130_fd_sc_hs__nand2b_2 _261_ (.A_N(\dpath.a_lt_b$in0[2] ),
    .B(\dpath.a_lt_b$in1[2] ),
    .Y(_044_));
 sky130_fd_sc_hs__nand2_2 _262_ (.A(_044_),
    .B(_043_),
    .Y(_045_));
 sky130_fd_sc_hs__nor2_2 _263_ (.A(_045_),
    .B(_042_),
    .Y(_046_));
 sky130_fd_sc_hs__nand2_2 _264_ (.A(_039_),
    .B(_046_),
    .Y(_047_));
 sky130_fd_sc_hs__inv_2 _265_ (.A(net1),
    .Y(_048_));
 sky130_fd_sc_hs__nor2_1 _266_ (.A(\dpath.a_lt_b$in0[3] ),
    .B(_048_),
    .Y(_049_));
 sky130_fd_sc_hs__o21a_1 _267_ (.A1(_043_),
    .A2(_049_),
    .B1(_040_),
    .X(_050_));
 sky130_fd_sc_hs__nand2_8 _268_ (.A(_050_),
    .B(_047_),
    .Y(_051_));
 sky130_fd_sc_hs__inv_1 _269_ (.A(\dpath.a_lt_b$in1[7] ),
    .Y(_052_));
 sky130_fd_sc_hs__nand2_1 _270_ (.A(_052_),
    .B(\dpath.a_lt_b$in0[7] ),
    .Y(_053_));
 sky130_fd_sc_hs__nand2b_1 _271_ (.A_N(\dpath.a_lt_b$in0[7] ),
    .B(\dpath.a_lt_b$in1[7] ),
    .Y(_054_));
 sky130_fd_sc_hs__and2_4 _272_ (.A(_054_),
    .B(_053_),
    .X(_055_));
 sky130_fd_sc_hs__xnor2_4 _273_ (.A(\dpath.a_lt_b$in0[6] ),
    .B(\dpath.a_lt_b$in1[6] ),
    .Y(_056_));
 sky130_fd_sc_hs__nand2_2 _274_ (.A(_055_),
    .B(_056_),
    .Y(_057_));
 sky130_fd_sc_hs__inv_1 _275_ (.A(\dpath.a_lt_b$in1[5] ),
    .Y(_058_));
 sky130_fd_sc_hs__nand2_2 _276_ (.A(_058_),
    .B(\dpath.a_lt_b$in0[5] ),
    .Y(_059_));
 sky130_fd_sc_hs__nand2b_2 _277_ (.A_N(\dpath.a_lt_b$in0[5] ),
    .B(\dpath.a_lt_b$in1[5] ),
    .Y(_060_));
 sky130_fd_sc_hs__and2_4 _278_ (.A(_059_),
    .B(_060_),
    .X(_061_));
 sky130_fd_sc_hs__xnor2_4 _279_ (.A(\dpath.a_lt_b$in1[4] ),
    .B(\dpath.a_lt_b$in0[4] ),
    .Y(_062_));
 sky130_fd_sc_hs__nand2_1 _280_ (.A(_061_),
    .B(_062_),
    .Y(_063_));
 sky130_fd_sc_hs__nor2_2 _281_ (.A(_057_),
    .B(_063_),
    .Y(_064_));
 sky130_fd_sc_hs__nand2_2 _282_ (.A(_051_),
    .B(_064_),
    .Y(_065_));
 sky130_fd_sc_hs__inv_2 _283_ (.A(\dpath.a_lt_b$in1[6] ),
    .Y(_066_));
 sky130_fd_sc_hs__nand2_1 _284_ (.A(_066_),
    .B(\dpath.a_lt_b$in0[6] ),
    .Y(_067_));
 sky130_fd_sc_hs__a21boi_1 _285_ (.A1(_053_),
    .A2(_067_),
    .B1_N(_054_),
    .Y(_068_));
 sky130_fd_sc_hs__inv_2 _286_ (.A(\dpath.a_lt_b$in1[4] ),
    .Y(_069_));
 sky130_fd_sc_hs__nand2_1 _287_ (.A(_069_),
    .B(\dpath.a_lt_b$in0[4] ),
    .Y(_070_));
 sky130_fd_sc_hs__nand2_1 _288_ (.A(_059_),
    .B(_070_),
    .Y(_071_));
 sky130_fd_sc_hs__nand2_1 _289_ (.A(_071_),
    .B(_060_),
    .Y(_072_));
 sky130_fd_sc_hs__nor2_2 _290_ (.A(_057_),
    .B(_072_),
    .Y(_073_));
 sky130_fd_sc_hs__nor2_4 _291_ (.A(_068_),
    .B(_073_),
    .Y(_074_));
 sky130_fd_sc_hs__nand2_8 _292_ (.A(_074_),
    .B(_065_),
    .Y(_075_));
 sky130_fd_sc_hs__inv_2 _293_ (.A(\dpath.a_lt_b$in0[9] ),
    .Y(_076_));
 sky130_fd_sc_hs__xnor2_4 _294_ (.A(\dpath.a_lt_b$in1[9] ),
    .B(_076_),
    .Y(_077_));
 sky130_fd_sc_hs__inv_2 _295_ (.A(\dpath.a_lt_b$in1[8] ),
    .Y(_078_));
 sky130_fd_sc_hs__nand2_4 _296_ (.A(_078_),
    .B(\dpath.a_lt_b$in0[8] ),
    .Y(_079_));
 sky130_fd_sc_hs__inv_2 _297_ (.A(\dpath.a_lt_b$in0[8] ),
    .Y(_080_));
 sky130_fd_sc_hs__nand2_1 _298_ (.A(_080_),
    .B(\dpath.a_lt_b$in1[8] ),
    .Y(_081_));
 sky130_fd_sc_hs__nand2_4 _299_ (.A(_079_),
    .B(_081_),
    .Y(_082_));
 sky130_fd_sc_hs__xnor2_4 _300_ (.A(\dpath.a_lt_b$in1[10] ),
    .B(\dpath.a_lt_b$in0[10] ),
    .Y(_083_));
 sky130_fd_sc_hs__inv_1 _301_ (.A(\dpath.a_lt_b$in1[11] ),
    .Y(_084_));
 sky130_fd_sc_hs__nand2_4 _302_ (.A(_084_),
    .B(\dpath.a_lt_b$in0[11] ),
    .Y(_085_));
 sky130_fd_sc_hs__inv_1 _303_ (.A(\dpath.a_lt_b$in0[11] ),
    .Y(_086_));
 sky130_fd_sc_hs__nand2_2 _304_ (.A(_086_),
    .B(\dpath.a_lt_b$in1[11] ),
    .Y(_087_));
 sky130_fd_sc_hs__nand3_4 _305_ (.A(_083_),
    .B(_085_),
    .C(_087_),
    .Y(_088_));
 sky130_fd_sc_hs__nor3_4 _306_ (.A(_077_),
    .B(_082_),
    .C(_088_),
    .Y(_089_));
 sky130_fd_sc_hs__nand2_2 _307_ (.A(_075_),
    .B(_089_),
    .Y(_090_));
 sky130_fd_sc_hs__inv_1 _308_ (.A(\dpath.a_lt_b$in1[10] ),
    .Y(_091_));
 sky130_fd_sc_hs__nand2_1 _309_ (.A(_091_),
    .B(\dpath.a_lt_b$in0[10] ),
    .Y(_092_));
 sky130_fd_sc_hs__nand2_4 _310_ (.A(_085_),
    .B(_087_),
    .Y(_093_));
 sky130_fd_sc_hs__o21ai_2 _311_ (.A1(_092_),
    .A2(_093_),
    .B1(_085_),
    .Y(_094_));
 sky130_fd_sc_hs__maj3_1 _312_ (.A(\dpath.a_lt_b$in1[9] ),
    .B(_079_),
    .C(_076_),
    .X(_095_));
 sky130_fd_sc_hs__nor2_1 _313_ (.A(_088_),
    .B(_095_),
    .Y(_096_));
 sky130_fd_sc_hs__nor2_1 _314_ (.A(_094_),
    .B(_096_),
    .Y(_097_));
 sky130_fd_sc_hs__nand2_2 _315_ (.A(_097_),
    .B(_090_),
    .Y(_098_));
 sky130_fd_sc_hs__inv_2 _316_ (.A(\dpath.a_lt_b$in0[12] ),
    .Y(_099_));
 sky130_fd_sc_hs__nor2_4 _317_ (.A(\dpath.a_lt_b$in1[12] ),
    .B(_099_),
    .Y(_100_));
 sky130_fd_sc_hs__clkinv_2 _318_ (.A(_100_),
    .Y(_101_));
 sky130_fd_sc_hs__nand2_2 _319_ (.A(_099_),
    .B(\dpath.a_lt_b$in1[12] ),
    .Y(_102_));
 sky130_fd_sc_hs__nand2_8 _320_ (.A(_101_),
    .B(_102_),
    .Y(_103_));
 sky130_fd_sc_hs__inv_2 _321_ (.A(\dpath.a_lt_b$in1[13] ),
    .Y(_104_));
 sky130_fd_sc_hs__nor2_1 _322_ (.A(\dpath.a_lt_b$in0[13] ),
    .B(_104_),
    .Y(_105_));
 sky130_fd_sc_hs__and2_1 _323_ (.A(_104_),
    .B(\dpath.a_lt_b$in0[13] ),
    .X(_106_));
 sky130_fd_sc_hs__nor2_4 _324_ (.A(_105_),
    .B(_106_),
    .Y(_107_));
 sky130_fd_sc_hs__inv_2 _325_ (.A(_107_),
    .Y(_108_));
 sky130_fd_sc_hs__nor2_1 _326_ (.A(_103_),
    .B(_108_),
    .Y(_109_));
 sky130_fd_sc_hs__nand2_2 _327_ (.A(_109_),
    .B(_098_),
    .Y(_110_));
 sky130_fd_sc_hs__a21oi_4 _328_ (.A1(_107_),
    .A2(_100_),
    .B1(_106_),
    .Y(_111_));
 sky130_fd_sc_hs__nand2_2 _329_ (.A(_110_),
    .B(_111_),
    .Y(_112_));
 sky130_fd_sc_hs__xnor2_4 _330_ (.A(\dpath.a_lt_b$in1[14] ),
    .B(\dpath.a_lt_b$in0[14] ),
    .Y(_113_));
 sky130_fd_sc_hs__nand2_2 _331_ (.A(_112_),
    .B(_113_),
    .Y(_114_));
 sky130_fd_sc_hs__inv_1 _332_ (.A(\dpath.a_lt_b$in0[14] ),
    .Y(_115_));
 sky130_fd_sc_hs__nor2_1 _333_ (.A(\dpath.a_lt_b$in1[14] ),
    .B(_115_),
    .Y(_116_));
 sky130_fd_sc_hs__inv_1 _334_ (.A(_116_),
    .Y(_117_));
 sky130_fd_sc_hs__nand2_1 _335_ (.A(_117_),
    .B(_114_),
    .Y(_118_));
 sky130_fd_sc_hs__inv_2 _336_ (.A(\dpath.a_lt_b$in1[15] ),
    .Y(_119_));
 sky130_fd_sc_hs__nor2_1 _337_ (.A(\dpath.a_lt_b$in0[15] ),
    .B(_119_),
    .Y(_120_));
 sky130_fd_sc_hs__and2_1 _338_ (.A(_119_),
    .B(\dpath.a_lt_b$in0[15] ),
    .X(_121_));
 sky130_fd_sc_hs__nor2_4 _339_ (.A(_120_),
    .B(_121_),
    .Y(_122_));
 sky130_fd_sc_hs__nand2_1 _340_ (.A(_118_),
    .B(_122_),
    .Y(_123_));
 sky130_fd_sc_hs__inv_1 _341_ (.A(_122_),
    .Y(_124_));
 sky130_fd_sc_hs__nand3_1 _342_ (.A(_114_),
    .B(_117_),
    .C(_124_),
    .Y(_125_));
 sky130_fd_sc_hs__and2_2 _343_ (.A(_123_),
    .B(_125_),
    .X(resp_msg[15]));
 sky130_fd_sc_hs__xnor2_4 _344_ (.A(\dpath.a_lt_b$in1[1] ),
    .B(\dpath.a_lt_b$in0[1] ),
    .Y(_126_));
 sky130_fd_sc_hs__xnor2_4 _345_ (.A(_035_),
    .B(_126_),
    .Y(resp_msg[1]));
 sky130_fd_sc_hs__xnor2_4 _346_ (.A(net31),
    .B(net4),
    .Y(resp_msg[2]));
 sky130_fd_sc_hs__a21boi_2 _347_ (.A1(net3),
    .A2(_044_),
    .B1_N(_043_),
    .Y(_127_));
 sky130_fd_sc_hs__xor2_4 _348_ (.A(net12),
    .B(_127_),
    .X(resp_msg[3]));
 sky130_fd_sc_hs__xor2_4 _349_ (.A(_062_),
    .B(net13),
    .X(resp_msg[4]));
 sky130_fd_sc_hs__nand2_1 _350_ (.A(_051_),
    .B(_062_),
    .Y(_128_));
 sky130_fd_sc_hs__nand2_2 _351_ (.A(_128_),
    .B(_070_),
    .Y(_129_));
 sky130_fd_sc_hs__xor2_4 _352_ (.A(_061_),
    .B(_129_),
    .X(resp_msg[5]));
 sky130_fd_sc_hs__nand3_1 _353_ (.A(_051_),
    .B(_061_),
    .C(_062_),
    .Y(_130_));
 sky130_fd_sc_hs__nand2_2 _354_ (.A(_130_),
    .B(_072_),
    .Y(_131_));
 sky130_fd_sc_hs__xor2_4 _355_ (.A(net21),
    .B(_131_),
    .X(resp_msg[6]));
 sky130_fd_sc_hs__nand2_1 _356_ (.A(_131_),
    .B(net20),
    .Y(_132_));
 sky130_fd_sc_hs__nand2_2 _357_ (.A(_132_),
    .B(_067_),
    .Y(_133_));
 sky130_fd_sc_hs__xor2_4 _358_ (.A(_055_),
    .B(_133_),
    .X(resp_msg[7]));
 sky130_fd_sc_hs__xnor2_4 _359_ (.A(_082_),
    .B(net9),
    .Y(resp_msg[8]));
 sky130_fd_sc_hs__nand3_1 _360_ (.A(_075_),
    .B(_079_),
    .C(_081_),
    .Y(_134_));
 sky130_fd_sc_hs__nand2_2 _361_ (.A(_134_),
    .B(_079_),
    .Y(_135_));
 sky130_fd_sc_hs__xnor2_4 _362_ (.A(_077_),
    .B(_135_),
    .Y(resp_msg[9]));
 sky130_fd_sc_hs__nor2_1 _363_ (.A(_082_),
    .B(_077_),
    .Y(_136_));
 sky130_fd_sc_hs__nand2_1 _364_ (.A(_075_),
    .B(_136_),
    .Y(_137_));
 sky130_fd_sc_hs__nand2_2 _365_ (.A(_095_),
    .B(_137_),
    .Y(_138_));
 sky130_fd_sc_hs__xor2_4 _366_ (.A(_083_),
    .B(net37),
    .X(resp_msg[10]));
 sky130_fd_sc_hs__nand2_1 _367_ (.A(_138_),
    .B(_083_),
    .Y(_139_));
 sky130_fd_sc_hs__nand2_2 _368_ (.A(_139_),
    .B(_092_),
    .Y(_140_));
 sky130_fd_sc_hs__xnor2_4 _369_ (.A(_093_),
    .B(_140_),
    .Y(resp_msg[11]));
 sky130_fd_sc_hs__xnor2_4 _370_ (.A(_103_),
    .B(_098_),
    .Y(resp_msg[12]));
 sky130_fd_sc_hs__inv_1 _371_ (.A(_103_),
    .Y(_141_));
 sky130_fd_sc_hs__nand2_1 _372_ (.A(_098_),
    .B(_141_),
    .Y(_142_));
 sky130_fd_sc_hs__nand2_2 _373_ (.A(_142_),
    .B(_101_),
    .Y(_143_));
 sky130_fd_sc_hs__xnor2_4 _374_ (.A(_143_),
    .B(_108_),
    .Y(resp_msg[13]));
 sky130_fd_sc_hs__xor2_4 _375_ (.A(_113_),
    .B(net10),
    .X(resp_msg[14]));
 sky130_fd_sc_hs__inv_2 _376_ (.A(\dpath.a_lt_b$in1[0] ),
    .Y(_144_));
 sky130_fd_sc_hs__xnor2_4 _377_ (.A(net33),
    .B(_144_),
    .Y(resp_msg[0]));
 sky130_fd_sc_hs__inv_1 _378_ (.A(\ctrl.state.out[2] ),
    .Y(_145_));
 sky130_fd_sc_hs__nor2_1 _379_ (.A(reset),
    .B(_145_),
    .Y(_146_));
 sky130_fd_sc_hs__nor4_4 _380_ (.A(\dpath.a_lt_b$in1[12] ),
    .B(\dpath.a_lt_b$in1[13] ),
    .C(\dpath.a_lt_b$in1[14] ),
    .D(\dpath.a_lt_b$in1[15] ),
    .Y(_147_));
 sky130_fd_sc_hs__nor4_4 _381_ (.A(\dpath.a_lt_b$in1[8] ),
    .B(\dpath.a_lt_b$in1[9] ),
    .C(\dpath.a_lt_b$in1[10] ),
    .D(\dpath.a_lt_b$in1[11] ),
    .Y(_148_));
 sky130_fd_sc_hs__nor4_4 _382_ (.A(net24),
    .B(net19),
    .C(net14),
    .D(net11),
    .Y(_149_));
 sky130_fd_sc_hs__nor4_4 _383_ (.A(net6),
    .B(net2),
    .C(net32),
    .D(\dpath.a_lt_b$in1[1] ),
    .Y(_150_));
 sky130_fd_sc_hs__nand4_2 _384_ (.A(_147_),
    .B(_148_),
    .C(_149_),
    .D(_150_),
    .Y(_151_));
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_0_8 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hs__nand2_1 _387_ (.A(req_rdy),
    .B(req_val),
    .Y(_154_));
 sky130_fd_sc_hs__o2bb2ai_1 _388_ (.A1_N(_146_),
    .A2_N(_151_),
    .B1(reset),
    .B2(_154_),
    .Y(_002_));
 sky130_fd_sc_hs__nor2_8 _389_ (.A(\ctrl.state.out[2] ),
    .B(req_rdy),
    .Y(_155_));
 sky130_fd_sc_hs__and2_1 _390_ (.A(_155_),
    .B(\ctrl.state.out[1] ),
    .X(resp_val));
 sky130_fd_sc_hs__clkinv_4 _391_ (.A(req_rdy),
    .Y(_156_));
 sky130_fd_sc_hs__a21oi_1 _392_ (.A1(resp_val),
    .A2(resp_rdy),
    .B1(reset),
    .Y(_157_));
 sky130_fd_sc_hs__o21ai_1 _393_ (.A1(_156_),
    .A2(req_val),
    .B1(_157_),
    .Y(_000_));
 sky130_fd_sc_hs__nand2_1 _394_ (.A(_157_),
    .B(\ctrl.state.out[1] ),
    .Y(_158_));
 sky130_fd_sc_hs__o31ai_1 _395_ (.A1(_145_),
    .A2(reset),
    .A3(_151_),
    .B1(_158_),
    .Y(_001_));
 sky130_fd_sc_hs__or2_1 _396_ (.A(_094_),
    .B(_096_),
    .X(_159_));
 sky130_fd_sc_hs__nand2_2 _397_ (.A(_122_),
    .B(_113_),
    .Y(_160_));
 sky130_fd_sc_hs__nor3_4 _398_ (.A(_103_),
    .B(_160_),
    .C(_108_),
    .Y(_161_));
 sky130_fd_sc_hs__a21oi_1 _399_ (.A1(_122_),
    .A2(_116_),
    .B1(_121_),
    .Y(_162_));
 sky130_fd_sc_hs__o21ai_2 _400_ (.A1(_160_),
    .A2(_111_),
    .B1(_162_),
    .Y(_163_));
 sky130_fd_sc_hs__a21oi_4 _401_ (.A1(_159_),
    .A2(_161_),
    .B1(_163_),
    .Y(_164_));
 sky130_fd_sc_hs__nand3_4 _402_ (.A(net8),
    .B(_161_),
    .C(_089_),
    .Y(_165_));
 sky130_fd_sc_hs__nand2_8 _403_ (.A(_164_),
    .B(_165_),
    .Y(_166_));
 sky130_fd_sc_hs__nor2_4 _404_ (.A(_145_),
    .B(_166_),
    .Y(_167_));
 sky130_fd_sc_hs__nor2_8 _405_ (.A(req_rdy),
    .B(_167_),
    .Y(_168_));
 sky130_fd_sc_hs__clkinv_8 _406_ (.A(_168_),
    .Y(_169_));
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hs__nand2_4 _408_ (.A(_156_),
    .B(\ctrl.state.out[2] ),
    .Y(_171_));
 sky130_fd_sc_hs__nor2_8 _409_ (.A(_166_),
    .B(_171_),
    .Y(_172_));
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hs__a22oi_1 _411_ (.A1(req_rdy),
    .A2(req_msg[0]),
    .B1(net38),
    .B2(net34),
    .Y(_174_));
 sky130_fd_sc_hs__o21ai_1 _412_ (.A1(_144_),
    .A2(_169_),
    .B1(_174_),
    .Y(_003_));
 sky130_fd_sc_hs__a22oi_1 _413_ (.A1(req_rdy),
    .A2(req_msg[1]),
    .B1(net43),
    .B2(\dpath.a_lt_b$in0[1] ),
    .Y(_175_));
 sky130_fd_sc_hs__o21ai_1 _414_ (.A1(_037_),
    .A2(_169_),
    .B1(_175_),
    .Y(_004_));
 sky130_fd_sc_hs__inv_1 _415_ (.A(net5),
    .Y(_176_));
 sky130_fd_sc_hs__a22oi_1 _416_ (.A1(req_rdy),
    .A2(req_msg[2]),
    .B1(net38),
    .B2(net23),
    .Y(_177_));
 sky130_fd_sc_hs__o21ai_1 _417_ (.A1(_176_),
    .A2(_169_),
    .B1(_177_),
    .Y(_005_));
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hs__a22oi_1 _419_ (.A1(req_rdy),
    .A2(req_msg[3]),
    .B1(net43),
    .B2(net7),
    .Y(_179_));
 sky130_fd_sc_hs__o21ai_1 _420_ (.A1(net26),
    .A2(_169_),
    .B1(_179_),
    .Y(_006_));
 sky130_fd_sc_hs__a22oi_1 _421_ (.A1(req_rdy),
    .A2(req_msg[4]),
    .B1(net43),
    .B2(\dpath.a_lt_b$in0[4] ),
    .Y(_180_));
 sky130_fd_sc_hs__o21ai_1 _422_ (.A1(_069_),
    .A2(_169_),
    .B1(_180_),
    .Y(_007_));
 sky130_fd_sc_hs__a22oi_1 _423_ (.A1(req_rdy),
    .A2(req_msg[5]),
    .B1(net38),
    .B2(\dpath.a_lt_b$in0[5] ),
    .Y(_181_));
 sky130_fd_sc_hs__o21ai_1 _424_ (.A1(_058_),
    .A2(_169_),
    .B1(_181_),
    .Y(_008_));
 sky130_fd_sc_hs__a22oi_1 _425_ (.A1(req_rdy),
    .A2(req_msg[6]),
    .B1(net38),
    .B2(\dpath.a_lt_b$in0[6] ),
    .Y(_182_));
 sky130_fd_sc_hs__o21ai_1 _426_ (.A1(_066_),
    .A2(_169_),
    .B1(_182_),
    .Y(_009_));
 sky130_fd_sc_hs__a22oi_1 _427_ (.A1(req_rdy),
    .A2(req_msg[7]),
    .B1(net38),
    .B2(\dpath.a_lt_b$in0[7] ),
    .Y(_183_));
 sky130_fd_sc_hs__o21ai_1 _428_ (.A1(_052_),
    .A2(_169_),
    .B1(_183_),
    .Y(_010_));
 sky130_fd_sc_hs__nor2_1 _429_ (.A(req_msg[8]),
    .B(_156_),
    .Y(_184_));
 sky130_fd_sc_hs__a21oi_1 _430_ (.A1(_156_),
    .A2(_080_),
    .B1(_184_),
    .Y(_185_));
 sky130_fd_sc_hs__nor2_1 _431_ (.A(_185_),
    .B(_168_),
    .Y(_186_));
 sky130_fd_sc_hs__a21oi_1 _432_ (.A1(_078_),
    .A2(_168_),
    .B1(_186_),
    .Y(_011_));
 sky130_fd_sc_hs__nand2_1 _433_ (.A(_168_),
    .B(\dpath.a_lt_b$in1[9] ),
    .Y(_187_));
 sky130_fd_sc_hs__nor2_1 _434_ (.A(req_msg[9]),
    .B(_156_),
    .Y(_188_));
 sky130_fd_sc_hs__a21oi_1 _435_ (.A1(_156_),
    .A2(_076_),
    .B1(_188_),
    .Y(_189_));
 sky130_fd_sc_hs__nand2_1 _436_ (.A(_169_),
    .B(_189_),
    .Y(_190_));
 sky130_fd_sc_hs__nand2_1 _437_ (.A(_187_),
    .B(_190_),
    .Y(_012_));
 sky130_fd_sc_hs__a22oi_1 _438_ (.A1(req_rdy),
    .A2(req_msg[10]),
    .B1(net44),
    .B2(\dpath.a_lt_b$in0[10] ),
    .Y(_191_));
 sky130_fd_sc_hs__o21ai_1 _439_ (.A1(_091_),
    .A2(_169_),
    .B1(_191_),
    .Y(_013_));
 sky130_fd_sc_hs__nor2_1 _440_ (.A(req_msg[11]),
    .B(_156_),
    .Y(_192_));
 sky130_fd_sc_hs__a21oi_1 _441_ (.A1(_156_),
    .A2(_086_),
    .B1(_192_),
    .Y(_193_));
 sky130_fd_sc_hs__nor2_1 _442_ (.A(_193_),
    .B(_168_),
    .Y(_194_));
 sky130_fd_sc_hs__a21oi_1 _443_ (.A1(_084_),
    .A2(_168_),
    .B1(_194_),
    .Y(_014_));
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hs__a22oi_1 _445_ (.A1(req_rdy),
    .A2(req_msg[12]),
    .B1(net38),
    .B2(\dpath.a_lt_b$in0[12] ),
    .Y(_196_));
 sky130_fd_sc_hs__nand2_1 _446_ (.A(_168_),
    .B(\dpath.a_lt_b$in1[12] ),
    .Y(_197_));
 sky130_fd_sc_hs__nand2_1 _447_ (.A(_196_),
    .B(_197_),
    .Y(_015_));
 sky130_fd_sc_hs__a22oi_1 _448_ (.A1(req_rdy),
    .A2(req_msg[13]),
    .B1(net38),
    .B2(\dpath.a_lt_b$in0[13] ),
    .Y(_198_));
 sky130_fd_sc_hs__o21ai_1 _449_ (.A1(_104_),
    .A2(_169_),
    .B1(_198_),
    .Y(_016_));
 sky130_fd_sc_hs__a22oi_1 _450_ (.A1(req_rdy),
    .A2(req_msg[14]),
    .B1(net38),
    .B2(\dpath.a_lt_b$in0[14] ),
    .Y(_199_));
 sky130_fd_sc_hs__nand2_1 _451_ (.A(_168_),
    .B(\dpath.a_lt_b$in1[14] ),
    .Y(_200_));
 sky130_fd_sc_hs__nand2_1 _452_ (.A(_199_),
    .B(_200_),
    .Y(_017_));
 sky130_fd_sc_hs__a22oi_1 _453_ (.A1(req_rdy),
    .A2(req_msg[15]),
    .B1(net38),
    .B2(\dpath.a_lt_b$in0[15] ),
    .Y(_201_));
 sky130_fd_sc_hs__o21ai_1 _454_ (.A1(_119_),
    .A2(_169_),
    .B1(_201_),
    .Y(_018_));
 sky130_fd_sc_hs__inv_4 _455_ (.A(_172_),
    .Y(_202_));
 sky130_fd_sc_hs__a21oi_4 _456_ (.A1(_165_),
    .A2(_164_),
    .B1(_171_),
    .Y(_203_));
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hs__nand2_1 _458_ (.A(net42),
    .B(resp_msg[0]),
    .Y(_205_));
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hs__a22oi_1 _460_ (.A1(req_rdy),
    .A2(req_msg[16]),
    .B1(_155_),
    .B2(net35),
    .Y(_207_));
 sky130_fd_sc_hs__o211ai_1 _461_ (.A1(_144_),
    .A2(_202_),
    .B1(_205_),
    .C1(_207_),
    .Y(_019_));
 sky130_fd_sc_hs__nand2_1 _462_ (.A(net42),
    .B(resp_msg[1]),
    .Y(_208_));
 sky130_fd_sc_hs__nand2_1 _463_ (.A(net43),
    .B(\dpath.a_lt_b$in1[1] ),
    .Y(_209_));
 sky130_fd_sc_hs__nand2_1 _464_ (.A(_155_),
    .B(\dpath.a_lt_b$in0[1] ),
    .Y(_210_));
 sky130_fd_sc_hs__nand2_1 _465_ (.A(req_rdy),
    .B(req_msg[17]),
    .Y(_211_));
 sky130_fd_sc_hs__nand4_1 _466_ (.A(_208_),
    .B(_209_),
    .C(_210_),
    .D(_211_),
    .Y(_020_));
 sky130_fd_sc_hs__nand2_1 _467_ (.A(net42),
    .B(resp_msg[2]),
    .Y(_212_));
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hs__a22oi_1 _469_ (.A1(req_msg[18]),
    .A2(req_rdy),
    .B1(_155_),
    .B2(net22),
    .Y(_214_));
 sky130_fd_sc_hs__o211ai_1 _470_ (.A1(_176_),
    .A2(_202_),
    .B1(_212_),
    .C1(_214_),
    .Y(_021_));
 sky130_fd_sc_hs__nand2_1 _471_ (.A(net40),
    .B(resp_msg[3]),
    .Y(_215_));
 sky130_fd_sc_hs__a22oi_1 _472_ (.A1(req_msg[19]),
    .A2(req_rdy),
    .B1(_155_),
    .B2(net7),
    .Y(_216_));
 sky130_fd_sc_hs__o211ai_1 _473_ (.A1(_048_),
    .A2(_202_),
    .B1(_215_),
    .C1(_216_),
    .Y(_022_));
 sky130_fd_sc_hs__nand2_1 _474_ (.A(net40),
    .B(resp_msg[4]),
    .Y(_217_));
 sky130_fd_sc_hs__a22oi_1 _475_ (.A1(req_msg[20]),
    .A2(req_rdy),
    .B1(_155_),
    .B2(\dpath.a_lt_b$in0[4] ),
    .Y(_218_));
 sky130_fd_sc_hs__o211ai_1 _476_ (.A1(_069_),
    .A2(_202_),
    .B1(_217_),
    .C1(_218_),
    .Y(_023_));
 sky130_fd_sc_hs__nand2_1 _477_ (.A(net40),
    .B(resp_msg[5]),
    .Y(_219_));
 sky130_fd_sc_hs__a22oi_1 _478_ (.A1(req_msg[21]),
    .A2(req_rdy),
    .B1(_155_),
    .B2(net36),
    .Y(_220_));
 sky130_fd_sc_hs__o211ai_1 _479_ (.A1(_058_),
    .A2(_202_),
    .B1(_219_),
    .C1(_220_),
    .Y(_024_));
 sky130_fd_sc_hs__nand2_1 _480_ (.A(net40),
    .B(resp_msg[6]),
    .Y(_221_));
 sky130_fd_sc_hs__a22oi_1 _481_ (.A1(req_msg[22]),
    .A2(req_rdy),
    .B1(_155_),
    .B2(\dpath.a_lt_b$in0[6] ),
    .Y(_222_));
 sky130_fd_sc_hs__o211ai_1 _482_ (.A1(_066_),
    .A2(_202_),
    .B1(_221_),
    .C1(_222_),
    .Y(_025_));
 sky130_fd_sc_hs__a22oi_1 _483_ (.A1(req_msg[23]),
    .A2(req_rdy),
    .B1(_155_),
    .B2(\dpath.a_lt_b$in0[7] ),
    .Y(_223_));
 sky130_fd_sc_hs__nand2_1 _484_ (.A(resp_msg[7]),
    .B(net40),
    .Y(_224_));
 sky130_fd_sc_hs__o211ai_1 _485_ (.A1(_052_),
    .A2(_202_),
    .B1(_223_),
    .C1(_224_),
    .Y(_026_));
 sky130_fd_sc_hs__nand2_1 _486_ (.A(net40),
    .B(resp_msg[8]),
    .Y(_225_));
 sky130_fd_sc_hs__nand2_1 _487_ (.A(net43),
    .B(\dpath.a_lt_b$in1[8] ),
    .Y(_226_));
 sky130_fd_sc_hs__nand2_4 _488_ (.A(req_msg[24]),
    .B(req_rdy),
    .Y(_227_));
 sky130_fd_sc_hs__nand2_1 _489_ (.A(_155_),
    .B(\dpath.a_lt_b$in0[8] ),
    .Y(_228_));
 sky130_fd_sc_hs__nand4_1 _490_ (.A(_225_),
    .B(_226_),
    .C(_227_),
    .D(_228_),
    .Y(_027_));
 sky130_fd_sc_hs__nand2_1 _491_ (.A(resp_msg[9]),
    .B(net40),
    .Y(_229_));
 sky130_fd_sc_hs__nand2_1 _492_ (.A(_172_),
    .B(\dpath.a_lt_b$in1[9] ),
    .Y(_230_));
 sky130_fd_sc_hs__nand2_1 _493_ (.A(req_msg[25]),
    .B(req_rdy),
    .Y(_231_));
 sky130_fd_sc_hs__nand2_1 _494_ (.A(_155_),
    .B(\dpath.a_lt_b$in0[9] ),
    .Y(_232_));
 sky130_fd_sc_hs__nand4_1 _495_ (.A(_229_),
    .B(_230_),
    .C(_231_),
    .D(_232_),
    .Y(_028_));
 sky130_fd_sc_hs__nand2_1 _496_ (.A(net41),
    .B(resp_msg[10]),
    .Y(_233_));
 sky130_fd_sc_hs__a22oi_1 _497_ (.A1(req_msg[26]),
    .A2(req_rdy),
    .B1(_155_),
    .B2(\dpath.a_lt_b$in0[10] ),
    .Y(_234_));
 sky130_fd_sc_hs__o211ai_1 _498_ (.A1(_091_),
    .A2(_202_),
    .B1(_233_),
    .C1(_234_),
    .Y(_029_));
 sky130_fd_sc_hs__nand2_1 _499_ (.A(resp_msg[11]),
    .B(net39),
    .Y(_235_));
 sky130_fd_sc_hs__nand2_1 _500_ (.A(net45),
    .B(\dpath.a_lt_b$in1[11] ),
    .Y(_236_));
 sky130_fd_sc_hs__nor3_1 _501_ (.A(\ctrl.state.out[2] ),
    .B(req_rdy),
    .C(_086_),
    .Y(_237_));
 sky130_fd_sc_hs__a21oi_1 _502_ (.A1(req_msg[27]),
    .A2(req_rdy),
    .B1(_237_),
    .Y(_238_));
 sky130_fd_sc_hs__nand3_1 _503_ (.A(_235_),
    .B(_236_),
    .C(_238_),
    .Y(_030_));
 sky130_fd_sc_hs__nand2_1 _504_ (.A(net42),
    .B(resp_msg[12]),
    .Y(_239_));
 sky130_fd_sc_hs__nand2_1 _505_ (.A(net45),
    .B(\dpath.a_lt_b$in1[12] ),
    .Y(_240_));
 sky130_fd_sc_hs__nand2_1 _506_ (.A(_155_),
    .B(\dpath.a_lt_b$in0[12] ),
    .Y(_241_));
 sky130_fd_sc_hs__nand2_4 _507_ (.A(req_msg[28]),
    .B(req_rdy),
    .Y(_242_));
 sky130_fd_sc_hs__nand4_1 _508_ (.A(_239_),
    .B(_240_),
    .C(_241_),
    .D(_242_),
    .Y(_031_));
 sky130_fd_sc_hs__nand2_1 _509_ (.A(resp_msg[13]),
    .B(net39),
    .Y(_243_));
 sky130_fd_sc_hs__nand2_1 _510_ (.A(net38),
    .B(\dpath.a_lt_b$in1[13] ),
    .Y(_244_));
 sky130_fd_sc_hs__a22oi_1 _511_ (.A1(req_msg[29]),
    .A2(req_rdy),
    .B1(_155_),
    .B2(\dpath.a_lt_b$in0[13] ),
    .Y(_245_));
 sky130_fd_sc_hs__nand3_1 _512_ (.A(_243_),
    .B(_244_),
    .C(_245_),
    .Y(_032_));
 sky130_fd_sc_hs__nand2_1 _513_ (.A(resp_msg[14]),
    .B(net42),
    .Y(_246_));
 sky130_fd_sc_hs__nand2_1 _514_ (.A(net38),
    .B(\dpath.a_lt_b$in1[14] ),
    .Y(_247_));
 sky130_fd_sc_hs__a22oi_1 _515_ (.A1(req_msg[30]),
    .A2(req_rdy),
    .B1(_155_),
    .B2(\dpath.a_lt_b$in0[14] ),
    .Y(_248_));
 sky130_fd_sc_hs__nand3_1 _516_ (.A(_246_),
    .B(_247_),
    .C(_248_),
    .Y(_033_));
 sky130_fd_sc_hs__nand3_1 _517_ (.A(_123_),
    .B(_125_),
    .C(net42),
    .Y(_249_));
 sky130_fd_sc_hs__a22o_1 _518_ (.A1(req_msg[31]),
    .A2(req_rdy),
    .B1(_155_),
    .B2(\dpath.a_lt_b$in0[15] ),
    .X(_250_));
 sky130_fd_sc_hs__a21oi_1 _519_ (.A1(net45),
    .A2(\dpath.a_lt_b$in1[15] ),
    .B1(_250_),
    .Y(_251_));
 sky130_fd_sc_hs__nand2_1 _520_ (.A(_249_),
    .B(_251_),
    .Y(_034_));
 sky130_fd_sc_hs__dfxtp_4 _521_ (.D(_000_),
    .Q(req_rdy),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hs__dfxtp_1 _522_ (.D(_001_),
    .Q(\ctrl.state.out[1] ),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hs__dfxtp_4 _523_ (.D(_002_),
    .Q(\ctrl.state.out[2] ),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _524_ (.D(_003_),
    .Q(\dpath.a_lt_b$in1[0] ),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hs__dfxtp_4 _525_ (.D(_004_),
    .Q(\dpath.a_lt_b$in1[1] ),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _526_ (.D(_005_),
    .Q(\dpath.a_lt_b$in1[2] ),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _527_ (.D(_006_),
    .Q(\dpath.a_lt_b$in1[3] ),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hs__dfxtp_4 _528_ (.D(_007_),
    .Q(\dpath.a_lt_b$in1[4] ),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _529_ (.D(_008_),
    .Q(\dpath.a_lt_b$in1[5] ),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _530_ (.D(_009_),
    .Q(\dpath.a_lt_b$in1[6] ),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _531_ (.D(_010_),
    .Q(\dpath.a_lt_b$in1[7] ),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _532_ (.D(_011_),
    .Q(\dpath.a_lt_b$in1[8] ),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hs__dfxtp_4 _533_ (.D(_012_),
    .Q(\dpath.a_lt_b$in1[9] ),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _534_ (.D(_013_),
    .Q(\dpath.a_lt_b$in1[10] ),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _535_ (.D(_014_),
    .Q(\dpath.a_lt_b$in1[11] ),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _536_ (.D(_015_),
    .Q(\dpath.a_lt_b$in1[12] ),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _537_ (.D(_016_),
    .Q(\dpath.a_lt_b$in1[13] ),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hs__dfxtp_4 _538_ (.D(_017_),
    .Q(\dpath.a_lt_b$in1[14] ),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _539_ (.D(_018_),
    .Q(\dpath.a_lt_b$in1[15] ),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _540_ (.D(_019_),
    .Q(\dpath.a_lt_b$in0[0] ),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _541_ (.D(_020_),
    .Q(\dpath.a_lt_b$in0[1] ),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _542_ (.D(_021_),
    .Q(\dpath.a_lt_b$in0[2] ),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _543_ (.D(_022_),
    .Q(\dpath.a_lt_b$in0[3] ),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _544_ (.D(_023_),
    .Q(\dpath.a_lt_b$in0[4] ),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _545_ (.D(_024_),
    .Q(\dpath.a_lt_b$in0[5] ),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _546_ (.D(_025_),
    .Q(\dpath.a_lt_b$in0[6] ),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _547_ (.D(_026_),
    .Q(\dpath.a_lt_b$in0[7] ),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hs__dfxtp_1 _548_ (.D(_027_),
    .Q(\dpath.a_lt_b$in0[8] ),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hs__dfxtp_1 _549_ (.D(_028_),
    .Q(\dpath.a_lt_b$in0[9] ),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _550_ (.D(_029_),
    .Q(\dpath.a_lt_b$in0[10] ),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hs__dfxtp_1 _551_ (.D(_030_),
    .Q(\dpath.a_lt_b$in0[11] ),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hs__dfxtp_1 _552_ (.D(_031_),
    .Q(\dpath.a_lt_b$in0[12] ),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hs__dfxtp_1 _553_ (.D(_032_),
    .Q(\dpath.a_lt_b$in0[13] ),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hs__dfxtp_2 _554_ (.D(_033_),
    .Q(\dpath.a_lt_b$in0[14] ),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hs__dfxtp_1 _555_ (.D(_034_),
    .Q(\dpath.a_lt_b$in0[15] ),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_0_9 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_0_10 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_0_11 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_0_12 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_0_13 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_0_14 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_0_15 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_0_16 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_0_17 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_0_18 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_0_19 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_1_20 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_1_21 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_1_22 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_1_23 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_1_24 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_1_25 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_1_26 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_1_27 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_1_28 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_1_29 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_2_30 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_2_31 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_2_32 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_2_33 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_2_34 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_2_35 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_2_36 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_2_37 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_2_38 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_2_39 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_3_40 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_3_41 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_3_42 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_3_43 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_3_44 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_3_45 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_3_46 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_3_47 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_3_48 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_3_49 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_4_50 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_4_51 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_4_52 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_4_53 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_4_54 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_4_55 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_4_56 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_4_57 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_4_58 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_4_59 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_5_60 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_5_61 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_5_62 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_5_63 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_5_64 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_5_65 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_5_66 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_5_67 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_5_68 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_5_69 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_6_70 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_6_71 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_6_72 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_6_73 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_6_74 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_6_75 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_6_76 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_6_77 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_6_78 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_6_79 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_7_80 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_7_81 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_7_82 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_7_83 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_7_84 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_7_85 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_7_86 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_7_87 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_7_88 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_7_89 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_8_90 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_8_91 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_8_92 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_8_93 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_8_94 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_8_95 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_8_96 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_8_97 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_8_98 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_8_99 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_9_100 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_9_101 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_9_102 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_9_103 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_9_104 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_9_105 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_9_106 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_9_107 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_9_108 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_9_109 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_10_110 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_10_111 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_10_112 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_10_113 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_10_114 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_10_115 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_10_116 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_10_117 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_10_118 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_10_119 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_11_120 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_11_121 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_11_122 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_11_123 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_11_124 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_11_125 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_11_126 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_11_127 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_11_128 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_11_129 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_12_130 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_12_131 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_12_132 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_12_133 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_12_134 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_12_135 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_12_136 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_12_137 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_12_138 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_12_139 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_13_140 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_13_141 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_13_142 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_13_143 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_13_144 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_13_145 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_13_146 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_13_147 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_13_148 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_13_149 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_14_150 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_14_151 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_14_152 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_14_153 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_14_154 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_14_155 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_14_156 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_14_157 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_14_158 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_14_159 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_15_160 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_15_161 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_15_162 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_15_163 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_15_164 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_15_165 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_15_166 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_15_167 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_15_168 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_15_169 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_16_170 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_16_171 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_16_172 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_16_173 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_16_174 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_16_175 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_16_176 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_16_177 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_16_178 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_16_179 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_17_180 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_17_181 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_17_182 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_17_183 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_17_184 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_17_185 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_17_186 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_17_187 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_17_188 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_17_189 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_18_190 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_18_191 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_18_192 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_18_193 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_18_194 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_18_195 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_18_196 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_18_197 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_18_198 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_18_199 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_19_200 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_19_201 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_19_202 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_19_203 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_19_204 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_19_205 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_19_206 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_19_207 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_19_208 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_19_209 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_20_210 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_20_211 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_20_212 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_20_213 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_20_214 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_20_215 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_20_216 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_20_217 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_20_218 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_20_219 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_21_220 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_21_221 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_21_222 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_21_223 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_21_224 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_21_225 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_21_226 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_21_227 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_21_228 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_21_229 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_22_230 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_22_231 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_22_232 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_22_233 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_22_234 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_22_235 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_22_236 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_22_237 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_22_238 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_22_239 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_23_240 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_23_241 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_23_242 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_23_243 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_23_244 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_23_245 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_23_246 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_23_247 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_23_248 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_23_249 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_24_250 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_24_251 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_24_252 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_24_253 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_24_254 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_24_255 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_24_256 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_24_257 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_24_258 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_24_259 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_25_260 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_25_261 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_25_262 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_25_263 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_25_264 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_25_265 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_25_266 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_25_267 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_25_268 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_25_269 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_26_270 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_26_271 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_26_272 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_26_273 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_26_274 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_26_275 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_26_276 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_26_277 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_26_278 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_26_279 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_27_280 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_27_281 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_27_282 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_27_283 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_27_284 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_27_285 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_27_286 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_27_287 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_27_288 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_27_289 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_28_290 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_28_291 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_28_292 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_28_293 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_28_294 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_28_295 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_28_296 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_28_297 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_28_298 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_28_299 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_29_300 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_29_301 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_29_302 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_29_303 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_29_304 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_29_305 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_29_306 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_29_307 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_29_308 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_29_309 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_30_310 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_30_311 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_30_312 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_30_313 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_30_314 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_30_315 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_30_316 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_30_317 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_30_318 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_30_319 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_31_320 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_31_321 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_31_322 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_31_323 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_31_324 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_31_325 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_31_326 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_31_327 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_31_328 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_31_329 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_32_330 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_32_331 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_32_332 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_32_333 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_32_334 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_32_335 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_32_336 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_32_337 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_32_338 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_32_339 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_33_340 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_33_341 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_33_342 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_33_343 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_33_344 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_33_345 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_33_346 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_33_347 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_33_348 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_33_349 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_34_350 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_34_351 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_34_352 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_34_353 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_34_354 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_34_355 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_34_356 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_34_357 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_34_358 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_34_359 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_35_360 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_35_361 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_35_362 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_35_363 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_35_364 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_35_365 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_35_366 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_35_367 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_35_368 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_35_369 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_36_370 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_36_371 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_36_372 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_36_373 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_36_374 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_36_375 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_36_376 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_36_377 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_36_378 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_36_379 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_37_380 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_37_381 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_37_382 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_37_383 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_37_384 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_37_385 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_37_386 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_37_387 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_37_388 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_37_389 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_38_390 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_38_391 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_38_392 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_38_393 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_38_394 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_38_395 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_38_396 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_38_397 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_38_398 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_38_399 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_39_400 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_39_401 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_39_402 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_39_403 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_39_404 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_39_405 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_39_406 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_39_407 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_39_408 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_39_409 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_40_410 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_40_411 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_40_412 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_40_413 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_40_414 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_40_415 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_40_416 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_40_417 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_40_418 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_40_419 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_41_420 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_41_421 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_41_422 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_41_423 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_41_424 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_41_425 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_41_426 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_41_427 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_41_428 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_41_429 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_42_430 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_42_431 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_42_432 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_42_433 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_42_434 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_42_435 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_42_436 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_42_437 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_42_438 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_42_439 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_43_440 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_43_441 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_43_442 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_43_443 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_43_444 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_43_445 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_43_446 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_43_447 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_43_448 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_43_449 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_44_450 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_44_451 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_44_452 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_44_453 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_44_454 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_44_455 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_44_456 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_44_457 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_44_458 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_44_459 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_45_460 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_45_461 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_45_462 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_45_463 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_45_464 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_45_465 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_45_466 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_45_467 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_45_468 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_45_469 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_46_470 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_46_471 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_46_472 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_46_473 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_46_474 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_46_475 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_46_476 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_46_477 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_46_478 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_46_479 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_47_480 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_47_481 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_47_482 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_47_483 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_47_484 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_47_485 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_47_486 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_47_487 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_47_488 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_47_489 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_48_490 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_48_491 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_48_492 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_48_493 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_48_494 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_48_495 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_48_496 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_48_497 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_48_498 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_48_499 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_49_500 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_49_501 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_49_502 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_49_503 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_49_504 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_49_505 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_49_506 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_49_507 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_49_508 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_49_509 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_50_510 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_50_511 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_50_512 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_50_513 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_50_514 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_50_515 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_50_516 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_50_517 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_50_518 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_50_519 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_51_520 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_51_521 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_51_522 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_51_523 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_51_524 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_51_525 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_51_526 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_51_527 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_51_528 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_51_529 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_52_530 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_52_531 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_52_532 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_52_533 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_52_534 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_52_535 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_52_536 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_52_537 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_52_538 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_52_539 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_53_540 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_53_541 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_53_542 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_53_543 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_53_544 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_53_545 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_53_546 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_53_547 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_53_548 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_53_549 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_54_550 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_54_551 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_54_552 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_54_553 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_54_554 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_54_555 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_54_556 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_54_557 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_54_558 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_54_559 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_55_560 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_55_561 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_55_562 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_55_563 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_55_564 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_55_565 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_55_566 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_55_567 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_55_568 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_55_569 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_56_570 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_56_571 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_56_572 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_56_573 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_56_574 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_56_575 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_56_576 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_56_577 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_56_578 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_56_579 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_57_580 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_57_581 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_57_582 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_57_583 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_57_584 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_57_585 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_57_586 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_57_587 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_57_588 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_57_589 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_58_590 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_58_591 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_58_592 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_58_593 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_58_594 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_58_595 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_58_596 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_58_597 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_58_598 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_58_599 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_59_600 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_59_601 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_59_602 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_59_603 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_59_604 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_59_605 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_59_606 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_59_607 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_59_608 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_59_609 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_60_610 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_60_611 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_60_612 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_60_613 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_60_614 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_60_615 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_60_616 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_60_617 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_60_618 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_60_619 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_61_620 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_61_621 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_61_622 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_61_623 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_61_624 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_61_625 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_61_626 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_61_627 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_61_628 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_61_629 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_62_630 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_62_631 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_62_632 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_62_633 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_62_634 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_62_635 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_62_636 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_62_637 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_62_638 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_62_639 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_63_640 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_63_641 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_63_642 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_63_643 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_63_644 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_63_645 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_63_646 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_63_647 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_63_648 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_63_649 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_64_650 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_64_651 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_64_652 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_64_653 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_64_654 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_64_655 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_64_656 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_64_657 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_64_658 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_64_659 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_65_660 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_65_661 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_65_662 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_65_663 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_65_664 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_65_665 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_65_666 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_65_667 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_65_668 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_65_669 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_66_670 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_66_671 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_66_672 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_66_673 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_66_674 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_66_675 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_66_676 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_66_677 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_66_678 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_66_679 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_67_680 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_67_681 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_67_682 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_67_683 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_67_684 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_67_685 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_67_686 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_67_687 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_67_688 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_67_689 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_68_690 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_68_691 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_68_692 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_68_693 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_68_694 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_68_695 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_68_696 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_68_697 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_68_698 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_68_699 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_69_700 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_69_701 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_69_702 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_69_703 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_69_704 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_69_705 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_69_706 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_69_707 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_69_708 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_69_709 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_70_710 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_70_711 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_70_712 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_70_713 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_70_714 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_70_715 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_70_716 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_70_717 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_70_718 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_70_719 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_71_720 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_71_721 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_71_722 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_71_723 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_71_724 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_71_725 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_71_726 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_71_727 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_71_728 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_71_729 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_72_730 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_72_731 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_72_732 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_72_733 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_72_734 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_72_735 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_72_736 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_72_737 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_72_738 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_72_739 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_73_740 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_73_741 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_73_742 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_73_743 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_73_744 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_73_745 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_73_746 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_73_747 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_73_748 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_73_749 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_74_750 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_74_751 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_74_752 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_74_753 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_74_754 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_74_755 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_74_756 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_74_757 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_74_758 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_74_759 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_75_760 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_75_761 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_75_762 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_75_763 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_75_764 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_75_765 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_75_766 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_75_767 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_75_768 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_75_769 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_76_770 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_76_771 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_76_772 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_76_773 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_76_774 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_76_775 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_76_776 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_76_777 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_76_778 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_76_779 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_77_780 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_77_781 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_77_782 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_77_783 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_77_784 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_77_785 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_77_786 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_77_787 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_77_788 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_77_789 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_78_790 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_78_791 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_78_792 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_78_793 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_78_794 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_78_795 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_78_796 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_78_797 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_78_798 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_78_799 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_79_800 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_79_801 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_79_802 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_79_803 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_79_804 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_79_805 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_79_806 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_79_807 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_79_808 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_79_809 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_80_810 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_80_811 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_80_812 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_80_813 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_80_814 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_80_815 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_80_816 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_80_817 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_80_818 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_80_819 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_81_820 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_81_821 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_81_822 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_81_823 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_81_824 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_81_825 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_81_826 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_81_827 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_81_828 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_81_829 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_82_830 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_82_831 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_82_832 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_82_833 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_82_834 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_82_835 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_82_836 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_82_837 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_82_838 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_82_839 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_82_840 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_82_841 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_82_842 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_82_843 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_82_844 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_82_845 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_82_846 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_82_847 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_82_848 ();
 sky130_fd_sc_hs__tap_1 TAP_TAPCELL_ROW_82_849 ();
 sky130_fd_sc_hs__clkbuf_4 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hs__clkbuf_4 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hs__clkbuf_4 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hs__clkbuf_4 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hs__clkbuf_4 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hs__bufinv_16 clkload0 (.A(clknet_2_0__leaf_clk));
 sky130_fd_sc_hs__clkinv_4 clkload1 (.A(clknet_2_1__leaf_clk));
 sky130_fd_sc_hs__clkinv_2 clkload2 (.A(clknet_2_2__leaf_clk));
 sky130_fd_sc_hs__clkbuf_2 rebuffer1 (.A(\dpath.a_lt_b$in1[3] ),
    .X(net1));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer2 (.A(net15),
    .X(net2));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer3 (.A(_039_),
    .X(net3));
 sky130_fd_sc_hs__dlymetal6s2s_1 rebuffer4 (.A(net3),
    .X(net4));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer5 (.A(\dpath.a_lt_b$in1[2] ),
    .X(net5));
 sky130_fd_sc_hs__buf_2 rebuffer6 (.A(net27),
    .X(net6));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer7 (.A(\dpath.a_lt_b$in0[3] ),
    .X(net7));
 sky130_fd_sc_hs__buf_1 rebuffer8 (.A(net25),
    .X(net8));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer9 (.A(_075_),
    .X(net9));
 sky130_fd_sc_hs__clkbuf_2 rebuffer10 (.A(_112_),
    .X(net10));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer11 (.A(\dpath.a_lt_b$in1[7] ),
    .X(net11));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer12 (.A(_042_),
    .X(net12));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer13 (.A(_051_),
    .X(net13));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer14 (.A(\dpath.a_lt_b$in1[6] ),
    .X(net14));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer15 (.A(net16),
    .X(net15));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer16 (.A(net17),
    .X(net16));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer17 (.A(\dpath.a_lt_b$in1[3] ),
    .X(net17));
 sky130_fd_sc_hs__buf_1 rebuffer18 (.A(\dpath.a_lt_b$in1[3] ),
    .X(net18));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer19 (.A(\dpath.a_lt_b$in1[5] ),
    .X(net19));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer20 (.A(_056_),
    .X(net20));
 sky130_fd_sc_hs__dlymetal6s2s_1 rebuffer21 (.A(net20),
    .X(net21));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer22 (.A(\dpath.a_lt_b$in0[2] ),
    .X(net22));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer23 (.A(\dpath.a_lt_b$in0[2] ),
    .X(net23));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer24 (.A(\dpath.a_lt_b$in1[4] ),
    .X(net24));
 sky130_fd_sc_hs__dlymetal6s2s_1 rebuffer25 (.A(_075_),
    .X(net25));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer26 (.A(_048_),
    .X(net26));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer27 (.A(net28),
    .X(net27));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer28 (.A(net29),
    .X(net28));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer29 (.A(net30),
    .X(net29));
 sky130_fd_sc_hs__buf_1 rebuffer30 (.A(\dpath.a_lt_b$in1[2] ),
    .X(net30));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer31 (.A(_045_),
    .X(net31));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer32 (.A(\dpath.a_lt_b$in1[0] ),
    .X(net32));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer33 (.A(\dpath.a_lt_b$in0[0] ),
    .X(net33));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer34 (.A(net33),
    .X(net34));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer35 (.A(\dpath.a_lt_b$in0[0] ),
    .X(net35));
 sky130_fd_sc_hs__dlygate4sd2_1 rebuffer36 (.A(\dpath.a_lt_b$in0[5] ),
    .X(net36));
 sky130_fd_sc_hs__buf_4 rebuffer37 (.A(_138_),
    .X(net37));
 sky130_fd_sc_hs__buf_8 split38 (.A(_172_),
    .X(net38));
 sky130_fd_sc_hs__dlymetal6s2s_1 rebuffer39 (.A(_203_),
    .X(net39));
 sky130_fd_sc_hs__buf_8 rebuffer40 (.A(_203_),
    .X(net40));
 sky130_fd_sc_hs__dlymetal6s2s_1 rebuffer41 (.A(_203_),
    .X(net41));
 sky130_fd_sc_hs__buf_8 rebuffer42 (.A(_203_),
    .X(net42));
 sky130_fd_sc_hs__buf_4 rebuffer43 (.A(_172_),
    .X(net43));
 sky130_fd_sc_hs__dlymetal6s2s_1 rebuffer44 (.A(_172_),
    .X(net44));
 sky130_fd_sc_hs__buf_4 rebuffer45 (.A(_172_),
    .X(net45));
endmodule
