VERSION 5.7 ;

MACRO digital_pll
  CLASS BLOCK ;
  FOREIGN digital_pll ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 75.000 ;
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 41.050 69.460 42.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 41.040 5.200 42.640 68.240 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 21.050 69.460 22.650 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 61.050 69.460 62.650 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.040 5.200 22.640 68.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 61.040 5.200 62.640 68.240 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 69.460 68.085 ;
      LAYER met1 ;
        RECT 2.830 5.200 72.150 68.980 ;
      LAYER met2 ;
        RECT 3.410 70.720 8.090 72.605 ;
        RECT 8.930 70.720 14.070 72.605 ;
        RECT 14.910 70.720 19.590 72.605 ;
        RECT 20.430 70.720 25.570 72.605 ;
        RECT 26.410 70.720 31.090 72.605 ;
        RECT 31.930 70.720 37.070 72.605 ;
        RECT 37.910 70.720 42.590 72.605 ;
        RECT 43.430 70.720 48.570 72.605 ;
        RECT 49.410 70.720 54.090 72.605 ;
        RECT 54.930 70.720 60.070 72.605 ;
        RECT 60.910 70.720 65.590 72.605 ;
        RECT 66.430 70.720 71.570 72.605 ;
        RECT 2.860 4.280 72.120 70.720 ;
        RECT 2.860 2.195 18.210 4.280 ;
        RECT 19.050 2.195 55.470 4.280 ;
        RECT 56.310 2.195 72.120 4.280 ;
      LAYER met3 ;
        RECT 4.400 71.720 71.000 72.585 ;
        RECT 4.000 69.040 71.000 71.720 ;
        RECT 4.000 68.360 70.600 69.040 ;
        RECT 4.400 67.640 70.600 68.360 ;
        RECT 4.400 66.960 71.000 67.640 ;
        RECT 4.000 63.600 71.000 66.960 ;
        RECT 4.400 62.200 71.000 63.600 ;
        RECT 4.000 58.840 71.000 62.200 ;
        RECT 4.400 57.440 71.000 58.840 ;
        RECT 4.000 56.800 71.000 57.440 ;
        RECT 4.000 55.400 70.600 56.800 ;
        RECT 4.000 54.080 71.000 55.400 ;
        RECT 4.400 52.680 71.000 54.080 ;
        RECT 4.000 49.320 71.000 52.680 ;
        RECT 4.400 47.920 71.000 49.320 ;
        RECT 4.000 44.560 71.000 47.920 ;
        RECT 4.400 43.160 70.600 44.560 ;
        RECT 4.000 40.480 71.000 43.160 ;
        RECT 4.400 39.080 71.000 40.480 ;
        RECT 4.000 35.720 71.000 39.080 ;
        RECT 4.400 34.320 71.000 35.720 ;
        RECT 4.000 31.640 71.000 34.320 ;
        RECT 4.000 30.960 70.600 31.640 ;
        RECT 4.400 30.240 70.600 30.960 ;
        RECT 4.400 29.560 71.000 30.240 ;
        RECT 4.000 26.200 71.000 29.560 ;
        RECT 4.400 24.800 71.000 26.200 ;
        RECT 4.000 21.440 71.000 24.800 ;
        RECT 4.400 20.040 71.000 21.440 ;
        RECT 4.000 19.400 71.000 20.040 ;
        RECT 4.000 18.000 70.600 19.400 ;
        RECT 4.000 16.680 71.000 18.000 ;
        RECT 4.400 15.280 71.000 16.680 ;
        RECT 4.000 11.920 71.000 15.280 ;
        RECT 4.400 10.520 71.000 11.920 ;
        RECT 4.000 7.160 71.000 10.520 ;
        RECT 4.400 5.760 70.600 7.160 ;
        RECT 4.000 3.080 71.000 5.760 ;
        RECT 4.400 2.215 71.000 3.080 ;
      LAYER met4 ;
        RECT 0 0 75.0 10.0 ;
        RECT 0 65.0 75.0 75.0 ;
  END
END digital_pll

END LIBRARY