module counter (out);
   output out;
   DFFPOSX1 d0 (.Q(out));
endmodule

