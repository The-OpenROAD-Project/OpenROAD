VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO h4
   CLASS BLOCK ;
   SIZE 166.8 BY 240 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   PIN FE_OCPN57649_FE_OFN47241_n_6273_bar
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 132.95 0.51 133.05 ;
      END
   END FE_OCPN57649_FE_OFN47241_n_6273_bar

   PIN FE_OCPN61274_n_33700_bar
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 17.15 166.8 17.25 ;
      END
   END FE_OCPN61274_n_33700_bar

   PIN FE_OCPN61430_n_31308
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 236.35 0.51 236.45 ;
      END
   END FE_OCPN61430_n_31308

   PIN FE_OCPN61542_FE_OFN47238_mux_k_ln251_z_5__4323813_bar
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 144.95 0.51 145.05 ;
      END
   END FE_OCPN61542_FE_OFN47238_mux_k_ln251_z_5__4323813_bar

   PIN FE_OCPN61544_n_35219
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 120.55 0.51 120.65 ;
      END
   END FE_OCPN61544_n_35219

   PIN FE_OCPN61546_n_35219
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 72.5 0.255 72.7 ;
      END
   END FE_OCPN61546_n_35219

   PIN FE_OCPN62339_n_65283
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 161.95 0.51 162.05 ;
      END
   END FE_OCPN62339_n_65283

   PIN FE_OCPN63165_n_34645
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 75.95 0.51 76.05 ;
      END
   END FE_OCPN63165_n_34645

   PIN FE_OCPN63166_n_34645
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 66.15 0.51 66.25 ;
      END
   END FE_OCPN63166_n_34645

   PIN FE_OCPN63167_n_34645
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 97.15 0.51 97.25 ;
      END
   END FE_OCPN63167_n_34645

   PIN FE_OCPN63170_n_34645
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 74.95 0.51 75.05 ;
      END
   END FE_OCPN63170_n_34645

   PIN FE_OCPN63172_n_34609
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 49.15 0.51 49.25 ;
      END
   END FE_OCPN63172_n_34609

   PIN FE_OCPN63184_n_34610
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 109.55 0.51 109.65 ;
      END
   END FE_OCPN63184_n_34610

   PIN FE_OCPN63185_n_34610
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 68.95 0.51 69.05 ;
      END
   END FE_OCPN63185_n_34610

   PIN FE_OCPN63189_FE_OFN47238_mux_k_ln251_z_5__4323813_bar
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 80.75 0.51 80.85 ;
      END
   END FE_OCPN63189_FE_OFN47238_mux_k_ln251_z_5__4323813_bar

   PIN FE_OCPN63285_n_35466
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 108.35 0.51 108.45 ;
      END
   END FE_OCPN63285_n_35466

   PIN FE_OCPN63376_FE_OFN38554_n_42605
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 188.55 0.51 188.65 ;
      END
   END FE_OCPN63376_FE_OFN38554_n_42605

   PIN FE_OCPN63733_n_34650
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 68.95 0.51 69.05 ;
      END
   END FE_OCPN63733_n_34650

   PIN FE_OCPN63744_n_34677
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 102.95 0.51 103.05 ;
      END
   END FE_OCPN63744_n_34677

   PIN FE_OFN27591_n_36720
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 207.55 0.51 207.65 ;
      END
   END FE_OFN27591_n_36720

   PIN FE_OFN27671_n_36750
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 222.95 0.51 223.05 ;
      END
   END FE_OFN27671_n_36750

   PIN FE_OFN27677_n_36830
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 225.55 0.51 225.65 ;
      END
   END FE_OFN27677_n_36830

   PIN FE_OFN27695_n_36869
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 137.55 166.8 137.65 ;
      END
   END FE_OFN27695_n_36869

   PIN FE_OFN27737_n_36719
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 214.95 0.51 215.05 ;
      END
   END FE_OFN27737_n_36719

   PIN FE_OFN27793_n_36739
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 226.15 0.51 226.25 ;
      END
   END FE_OFN27793_n_36739

   PIN FE_OFN27858_n_36176
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 236.55 0.51 236.65 ;
      END
   END FE_OFN27858_n_36176

   PIN FE_OFN27943_n_36631
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 112.05 0 112.15 0.51 ;
      END
   END FE_OFN27943_n_36631

   PIN FE_OFN27945_n_36632
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 110.65 0 110.75 0.51 ;
      END
   END FE_OFN27945_n_36632

   PIN FE_OFN28066_n_36155
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 109.05 0 109.15 0.51 ;
      END
   END FE_OFN28066_n_36155

   PIN FE_OFN28109_n_36231
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 99.35 166.8 99.45 ;
      END
   END FE_OFN28109_n_36231

   PIN FE_OFN28150_n_36991
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 170.95 166.8 171.05 ;
      END
   END FE_OFN28150_n_36991

   PIN FE_OFN28264_n_36480
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 152.95 166.8 153.05 ;
      END
   END FE_OFN28264_n_36480

   PIN FE_OFN30064_n_39931
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 90.55 166.8 90.65 ;
      END
   END FE_OFN30064_n_39931

   PIN FE_OFN32324_g2_n_3744391
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 151.75 166.8 151.85 ;
      END
   END FE_OFN32324_g2_n_3744391

   PIN FE_OFN32385_n_21110
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 135.15 166.8 135.25 ;
      END
   END FE_OFN32385_n_21110

   PIN FE_OFN32386_n_21110
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 164.15 0.51 164.25 ;
      END
   END FE_OFN32386_n_21110

   PIN FE_OFN32390_n_59356
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 160.9 0.255 161.1 ;
      END
   END FE_OFN32390_n_59356

   PIN FE_OFN34192_n_82
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 138.95 166.8 139.05 ;
      END
   END FE_OFN34192_n_82

   PIN FE_OFN34385_n_7916
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 215.55 0.51 215.65 ;
      END
   END FE_OFN34385_n_7916

   PIN FE_OFN35296_n_5226969_bar
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 95.35 166.8 95.45 ;
      END
   END FE_OFN35296_n_5226969_bar

   PIN FE_OFN35387_eq_15876_46_n_18
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 122.95 0.51 123.05 ;
      END
   END FE_OFN35387_eq_15876_46_n_18

   PIN FE_OFN35405_eq_15784_44_n_18
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 55.65 239.49 55.75 240 ;
      END
   END FE_OFN35405_eq_15784_44_n_18

   PIN FE_OFN35416_eq_15782_44_n_18
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 20.05 239.49 20.15 240 ;
      END
   END FE_OFN35416_eq_15782_44_n_18

   PIN FE_OFN35557_n_48868
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 173.15 0.51 173.25 ;
      END
   END FE_OFN35557_n_48868

   PIN FE_OFN35566_n_48307
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 143.75 0.51 143.85 ;
      END
   END FE_OFN35566_n_48307

   PIN FE_OFN35724_n_49478
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 19.25 239.49 19.35 240 ;
      END
   END FE_OFN35724_n_49478

   PIN FE_OFN35827_n_43179
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 38.95 0.51 39.05 ;
      END
   END FE_OFN35827_n_43179

   PIN FE_OFN35833_n_41388
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 17.95 0.51 18.05 ;
      END
   END FE_OFN35833_n_41388

   PIN FE_OFN35980_n_51064
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 183.15 0.51 183.25 ;
      END
   END FE_OFN35980_n_51064

   PIN FE_OFN35982_n_51575
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 180.95 0.51 181.05 ;
      END
   END FE_OFN35982_n_51575

   PIN FE_OFN36039_n_49324
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 176.95 0.51 177.05 ;
      END
   END FE_OFN36039_n_49324

   PIN FE_OFN36056_n_43053
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 29.05 0 29.15 0.51 ;
      END
   END FE_OFN36056_n_43053

   PIN FE_OFN36062_n_40128
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 35.55 0.51 35.65 ;
      END
   END FE_OFN36062_n_40128

   PIN FE_OFN36065_n_48779
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 153.55 0.51 153.65 ;
      END
   END FE_OFN36065_n_48779

   PIN FE_OFN36096_n_48764
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 136.65 0 136.75 0.51 ;
      END
   END FE_OFN36096_n_48764

   PIN FE_OFN36240_n_48902
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 151.35 0.51 151.45 ;
      END
   END FE_OFN36240_n_48902

   PIN FE_OFN36242_n_49413
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 143.35 0.51 143.45 ;
      END
   END FE_OFN36242_n_49413

   PIN FE_OFN36289_n_35472
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 59.95 0.51 60.05 ;
      END
   END FE_OFN36289_n_35472

   PIN FE_OFN36290_n_35472
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 53.75 0.51 53.85 ;
      END
   END FE_OFN36290_n_35472

   PIN FE_OFN36305_sub_ln263_unr88_z_4__4328191
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 90.15 0.51 90.25 ;
      END
   END FE_OFN36305_sub_ln263_unr88_z_4__4328191

   PIN FE_OFN36306_sub_ln263_unr88_z_4__4328191
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 90.35 0.51 90.45 ;
      END
   END FE_OFN36306_sub_ln263_unr88_z_4__4328191

   PIN FE_OFN36312_n_41464
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 99.75 0.51 99.85 ;
      END
   END FE_OFN36312_n_41464

   PIN FE_OFN36434_n_51052
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 20.05 239.49 20.15 240 ;
      END
   END FE_OFN36434_n_51052

   PIN FE_OFN36478_n_39632
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 144.15 0.51 144.25 ;
      END
   END FE_OFN36478_n_39632

   PIN FE_OFN36488_n_35474
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 57.15 0.51 57.25 ;
      END
   END FE_OFN36488_n_35474

   PIN FE_OFN36489_n_35474
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 109.1 0.255 109.3 ;
      END
   END FE_OFN36489_n_35474

   PIN FE_OFN36543_n_49063
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 117.15 0.51 117.25 ;
      END
   END FE_OFN36543_n_49063

   PIN FE_OFN36564_n_48859
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 195.15 0.51 195.25 ;
      END
   END FE_OFN36564_n_48859

   PIN FE_OFN36573_n_48806
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 124.05 0 124.15 0.51 ;
      END
   END FE_OFN36573_n_48806

   PIN FE_OFN36582_n_34613
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 52.9 0.255 53.1 ;
      END
   END FE_OFN36582_n_34613

   PIN FE_OFN36613_n_49060
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 16.95 0.51 17.05 ;
      END
   END FE_OFN36613_n_49060

   PIN FE_OFN36690_n_34610
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 47.55 0.51 47.65 ;
      END
   END FE_OFN36690_n_34610

   PIN FE_OFN36698_n_43262
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 63.35 0.51 63.45 ;
      END
   END FE_OFN36698_n_43262

   PIN FE_OFN36710_n_39974
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 18.75 0.51 18.85 ;
      END
   END FE_OFN36710_n_39974

   PIN FE_OFN36729_n_35568
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 79.95 0.51 80.05 ;
      END
   END FE_OFN36729_n_35568

   PIN FE_OFN36733_n_35568
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 66.95 0.51 67.05 ;
      END
   END FE_OFN36733_n_35568

   PIN FE_OFN36770_n_40005
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 17.35 0.51 17.45 ;
      END
   END FE_OFN36770_n_40005

   PIN FE_OFN36771_n_41490
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 106.95 0.51 107.05 ;
      END
   END FE_OFN36771_n_41490

   PIN FE_OFN36774_n_39746
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 101.35 0.51 101.45 ;
      END
   END FE_OFN36774_n_39746

   PIN FE_OFN36787_sub_14956_48_n_104
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 28.35 0.51 28.45 ;
      END
   END FE_OFN36787_sub_14956_48_n_104

   PIN FE_OFN37075_sub_15040_54_n_115
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 113.35 0.51 113.45 ;
      END
   END FE_OFN37075_sub_15040_54_n_115

   PIN FE_OFN37708_n_42708
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 6.15 166.8 6.25 ;
      END
   END FE_OFN37708_n_42708

   PIN FE_OFN38237_sub_15041_54_n_115
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 125.75 0.51 125.85 ;
      END
   END FE_OFN38237_sub_15041_54_n_115

   PIN FE_OFN38498_n_42702
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 143.95 0.51 144.05 ;
      END
   END FE_OFN38498_n_42702

   PIN FE_OFN38572_n_35480
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 43.9 0.255 44.1 ;
      END
   END FE_OFN38572_n_35480

   PIN FE_OFN41497_sub_15040_54_n_63
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 53.95 0.51 54.05 ;
      END
   END FE_OFN41497_sub_15040_54_n_63

   PIN FE_OFN41895_n_226
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 151.95 166.8 152.05 ;
      END
   END FE_OFN41895_n_226

   PIN FE_OFN41977_n_228
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 148.75 166.8 148.85 ;
      END
   END FE_OFN41977_n_228

   PIN FE_OFN43137_n_35287
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 200.9 0.255 201.1 ;
      END
   END FE_OFN43137_n_35287

   PIN FE_OFN43147_n_35287
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.545 127.7 166.8 127.9 ;
      END
   END FE_OFN43147_n_35287

   PIN FE_OFN44003_n_35331
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 222.95 166.8 223.05 ;
      END
   END FE_OFN44003_n_35331

   PIN FE_OFN46305_n_35331
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 127.35 166.8 127.45 ;
      END
   END FE_OFN46305_n_35331

   PIN FE_OFN46746_n_57645
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 198.55 0.51 198.65 ;
      END
   END FE_OFN46746_n_57645

   PIN FE_OFN46835_n_18055
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.545 196.9 166.8 197.1 ;
      END
   END FE_OFN46835_n_18055

   PIN FE_OFN46837_n_5223349_bar
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.545 206.1 166.8 206.3 ;
      END
   END FE_OFN46837_n_5223349_bar

   PIN FE_OFN47466_sub_15040_54_n_63
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 69.35 0.51 69.45 ;
      END
   END FE_OFN47466_sub_15040_54_n_63

   PIN FE_OFN47467_sub_15040_54_n_63
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 71.35 0.51 71.45 ;
      END
   END FE_OFN47467_sub_15040_54_n_63

   PIN FE_OFN47469_sub_15027_54_n_55
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 108.55 0.51 108.65 ;
      END
   END FE_OFN47469_sub_15027_54_n_55

   PIN FE_OFN48512_n_59356
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 72.15 0.51 72.25 ;
      END
   END FE_OFN48512_n_59356

   PIN FE_OFN49008_n_39642
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 47.15 0.51 47.25 ;
      END
   END FE_OFN49008_n_39642

   PIN FE_OFN49020_n_42611
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 148.55 0.51 148.65 ;
      END
   END FE_OFN49020_n_42611

   PIN FE_OFN49964_n_48908
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 225.95 0.51 226.05 ;
      END
   END FE_OFN49964_n_48908

   PIN FE_OFN49999_n_49354
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 173.35 0.51 173.45 ;
      END
   END FE_OFN49999_n_49354

   PIN FE_OFN50041_n_49465
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 126.75 0.51 126.85 ;
      END
   END FE_OFN50041_n_49465

   PIN FE_OFN50111_n_49480
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 153.55 0.51 153.65 ;
      END
   END FE_OFN50111_n_49480

   PIN FE_OFN50218_n_51418
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 153.75 0.51 153.85 ;
      END
   END FE_OFN50218_n_51418

   PIN FE_OFN50523_n_57647
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 225.75 0.51 225.85 ;
      END
   END FE_OFN50523_n_57647

   PIN FE_OFN50623_n_57653
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 150.15 0.51 150.25 ;
      END
   END FE_OFN50623_n_57653

   PIN FE_OFN54179_n_57047
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 92.05 239.49 92.15 240 ;
      END
   END FE_OFN54179_n_57047

   PIN FE_OFN54264_n_57053
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 81.45 239.49 81.55 240 ;
      END
   END FE_OFN54264_n_57053

   PIN FE_OFN70124_n_36963
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 235.15 0.51 235.25 ;
      END
   END FE_OFN70124_n_36963

   PIN FE_OFN71221_n_51388
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 126.95 0.51 127.05 ;
      END
   END FE_OFN71221_n_51388

   PIN FE_OFN71870_n_49472
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 222.95 0.51 223.05 ;
      END
   END FE_OFN71870_n_49472

   PIN FE_OFN71874_n_48941
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 198.95 0.51 199.05 ;
      END
   END FE_OFN71874_n_48941

   PIN FE_OFN71876_n_49492
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 210.95 0.51 211.05 ;
      END
   END FE_OFN71876_n_49492

   PIN FE_OFN71880_n_48888
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 6.65 239.49 6.75 240 ;
      END
   END FE_OFN71880_n_48888

   PIN FE_OFN71884_n_49381
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 6.65 239.49 6.75 240 ;
      END
   END FE_OFN71884_n_49381

   PIN FE_OFN71898_n_49468
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 193.15 0.51 193.25 ;
      END
   END FE_OFN71898_n_49468

   PIN FE_OFN71900_n_48857
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 171.55 0.51 171.65 ;
      END
   END FE_OFN71900_n_48857

   PIN FE_OFN71903_n_48879
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 193.35 0.51 193.45 ;
      END
   END FE_OFN71903_n_48879

   PIN FE_OFN71950_n_49434
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 173.55 0.51 173.65 ;
      END
   END FE_OFN71950_n_49434

   PIN FE_OFN72307_n_35478
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 108.15 0.51 108.25 ;
      END
   END FE_OFN72307_n_35478

   PIN FE_OFN72308_n_35478
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 71.75 0.51 71.85 ;
      END
   END FE_OFN72308_n_35478

   PIN FE_OFN72343_n_40157
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 127.15 0.51 127.25 ;
      END
   END FE_OFN72343_n_40157

   PIN FE_OFN72353_n_34646
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 54.95 0.51 55.05 ;
      END
   END FE_OFN72353_n_34646

   PIN FE_OFN72354_n_34646
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 66.35 0.51 66.45 ;
      END
   END FE_OFN72354_n_34646

   PIN FE_OFN73017_n_35230
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 98.15 0.51 98.25 ;
      END
   END FE_OFN73017_n_35230

   PIN FE_OFN74845_n_34783
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 46.95 0.51 47.05 ;
      END
   END FE_OFN74845_n_34783

   PIN FE_OFN74988_n_34728
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 138.25 0 138.35 0.51 ;
      END
   END FE_OFN74988_n_34728

   PIN FE_OFN75036_n_39918
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 188.75 166.8 188.85 ;
      END
   END FE_OFN75036_n_39918

   PIN FE_OFN83546_n_36628
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 170.75 0.51 170.85 ;
      END
   END FE_OFN83546_n_36628

   PIN FE_OFN83569_n_36967
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 28.85 239.49 28.95 240 ;
      END
   END FE_OFN83569_n_36967

   PIN FE_OFN83591_n_36801
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 72.15 0.51 72.25 ;
      END
   END FE_OFN83591_n_36801

   PIN FE_OFN84427_n_48865
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 99.95 0.51 100.05 ;
      END
   END FE_OFN84427_n_48865

   PIN FE_OFN84447_eq_15948_66_n_18
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 152.45 0 152.55 0.51 ;
      END
   END FE_OFN84447_eq_15948_66_n_18

   PIN FE_OFN84485_n_45279
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 145.15 0.51 145.25 ;
      END
   END FE_OFN84485_n_45279

   PIN FE_OFN84520_n_51062
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 10.45 239.49 10.55 240 ;
      END
   END FE_OFN84520_n_51062

   PIN FE_OFN84522_n_51648
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 19.65 239.49 19.75 240 ;
      END
   END FE_OFN84522_n_51648

   PIN FE_OFN84525_n_51588
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 6.45 239.49 6.55 240 ;
      END
   END FE_OFN84525_n_51588

   PIN FE_OFN84528_n_48932
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 13.05 239.49 13.15 240 ;
      END
   END FE_OFN84528_n_48932

   PIN FE_OFN84547_n_51122
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 9.25 239.49 9.35 240 ;
      END
   END FE_OFN84547_n_51122

   PIN FE_OFN84549_n_51605
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 183.35 0.51 183.45 ;
      END
   END FE_OFN84549_n_51605

   PIN FE_OFN84711_n_48951
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 188.95 0.51 189.05 ;
      END
   END FE_OFN84711_n_48951

   PIN FE_OFN84743_n_61607
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 167.35 166.8 167.45 ;
      END
   END FE_OFN84743_n_61607

   PIN FE_OFN86863_n_34728
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 45.35 0.51 45.45 ;
      END
   END FE_OFN86863_n_34728

   PIN FE_OFN87003_n_36103
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 180.95 166.8 181.05 ;
      END
   END FE_OFN87003_n_36103

   PIN FE_OFN97682_n_36483
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 162.95 166.8 163.05 ;
      END
   END FE_OFN97682_n_36483

   PIN FE_OFN97790_n_7079
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 92.05 239.49 92.15 240 ;
      END
   END FE_OFN97790_n_7079

   PIN FE_OFN98056_n_43238
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 180.15 0.51 180.25 ;
      END
   END FE_OFN98056_n_43238

   PIN FE_OFN98707_n_35230
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 96.95 0.51 97.05 ;
      END
   END FE_OFN98707_n_35230

   PIN FE_RN_1121_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 162.15 0.51 162.25 ;
      END
   END FE_RN_1121_0

   PIN FE_RN_1136_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 82.65 0 82.75 0.51 ;
      END
   END FE_RN_1136_0

   PIN FE_RN_1694_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 90.55 0.51 90.65 ;
      END
   END FE_RN_1694_0

   PIN add_85566_69_n_36
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 191.35 166.8 191.45 ;
      END
   END add_85566_69_n_36

   PIN eq_15818_44_n_18
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 130.35 0.51 130.45 ;
      END
   END eq_15818_44_n_18

   PIN eq_15822_44_n_18
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 100.15 0.51 100.25 ;
      END
   END eq_15822_44_n_18

   PIN eq_15848_46_n_18
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 27.15 0.51 27.25 ;
      END
   END eq_15848_46_n_18

   PIN eq_15858_46_n_18
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 133.55 0.51 133.65 ;
      END
   END eq_15858_46_n_18

   PIN eq_15862_46_n_18
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 136.55 0.51 136.65 ;
      END
   END eq_15862_46_n_18

   PIN eq_15866_46_n_18
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 102.25 0 102.35 0.51 ;
      END
   END eq_15866_46_n_18

   PIN g2_m_5__3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 193.55 0.51 193.65 ;
      END
   END g2_m_5__3_

   PIN memread_edit_dist_g2_ln254_unr6_q_0_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 87.05 239.49 87.15 240 ;
      END
   END memread_edit_dist_g2_ln254_unr6_q_0_

   PIN memread_edit_dist_g2_ln254_unr6_q_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 143.65 239.49 143.75 240 ;
      END
   END memread_edit_dist_g2_ln254_unr6_q_3_

   PIN mux_g_ln477_q_117_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 147.95 166.8 148.05 ;
      END
   END mux_g_ln477_q_117_

   PIN mux_g_ln477_q_128_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 125.95 166.8 126.05 ;
      END
   END mux_g_ln477_q_128_

   PIN n_10566
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 57.45 239.49 57.55 240 ;
      END
   END n_10566

   PIN n_11993
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 181.95 0.51 182.05 ;
      END
   END n_11993

   PIN n_11994
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 206.55 0.51 206.65 ;
      END
   END n_11994

   PIN n_11995
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 204.95 166.8 205.05 ;
      END
   END n_11995

   PIN n_11997
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 197.95 0.51 198.05 ;
      END
   END n_11997

   PIN n_11998
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 212.95 0.51 213.05 ;
      END
   END n_11998

   PIN n_11999
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 207.75 166.8 207.85 ;
      END
   END n_11999

   PIN n_12000
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 235.55 0.51 235.65 ;
      END
   END n_12000

   PIN n_12001
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 194.95 166.8 195.05 ;
      END
   END n_12001

   PIN n_12002
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 206.75 0.51 206.85 ;
      END
   END n_12002

   PIN n_12003
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 224.35 166.8 224.45 ;
      END
   END n_12003

   PIN n_12004
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 207.75 0.51 207.85 ;
      END
   END n_12004

   PIN n_12005
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 166.29 207.55 166.8 207.65 ;
      END
   END n_12005

   PIN n_12006
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 225.15 0.51 225.25 ;
      END
   END n_12006

   PIN n_12026
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 206.95 0.51 207.05 ;
      END
   END n_12026

   PIN n_12027
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 190.35 0.51 190.45 ;
      END
   END n_12027

   PIN n_12345
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 197.95 166.8 198.05 ;
      END
   END n_12345

   PIN n_12353
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 207.35 0.51 207.45 ;
      END
   END n_12353

   PIN n_12926
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 236.75 0.51 236.85 ;
      END
   END n_12926

   PIN n_12932
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 236.95 0.51 237.05 ;
      END
   END n_12932

   PIN n_14365
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 192.15 166.8 192.25 ;
      END
   END n_14365

   PIN n_14987
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 237.15 0.51 237.25 ;
      END
   END n_14987

   PIN n_15857
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 214.95 166.8 215.05 ;
      END
   END n_15857

   PIN n_15877
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 216.15 166.8 216.25 ;
      END
   END n_15877

   PIN n_17531
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 206.55 166.8 206.65 ;
      END
   END n_17531

   PIN n_17902
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 202.55 166.8 202.65 ;
      END
   END n_17902

   PIN n_18259
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 197.35 166.8 197.45 ;
      END
   END n_18259

   PIN n_18380
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 206.95 166.8 207.05 ;
      END
   END n_18380

   PIN n_18657
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 214.1 0.255 214.3 ;
      END
   END n_18657

   PIN n_18826
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 25.85 0 25.95 0.51 ;
      END
   END n_18826

   PIN n_21936
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 191.75 166.8 191.85 ;
      END
   END n_21936

   PIN n_2287
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 223.15 0.51 223.25 ;
      END
   END n_2287

   PIN n_25366
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 98.55 0.51 98.65 ;
      END
   END n_25366

   PIN n_25372
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 80.95 0.51 81.05 ;
      END
   END n_25372

   PIN n_31455
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 181.15 166.8 181.25 ;
      END
   END n_31455

   PIN n_3429
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 145.85 239.49 145.95 240 ;
      END
   END n_3429

   PIN n_34414
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 136.15 0.51 136.25 ;
      END
   END n_34414

   PIN n_34611
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 47.5 0.255 47.7 ;
      END
   END n_34611

   PIN n_34613
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 70.9 0.255 71.1 ;
      END
   END n_34613

   PIN n_34614
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 44.9 0.255 45.1 ;
      END
   END n_34614

   PIN n_34647
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 57.3 0.255 57.5 ;
      END
   END n_34647

   PIN n_34648
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 108.7 0.255 108.9 ;
      END
   END n_34648

   PIN n_34649
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 90.75 0.51 90.85 ;
      END
   END n_34649

   PIN n_34684
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 105.95 0.51 106.05 ;
      END
   END n_34684

   PIN n_35083
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 116.75 0.51 116.85 ;
      END
   END n_35083

   PIN n_35219
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 123.15 0.51 123.25 ;
      END
   END n_35219

   PIN n_35229
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 100.9 0.255 101.1 ;
      END
   END n_35229

   PIN n_35231
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 79.3 0.255 79.5 ;
      END
   END n_35231

   PIN n_35232
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 27.3 0.255 27.5 ;
      END
   END n_35232

   PIN n_35448
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 94.75 0.51 94.85 ;
      END
   END n_35448

   PIN n_35471
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 44.3 0.255 44.5 ;
      END
   END n_35471

   PIN n_35472
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 71.55 0.51 71.65 ;
      END
   END n_35472

   PIN n_35475
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 17.15 0.51 17.25 ;
      END
   END n_35475

   PIN n_35476
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 98.95 0.51 99.05 ;
      END
   END n_35476

   PIN n_35477
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 116.1 0.255 116.3 ;
      END
   END n_35477

   PIN n_35479
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 63.55 0.51 63.65 ;
      END
   END n_35479

   PIN n_35507
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 58.75 0.51 58.85 ;
      END
   END n_35507

   PIN n_35515
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 6.95 0.51 7.05 ;
      END
   END n_35515

   PIN n_35563
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 73.3 0.255 73.5 ;
      END
   END n_35563

   PIN n_35567
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 57.5 0.255 57.7 ;
      END
   END n_35567

   PIN n_35590
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 90.95 0.51 91.05 ;
      END
   END n_35590

   PIN n_35722
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 49.95 0.51 50.05 ;
      END
   END n_35722

   PIN n_35728
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 37.35 0.51 37.45 ;
      END
   END n_35728

   PIN n_35774
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 59.35 166.8 59.45 ;
      END
   END n_35774

   PIN n_35775
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 80.35 0.51 80.45 ;
      END
   END n_35775

   PIN n_3604
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 44.85 239.49 44.95 240 ;
      END
   END n_3604

   PIN n_3608
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 57.65 239.49 57.75 240 ;
      END
   END n_3608

   PIN n_36089
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 188.95 166.8 189.05 ;
      END
   END n_36089

   PIN n_3612
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 220.15 0.51 220.25 ;
      END
   END n_3612

   PIN n_36199
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 99.55 166.8 99.65 ;
      END
   END n_36199

   PIN n_36776
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 145.85 0 145.95 0.51 ;
      END
   END n_36776

   PIN n_36959
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 29.05 239.49 29.15 240 ;
      END
   END n_36959

   PIN n_37013
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 100.65 239.49 100.75 240 ;
      END
   END n_37013

   PIN n_37017
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 234.95 0.51 235.05 ;
      END
   END n_37017

   PIN n_37026
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 168.95 166.8 169.05 ;
      END
   END n_37026

   PIN n_37033
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 180.55 166.8 180.65 ;
      END
   END n_37033

   PIN n_39567
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 135.15 0.51 135.25 ;
      END
   END n_39567

   PIN n_39579
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 128.95 0.51 129.05 ;
      END
   END n_39579

   PIN n_39580
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 126.35 0.51 126.45 ;
      END
   END n_39580

   PIN n_39675
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 48.75 0.51 48.85 ;
      END
   END n_39675

   PIN n_39833
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 80.15 0.51 80.25 ;
      END
   END n_39833

   PIN n_39839
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 89.15 0.51 89.25 ;
      END
   END n_39839

   PIN n_39854
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 57.15 166.8 57.25 ;
      END
   END n_39854

   PIN n_39882
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 197.55 0.51 197.65 ;
      END
   END n_39882

   PIN n_39911
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 158.95 166.8 159.05 ;
      END
   END n_39911

   PIN n_39920
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 108.35 166.8 108.45 ;
      END
   END n_39920

   PIN n_39965
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 103.35 0.51 103.45 ;
      END
   END n_39965

   PIN n_40114
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 109.75 0.51 109.85 ;
      END
   END n_40114

   PIN n_41399
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 72.35 0.51 72.45 ;
      END
   END n_41399

   PIN n_41410
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 119.95 0.51 120.05 ;
      END
   END n_41410

   PIN n_41424
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 134.55 0.51 134.65 ;
      END
   END n_41424

   PIN n_42305
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 58.55 0.51 58.65 ;
      END
   END n_42305

   PIN n_42524
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 100.65 0 100.75 0.51 ;
      END
   END n_42524

   PIN n_42707
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 6.35 166.8 6.45 ;
      END
   END n_42707

   PIN n_42987
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 118.95 0.51 119.05 ;
      END
   END n_42987

   PIN n_43058
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 99.15 0.51 99.25 ;
      END
   END n_43058

   PIN n_43098
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 99.35 0.51 99.45 ;
      END
   END n_43098

   PIN n_43116
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 98.75 0.51 98.85 ;
      END
   END n_43116

   PIN n_43142
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 128.95 0.51 129.05 ;
      END
   END n_43142

   PIN n_43174
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 9.75 0.51 9.85 ;
      END
   END n_43174

   PIN n_45172
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 28.15 0.51 28.25 ;
      END
   END n_45172

   PIN n_45277
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 120.15 0.51 120.25 ;
      END
   END n_45277

   PIN n_45524
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 89.55 0.51 89.65 ;
      END
   END n_45524

   PIN n_45825
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 18.75 166.8 18.85 ;
      END
   END n_45825

   PIN n_45972
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 58.35 0.51 58.45 ;
      END
   END n_45972

   PIN n_46005
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 80.55 0.51 80.65 ;
      END
   END n_46005

   PIN n_46166
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 35.75 0.51 35.85 ;
      END
   END n_46166

   PIN n_46167
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 35.95 0.51 36.05 ;
      END
   END n_46167

   PIN n_46192
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 73.45 0 73.55 0.51 ;
      END
   END n_46192

   PIN n_46540
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 90.95 166.8 91.05 ;
      END
   END n_46540

   PIN n_46555
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 18.95 166.8 19.05 ;
      END
   END n_46555

   PIN n_46557
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 55.85 0 55.95 0.51 ;
      END
   END n_46557

   PIN n_48369
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 180.35 0.51 180.45 ;
      END
   END n_48369

   PIN n_48630
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 136.35 0.51 136.45 ;
      END
   END n_48630

   PIN n_48760
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 100.85 0 100.95 0.51 ;
      END
   END n_48760

   PIN n_48784
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 19.15 166.8 19.25 ;
      END
   END n_48784

   PIN n_48790
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 45.35 166.8 45.45 ;
      END
   END n_48790

   PIN n_48801
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 45.55 166.8 45.65 ;
      END
   END n_48801

   PIN n_48882
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 58.65 0 58.75 0.51 ;
      END
   END n_48882

   PIN n_48894
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 144.55 0.51 144.65 ;
      END
   END n_48894

   PIN n_48907
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 225.95 0.51 226.05 ;
      END
   END n_48907

   PIN n_48913
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 162.35 0.51 162.45 ;
      END
   END n_48913

   PIN n_48927
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 164.35 0.51 164.45 ;
      END
   END n_48927

   PIN n_49353
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 47.75 0.51 47.85 ;
      END
   END n_49353

   PIN n_49364
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 151.55 0.51 151.65 ;
      END
   END n_49364

   PIN n_49837
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 207.35 0.51 207.45 ;
      END
   END n_49837

   PIN n_5042
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 100.95 0.51 101.05 ;
      END
   END n_5042

   PIN n_51039
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 188.75 0.51 188.85 ;
      END
   END n_51039

   PIN n_51043
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 171.75 0.51 171.85 ;
      END
   END n_51043

   PIN n_51046
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 56.45 239.49 56.55 240 ;
      END
   END n_51046

   PIN n_51219
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 171.35 0.51 171.45 ;
      END
   END n_51219

   PIN n_51577
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 198.75 0.51 198.85 ;
      END
   END n_51577

   PIN n_51584
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 226.15 0.51 226.25 ;
      END
   END n_51584

   PIN n_51600
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 198.15 0.51 198.25 ;
      END
   END n_51600

   PIN n_51640
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 103.45 239.49 103.55 240 ;
      END
   END n_51640

   PIN n_51655
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 234.75 0.51 234.85 ;
      END
   END n_51655

   PIN n_51678
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 6.75 0.51 6.85 ;
      END
   END n_51678

   PIN n_51711
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 189.15 0.51 189.25 ;
      END
   END n_51711

   PIN n_5226968_bar
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 118.95 166.8 119.05 ;
      END
   END n_5226968_bar

   PIN n_58231
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 115.35 166.8 115.45 ;
      END
   END n_58231

   PIN n_58248
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 117.15 166.8 117.25 ;
      END
   END n_58248

   PIN n_58255
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 119.35 166.8 119.45 ;
      END
   END n_58255

   PIN n_58274
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 36.75 166.8 36.85 ;
      END
   END n_58274

   PIN n_58468
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 99.75 166.8 99.85 ;
      END
   END n_58468

   PIN n_58771
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 120.95 166.8 121.05 ;
      END
   END n_58771

   PIN n_60940
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 107.35 0.51 107.45 ;
      END
   END n_60940

   PIN n_61
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 37.65 239.49 37.75 240 ;
      END
   END n_61

   PIN n_61009
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 143.55 0.51 143.65 ;
      END
   END n_61009

   PIN n_61819
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 99.55 0.51 99.65 ;
      END
   END n_61819

   PIN n_65255
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 37.55 0.51 37.65 ;
      END
   END n_65255

   PIN n_65263
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 103.45 0 103.55 0.51 ;
      END
   END n_65263

   PIN n_65290
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 100.45 239.49 100.55 240 ;
      END
   END n_65290

   PIN n_65302
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 109.65 239.49 109.75 240 ;
      END
   END n_65302

   PIN n_8376
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 202.75 0.51 202.85 ;
      END
   END n_8376

   PIN n_9348
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 207.15 166.8 207.25 ;
      END
   END n_9348

   PIN n_9349
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 216.35 166.8 216.45 ;
      END
   END n_9349

   PIN n_9350
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 212.95 166.8 213.05 ;
      END
   END n_9350

   PIN n_9351
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 213.15 166.8 213.25 ;
      END
   END n_9351

   PIN n_9353
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 213.95 166.8 214.05 ;
      END
   END n_9353

   PIN sub_14960_49_n_107
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 45.15 0.51 45.25 ;
      END
   END sub_14960_49_n_107

   PIN sub_14970_49_n_107
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 81.15 0.51 81.25 ;
      END
   END sub_14970_49_n_107

   PIN sub_14999_49_n_108
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 116.95 0.51 117.05 ;
      END
   END sub_14999_49_n_108

   PIN sub_15894_74_n_2572416
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 111.15 0.51 111.25 ;
      END
   END sub_15894_74_n_2572416

   PIN sub_ln263_unr104_z_3__4326697
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 108.75 0.51 108.85 ;
      END
   END sub_ln263_unr104_z_3__4326697

   PIN sub_ln263_unr36_z_6_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 120.35 0.51 120.45 ;
      END
   END sub_ln263_unr36_z_6_

   PIN sub_ln263_unr52_z_6_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 114.95 0.51 115.05 ;
      END
   END sub_ln263_unr52_z_6_

   PIN ternarymux_ln49_0_unr7_z_0__4472252
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 169.95 166.8 170.05 ;
      END
   END ternarymux_ln49_0_unr7_z_0__4472252

   PIN ternarymux_ln49_0_unr7_z_1__4472242
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 162.35 166.8 162.45 ;
      END
   END ternarymux_ln49_0_unr7_z_1__4472242

   PIN ternarymux_ln49_0_unr7_z_2__4472244
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 171.95 166.8 172.05 ;
      END
   END ternarymux_ln49_0_unr7_z_2__4472244

   PIN FE_OCPN57641_sub_14990_49_n_2572016
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 93.15 0.51 93.25 ;
      END
   END FE_OCPN57641_sub_14990_49_n_2572016

   PIN FE_OCPN57647_FE_OFN47241_n_6273_bar
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 133.35 0.51 133.45 ;
      END
   END FE_OCPN57647_FE_OFN47241_n_6273_bar

   PIN FE_OCPN57979_FE_OFN47238_mux_k_ln251_z_5__4323813_bar
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 130.55 0.51 130.65 ;
      END
   END FE_OCPN57979_FE_OFN47238_mux_k_ln251_z_5__4323813_bar

   PIN FE_OCPN58925_n_35465
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 141.15 0.51 141.25 ;
      END
   END FE_OCPN58925_n_35465

   PIN FE_OCPN59173_add_15054_37_n_30
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 80.95 0.51 81.05 ;
      END
   END FE_OCPN59173_add_15054_37_n_30

   PIN FE_OCPN61716_n_25369
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 107.95 0.51 108.05 ;
      END
   END FE_OCPN61716_n_25369

   PIN FE_OCPN62290_FE_OFN54291_sub_15040_54_n_2572501
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 80.15 0.51 80.25 ;
      END
   END FE_OCPN62290_FE_OFN54291_sub_15040_54_n_2572501

   PIN FE_OCPN62338_n_65283
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 90.35 166.8 90.45 ;
      END
   END FE_OCPN62338_n_65283

   PIN FE_OCPN63182_n_34649
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 89.5 0.255 89.7 ;
      END
   END FE_OCPN63182_n_34649

   PIN FE_OCPN63193_n_35226
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 114.95 0.51 115.05 ;
      END
   END FE_OCPN63193_n_35226

   PIN FE_OCPN63292_sub_15039_54_n_48
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 91.15 0.51 91.25 ;
      END
   END FE_OCPN63292_sub_15039_54_n_48

   PIN FE_OCPN63324_n_35588
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 82.95 0.51 83.05 ;
      END
   END FE_OCPN63324_n_35588

   PIN FE_OCPN63391_FE_OFN37146_sub_15016_49_n_98_bar
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 63.15 0.51 63.25 ;
      END
   END FE_OCPN63391_FE_OFN37146_sub_15016_49_n_98_bar

   PIN FE_OCPN63717_FE_OFN38588_mux_k_ln251_z_6__4323808_bar
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 126.55 0.51 126.65 ;
      END
   END FE_OCPN63717_FE_OFN38588_mux_k_ln251_z_6__4323808_bar

   PIN FE_OCPN63732_n_34650
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 69.15 0.51 69.25 ;
      END
   END FE_OCPN63732_n_34650

   PIN FE_OCPN63734_n_34650
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 49.5 0.255 49.7 ;
      END
   END FE_OCPN63734_n_34650

   PIN FE_OCPN63741_n_34677
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 88.95 0.51 89.05 ;
      END
   END FE_OCPN63741_n_34677

   PIN FE_OCPN99275_n_31308
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 154.85 239.49 154.95 240 ;
      END
   END FE_OCPN99275_n_31308

   PIN FE_OCP_RBN77513_n_58100
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 27.35 166.8 27.45 ;
      END
   END FE_OCP_RBN77513_n_58100

   PIN FE_OFN27525_n_36175
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 198.35 0.51 198.45 ;
      END
   END FE_OFN27525_n_36175

   PIN FE_OFN27527_n_36461
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 118.65 239.49 118.75 240 ;
      END
   END FE_OFN27527_n_36461

   PIN FE_OFN27529_n_36817
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 180.35 0.51 180.45 ;
      END
   END FE_OFN27529_n_36817

   PIN FE_OFN27719_n_36831
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 134.95 166.8 135.05 ;
      END
   END FE_OFN27719_n_36831

   PIN FE_OFN27721_n_36822
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 115.95 166.8 116.05 ;
      END
   END FE_OFN27721_n_36822

   PIN FE_OFN27723_n_36770
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 131.35 166.8 131.45 ;
      END
   END FE_OFN27723_n_36770

   PIN FE_OFN27736_n_36719
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 207.55 166.8 207.65 ;
      END
   END FE_OFN27736_n_36719

   PIN FE_OFN27941_n_36634
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 139.45 239.49 139.55 240 ;
      END
   END FE_OFN27941_n_36634

   PIN FE_OFN27988_n_36594
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 136.85 239.49 136.95 240 ;
      END
   END FE_OFN27988_n_36594

   PIN FE_OFN28005_n_36578
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 82.85 239.49 82.95 240 ;
      END
   END FE_OFN28005_n_36578

   PIN FE_OFN28007_n_36087
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 46.85 239.49 46.95 240 ;
      END
   END FE_OFN28007_n_36087

   PIN FE_OFN28009_n_36576
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 46.65 239.49 46.75 240 ;
      END
   END FE_OFN28009_n_36576

   PIN FE_OFN28011_n_36573
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 76.65 239.49 76.75 240 ;
      END
   END FE_OFN28011_n_36573

   PIN FE_OFN28149_n_36991
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 6.85 239.49 6.95 240 ;
      END
   END FE_OFN28149_n_36991

   PIN FE_OFN28263_n_36480
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 19.85 239.49 19.95 240 ;
      END
   END FE_OFN28263_n_36480

   PIN FE_OFN28266_n_37062
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 153.35 0.51 153.45 ;
      END
   END FE_OFN28266_n_37062

   PIN FE_OFN28302_n_36267
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 155.05 239.49 155.15 240 ;
      END
   END FE_OFN28302_n_36267

   PIN FE_OFN29813_n_59339
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 99.2 239.745 99.4 240 ;
      END
   END FE_OFN29813_n_59339

   PIN FE_OFN30059_n_34783
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 108.15 166.8 108.25 ;
      END
   END FE_OFN30059_n_34783

   PIN FE_OFN30063_n_39931
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 180.55 0.51 180.65 ;
      END
   END FE_OFN30063_n_39931

   PIN FE_OFN30374_n_34771
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 145.8 239.745 146 240 ;
      END
   END FE_OFN30374_n_34771

   PIN FE_OFN30391_n_34771
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.545 147.3 166.8 147.5 ;
      END
   END FE_OFN30391_n_34771

   PIN FE_OFN30393_n_34771
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 108.6 239.745 108.8 240 ;
      END
   END FE_OFN30393_n_34771

   PIN FE_OFN30500_n_34778
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.545 128.1 166.8 128.3 ;
      END
   END FE_OFN30500_n_34778

   PIN FE_OFN30777_n_34754
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 118 239.745 118.2 240 ;
      END
   END FE_OFN30777_n_34754

   PIN FE_OFN33694_n_871
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 64.85 239.49 64.95 240 ;
      END
   END FE_OFN33694_n_871

   PIN FE_OFN33863_n_71
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 236.15 0.51 236.25 ;
      END
   END FE_OFN33863_n_71

   PIN FE_OFN33942_n_93
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 19.85 239.49 19.95 240 ;
      END
   END FE_OFN33942_n_93

   PIN FE_OFN34078_n_87
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 28.85 239.49 28.95 240 ;
      END
   END FE_OFN34078_n_87

   PIN FE_OFN34099_n_86
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 77.85 239.49 77.95 240 ;
      END
   END FE_OFN34099_n_86

   PIN FE_OFN34189_n_82
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 138.95 0.51 139.05 ;
      END
   END FE_OFN34189_n_82

   PIN FE_OFN34490_n_224
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 158.95 0.51 159.05 ;
      END
   END FE_OFN34490_n_224

   PIN FE_OFN34615_n_223
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.545 126.9 166.8 127.1 ;
      END
   END FE_OFN34615_n_223

   PIN FE_OFN35134_n_61599
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 170.95 0.51 171.05 ;
      END
   END FE_OFN35134_n_61599

   PIN FE_OFN35392_n_43250
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 116.95 0.51 117.05 ;
      END
   END FE_OFN35392_n_43250

   PIN FE_OFN35421_eq_15766_42_n_18
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 65.05 0 65.15 0.51 ;
      END
   END FE_OFN35421_eq_15766_42_n_18

   PIN FE_OFN35722_n_49478
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 22.25 0 22.35 0.51 ;
      END
   END FE_OFN35722_n_49478

   PIN FE_OFN35745_n_60966
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 39.05 0 39.15 0.51 ;
      END
   END FE_OFN35745_n_60966

   PIN FE_OFN36439_n_43089
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 9.95 0.51 10.05 ;
      END
   END FE_OFN36439_n_43089

   PIN FE_OFN36449_n_39997
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 58.75 0.51 58.85 ;
      END
   END FE_OFN36449_n_39997

   PIN FE_OFN36464_n_43125
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 73.05 0 73.15 0.51 ;
      END
   END FE_OFN36464_n_43125

   PIN FE_OFN36476_n_39651
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 17.15 0.51 17.25 ;
      END
   END FE_OFN36476_n_39651

   PIN FE_OFN36503_n_48575
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 16.95 166.8 17.05 ;
      END
   END FE_OFN36503_n_48575

   PIN FE_OFN36505_n_43150
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 48.25 0 48.35 0.51 ;
      END
   END FE_OFN36505_n_43150

   PIN FE_OFN36515_n_45481
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 14.95 0.51 15.05 ;
      END
   END FE_OFN36515_n_45481

   PIN FE_OFN36569_n_34614
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 50.95 0.51 51.05 ;
      END
   END FE_OFN36569_n_34614

   PIN FE_OFN36584_n_51062
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 11.25 0 11.35 0.51 ;
      END
   END FE_OFN36584_n_51062

   PIN FE_OFN36712_n_35722
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 48.95 0.51 49.05 ;
      END
   END FE_OFN36712_n_35722

   PIN FE_OFN36738_n_45529
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 6.15 0.51 6.25 ;
      END
   END FE_OFN36738_n_45529

   PIN FE_OFN36754_n_35564
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 72.95 0.51 73.05 ;
      END
   END FE_OFN36754_n_35564

   PIN FE_OFN36782_n_43330
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 28.85 0 28.95 0.51 ;
      END
   END FE_OFN36782_n_43330

   PIN FE_OFN36821_n_48932
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 11.05 0 11.15 0.51 ;
      END
   END FE_OFN36821_n_48932

   PIN FE_OFN37107_n_39853
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 19.35 166.8 19.45 ;
      END
   END FE_OFN37107_n_39853

   PIN FE_OFN37260_n_45839
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 26.95 0.51 27.05 ;
      END
   END FE_OFN37260_n_45839

   PIN FE_OFN37689_n_45290
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 100.85 0 100.95 0.51 ;
      END
   END FE_OFN37689_n_45290

   PIN FE_OFN37713_n_45400
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 74.85 0 74.95 0.51 ;
      END
   END FE_OFN37713_n_45400

   PIN FE_OFN37718_n_39688
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 36.95 0.51 37.05 ;
      END
   END FE_OFN37718_n_39688

   PIN FE_OFN38279_sub_15035_54_n_74
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 80.35 0.51 80.45 ;
      END
   END FE_OFN38279_sub_15035_54_n_74

   PIN FE_OFN38497_n_42702
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 56.95 0.51 57.05 ;
      END
   END FE_OFN38497_n_42702

   PIN FE_OFN40808_n_35230
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 94.3 0.255 94.5 ;
      END
   END FE_OFN40808_n_35230

   PIN FE_OFN40809_n_35230
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 91.35 0.51 91.45 ;
      END
   END FE_OFN40809_n_35230

   PIN FE_OFN41487_sub_15027_54_n_55
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 129.95 0.51 130.05 ;
      END
   END FE_OFN41487_sub_15027_54_n_55

   PIN FE_OFN41911_n_227
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 235.95 0.51 236.05 ;
      END
   END FE_OFN41911_n_227

   PIN FE_OFN41974_n_228
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 148.75 0.51 148.85 ;
      END
   END FE_OFN41974_n_228

   PIN FE_OFN41984_n_228
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 152.75 166.8 152.85 ;
      END
   END FE_OFN41984_n_228

   PIN FE_OFN42379_n_44
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 64.85 239.49 64.95 240 ;
      END
   END FE_OFN42379_n_44

   PIN FE_OFN42673_n_16
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 136.85 239.49 136.95 240 ;
      END
   END FE_OFN42673_n_16

   PIN FE_OFN42800_n_11
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 100.25 239.49 100.35 240 ;
      END
   END FE_OFN42800_n_11

   PIN FE_OFN42823_n_10
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 117.45 239.49 117.55 240 ;
      END
   END FE_OFN42823_n_10

   PIN FE_OFN43021_n_35315
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 235.15 166.8 235.25 ;
      END
   END FE_OFN43021_n_35315

   PIN FE_OFN43045_n_35324
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.545 146.9 166.8 147.1 ;
      END
   END FE_OFN43045_n_35324

   PIN FE_OFN43227_n_35284
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 100.05 239.49 100.15 240 ;
      END
   END FE_OFN43227_n_35284

   PIN FE_OFN43246_n_35279
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 109.65 239.49 109.75 240 ;
      END
   END FE_OFN43246_n_35279

   PIN FE_OFN43814_n_67218
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 38 239.745 38.2 240 ;
      END
   END FE_OFN43814_n_67218

   PIN FE_OFN47463_sub_14941_55_n_80
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 80.75 0.51 80.85 ;
      END
   END FE_OFN47463_sub_14941_55_n_80

   PIN FE_OFN47468_sub_15027_54_n_55
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 125.15 0.51 125.25 ;
      END
   END FE_OFN47468_sub_15027_54_n_55

   PIN FE_OFN48046_sub_14960_49_n_142
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 37.15 0.51 37.25 ;
      END
   END FE_OFN48046_sub_14960_49_n_142

   PIN FE_OFN48509_n_59356
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 78.95 166.8 79.05 ;
      END
   END FE_OFN48509_n_59356

   PIN FE_OFN49847_n_77
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 88.85 239.49 88.95 240 ;
      END
   END FE_OFN49847_n_77

   PIN FE_OFN49963_n_48908
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 215.15 0.51 215.25 ;
      END
   END FE_OFN49963_n_48908

   PIN FE_OFN50044_n_49472
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 198.55 0.51 198.65 ;
      END
   END FE_OFN50044_n_49472

   PIN FE_OFN50045_n_51588
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 18.55 0.51 18.65 ;
      END
   END FE_OFN50045_n_51588

   PIN FE_OFN50048_n_51648
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 19.85 0 19.95 0.51 ;
      END
   END FE_OFN50048_n_51648

   PIN FE_OFN50217_n_51418
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 64.85 0 64.95 0.51 ;
      END
   END FE_OFN50217_n_51418

   PIN FE_OFN50653_n_58010
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 18.55 166.8 18.65 ;
      END
   END FE_OFN50653_n_58010

   PIN FE_OFN50871_n_35287
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.545 150.9 166.8 151.1 ;
      END
   END FE_OFN50871_n_35287

   PIN FE_OFN54182_n_57313
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 141.85 0 141.95 0.51 ;
      END
   END FE_OFN54182_n_57313

   PIN FE_OFN54227_n_57317
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 27.15 166.8 27.25 ;
      END
   END FE_OFN54227_n_57317

   PIN FE_OFN54578_n_21110
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 148.55 166.8 148.65 ;
      END
   END FE_OFN54578_n_21110

   PIN FE_OFN64099_n_55937
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 152.75 0.51 152.85 ;
      END
   END FE_OFN64099_n_55937

   PIN FE_OFN71220_n_51388
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 136.25 0 136.35 0.51 ;
      END
   END FE_OFN71220_n_51388

   PIN FE_OFN71873_n_48941
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 180.55 0.51 180.65 ;
      END
   END FE_OFN71873_n_48941

   PIN FE_OFN71875_n_49492
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 189.55 0.51 189.65 ;
      END
   END FE_OFN71875_n_49492

   PIN FE_OFN71879_n_48888
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 189.35 0.51 189.45 ;
      END
   END FE_OFN71879_n_48888

   PIN FE_OFN71883_n_49381
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 198.35 0.51 198.45 ;
      END
   END FE_OFN71883_n_49381

   PIN FE_OFN71949_n_49434
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 172.95 0.51 173.05 ;
      END
   END FE_OFN71949_n_49434

   PIN FE_OFN72112_n_45317
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 6.55 166.8 6.65 ;
      END
   END FE_OFN72112_n_45317

   PIN FE_OFN72158_n_43112
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 65.85 0 65.95 0.51 ;
      END
   END FE_OFN72158_n_43112

   PIN FE_OFN72170_n_42489
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 48.95 166.8 49.05 ;
      END
   END FE_OFN72170_n_42489

   PIN FE_OFN72809_sub_14939_54_n_87
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 59.75 0.51 59.85 ;
      END
   END FE_OFN72809_sub_14939_54_n_87

   PIN FE_OFN73560_n_50
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 123.85 239.49 123.95 240 ;
      END
   END FE_OFN73560_n_50

   PIN FE_OFN73816_n_234
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 91.85 239.49 91.95 240 ;
      END
   END FE_OFN73816_n_234

   PIN FE_OFN74055_ternarymux_ln49_0_unr7_z_3__4472243
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 197.75 166.8 197.85 ;
      END
   END FE_OFN74055_ternarymux_ln49_0_unr7_z_3__4472243

   PIN FE_OFN74157_n_883
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 171.15 0.51 171.25 ;
      END
   END FE_OFN74157_n_883

   PIN FE_OFN74165_n_876
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 36.65 0 36.75 0.51 ;
      END
   END FE_OFN74165_n_876

   PIN FE_OFN74186_n_875
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 28.65 0 28.75 0.51 ;
      END
   END FE_OFN74186_n_875

   PIN FE_OFN74237_n_223
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 226.5 0.255 226.7 ;
      END
   END FE_OFN74237_n_223

   PIN FE_OFN74738_n_526
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 37.85 239.49 37.95 240 ;
      END
   END FE_OFN74738_n_526

   PIN FE_OFN74885_n_34782
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 126.45 239.49 126.55 240 ;
      END
   END FE_OFN74885_n_34782

   PIN FE_OFN74896_n_34780
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 137.15 166.8 137.25 ;
      END
   END FE_OFN74896_n_34780

   PIN FE_OFN74982_n_34728
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 171.75 166.8 171.85 ;
      END
   END FE_OFN74982_n_34728

   PIN FE_OFN75096_n_34784
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 28.65 239.49 28.75 240 ;
      END
   END FE_OFN75096_n_34784

   PIN FE_OFN75341_n_35324
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 100.85 239.49 100.95 240 ;
      END
   END FE_OFN75341_n_35324

   PIN FE_OFN75380_n_35283
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 91.65 239.49 91.75 240 ;
      END
   END FE_OFN75380_n_35283

   PIN FE_OFN75718_FE_OCPN56136_n_35331
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 126.95 0.51 127.05 ;
      END
   END FE_OFN75718_FE_OCPN56136_n_35331

   PIN FE_OFN75726_n_35331
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 223.15 0.51 223.25 ;
      END
   END FE_OFN75726_n_35331

   PIN FE_OFN79437_n_57254
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 127.85 0 127.95 0.51 ;
      END
   END FE_OFN79437_n_57254

   PIN FE_OFN83573_n_36956
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 144.95 166.8 145.05 ;
      END
   END FE_OFN83573_n_36956

   PIN FE_OFN84709_n_43175
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 125.75 0.51 125.85 ;
      END
   END FE_OFN84709_n_43175

   PIN FE_OFN84938_n_7043
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 163.35 0.51 163.45 ;
      END
   END FE_OFN84938_n_7043

   PIN FE_OFN85149_n_222
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 73.65 239.49 73.75 240 ;
      END
   END FE_OFN85149_n_222

   PIN FE_OFN85189_n_226
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 112.75 166.8 112.85 ;
      END
   END FE_OFN85189_n_226

   PIN FE_OFN86333_n_4990
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 224.95 0.51 225.05 ;
      END
   END FE_OFN86333_n_4990

   PIN FE_OFN86459_n_7776
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 234.55 0.51 234.65 ;
      END
   END FE_OFN86459_n_7776

   PIN FE_OFN86874_n_34728
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 170.75 166.8 170.85 ;
      END
   END FE_OFN86874_n_34728

   PIN FE_OFN86916_n_34778
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.545 151.3 166.8 151.5 ;
      END
   END FE_OFN86916_n_34778

   PIN FE_OFN87971_n_35278
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 118.65 239.49 118.75 240 ;
      END
   END FE_OFN87971_n_35278

   PIN FE_OFN90264_n_57193
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 72.95 166.8 73.05 ;
      END
   END FE_OFN90264_n_57193

   PIN FE_OFN93509_n_57220
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 106.95 166.8 107.05 ;
      END
   END FE_OFN93509_n_57220

   PIN FE_OFN95954_n_57193
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 81.55 166.8 81.65 ;
      END
   END FE_OFN95954_n_57193

   PIN FE_OFN97666_n_36632
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 115.45 239.49 115.55 240 ;
      END
   END FE_OFN97666_n_36632

   PIN FE_OFN97681_n_36483
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 171.55 0.51 171.65 ;
      END
   END FE_OFN97681_n_36483

   PIN FE_OFN98055_n_43238
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 107.75 0.51 107.85 ;
      END
   END FE_OFN98055_n_43238

   PIN FE_OFN98229_n_865
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 161.75 0.51 161.85 ;
      END
   END FE_OFN98229_n_865

   PIN FE_RN_1119_0
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 144.15 0.51 144.25 ;
      END
   END FE_RN_1119_0

   PIN FE_RN_1120_0
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 154.95 0.51 155.05 ;
      END
   END FE_RN_1120_0

   PIN b_in_16_2
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 234.95 166.8 235.05 ;
      END
   END b_in_16_2

   PIN b_in_16_3
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 166.29 153.55 166.8 153.65 ;
      END
   END b_in_16_3

   PIN b_in_18_1
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 189.75 166.8 189.85 ;
      END
   END b_in_18_1

   PIN b_in_18_2
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 110.65 239.49 110.75 240 ;
      END
   END b_in_18_2

   PIN b_in_22_0
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 166.29 144.55 166.8 144.65 ;
      END
   END b_in_22_0

   PIN b_in_22_2
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 166.29 198.55 166.8 198.65 ;
      END
   END b_in_22_2

   PIN b_in_22_3
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 144.35 166.8 144.45 ;
      END
   END b_in_22_3

   PIN b_in_26_1
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 166.29 220.15 166.8 220.25 ;
      END
   END b_in_26_1

   PIN b_in_26_3
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 166.29 136.15 166.8 136.25 ;
      END
   END b_in_26_3

   PIN b_in_29_1
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 166.29 144.15 166.8 144.25 ;
      END
   END b_in_29_1

   PIN b_in_32_0
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 166.29 126.55 166.8 126.65 ;
      END
   END b_in_32_0

   PIN eq_15778_44_n_18
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 153.75 0.51 153.85 ;
      END
   END eq_15778_44_n_18

   PIN eq_15782_44_n_18
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 37.65 0 37.75 0.51 ;
      END
   END eq_15782_44_n_18

   PIN eq_15784_44_n_18
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 140.95 166.8 141.05 ;
      END
   END eq_15784_44_n_18

   PIN g2_q8_2_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 191.95 166.8 192.05 ;
      END
   END g2_q8_2_

   PIN g2_q8_3_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 207.35 166.8 207.45 ;
      END
   END g2_q8_3_

   PIN gt_16017_52_n_89
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 119.75 0.51 119.85 ;
      END
   END gt_16017_52_n_89

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 159.9 0.255 160.1 ;
      END
   END ispd_clk

   PIN memread_edit_dist_g2_ln254_unr7_q_4_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 180.35 166.8 180.45 ;
      END
   END memread_edit_dist_g2_ln254_unr7_q_4_

   PIN memread_edit_dist_g2_ln254_unr7_q_6_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 180.75 166.8 180.85 ;
      END
   END memread_edit_dist_g2_ln254_unr7_q_6_

   PIN memread_edit_dist_g2_ln254_unr7_q_7_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 180.15 166.8 180.25 ;
      END
   END memread_edit_dist_g2_ln254_unr7_q_7_

   PIN memread_edit_dist_g2_ln254_unr8_q_11_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 137.35 166.8 137.45 ;
      END
   END memread_edit_dist_g2_ln254_unr8_q_11_

   PIN memread_edit_dist_g2_ln254_unr8_q_9_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 108.55 166.8 108.65 ;
      END
   END memread_edit_dist_g2_ln254_unr8_q_9_

   PIN mux_g_ln477_q_65_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 213.55 0.51 213.65 ;
      END
   END mux_g_ln477_q_65_

   PIN mux_k_ln251_z_7__4323810
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 71.55 0.51 71.65 ;
      END
   END mux_k_ln251_z_7__4323810

   PIN n_11915
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 235.1 0.255 235.3 ;
      END
   END n_11915

   PIN n_12782
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 197.55 166.8 197.65 ;
      END
   END n_12782

   PIN n_14602
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 235.75 0.51 235.85 ;
      END
   END n_14602

   PIN n_15146
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.545 203.7 166.8 203.9 ;
      END
   END n_15146

   PIN n_15147
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.545 203.3 166.8 203.5 ;
      END
   END n_15147

   PIN n_18127
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 215.95 166.8 216.05 ;
      END
   END n_18127

   PIN n_18128
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 206.75 166.8 206.85 ;
      END
   END n_18128

   PIN n_18558
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 224.95 0.51 225.05 ;
      END
   END n_18558

   PIN n_18559
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 203.75 0.51 203.85 ;
      END
   END n_18559

   PIN n_18725
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 225.75 0.51 225.85 ;
      END
   END n_18725

   PIN n_18732
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 215.75 0.51 215.85 ;
      END
   END n_18732

   PIN n_18789
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 197.75 0.51 197.85 ;
      END
   END n_18789

   PIN n_18799
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 207.15 0.51 207.25 ;
      END
   END n_18799

   PIN n_18800
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 225.55 0.51 225.65 ;
      END
   END n_18800

   PIN n_18801
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 203.55 0.51 203.65 ;
      END
   END n_18801

   PIN n_18802
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 214.95 0.51 215.05 ;
      END
   END n_18802

   PIN n_18803
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 203.35 0.51 203.45 ;
      END
   END n_18803

   PIN n_18804
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 213.35 0.51 213.45 ;
      END
   END n_18804

   PIN n_18805
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 179.95 0.51 180.05 ;
      END
   END n_18805

   PIN n_2103
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 136.95 166.8 137.05 ;
      END
   END n_2103

   PIN n_21081
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 20.85 0 20.95 0.51 ;
      END
   END n_21081

   PIN n_21433
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 142.95 0.51 143.05 ;
      END
   END n_21433

   PIN n_22021
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 191.55 166.8 191.65 ;
      END
   END n_22021

   PIN n_25369
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 92.95 0.51 93.05 ;
      END
   END n_25369

   PIN n_25529
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 44.95 0.51 45.05 ;
      END
   END n_25529

   PIN n_31306
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.545 171.3 166.8 171.5 ;
      END
   END n_31306

   PIN n_3207
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 125.75 166.8 125.85 ;
      END
   END n_3207

   PIN n_34362
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 124.95 0.51 125.05 ;
      END
   END n_34362

   PIN n_34472
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 79.75 0.51 79.85 ;
      END
   END n_34472

   PIN n_34609
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 62.75 0.51 62.85 ;
      END
   END n_34609

   PIN n_34612
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 89.1 0.255 89.3 ;
      END
   END n_34612

   PIN n_34634
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 59.55 0.51 59.65 ;
      END
   END n_34634

   PIN n_34645
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 125.35 0.51 125.45 ;
      END
   END n_34645

   PIN n_34646
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 84.95 0.51 85.05 ;
      END
   END n_34646

   PIN n_35217
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 122.95 0.51 123.05 ;
      END
   END n_35217

   PIN n_35218
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 119.55 0.51 119.65 ;
      END
   END n_35218

   PIN n_35228
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 53.95 0.51 54.05 ;
      END
   END n_35228

   PIN n_35247
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 27.7 0.255 27.9 ;
      END
   END n_35247

   PIN n_35259
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 108.15 0.51 108.25 ;
      END
   END n_35259

   PIN n_35458
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 108.35 0.51 108.45 ;
      END
   END n_35458

   PIN n_35468
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 6.55 0.51 6.65 ;
      END
   END n_35468

   PIN n_35499
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 60.95 0.51 61.05 ;
      END
   END n_35499

   PIN n_35514
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 17.75 0.51 17.85 ;
      END
   END n_35514

   PIN n_35556
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 109.15 0.51 109.25 ;
      END
   END n_35556

   PIN n_35613
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 18.55 0.51 18.65 ;
      END
   END n_35613

   PIN n_35675
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 110.95 0.51 111.05 ;
      END
   END n_35675

   PIN n_3606
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 161.55 0.51 161.65 ;
      END
   END n_3606

   PIN n_3607
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 36.15 0.51 36.25 ;
      END
   END n_3607

   PIN n_3610
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 66.65 0 66.75 0.51 ;
      END
   END n_3610

   PIN n_36155
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 75.05 239.49 75.15 240 ;
      END
   END n_36155

   PIN n_36176
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 41.85 239.49 41.95 240 ;
      END
   END n_36176

   PIN n_36231
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 43.85 239.49 43.95 240 ;
      END
   END n_36231

   PIN n_36631
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 111.45 239.49 111.55 240 ;
      END
   END n_36631

   PIN n_36739
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 136.65 239.49 136.75 240 ;
      END
   END n_36739

   PIN n_36801
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 104.95 166.8 105.05 ;
      END
   END n_36801

   PIN n_39564
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 59.35 0.51 59.45 ;
      END
   END n_39564

   PIN n_39617
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 126.35 0.51 126.45 ;
      END
   END n_39617

   PIN n_39641
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 16.95 0.51 17.05 ;
      END
   END n_39641

   PIN n_39644
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 6.35 0.51 6.45 ;
      END
   END n_39644

   PIN n_39646
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 83.15 0.51 83.25 ;
      END
   END n_39646

   PIN n_39648
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 17.55 0.51 17.65 ;
      END
   END n_39648

   PIN n_39682
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 44.75 0.51 44.85 ;
      END
   END n_39682

   PIN n_39687
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 27.5 0.255 27.7 ;
      END
   END n_39687

   PIN n_39918
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 133.65 239.49 133.75 240 ;
      END
   END n_39918

   PIN n_40005
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 62.95 0.51 63.05 ;
      END
   END n_40005

   PIN n_40121
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 58.55 0.51 58.65 ;
      END
   END n_40121

   PIN n_40134
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 53.35 0.51 53.45 ;
      END
   END n_40134

   PIN n_40243
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 89.95 0.51 90.05 ;
      END
   END n_40243

   PIN n_41327
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 46.95 0.51 47.05 ;
      END
   END n_41327

   PIN n_42466
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 71.75 0.51 71.85 ;
      END
   END n_42466

   PIN n_42535
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 71.95 0.51 72.05 ;
      END
   END n_42535

   PIN n_42576
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 152.55 0.51 152.65 ;
      END
   END n_42576

   PIN n_43051
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 39.35 0.51 39.45 ;
      END
   END n_43051

   PIN n_43053
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 86.85 0 86.95 0.51 ;
      END
   END n_43053

   PIN n_43108
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 153.35 0.51 153.45 ;
      END
   END n_43108

   PIN n_43183
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 125.55 0.51 125.65 ;
      END
   END n_43183

   PIN n_43245
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 70.05 0 70.15 0.51 ;
      END
   END n_43245

   PIN n_43247
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 125.95 0.51 126.05 ;
      END
   END n_43247

   PIN n_43262
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 80.55 0.51 80.65 ;
      END
   END n_43262

   PIN n_45279
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 143.15 0.51 143.25 ;
      END
   END n_45279

   PIN n_45298
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 73.65 0 73.75 0.51 ;
      END
   END n_45298

   PIN n_45350
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 26.95 0.51 27.05 ;
      END
   END n_45350

   PIN n_45382
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 142.95 0.51 143.05 ;
      END
   END n_45382

   PIN n_45483
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 56.95 166.8 57.05 ;
      END
   END n_45483

   PIN n_45488
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 56.95 0.51 57.05 ;
      END
   END n_45488

   PIN n_46118
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 64.65 0 64.75 0.51 ;
      END
   END n_46118

   PIN n_46120
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 153.15 0.51 153.25 ;
      END
   END n_46120

   PIN n_46121
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 146.95 0.51 147.05 ;
      END
   END n_46121

   PIN n_46176
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 117.75 0.51 117.85 ;
      END
   END n_46176

   PIN n_46186
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 139.15 0.51 139.25 ;
      END
   END n_46186

   PIN n_468
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 166.75 166.8 166.85 ;
      END
   END n_468

   PIN n_48346
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 133.15 0.51 133.25 ;
      END
   END n_48346

   PIN n_48398
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 130.75 0.51 130.85 ;
      END
   END n_48398

   PIN n_48568
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 152.95 0.51 153.05 ;
      END
   END n_48568

   PIN n_48648
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 119.35 0.51 119.45 ;
      END
   END n_48648

   PIN n_48764
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 71.95 0.51 72.05 ;
      END
   END n_48764

   PIN n_48806
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 126.15 0.51 126.25 ;
      END
   END n_48806

   PIN n_48859
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 194.95 0.51 195.05 ;
      END
   END n_48859

   PIN n_48865
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 53.55 0.51 53.65 ;
      END
   END n_48865

   PIN n_48868
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 163.15 0.51 163.25 ;
      END
   END n_48868

   PIN n_48879
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 134.95 0.51 135.05 ;
      END
   END n_48879

   PIN n_48902
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 151.15 0.51 151.25 ;
      END
   END n_48902

   PIN n_48951
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 107.55 0.51 107.65 ;
      END
   END n_48951

   PIN n_49060
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 27.95 0.51 28.05 ;
      END
   END n_49060

   PIN n_49063
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 39.15 0.51 39.25 ;
      END
   END n_49063

   PIN n_49214
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 134.75 0.51 134.85 ;
      END
   END n_49214

   PIN n_49324
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 107.15 0.51 107.25 ;
      END
   END n_49324

   PIN n_49413
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 116.75 0.51 116.85 ;
      END
   END n_49413

   PIN n_49468
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 164.95 0.51 165.05 ;
      END
   END n_49468

   PIN n_49480
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 40.75 0.51 40.85 ;
      END
   END n_49480

   PIN n_4992
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 85.45 239.49 85.55 240 ;
      END
   END n_4992

   PIN n_4999
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 192.95 0.51 193.05 ;
      END
   END n_4999

   PIN n_51064
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 182.95 0.51 183.05 ;
      END
   END n_51064

   PIN n_51122
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 99.15 0.51 99.25 ;
      END
   END n_51122

   PIN n_51575
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 9.55 0.51 9.65 ;
      END
   END n_51575

   PIN n_51605
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 98.95 0.51 99.05 ;
      END
   END n_51605

   PIN n_5223120_bar
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 150.95 0.51 151.05 ;
      END
   END n_5223120_bar

   PIN n_5226969_bar
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 116.55 0.51 116.65 ;
      END
   END n_5226969_bar

   PIN n_55934
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 153.15 0.51 153.25 ;
      END
   END n_55934

   PIN n_55936
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 140.95 0.51 141.05 ;
      END
   END n_55936

   PIN n_56252
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 144.35 0.51 144.45 ;
      END
   END n_56252

   PIN n_57047
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 77.45 0 77.55 0.51 ;
      END
   END n_57047

   PIN n_57053
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 38.15 0.51 38.25 ;
      END
   END n_57053

   PIN n_57311
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 36.95 166.8 37.05 ;
      END
   END n_57311

   PIN n_57315
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 26.95 166.8 27.05 ;
      END
   END n_57315

   PIN n_57327
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 27.55 166.8 27.65 ;
      END
   END n_57327

   PIN n_57353
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 82.85 0 82.95 0.51 ;
      END
   END n_57353

   PIN n_57645
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 46.85 0 46.95 0.51 ;
      END
   END n_57645

   PIN n_57647
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 79.45 0 79.55 0.51 ;
      END
   END n_57647

   PIN n_57653
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 64.85 0 64.95 0.51 ;
      END
   END n_57653

   PIN n_58064
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 72.55 166.8 72.65 ;
      END
   END n_58064

   PIN n_58080
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 10.85 0 10.95 0.51 ;
      END
   END n_58080

   PIN n_58240
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 192.15 0.51 192.25 ;
      END
   END n_58240

   PIN n_58241
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 171.35 0.51 171.45 ;
      END
   END n_58241

   PIN n_58283
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 108.65 0 108.75 0.51 ;
      END
   END n_58283

   PIN n_58284
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 112.45 0 112.55 0.51 ;
      END
   END n_58284

   PIN n_58286
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 102.65 239.49 102.75 240 ;
      END
   END n_58286

   PIN n_58527
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 134.75 166.8 134.85 ;
      END
   END n_58527

   PIN n_58659
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 120.65 0 120.75 0.51 ;
      END
   END n_58659

   PIN n_58718
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 127.65 239.49 127.75 240 ;
      END
   END n_58718

   PIN n_58790
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 22.65 0 22.75 0.51 ;
      END
   END n_58790

   PIN n_58825
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 179.75 0.51 179.85 ;
      END
   END n_58825

   PIN n_60890
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 202.75 166.8 202.85 ;
      END
   END n_60890

   PIN n_61607
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 162.95 0.51 163.05 ;
      END
   END n_61607

   PIN n_61644
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 119.15 0.51 119.25 ;
      END
   END n_61644

   PIN n_61668
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 161.35 0.51 161.45 ;
      END
   END n_61668

   PIN n_6483
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 37.65 239.49 37.75 240 ;
      END
   END n_6483

   PIN n_65339
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.545 190.9 166.8 191.1 ;
      END
   END n_65339

   PIN n_67179
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 225.55 166.8 225.65 ;
      END
   END n_67179

   PIN n_7530
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 213.75 0.51 213.85 ;
      END
   END n_7530

   PIN n_7532
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 207.55 0.51 207.65 ;
      END
   END n_7532

   PIN n_7534
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 213.15 0.51 213.25 ;
      END
   END n_7534

   PIN n_7535
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 223.95 0.51 224.05 ;
      END
   END n_7535

   PIN n_7538
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 234.55 0.51 234.65 ;
      END
   END n_7538

   PIN n_8012
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 237.35 0.51 237.45 ;
      END
   END n_8012

   PIN n_8483
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 110.05 239.49 110.15 240 ;
      END
   END n_8483

   PIN sub_14999_49_n_82
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 58.15 0.51 58.25 ;
      END
   END sub_14999_49_n_82

   PIN sub_15028_54_n_56
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 136.95 0.51 137.05 ;
      END
   END sub_15028_54_n_56

   PIN sub_15040_54_n_63
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 78.95 0.51 79.05 ;
      END
   END sub_15040_54_n_63

   PIN ternarymux_ln49_0_unr5_z_7__4471875
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 225.35 0.51 225.45 ;
      END
   END ternarymux_ln49_0_unr5_z_7__4471875

   PIN ternarymux_ln49_0_unr7_z_3__4472243
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 202.35 166.8 202.45 ;
      END
   END ternarymux_ln49_0_unr7_z_3__4472243

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 166.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 166.8 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 166.8 8.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 11.745 166.8 12.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 15.745 166.8 16.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 19.745 166.8 20.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 23.745 166.8 24.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 27.745 166.8 28.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 31.745 166.8 32.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 35.745 166.8 36.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 39.745 166.8 40.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 43.745 166.8 44.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 47.745 166.8 48.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 51.745 166.8 52.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 55.745 166.8 56.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 59.745 166.8 60.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 63.745 166.8 64.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 67.745 166.8 68.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 71.745 166.8 72.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 75.745 166.8 76.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 79.745 166.8 80.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 83.745 166.8 84.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 87.745 166.8 88.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 91.745 166.8 92.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 95.745 166.8 96.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 99.745 166.8 100.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 103.745 166.8 104.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 107.745 166.8 108.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 111.745 166.8 112.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 115.745 166.8 116.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 119.745 166.8 120.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 123.745 166.8 124.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 127.745 166.8 128.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 131.745 166.8 132.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 135.745 166.8 136.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 139.745 166.8 140.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 143.745 166.8 144.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 147.745 166.8 148.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 151.745 166.8 152.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 155.745 166.8 156.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 159.745 166.8 160.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 163.745 166.8 164.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 167.745 166.8 168.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 171.745 166.8 172.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 175.745 166.8 176.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 179.745 166.8 180.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 183.745 166.8 184.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 187.745 166.8 188.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 191.745 166.8 192.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 195.745 166.8 196.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 199.745 166.8 200.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 203.745 166.8 204.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 207.745 166.8 208.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 211.745 166.8 212.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 215.745 166.8 216.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 219.745 166.8 220.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 223.745 166.8 224.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 227.745 166.8 228.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 231.745 166.8 232.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 235.745 166.8 236.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 239.745 166.8 240.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 166.8 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 166.8 6.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 9.745 166.8 10.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 13.745 166.8 14.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 17.745 166.8 18.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 21.745 166.8 22.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 25.745 166.8 26.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 29.745 166.8 30.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 33.745 166.8 34.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 37.745 166.8 38.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 41.745 166.8 42.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 45.745 166.8 46.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 49.745 166.8 50.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 53.745 166.8 54.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 57.745 166.8 58.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 61.745 166.8 62.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 65.745 166.8 66.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 69.745 166.8 70.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 73.745 166.8 74.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 77.745 166.8 78.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 81.745 166.8 82.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 85.745 166.8 86.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 89.745 166.8 90.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 93.745 166.8 94.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 97.745 166.8 98.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 101.745 166.8 102.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 105.745 166.8 106.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 109.745 166.8 110.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 113.745 166.8 114.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 117.745 166.8 118.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 121.745 166.8 122.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 125.745 166.8 126.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 129.745 166.8 130.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 133.745 166.8 134.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 137.745 166.8 138.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 141.745 166.8 142.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 145.745 166.8 146.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 149.745 166.8 150.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 153.745 166.8 154.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 157.745 166.8 158.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 161.745 166.8 162.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 165.745 166.8 166.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 169.745 166.8 170.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 173.745 166.8 174.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 177.745 166.8 178.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 181.745 166.8 182.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 185.745 166.8 186.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 189.745 166.8 190.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 193.745 166.8 194.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 197.745 166.8 198.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 201.745 166.8 202.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 205.745 166.8 206.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 209.745 166.8 210.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 213.745 166.8 214.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 217.745 166.8 218.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 221.745 166.8 222.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 225.745 166.8 226.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 229.745 166.8 230.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 233.745 166.8 234.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 237.745 166.8 238.255 ;
      END
   END vdd

   OBS
      LAYER metal1 ;
         RECT 0 0 166.8 240 ;
   END
   OBS
      LAYER metal2 ;
         RECT 0 0 166.8 240 ;
   END
   OBS
      LAYER metal3 ;
         RECT 0 0 166.8 240 ;
   END
   OBS
      LAYER metal4 ;
         RECT 0 0 166.8 240 ;
   END
   OBS
      LAYER metal5 ;
         RECT 0 0 166.8 240 ;
   END
END h4

MACRO h5
   CLASS BLOCK ;
   SIZE 166.8 BY 106 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   PIN FE_OFN37857_n_42354
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 79.35 0.51 79.45 ;
      END
   END FE_OFN37857_n_42354

   PIN FE_OFN38247_n_35860
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 66.35 166.8 66.45 ;
      END
   END FE_OFN38247_n_35860

   PIN FE_OFN38253_n_35857
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.545 56.3 166.8 56.5 ;
      END
   END FE_OFN38253_n_35857

   PIN FE_OFN52040_n_35867
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 78.95 166.8 79.05 ;
      END
   END FE_OFN52040_n_35867

   PIN FE_OFN52045_n_35865
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.545 65.1 166.8 65.3 ;
      END
   END FE_OFN52045_n_35865

   PIN FE_OFN52558_n_35866
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 47.55 166.8 47.65 ;
      END
   END FE_OFN52558_n_35866

   PIN FE_OFN53041_n_35859
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 65.95 166.8 66.05 ;
      END
   END FE_OFN53041_n_35859

   PIN FE_OFN53042_n_35859
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 79.15 166.8 79.25 ;
      END
   END FE_OFN53042_n_35859

   PIN FE_OFN54030_n_50641
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 28.95 166.8 29.05 ;
      END
   END FE_OFN54030_n_50641

   PIN FE_OFN54849_n_35866
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 66.55 166.8 66.65 ;
      END
   END FE_OFN54849_n_35866

   PIN FE_OFN69501_n_50570
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 84.75 166.8 84.85 ;
      END
   END FE_OFN69501_n_50570

   PIN FE_OFN69852_n_50569
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 84.95 166.8 85.05 ;
      END
   END FE_OFN69852_n_50569

   PIN FE_OFN72698_n_34489
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 4.05 105.49 4.15 106 ;
      END
   END FE_OFN72698_n_34489

   PIN FE_OFN87330_n_42357
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 44.05 105.49 44.15 106 ;
      END
   END FE_OFN87330_n_42357

   PIN FE_OFN87336_n_42354
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 84.5 0.255 84.7 ;
      END
   END FE_OFN87336_n_42354

   PIN FE_OFN89085_n_34489
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 42.95 0.51 43.05 ;
      END
   END FE_OFN89085_n_34489

   PIN FE_OFN89086_n_34489
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 54.95 0.51 55.05 ;
      END
   END FE_OFN89086_n_34489

   PIN FE_OFN90160_n_57651
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 61.05 105.49 61.15 106 ;
      END
   END FE_OFN90160_n_57651

   PIN FE_OFN97083_n_50558
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 67.35 166.8 67.45 ;
      END
   END FE_OFN97083_n_50558

   PIN FE_RN_1854_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 38.95 166.8 39.05 ;
      END
   END FE_RN_1854_0

   PIN FE_RN_2772_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 84.55 166.8 84.65 ;
      END
   END FE_RN_2772_0

   PIN n_35857
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.545 65.5 166.8 65.7 ;
      END
   END n_35857

   PIN n_35859
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.545 61.7 166.8 61.9 ;
      END
   END n_35859

   PIN n_35860
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.545 74.7 166.8 74.9 ;
      END
   END n_35860

   PIN n_35861
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.545 46.5 166.8 46.7 ;
      END
   END n_35861

   PIN n_42357
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 97.15 0.51 97.25 ;
      END
   END n_42357

   PIN n_49961
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 49.05 105.49 49.15 106 ;
      END
   END n_49961

   PIN n_49962
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 38.25 105.49 38.35 106 ;
      END
   END n_49962

   PIN n_50542
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 85.15 166.8 85.25 ;
      END
   END n_50542

   PIN n_50543
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 98.35 166.8 98.45 ;
      END
   END n_50543

   PIN n_50544
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 85.35 166.8 85.45 ;
      END
   END n_50544

   PIN n_50552
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 45.95 166.8 46.05 ;
      END
   END n_50552

   PIN n_50559
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 85.55 166.8 85.65 ;
      END
   END n_50559

   PIN n_50561
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 75.15 166.8 75.25 ;
      END
   END n_50561

   PIN n_50565
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 97.95 166.8 98.05 ;
      END
   END n_50565

   PIN n_50566
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 85.75 166.8 85.85 ;
      END
   END n_50566

   PIN n_50571
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 98.15 166.8 98.25 ;
      END
   END n_50571

   PIN n_50588
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 85.95 166.8 86.05 ;
      END
   END n_50588

   PIN n_50664
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 97.55 166.8 97.65 ;
      END
   END n_50664

   PIN n_50670
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 55.25 105.49 55.35 106 ;
      END
   END n_50670

   PIN n_50675
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 42.95 166.8 43.05 ;
      END
   END n_50675

   PIN n_50676
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 27.35 166.8 27.45 ;
      END
   END n_50676

   PIN n_50685
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 9.75 166.8 9.85 ;
      END
   END n_50685

   PIN n_50688
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 147.05 105.49 147.15 106 ;
      END
   END n_50688

   PIN n_50692
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 9.95 166.8 10.05 ;
      END
   END n_50692

   PIN n_50693
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 80.45 105.49 80.55 106 ;
      END
   END n_50693

   PIN n_50695
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 135.85 105.49 135.95 106 ;
      END
   END n_50695

   PIN n_50696
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 17.85 105.49 17.95 106 ;
      END
   END n_50696

   PIN n_50698
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 83.25 105.49 83.35 106 ;
      END
   END n_50698

   PIN n_50699
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 63.15 166.8 63.25 ;
      END
   END n_50699

   PIN n_50700
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 160.25 105.49 160.35 106 ;
      END
   END n_50700

   PIN n_50701
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 10.15 166.8 10.25 ;
      END
   END n_50701

   PIN n_50702
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 92.85 105.49 92.95 106 ;
      END
   END n_50702

   PIN n_50703
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 93.85 105.49 93.95 106 ;
      END
   END n_50703

   PIN n_50704
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 53.65 105.49 53.75 106 ;
      END
   END n_50704

   PIN n_50705
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 27.55 166.8 27.65 ;
      END
   END n_50705

   PIN n_50706
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 10.35 166.8 10.45 ;
      END
   END n_50706

   PIN n_50708
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 66.65 105.49 66.75 106 ;
      END
   END n_50708

   PIN n_50709
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 106.65 105.49 106.75 106 ;
      END
   END n_50709

   PIN n_50711
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 46.15 166.8 46.25 ;
      END
   END n_50711

   PIN n_50712
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 22.25 105.49 22.35 106 ;
      END
   END n_50712

   PIN n_52622
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 161.65 105.49 161.75 106 ;
      END
   END n_52622

   PIN n_52631
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 10.45 105.49 10.55 106 ;
      END
   END n_52631

   PIN n_52632
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 122.65 105.49 122.75 106 ;
      END
   END n_52632

   PIN n_52633
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 110.05 105.49 110.15 106 ;
      END
   END n_52633

   PIN n_52634
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 48.05 105.49 48.15 106 ;
      END
   END n_52634

   PIN n_52635
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 129.05 105.49 129.15 106 ;
      END
   END n_52635

   PIN n_52639
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 136.05 105.49 136.15 106 ;
      END
   END n_52639

   PIN n_52641
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 120.25 105.49 120.35 106 ;
      END
   END n_52641

   PIN n_52661
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 76.05 105.49 76.15 106 ;
      END
   END n_52661

   PIN n_62553
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 19.65 105.49 19.75 106 ;
      END
   END n_62553

   PIN n_62555
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 63.25 105.49 63.35 106 ;
      END
   END n_62555

   PIN n_62557
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 79.75 166.8 79.85 ;
      END
   END n_62557

   PIN n_62559
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 6.65 105.49 6.75 106 ;
      END
   END n_62559

   PIN n_62567
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 101.65 105.49 101.75 106 ;
      END
   END n_62567

   PIN n_62579
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 28.85 105.49 28.95 106 ;
      END
   END n_62579

   PIN n_62581
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 31.05 105.49 31.15 106 ;
      END
   END n_62581

   PIN n_62582
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 82.25 105.49 82.35 106 ;
      END
   END n_62582

   PIN FE_OFN49462_n_35858
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 56.95 166.8 57.05 ;
      END
   END FE_OFN49462_n_35858

   PIN FE_OFN49464_n_35858
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 46.95 166.8 47.05 ;
      END
   END FE_OFN49464_n_35858

   PIN FE_OFN49465_n_35858
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 26.95 166.8 27.05 ;
      END
   END FE_OFN49465_n_35858

   PIN FE_OFN49995_n_42354
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 55.45 105.49 55.55 106 ;
      END
   END FE_OFN49995_n_42354

   PIN FE_OFN52037_n_35867
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.545 44.9 166.8 45.1 ;
      END
   END FE_OFN52037_n_35867

   PIN FE_OFN52042_n_35865
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 47.35 166.8 47.45 ;
      END
   END FE_OFN52042_n_35865

   PIN FE_OFN52416_n_35863
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.545 9.3 166.8 9.5 ;
      END
   END FE_OFN52416_n_35863

   PIN FE_OFN52418_n_35863
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 61.35 166.8 61.45 ;
      END
   END FE_OFN52418_n_35863

   PIN FE_OFN54846_n_35866
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 66.15 166.8 66.25 ;
      END
   END FE_OFN54846_n_35866

   PIN FE_OFN69978_n_46751
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 78.95 0.51 79.05 ;
      END
   END FE_OFN69978_n_46751

   PIN FE_OFN79654_n_47488
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 116.25 105.49 116.35 106 ;
      END
   END FE_OFN79654_n_47488

   PIN FE_OFN87240_n_42521
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 86.15 166.8 86.25 ;
      END
   END FE_OFN87240_n_42521

   PIN FE_OFN87249_n_35860
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 67.15 166.8 67.25 ;
      END
   END FE_OFN87249_n_35860

   PIN FE_OFN87331_n_42357
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 44.25 105.49 44.35 106 ;
      END
   END FE_OFN87331_n_42357

   PIN FE_OFN90096_n_47429
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 118.25 0 118.35 0.51 ;
      END
   END FE_OFN90096_n_47429

   PIN FE_OFN90159_n_57651
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 107.05 105.49 107.15 106 ;
      END
   END FE_OFN90159_n_57651

   PIN FE_OFN95252_n_47584
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 96.95 0.51 97.05 ;
      END
   END FE_OFN95252_n_47584

   PIN FE_RN_1856_0
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 39.35 166.8 39.45 ;
      END
   END FE_RN_1856_0

   PIN FE_RN_5578_0
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 62.95 166.8 63.05 ;
      END
   END FE_RN_5578_0

   PIN n_34489
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 22.75 0.51 22.85 ;
      END
   END n_34489

   PIN n_35863
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 8.95 166.8 9.05 ;
      END
   END n_35863

   PIN n_35865
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 45.35 166.8 45.45 ;
      END
   END n_35865

   PIN n_42516
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.545 78.5 166.8 78.7 ;
      END
   END n_42516

   PIN n_42517
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.545 60.3 166.8 60.5 ;
      END
   END n_42517

   PIN n_42518
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.545 96.5 166.8 96.7 ;
      END
   END n_42518

   PIN n_42520
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 97.35 166.8 97.45 ;
      END
   END n_42520

   PIN n_42522
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.545 96.9 166.8 97.1 ;
      END
   END n_42522

   PIN n_46750
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 84.95 0.51 85.05 ;
      END
   END n_46750

   PIN n_46752
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 75.15 0.51 75.25 ;
      END
   END n_46752

   PIN n_46753
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 66.55 0.51 66.65 ;
      END
   END n_46753

   PIN n_47344
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 25.35 0.51 25.45 ;
      END
   END n_47344

   PIN n_47346
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 48.55 0.51 48.65 ;
      END
   END n_47346

   PIN n_47348
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 48.35 0.51 48.45 ;
      END
   END n_47348

   PIN n_47357
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 66.95 166.8 67.05 ;
      END
   END n_47357

   PIN n_47360
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 79.55 166.8 79.65 ;
      END
   END n_47360

   PIN n_47361
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 9.55 0.51 9.65 ;
      END
   END n_47361

   PIN n_47365
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 30.55 0.51 30.65 ;
      END
   END n_47365

   PIN n_47366
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 79.15 0.51 79.25 ;
      END
   END n_47366

   PIN n_47369
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 45.15 0.51 45.25 ;
      END
   END n_47369

   PIN n_47370
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 61.15 166.8 61.25 ;
      END
   END n_47370

   PIN n_47371
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 22.55 0.51 22.65 ;
      END
   END n_47371

   PIN n_47372
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 9.75 0.51 9.85 ;
      END
   END n_47372

   PIN n_47373
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 25.15 0.51 25.25 ;
      END
   END n_47373

   PIN n_47374
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 61.35 0.51 61.45 ;
      END
   END n_47374

   PIN n_47375
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 22.35 0.51 22.45 ;
      END
   END n_47375

   PIN n_47376
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 27.35 0.51 27.45 ;
      END
   END n_47376

   PIN n_47377
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 27.15 0.51 27.25 ;
      END
   END n_47377

   PIN n_47378
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 48.15 0.51 48.25 ;
      END
   END n_47378

   PIN n_47379
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 39.55 0.51 39.65 ;
      END
   END n_47379

   PIN n_47380
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 9.35 0.51 9.45 ;
      END
   END n_47380

   PIN n_47383
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 61.15 0.51 61.25 ;
      END
   END n_47383

   PIN n_47384
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 39.95 0.51 40.05 ;
      END
   END n_47384

   PIN n_47385
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 66.75 0.51 66.85 ;
      END
   END n_47385

   PIN n_47386
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 75.35 0.51 75.45 ;
      END
   END n_47386

   PIN n_47389
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 30.35 0.51 30.45 ;
      END
   END n_47389

   PIN n_47390
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 44.95 0.51 45.05 ;
      END
   END n_47390

   PIN n_47391
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 22.15 0.51 22.25 ;
      END
   END n_47391

   PIN n_47416
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 46.95 0.51 47.05 ;
      END
   END n_47416

   PIN n_47419
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 46.95 0.51 47.05 ;
      END
   END n_47419

   PIN n_47427
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 21.75 0.51 21.85 ;
      END
   END n_47427

   PIN n_47431
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 30.15 0.51 30.25 ;
      END
   END n_47431

   PIN n_47437
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 45.75 166.8 45.85 ;
      END
   END n_47437

   PIN n_47438
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 45.55 166.8 45.65 ;
      END
   END n_47438

   PIN n_47441
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 39.35 0.51 39.45 ;
      END
   END n_47441

   PIN n_47442
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 39.75 0.51 39.85 ;
      END
   END n_47442

   PIN n_47445
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 21.95 0.51 22.05 ;
      END
   END n_47445

   PIN n_47472
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 12.55 0.51 12.65 ;
      END
   END n_47472

   PIN n_47489
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 26.95 0.51 27.05 ;
      END
   END n_47489

   PIN n_47507
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 60.95 0.51 61.05 ;
      END
   END n_47507

   PIN n_47510
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 57.15 0.51 57.25 ;
      END
   END n_47510

   PIN n_47557
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 21.55 0.51 21.65 ;
      END
   END n_47557

   PIN n_47573
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 39.15 0.51 39.25 ;
      END
   END n_47573

   PIN n_47577
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 9.15 0.51 9.25 ;
      END
   END n_47577

   PIN n_47580
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 24.95 0.51 25.05 ;
      END
   END n_47580

   PIN n_47581
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 8.95 0.51 9.05 ;
      END
   END n_47581

   PIN n_47587
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 148.65 105.49 148.75 106 ;
      END
   END n_47587

   PIN n_47589
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 66.75 166.8 66.85 ;
      END
   END n_47589

   PIN n_47591
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 97.75 166.8 97.85 ;
      END
   END n_47591

   PIN n_50557
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 27.15 166.8 27.25 ;
      END
   END n_50557

   PIN n_50558
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 47.15 166.8 47.25 ;
      END
   END n_50558

   PIN n_50569
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 56.75 166.8 56.85 ;
      END
   END n_50569

   PIN n_50589
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 60.95 166.8 61.05 ;
      END
   END n_50589

   PIN n_50591
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 47.75 166.8 47.85 ;
      END
   END n_50591

   PIN n_50662
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 60.75 166.8 60.85 ;
      END
   END n_50662

   PIN n_50667
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 166.29 79.35 166.8 79.45 ;
      END
   END n_50667

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 166.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 166.8 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 166.8 8.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 11.745 166.8 12.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 15.745 166.8 16.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 19.745 166.8 20.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 23.745 166.8 24.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 27.745 166.8 28.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 31.745 166.8 32.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 35.745 166.8 36.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 39.745 166.8 40.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 43.745 166.8 44.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 47.745 166.8 48.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 51.745 166.8 52.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 55.745 166.8 56.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 59.745 166.8 60.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 63.745 166.8 64.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 67.745 166.8 68.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 71.745 166.8 72.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 75.745 166.8 76.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 79.745 166.8 80.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 83.745 166.8 84.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 87.745 166.8 88.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 91.745 166.8 92.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 95.745 166.8 96.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 99.745 166.8 100.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 103.745 166.8 104.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 166.8 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 166.8 6.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 9.745 166.8 10.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 13.745 166.8 14.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 17.745 166.8 18.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 21.745 166.8 22.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 25.745 166.8 26.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 29.745 166.8 30.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 33.745 166.8 34.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 37.745 166.8 38.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 41.745 166.8 42.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 45.745 166.8 46.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 49.745 166.8 50.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 53.745 166.8 54.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 57.745 166.8 58.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 61.745 166.8 62.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 65.745 166.8 66.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 69.745 166.8 70.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 73.745 166.8 74.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 77.745 166.8 78.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 81.745 166.8 82.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 85.745 166.8 86.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 89.745 166.8 90.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 93.745 166.8 94.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 97.745 166.8 98.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 101.745 166.8 102.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 105.745 166.8 106.255 ;
      END
   END vdd

   OBS
      LAYER metal1 ;
         RECT 0 0 166.8 106 ;
   END
   OBS
      LAYER metal2 ;
         RECT 0 0 166.8 106 ;
   END
   OBS
      LAYER metal3 ;
         RECT 0 0 166.8 106 ;
   END
   OBS
      LAYER metal4 ;
         RECT 0 0 166.8 106 ;
   END
   OBS
      LAYER metal5 ;
         RECT 0 0 166.8 106 ;
   END
END h5

MACRO h6
   CLASS BLOCK ;
   SIZE 161.4 BY 186 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   PIN FE_OCPN58665_n_40293
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 23.45 185.49 23.55 186 ;
      END
   END FE_OCPN58665_n_40293

   PIN FE_OCPN58699_n_40977
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 95.75 0.51 95.85 ;
      END
   END FE_OCPN58699_n_40977

   PIN FE_OCPN59731_n_40871
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 95.95 0.51 96.05 ;
      END
   END FE_OCPN59731_n_40871

   PIN FE_OCPN59829_FE_OFN27411_n_40407
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 141.55 161.4 141.65 ;
      END
   END FE_OCPN59829_FE_OFN27411_n_40407

   PIN FE_OCPN60004_n_40991
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 91.55 0.51 91.65 ;
      END
   END FE_OCPN60004_n_40991

   PIN FE_OCPN60013_n_40453
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 149.45 185.49 149.55 186 ;
      END
   END FE_OCPN60013_n_40453

   PIN FE_OCPN60445_n_40884
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 93.75 0.51 93.85 ;
      END
   END FE_OCPN60445_n_40884

   PIN FE_OCPN60817_FE_OFN50247_n_40462
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 77.15 161.4 77.25 ;
      END
   END FE_OCPN60817_FE_OFN50247_n_40462

   PIN FE_OCPN60825_n_40739
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 107.15 0.51 107.25 ;
      END
   END FE_OCPN60825_n_40739

   PIN FE_OCPN60829_n_40773
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 134.95 161.4 135.05 ;
      END
   END FE_OCPN60829_n_40773

   PIN FE_OCPN60889_n_40624
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 96.55 161.4 96.65 ;
      END
   END FE_OCPN60889_n_40624

   PIN FE_OCPN60892_n_40626
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 92.95 161.4 93.05 ;
      END
   END FE_OCPN60892_n_40626

   PIN FE_OCPN60896_n_40916
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 122.75 0.51 122.85 ;
      END
   END FE_OCPN60896_n_40916

   PIN FE_OCPN61157_n_40452
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 94.95 0.51 95.05 ;
      END
   END FE_OCPN61157_n_40452

   PIN FE_OCPN61165_n_40736
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 114.95 0.51 115.05 ;
      END
   END FE_OCPN61165_n_40736

   PIN FE_OCPN61186_n_40442
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 96.35 161.4 96.45 ;
      END
   END FE_OCPN61186_n_40442

   PIN FE_OCPN61190_n_40385
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 104.35 0.51 104.45 ;
      END
   END FE_OCPN61190_n_40385

   PIN FE_OCPN61194_n_40543
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 95.15 0.51 95.25 ;
      END
   END FE_OCPN61194_n_40543

   PIN FE_OCPN61198_FE_OFN4340_n_40574
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 67.85 185.49 67.95 186 ;
      END
   END FE_OCPN61198_FE_OFN4340_n_40574

   PIN FE_OCPN61200_FE_OFN26050_n_40461
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 150.55 161.4 150.65 ;
      END
   END FE_OCPN61200_FE_OFN26050_n_40461

   PIN FE_OCPN61205_n_40748
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 96.15 0.51 96.25 ;
      END
   END FE_OCPN61205_n_40748

   PIN FE_OCPN61340_n_40638
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 113.45 185.49 113.55 186 ;
      END
   END FE_OCPN61340_n_40638

   PIN FE_OCPN61708_n_40671
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 168.95 0.51 169.05 ;
      END
   END FE_OCPN61708_n_40671

   PIN FE_OCPN62299_FE_OFN53822_n_40455
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 114.55 0.51 114.65 ;
      END
   END FE_OCPN62299_FE_OFN53822_n_40455

   PIN FE_OCPN62464_n_40460
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 63.95 0.51 64.05 ;
      END
   END FE_OCPN62464_n_40460

   PIN FE_OCPN62757_n_40522
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 150.15 0.51 150.25 ;
      END
   END FE_OCPN62757_n_40522

   PIN FE_OCPN62762_n_40389
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 162.95 161.4 163.05 ;
      END
   END FE_OCPN62762_n_40389

   PIN FE_OCPN62778_n_40539
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 167.95 0.51 168.05 ;
      END
   END FE_OCPN62778_n_40539

   PIN FE_OCPN63314_n_40689
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 35.75 0.51 35.85 ;
      END
   END FE_OCPN63314_n_40689

   PIN FE_OCPN63402_n_40695
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 77.05 185.49 77.15 186 ;
      END
   END FE_OCPN63402_n_40695

   PIN FE_OCPN63686_n_40655
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 68.25 185.49 68.35 186 ;
      END
   END FE_OCPN63686_n_40655

   PIN FE_OCPN63879_n_40667
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 100.25 185.49 100.35 186 ;
      END
   END FE_OCPN63879_n_40667

   PIN FE_OCPN76175_n_40685
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 31.85 185.49 31.95 186 ;
      END
   END FE_OCPN76175_n_40685

   PIN FE_OCPN76176_n_40685
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 131.45 185.49 131.55 186 ;
      END
   END FE_OCPN76176_n_40685

   PIN FE_OCPN76225_n_40728
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 49.55 0.51 49.65 ;
      END
   END FE_OCPN76225_n_40728

   PIN FE_OCPN76871_n_40344
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 140.15 0.51 140.25 ;
      END
   END FE_OCPN76871_n_40344

   PIN FE_OCPN76899_n_40732
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 21.15 0.51 21.25 ;
      END
   END FE_OCPN76899_n_40732

   PIN FE_OCPN77057_n_40646
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 64.75 0.51 64.85 ;
      END
   END FE_OCPN77057_n_40646

   PIN FE_OCPN77058_n_40646
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 77.55 0.51 77.65 ;
      END
   END FE_OCPN77058_n_40646

   PIN FE_OCPN78169_n_40634
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 104.25 185.49 104.35 186 ;
      END
   END FE_OCPN78169_n_40634

   PIN FE_OCPN78237_FE_OFN3733_n_40730
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 50.75 0.51 50.85 ;
      END
   END FE_OCPN78237_FE_OFN3733_n_40730

   PIN FE_OCPN95535_n_40744
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 132.35 161.4 132.45 ;
      END
   END FE_OCPN95535_n_40744

   PIN FE_OCPN95538_FE_OFN90000_n_40684
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 59.55 0.51 59.65 ;
      END
   END FE_OCPN95538_FE_OFN90000_n_40684

   PIN FE_OCPN95613_FE_OFN89862_n_40309
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 123.15 161.4 123.25 ;
      END
   END FE_OCPN95613_FE_OFN89862_n_40309

   PIN FE_OCPN95619_n_40607
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 148.95 161.4 149.05 ;
      END
   END FE_OCPN95619_n_40607

   PIN FE_OCPN95761_n_40465
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 122.25 185.49 122.35 186 ;
      END
   END FE_OCPN95761_n_40465

   PIN FE_OCPN95853_FE_OFN90041_n_40381
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 160.89 178.95 161.4 179.05 ;
      END
   END FE_OCPN95853_FE_OFN90041_n_40381

   PIN FE_OCP_DRV_N76452_FE_OFN67430_n_40505
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 86.55 0.51 86.65 ;
      END
   END FE_OCP_DRV_N76452_FE_OFN67430_n_40505

   PIN FE_OCP_DRV_N76464_FE_OFN66917_n_40672
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 141.75 161.4 141.85 ;
      END
   END FE_OCP_DRV_N76464_FE_OFN66917_n_40672

   PIN FE_OCP_DRV_N78200_FE_OFN37047_n_35919
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 35.15 0.51 35.25 ;
      END
   END FE_OCP_DRV_N78200_FE_OFN37047_n_35919

   PIN FE_OFN3336_n_57614
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 6.25 185.49 6.35 186 ;
      END
   END FE_OFN3336_n_57614

   PIN FE_OFN35849_n_52031
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 59.85 185.49 59.95 186 ;
      END
   END FE_OFN35849_n_52031

   PIN FE_OFN35858_n_52027
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 69.85 185.49 69.95 186 ;
      END
   END FE_OFN35858_n_52027

   PIN FE_OFN35873_n_52030
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 41.05 185.49 41.15 186 ;
      END
   END FE_OFN35873_n_52030

   PIN FE_OFN35875_n_52030
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 15.25 185.49 15.35 186 ;
      END
   END FE_OFN35875_n_52030

   PIN FE_OFN35909_n_52083
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 42.35 0.51 42.45 ;
      END
   END FE_OFN35909_n_52083

   PIN FE_OFN35925_n_52086
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 62.95 0.51 63.05 ;
      END
   END FE_OFN35925_n_52086

   PIN FE_OFN35933_n_52028
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 112.65 185.49 112.75 186 ;
      END
   END FE_OFN35933_n_52028

   PIN FE_OFN35937_n_52028
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 17.2 185.745 17.4 186 ;
      END
   END FE_OFN35937_n_52028

   PIN FE_OFN36907_n_35904
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 148.95 0.51 149.05 ;
      END
   END FE_OFN36907_n_35904

   PIN FE_OFN36908_n_35904
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 59.8 185.745 60 186 ;
      END
   END FE_OFN36908_n_35904

   PIN FE_OFN36982_n_45345
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 41.85 185.49 41.95 186 ;
      END
   END FE_OFN36982_n_45345

   PIN FE_OFN37047_n_35919
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 41.75 0.51 41.85 ;
      END
   END FE_OFN37047_n_35919

   PIN FE_OFN4914_n_56419
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 141.75 0.51 141.85 ;
      END
   END FE_OFN4914_n_56419

   PIN FE_OFN50279_n_52028
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 76.95 0.51 77.05 ;
      END
   END FE_OFN50279_n_52028

   PIN FE_OFN50280_n_52028
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 132.55 0.51 132.65 ;
      END
   END FE_OFN50280_n_52028

   PIN FE_OFN50334_n_52030
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 60.05 185.49 60.15 186 ;
      END
   END FE_OFN50334_n_52030

   PIN FE_OFN50335_n_52030
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 86.15 0.51 86.25 ;
      END
   END FE_OFN50335_n_52030

   PIN FE_OFN53021_n_40337
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 121.75 0.51 121.85 ;
      END
   END FE_OFN53021_n_40337

   PIN FE_OFN53588_n_40797
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 60.55 161.4 60.65 ;
      END
   END FE_OFN53588_n_40797

   PIN FE_OFN53589_n_40797
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 69.75 0.51 69.85 ;
      END
   END FE_OFN53589_n_40797

   PIN FE_OFN53785_n_52084
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 50.35 0.51 50.45 ;
      END
   END FE_OFN53785_n_52084

   PIN FE_OFN53787_n_52080
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 27.05 185.49 27.15 186 ;
      END
   END FE_OFN53787_n_52080

   PIN FE_OFN53788_n_52080
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 141.95 0.51 142.05 ;
      END
   END FE_OFN53788_n_52080

   PIN FE_OFN53789_n_52080
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 40.45 185.49 40.55 186 ;
      END
   END FE_OFN53789_n_52080

   PIN FE_OFN53790_n_52080
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 96.75 0.51 96.85 ;
      END
   END FE_OFN53790_n_52080

   PIN FE_OFN53791_n_52027
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 43.75 0.51 43.85 ;
      END
   END FE_OFN53791_n_52027

   PIN FE_OFN53792_n_52027
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 77.45 185.49 77.55 186 ;
      END
   END FE_OFN53792_n_52027

   PIN FE_OFN53795_n_52027
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 42.05 185.49 42.15 186 ;
      END
   END FE_OFN53795_n_52027

   PIN FE_OFN53796_n_52087
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 85.95 0.51 86.05 ;
      END
   END FE_OFN53796_n_52087

   PIN FE_OFN53797_n_52087
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 41.6 185.745 41.8 186 ;
      END
   END FE_OFN53797_n_52087

   PIN FE_OFN53798_n_52087
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 41.25 185.49 41.35 186 ;
      END
   END FE_OFN53798_n_52087

   PIN FE_OFN53806_n_52029
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 17.85 185.49 17.95 186 ;
      END
   END FE_OFN53806_n_52029

   PIN FE_OFN53807_n_52029
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 105.95 0.51 106.05 ;
      END
   END FE_OFN53807_n_52029

   PIN FE_OFN53808_n_52029
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 77.8 185.745 78 186 ;
      END
   END FE_OFN53808_n_52029

   PIN FE_OFN53810_n_52029
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 120.05 185.49 120.15 186 ;
      END
   END FE_OFN53810_n_52029

   PIN FE_OFN53813_n_52029
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 107.35 0.51 107.45 ;
      END
   END FE_OFN53813_n_52029

   PIN FE_OFN53847_n_52031
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 32.85 185.49 32.95 186 ;
      END
   END FE_OFN53847_n_52031

   PIN FE_OFN53848_n_52031
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 62.95 0.51 63.05 ;
      END
   END FE_OFN53848_n_52031

   PIN FE_OFN53852_n_52081
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 168.55 0.51 168.65 ;
      END
   END FE_OFN53852_n_52081

   PIN FE_OFN53929_n_52024
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 142.55 0.51 142.65 ;
      END
   END FE_OFN53929_n_52024

   PIN FE_OFN53930_n_52024
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 14.85 185.49 14.95 186 ;
      END
   END FE_OFN53930_n_52024

   PIN FE_OFN53951_n_40618
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 76.95 161.4 77.05 ;
      END
   END FE_OFN53951_n_40618

   PIN FE_OFN53970_n_40476
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 49.75 0.51 49.85 ;
      END
   END FE_OFN53970_n_40476

   PIN FE_OFN53975_n_52082
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 93.95 0.51 94.05 ;
      END
   END FE_OFN53975_n_52082

   PIN FE_OFN53976_n_52082
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 122.95 0.51 123.05 ;
      END
   END FE_OFN53976_n_52082

   PIN FE_OFN54053_n_53997
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 7.75 0.51 7.85 ;
      END
   END FE_OFN54053_n_53997

   PIN FE_OFN55531_n_45338
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 32.45 185.49 32.55 186 ;
      END
   END FE_OFN55531_n_45338

   PIN FE_OFN55721_n_52025
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 129.45 185.49 129.55 186 ;
      END
   END FE_OFN55721_n_52025

   PIN FE_OFN55722_n_52025
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 77.95 0.51 78.05 ;
      END
   END FE_OFN55722_n_52025

   PIN FE_OFN55723_n_52025
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 158.75 0.51 158.85 ;
      END
   END FE_OFN55723_n_52025

   PIN FE_OFN55724_n_52025
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 49.85 185.49 49.95 186 ;
      END
   END FE_OFN55724_n_52025

   PIN FE_OFN55763_n_52086
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 23.25 185.49 23.35 186 ;
      END
   END FE_OFN55763_n_52086

   PIN FE_OFN55765_n_52086
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 59.4 185.745 59.6 186 ;
      END
   END FE_OFN55765_n_52086

   PIN FE_OFN55829_n_52085
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 6.65 185.49 6.75 186 ;
      END
   END FE_OFN55829_n_52085

   PIN FE_OFN55830_n_52085
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 42.25 185.49 42.35 186 ;
      END
   END FE_OFN55830_n_52085

   PIN FE_OFN55832_n_52085
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 51.75 0.51 51.85 ;
      END
   END FE_OFN55832_n_52085

   PIN FE_OFN64709_n_40441
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 149.65 185.49 149.75 186 ;
      END
   END FE_OFN64709_n_40441

   PIN FE_OFN64798_n_40578
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 66.85 185.49 66.95 186 ;
      END
   END FE_OFN64798_n_40578

   PIN FE_OFN64923_n_40587
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 77.25 185.49 77.35 186 ;
      END
   END FE_OFN64923_n_40587

   PIN FE_OFN67632_n_40380
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 69.95 0.51 70.05 ;
      END
   END FE_OFN67632_n_40380

   PIN FE_OFN67675_n_41246
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 41.95 0.51 42.05 ;
      END
   END FE_OFN67675_n_41246

   PIN FE_OFN68512_n_40584
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 59.05 185.49 59.15 186 ;
      END
   END FE_OFN68512_n_40584

   PIN FE_OFN68513_n_40584
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 64.15 0.51 64.25 ;
      END
   END FE_OFN68513_n_40584

   PIN FE_OFN68659_n_41001
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 177.75 0.51 177.85 ;
      END
   END FE_OFN68659_n_41001

   PIN FE_OFN68752_n_40468
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 59.25 185.49 59.35 186 ;
      END
   END FE_OFN68752_n_40468

   PIN FE_OFN69011_n_40742
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 135.15 161.4 135.25 ;
      END
   END FE_OFN69011_n_40742

   PIN FE_OFN69206_n_40725
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 68.35 0.51 68.45 ;
      END
   END FE_OFN69206_n_40725

   PIN FE_OFN69664_n_40499
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 77.35 0.51 77.45 ;
      END
   END FE_OFN69664_n_40499

   PIN FE_OFN69889_n_40422
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 96.95 0.51 97.05 ;
      END
   END FE_OFN69889_n_40422

   PIN FE_OFN70042_n_40615
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 77.25 185.49 77.35 186 ;
      END
   END FE_OFN70042_n_40615

   PIN FE_OFN79586_n_40690
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 50.25 185.49 50.35 186 ;
      END
   END FE_OFN79586_n_40690

   PIN FE_OFN79626_n_40616
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 160.89 159.55 161.4 159.65 ;
      END
   END FE_OFN79626_n_40616

   PIN FE_OFN80551_n_41085
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 150.35 161.4 150.45 ;
      END
   END FE_OFN80551_n_41085

   PIN FE_OFN81546_n_40579
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 114.55 161.4 114.65 ;
      END
   END FE_OFN81546_n_40579

   PIN FE_OFN82254_n_40562
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 65.35 0.51 65.45 ;
      END
   END FE_OFN82254_n_40562

   PIN FE_OFN82720_n_40745
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 159.35 0.51 159.45 ;
      END
   END FE_OFN82720_n_40745

   PIN FE_OFN84632_n_45520
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 167.55 161.4 167.65 ;
      END
   END FE_OFN84632_n_45520

   PIN FE_OFN89562_n_40600
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 159.55 0.51 159.65 ;
      END
   END FE_OFN89562_n_40600

   PIN FE_OFN89690_n_40666
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 121.15 161.4 121.25 ;
      END
   END FE_OFN89690_n_40666

   PIN FE_OFN89775_n_40818
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 132.75 0.51 132.85 ;
      END
   END FE_OFN89775_n_40818

   PIN FE_OFN89783_n_41094
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 79.95 0.51 80.05 ;
      END
   END FE_OFN89783_n_41094

   PIN FE_OFN89834_n_40765
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 22.05 185.49 22.15 186 ;
      END
   END FE_OFN89834_n_40765

   PIN FE_OFN89889_n_40579
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 78.35 161.4 78.45 ;
      END
   END FE_OFN89889_n_40579

   PIN FE_OFN89896_n_40690
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 95.25 185.49 95.35 186 ;
      END
   END FE_OFN89896_n_40690

   PIN FE_OFN89931_n_41129
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 123.25 185.49 123.35 186 ;
      END
   END FE_OFN89931_n_41129

   PIN FE_OFN89946_n_40368
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 70.15 0.51 70.25 ;
      END
   END FE_OFN89946_n_40368

   PIN FE_OFN89969_n_40791
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 151.25 185.49 151.35 186 ;
      END
   END FE_OFN89969_n_40791

   PIN FE_OFN89991_n_40449
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 42.55 0.51 42.65 ;
      END
   END FE_OFN89991_n_40449

   PIN FE_OFN89995_n_40526
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 131.65 185.49 131.75 186 ;
      END
   END FE_OFN89995_n_40526

   PIN FE_OFN89996_n_40526
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 121.35 161.4 121.45 ;
      END
   END FE_OFN89996_n_40526

   PIN FE_OFN90072_FE_OCPN57974_n_40531
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 132.55 161.4 132.65 ;
      END
   END FE_OFN90072_FE_OCPN57974_n_40531

   PIN FE_OFN90077_n_40436
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 76.85 185.49 76.95 186 ;
      END
   END FE_OFN90077_n_40436

   PIN FE_OFN90083_n_40637
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 142.15 0.51 142.25 ;
      END
   END FE_OFN90083_n_40637

   PIN FE_OFN92416_n_40768
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 132.95 0.51 133.05 ;
      END
   END FE_OFN92416_n_40768

   PIN FE_OFN92692_n_40849
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 42.75 0.51 42.85 ;
      END
   END FE_OFN92692_n_40849

   PIN FE_OFN92693_n_40849
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 42.95 0.51 43.05 ;
      END
   END FE_OFN92693_n_40849

   PIN FE_OFN92898_n_40770
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 119.55 0.51 119.65 ;
      END
   END FE_OFN92898_n_40770

   PIN FE_OFN93228_n_40835
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 77.75 0.51 77.85 ;
      END
   END FE_OFN93228_n_40835

   PIN FE_OFN95235_n_40680
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 78.15 0.51 78.25 ;
      END
   END FE_OFN95235_n_40680

   PIN FE_OFN95251_n_40692
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 97.65 185.49 97.75 186 ;
      END
   END FE_OFN95251_n_40692

   PIN FE_OFN95268_n_40689
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 35.95 0.51 36.05 ;
      END
   END FE_OFN95268_n_40689

   PIN FE_OFN96061_FE_OCPN59260_n_40732
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 59.15 0.51 59.25 ;
      END
   END FE_OFN96061_FE_OCPN59260_n_40732

   PIN FE_OFN96635_n_41231
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 114.75 0.51 114.85 ;
      END
   END FE_OFN96635_n_41231

   PIN FE_OFN96853_FE_OCPN61163_n_40472
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 96.35 0.51 96.45 ;
      END
   END FE_OFN96853_FE_OCPN61163_n_40472

   PIN FE_OFN96935_n_40586
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 151.15 0.51 151.25 ;
      END
   END FE_OFN96935_n_40586

   PIN FE_OFN96959_n_40592
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 86.25 185.49 86.35 186 ;
      END
   END FE_OFN96959_n_40592

   PIN FE_OFN97148_n_41111
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 106.15 0.51 106.25 ;
      END
   END FE_OFN97148_n_41111

   PIN FE_OFN97292_n_40798
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 86.45 185.49 86.55 186 ;
      END
   END FE_OFN97292_n_40798

   PIN FE_OFN97614_FE_OCPN61281_n_40613
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 86.45 185.49 86.55 186 ;
      END
   END FE_OFN97614_FE_OCPN61281_n_40613

   PIN FE_RN_3275_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 77.45 185.49 77.55 186 ;
      END
   END FE_RN_3275_0

   PIN FE_RN_3761_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 78.35 0.51 78.45 ;
      END
   END FE_RN_3761_0

   PIN FE_RN_541_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 31.25 185.49 31.35 186 ;
      END
   END FE_RN_541_0

   PIN n_44333
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 159.55 161.4 159.65 ;
      END
   END n_44333

   PIN n_44349
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 159.75 161.4 159.85 ;
      END
   END n_44349

   PIN n_44353
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 19.85 185.49 19.95 186 ;
      END
   END n_44353

   PIN n_44354
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 140.45 185.49 140.55 186 ;
      END
   END n_44354

   PIN n_44355
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 20.95 161.4 21.05 ;
      END
   END n_44355

   PIN n_44356
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 6.95 161.4 7.05 ;
      END
   END n_44356

   PIN n_44359
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 149.15 161.4 149.25 ;
      END
   END n_44359

   PIN n_44383
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 107.15 161.4 107.25 ;
      END
   END n_44383

   PIN n_44384
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 116.85 185.49 116.95 186 ;
      END
   END n_44384

   PIN n_45336
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 41.45 185.49 41.55 186 ;
      END
   END n_45336

   PIN n_45339
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 23.45 185.49 23.55 186 ;
      END
   END n_45339

   PIN n_45342
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 106.65 185.49 106.75 186 ;
      END
   END n_45342

   PIN n_45343
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 24.85 185.49 24.95 186 ;
      END
   END n_45343

   PIN n_45344
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 142.95 0.51 143.05 ;
      END
   END n_45344

   PIN n_45346
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 41.65 185.49 41.75 186 ;
      END
   END n_45346

   PIN n_52024
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 59.45 185.49 59.55 186 ;
      END
   END n_52024

   PIN n_52082
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 78.05 185.49 78.15 186 ;
      END
   END n_52082

   PIN n_53966
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 70.75 0.51 70.85 ;
      END
   END n_53966

   PIN n_53968
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 88.15 0.51 88.25 ;
      END
   END n_53968

   PIN n_53995
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 80.15 0.51 80.25 ;
      END
   END n_53995

   PIN n_53996
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 78.55 0.51 78.65 ;
      END
   END n_53996

   PIN n_54003
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 50.45 185.49 50.55 186 ;
      END
   END n_54003

   PIN n_54014
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 41.25 185.49 41.35 186 ;
      END
   END n_54014

   PIN n_54043
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 51.55 0.51 51.65 ;
      END
   END n_54043

   PIN n_54057
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 64.35 0.51 64.45 ;
      END
   END n_54057

   PIN n_54098
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 135.55 0.51 135.65 ;
      END
   END n_54098

   PIN n_54186
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 22.65 185.49 22.75 186 ;
      END
   END n_54186

   PIN n_54198
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 15.05 185.49 15.15 186 ;
      END
   END n_54198

   PIN n_54215
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 15.65 185.49 15.75 186 ;
      END
   END n_54215

   PIN n_54238
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 22.85 185.49 22.95 186 ;
      END
   END n_54238

   PIN n_54239
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 23.05 185.49 23.15 186 ;
      END
   END n_54239

   PIN n_56417
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 58.85 185.49 58.95 186 ;
      END
   END n_56417

   PIN n_56423
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 6.45 185.49 6.55 186 ;
      END
   END n_56423

   PIN n_56424
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 5.45 185.49 5.55 186 ;
      END
   END n_56424

   PIN n_56425
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 114.55 0.51 114.65 ;
      END
   END n_56425

   PIN n_56426
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 123.15 0.51 123.25 ;
      END
   END n_56426

   PIN n_56429
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 34.95 0.51 35.05 ;
      END
   END n_56429

   PIN n_57591
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 77.85 185.49 77.95 186 ;
      END
   END n_57591

   PIN n_58389
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 121.95 0.51 122.05 ;
      END
   END n_58389

   PIN n_58593
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 5.65 185.49 5.75 186 ;
      END
   END n_58593

   PIN n_58665
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 178.95 0.51 179.05 ;
      END
   END n_58665

   PIN FE_OCPN57928_n_40786
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 63.75 0.51 63.85 ;
      END
   END FE_OCPN57928_n_40786

   PIN FE_OCPN57974_n_40531
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 22.15 0.51 22.25 ;
      END
   END FE_OCPN57974_n_40531

   PIN FE_OCPN58664_n_40293
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 49.95 0.51 50.05 ;
      END
   END FE_OCPN58664_n_40293

   PIN FE_OCPN58691_n_40304
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 60.55 0.51 60.65 ;
      END
   END FE_OCPN58691_n_40304

   PIN FE_OCPN58698_n_40977
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 51.35 0.51 51.45 ;
      END
   END FE_OCPN58698_n_40977

   PIN FE_OCPN59256_n_40667
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 179.15 0.51 179.25 ;
      END
   END FE_OCPN59256_n_40667

   PIN FE_OCPN59258_n_40370
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 87.55 0.51 87.65 ;
      END
   END FE_OCPN59258_n_40370

   PIN FE_OCPN59262_n_40728
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 41.55 0.51 41.65 ;
      END
   END FE_OCPN59262_n_40728

   PIN FE_OCPN59729_n_40871
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 91.35 0.51 91.45 ;
      END
   END FE_OCPN59729_n_40871

   PIN FE_OCPN59744_n_40606
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 7.55 0.51 7.65 ;
      END
   END FE_OCPN59744_n_40606

   PIN FE_OCPN59823_n_40673
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 52.25 185.49 52.35 186 ;
      END
   END FE_OCPN59823_n_40673

   PIN FE_OCPN59828_FE_OFN27411_n_40407
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 115.55 0.51 115.65 ;
      END
   END FE_OCPN59828_FE_OFN27411_n_40407

   PIN FE_OCPN59987_n_40388
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 72.15 0.51 72.25 ;
      END
   END FE_OCPN59987_n_40388

   PIN FE_OCPN60002_n_40991
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 91.15 0.51 91.25 ;
      END
   END FE_OCPN60002_n_40991

   PIN FE_OCPN60011_n_40453
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 82.05 185.49 82.15 186 ;
      END
   END FE_OCPN60011_n_40453

   PIN FE_OCPN60444_n_40884
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 93.55 0.51 93.65 ;
      END
   END FE_OCPN60444_n_40884

   PIN FE_OCPN60815_FE_OFN50247_n_40462
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 93.15 0.51 93.25 ;
      END
   END FE_OCPN60815_FE_OFN50247_n_40462

   PIN FE_OCPN60824_n_40739
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 114.35 0.51 114.45 ;
      END
   END FE_OCPN60824_n_40739

   PIN FE_OCPN60827_n_40753
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 120.95 161.4 121.05 ;
      END
   END FE_OCPN60827_n_40753

   PIN FE_OCPN60828_n_40773
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 135.35 0.51 135.45 ;
      END
   END FE_OCPN60828_n_40773

   PIN FE_OCPN60887_n_40624
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 107.35 0.51 107.45 ;
      END
   END FE_OCPN60887_n_40624

   PIN FE_OCPN60890_n_40626
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 92.95 0.51 93.05 ;
      END
   END FE_OCPN60890_n_40626

   PIN FE_OCPN60895_n_40916
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 106.95 0.51 107.05 ;
      END
   END FE_OCPN60895_n_40916

   PIN FE_OCPN60898_FE_OFN3733_n_40730
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 7.35 0.51 7.45 ;
      END
   END FE_OCPN60898_FE_OFN3733_n_40730

   PIN FE_OCPN61161_n_40733
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 50.55 0.51 50.65 ;
      END
   END FE_OCPN61161_n_40733

   PIN FE_OCPN61163_n_40472
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 90.95 0.51 91.05 ;
      END
   END FE_OCPN61163_n_40472

   PIN FE_OCPN61164_n_40736
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 105.35 0.51 105.45 ;
      END
   END FE_OCPN61164_n_40736

   PIN FE_OCPN61170_n_40664
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 14.65 185.49 14.75 186 ;
      END
   END FE_OCPN61170_n_40664

   PIN FE_OCPN61178_n_40494
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 79.15 0.51 79.25 ;
      END
   END FE_OCPN61178_n_40494

   PIN FE_OCPN61180_FE_OFN26782_n_40493
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 106.95 161.4 107.05 ;
      END
   END FE_OCPN61180_FE_OFN26782_n_40493

   PIN FE_OCPN61184_n_40665
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 167.75 0.51 167.85 ;
      END
   END FE_OCPN61184_n_40665

   PIN FE_OCPN61188_n_40458
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 105.75 0.51 105.85 ;
      END
   END FE_OCPN61188_n_40458

   PIN FE_OCPN61189_n_40385
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 49.35 0.51 49.45 ;
      END
   END FE_OCPN61189_n_40385

   PIN FE_OCPN61193_n_40543
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 59.35 0.51 59.45 ;
      END
   END FE_OCPN61193_n_40543

   PIN FE_OCPN61197_FE_OFN4340_n_40574
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 22.95 0.51 23.05 ;
      END
   END FE_OCPN61197_FE_OFN4340_n_40574

   PIN FE_OCPN61199_FE_OFN26050_n_40461
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 135.15 0.51 135.25 ;
      END
   END FE_OCPN61199_FE_OFN26050_n_40461

   PIN FE_OCPN61202_n_40700
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 141.55 0.51 141.65 ;
      END
   END FE_OCPN61202_n_40700

   PIN FE_OCPN61281_n_40613
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 169.15 0.51 169.25 ;
      END
   END FE_OCPN61281_n_40613

   PIN FE_OCPN61334_n_40487
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 77.15 0.51 77.25 ;
      END
   END FE_OCPN61334_n_40487

   PIN FE_OCPN61703_n_40614
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 87.35 0.51 87.45 ;
      END
   END FE_OCPN61703_n_40614

   PIN FE_OCPN61705_n_40652
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 87.15 0.51 87.25 ;
      END
   END FE_OCPN61705_n_40652

   PIN FE_OCPN61706_n_40671
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 168.75 0.51 168.85 ;
      END
   END FE_OCPN61706_n_40671

   PIN FE_OCPN61855_FE_OFN53951_n_40618
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 78.55 161.4 78.65 ;
      END
   END FE_OCPN61855_FE_OFN53951_n_40618

   PIN FE_OCPN61880_FE_OFN21562_n_40405
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 160.15 0.51 160.25 ;
      END
   END FE_OCPN61880_FE_OFN21562_n_40405

   PIN FE_OCPN61918_FE_OFN53968_n_40476
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 49.15 0.51 49.25 ;
      END
   END FE_OCPN61918_FE_OFN53968_n_40476

   PIN FE_OCPN62235_n_40789
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 93.35 0.51 93.45 ;
      END
   END FE_OCPN62235_n_40789

   PIN FE_OCPN62246_n_40447
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 7.15 0.51 7.25 ;
      END
   END FE_OCPN62246_n_40447

   PIN FE_OCPN62248_n_40471
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 32.25 185.49 32.35 186 ;
      END
   END FE_OCPN62248_n_40471

   PIN FE_OCPN62288_FE_OFN53950_n_40618
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 92.95 0.51 93.05 ;
      END
   END FE_OCPN62288_FE_OFN53950_n_40618

   PIN FE_OCPN62466_n_40460
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 15.55 0.51 15.65 ;
      END
   END FE_OCPN62466_n_40460

   PIN FE_OCPN62755_n_40522
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 114.15 0.51 114.25 ;
      END
   END FE_OCPN62755_n_40522

   PIN FE_OCPN62760_n_40389
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 163.15 0.51 163.25 ;
      END
   END FE_OCPN62760_n_40389

   PIN FE_OCPN62777_n_40539
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 159.95 0.51 160.05 ;
      END
   END FE_OCPN62777_n_40539

   PIN FE_OCPN63398_n_41185
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 159.15 0.51 159.25 ;
      END
   END FE_OCPN63398_n_41185

   PIN FE_OCPN63401_n_40695
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 121.55 0.51 121.65 ;
      END
   END FE_OCPN63401_n_40695

   PIN FE_OCPN63684_n_40655
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 146.95 0.51 147.05 ;
      END
   END FE_OCPN63684_n_40655

   PIN FE_OCPN63702_n_40513
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 21.95 0.51 22.05 ;
      END
   END FE_OCPN63702_n_40513

   PIN FE_OCPN63974_n_40634
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 34.65 185.49 34.75 186 ;
      END
   END FE_OCPN63974_n_40634

   PIN FE_OCPN76163_n_40638
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 113.05 185.49 113.15 186 ;
      END
   END FE_OCPN76163_n_40638

   PIN FE_OCPN76302_FE_OFN67600_n_40588
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 69.55 0.51 69.65 ;
      END
   END FE_OCPN76302_FE_OFN67600_n_40588

   PIN FE_OCPN76722_n_40452
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 15.75 0.51 15.85 ;
      END
   END FE_OCPN76722_n_40452

   PIN FE_OCPN76870_n_40344
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 63.55 0.51 63.65 ;
      END
   END FE_OCPN76870_n_40344

   PIN FE_OCPN77056_n_40657
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 167.55 0.51 167.65 ;
      END
   END FE_OCPN77056_n_40657

   PIN FE_OCPN95432_FE_OFN89660_n_40792
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 113.95 0.51 114.05 ;
      END
   END FE_OCPN95432_FE_OFN89660_n_40792

   PIN FE_OCPN95534_n_40744
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 121.15 0.51 121.25 ;
      END
   END FE_OCPN95534_n_40744

   PIN FE_OCPN95536_FE_OFN90000_n_40684
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 36.55 0.51 36.65 ;
      END
   END FE_OCPN95536_FE_OFN90000_n_40684

   PIN FE_OCPN95612_FE_OFN89862_n_40309
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 142.75 0.51 142.85 ;
      END
   END FE_OCPN95612_FE_OFN89862_n_40309

   PIN FE_OCPN95618_n_40607
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 141.35 0.51 141.45 ;
      END
   END FE_OCPN95618_n_40607

   PIN FE_OCPN95760_n_40465
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 181.55 0.51 181.65 ;
      END
   END FE_OCPN95760_n_40465

   PIN FE_OCPN99043_n_40638
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 159.75 0.51 159.85 ;
      END
   END FE_OCPN99043_n_40638

   PIN FE_OCP_DRV_N78196_n_40785
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 116.65 185.49 116.75 186 ;
      END
   END FE_OCP_DRV_N78196_n_40785

   PIN FE_OCP_DRV_N78718_FE_OFN69107_n_40425
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 51.55 0.51 51.65 ;
      END
   END FE_OCP_DRV_N78718_FE_OFN69107_n_40425

   PIN FE_OCP_DRV_N99398_FE_OFN98007_n_35906
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 95.45 185.49 95.55 186 ;
      END
   END FE_OCP_DRV_N99398_FE_OFN98007_n_35906

   PIN FE_OFN11400_n_40826
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 51.35 0.51 51.45 ;
      END
   END FE_OFN11400_n_40826

   PIN FE_OFN36963_n_35917
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 86.65 185.49 86.75 186 ;
      END
   END FE_OFN36963_n_35917

   PIN FE_OFN36981_n_45345
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 79.65 185.49 79.75 186 ;
      END
   END FE_OFN36981_n_45345

   PIN FE_OFN37043_n_35919
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 87.75 0.51 87.85 ;
      END
   END FE_OFN37043_n_35919

   PIN FE_OFN37045_n_35919
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 79.75 0.51 79.85 ;
      END
   END FE_OFN37045_n_35919

   PIN FE_OFN37046_n_35919
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 132.35 0.51 132.45 ;
      END
   END FE_OFN37046_n_35919

   PIN FE_OFN37067_n_35921
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 41.35 0.51 41.45 ;
      END
   END FE_OFN37067_n_35921

   PIN FE_OFN46443_n_35921
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 79.55 0.51 79.65 ;
      END
   END FE_OFN46443_n_35921

   PIN FE_OFN46639_n_35902
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 100.05 185.49 100.15 186 ;
      END
   END FE_OFN46639_n_35902

   PIN FE_OFN46654_n_35904
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 32.65 185.49 32.75 186 ;
      END
   END FE_OFN46654_n_35904

   PIN FE_OFN49989_n_40350
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 142.55 0.51 142.65 ;
      END
   END FE_OFN49989_n_40350

   PIN FE_OFN49990_n_40689
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 34.95 0.51 35.05 ;
      END
   END FE_OFN49990_n_40689

   PIN FE_OFN50159_n_51368
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 149.85 185.49 149.95 186 ;
      END
   END FE_OFN50159_n_51368

   PIN FE_OFN50261_n_51366
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 153.45 185.49 153.55 186 ;
      END
   END FE_OFN50261_n_51366

   PIN FE_OFN50310_n_40737
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 113.75 0.51 113.85 ;
      END
   END FE_OFN50310_n_40737

   PIN FE_OFN52335_n_45520
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 153.85 185.49 153.95 186 ;
      END
   END FE_OFN52335_n_45520

   PIN FE_OFN5281_n_40391
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 132.55 0.51 132.65 ;
      END
   END FE_OFN5281_n_40391

   PIN FE_OFN53002_n_40279
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 141.15 0.51 141.25 ;
      END
   END FE_OFN53002_n_40279

   PIN FE_OFN53022_n_40337
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 105.55 0.51 105.65 ;
      END
   END FE_OFN53022_n_40337

   PIN FE_OFN53283_n_40791
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 149.95 0.51 150.05 ;
      END
   END FE_OFN53283_n_40791

   PIN FE_OFN53291_n_41258
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 35.55 0.51 35.65 ;
      END
   END FE_OFN53291_n_41258

   PIN FE_OFN53587_n_40797
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 43.55 0.51 43.65 ;
      END
   END FE_OFN53587_n_40797

   PIN FE_OFN53642_n_40692
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 40.85 185.49 40.95 186 ;
      END
   END FE_OFN53642_n_40692

   PIN FE_OFN53722_n_40501
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 64.55 0.51 64.65 ;
      END
   END FE_OFN53722_n_40501

   PIN FE_OFN53780_n_52084
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 37.85 185.49 37.95 186 ;
      END
   END FE_OFN53780_n_52084

   PIN FE_OFN53782_n_52084
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 32.05 185.49 32.15 186 ;
      END
   END FE_OFN53782_n_52084

   PIN FE_OFN53783_n_52084
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 70.45 185.49 70.55 186 ;
      END
   END FE_OFN53783_n_52084

   PIN FE_OFN53822_n_40455
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 105.15 0.51 105.25 ;
      END
   END FE_OFN53822_n_40455

   PIN FE_OFN53850_n_52081
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 50.65 185.49 50.75 186 ;
      END
   END FE_OFN53850_n_52081

   PIN FE_OFN53963_n_40967
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 96.55 0.51 96.65 ;
      END
   END FE_OFN53963_n_40967

   PIN FE_OFN53973_n_52082
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 85.65 185.49 85.75 186 ;
      END
   END FE_OFN53973_n_52082

   PIN FE_OFN54887_n_45508
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 181.55 161.4 181.65 ;
      END
   END FE_OFN54887_n_45508

   PIN FE_OFN55725_n_52027
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 159.35 161.4 159.45 ;
      END
   END FE_OFN55725_n_52027

   PIN FE_OFN55732_n_52083
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 68.05 185.49 68.15 186 ;
      END
   END FE_OFN55732_n_52083

   PIN FE_OFN55733_n_52083
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 17.65 185.49 17.75 186 ;
      END
   END FE_OFN55733_n_52083

   PIN FE_OFN55736_n_52083
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 38.05 185.49 38.15 186 ;
      END
   END FE_OFN55736_n_52083

   PIN FE_OFN55761_n_52081
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 104.45 185.49 104.55 186 ;
      END
   END FE_OFN55761_n_52081

   PIN FE_OFN55822_n_52026
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 37.65 185.49 37.75 186 ;
      END
   END FE_OFN55822_n_52026

   PIN FE_OFN55823_n_52026
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 50.85 185.49 50.95 186 ;
      END
   END FE_OFN55823_n_52026

   PIN FE_OFN65159_n_57599
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 148.95 0.51 149.05 ;
      END
   END FE_OFN65159_n_57599

   PIN FE_OFN65264_n_40386
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 23.65 185.49 23.75 186 ;
      END
   END FE_OFN65264_n_40386

   PIN FE_OFN66190_n_40803
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 69.55 161.4 69.65 ;
      END
   END FE_OFN66190_n_40803

   PIN FE_OFN66462_n_41242
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 78.95 0.51 79.05 ;
      END
   END FE_OFN66462_n_41242

   PIN FE_OFN68662_n_41001
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 51.15 0.51 51.25 ;
      END
   END FE_OFN68662_n_41001

   PIN FE_OFN69662_n_40499
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 70.55 0.51 70.65 ;
      END
   END FE_OFN69662_n_40499

   PIN FE_OFN72075_n_35884
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 35.45 185.49 35.55 186 ;
      END
   END FE_OFN72075_n_35884

   PIN FE_OFN7415_n_57598
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 123.35 0.51 123.45 ;
      END
   END FE_OFN7415_n_57598

   PIN FE_OFN79894_n_53976
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 40.65 185.49 40.75 186 ;
      END
   END FE_OFN79894_n_53976

   PIN FE_OFN80051_n_54052
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 159.55 0.51 159.65 ;
      END
   END FE_OFN80051_n_54052

   PIN FE_OFN80076_n_57600
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 150.35 0.51 150.45 ;
      END
   END FE_OFN80076_n_57600

   PIN FE_OFN80128_n_40881
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 122.55 0.51 122.65 ;
      END
   END FE_OFN80128_n_40881

   PIN FE_OFN81050_n_40677
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 63.35 0.51 63.45 ;
      END
   END FE_OFN81050_n_40677

   PIN FE_OFN82374_n_40595
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 6.95 0.51 7.05 ;
      END
   END FE_OFN82374_n_40595

   PIN FE_OFN89560_n_40600
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 135.15 0.51 135.25 ;
      END
   END FE_OFN89560_n_40600

   PIN FE_OFN89563_n_40669
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 105.35 0.51 105.45 ;
      END
   END FE_OFN89563_n_40669

   PIN FE_OFN89691_n_40666
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 115.35 0.51 115.45 ;
      END
   END FE_OFN89691_n_40666

   PIN FE_OFN89714_n_40740
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 95.55 0.51 95.65 ;
      END
   END FE_OFN89714_n_40740

   PIN FE_OFN89774_n_40818
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 120.95 0.51 121.05 ;
      END
   END FE_OFN89774_n_40818

   PIN FE_OFN89904_n_41210
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 149.75 0.51 149.85 ;
      END
   END FE_OFN89904_n_41210

   PIN FE_OFN89935_n_40583
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 32.75 0.51 32.85 ;
      END
   END FE_OFN89935_n_40583

   PIN FE_OFN89944_n_40368
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 50.95 0.51 51.05 ;
      END
   END FE_OFN89944_n_40368

   PIN FE_OFN89967_n_40639
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 149.55 0.51 149.65 ;
      END
   END FE_OFN89967_n_40639

   PIN FE_OFN89998_n_40672
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 77.65 185.49 77.75 186 ;
      END
   END FE_OFN89998_n_40672

   PIN FE_OFN90003_n_41246
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 20.95 0.51 21.05 ;
      END
   END FE_OFN90003_n_41246

   PIN FE_OFN90026_n_40748
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 76.95 0.51 77.05 ;
      END
   END FE_OFN90026_n_40748

   PIN FE_OFN90039_n_40717
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 21.75 0.51 21.85 ;
      END
   END FE_OFN90039_n_40717

   PIN FE_OFN90040_n_40372
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 63.15 0.51 63.25 ;
      END
   END FE_OFN90040_n_40372

   PIN FE_OFN90041_n_40381
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 11.65 185.49 11.75 186 ;
      END
   END FE_OFN90041_n_40381

   PIN FE_OFN90067_n_40724
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 140.95 0.51 141.05 ;
      END
   END FE_OFN90067_n_40724

   PIN FE_OFN90075_n_40436
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 50.05 185.49 50.15 186 ;
      END
   END FE_OFN90075_n_40436

   PIN FE_OFN90079_n_40674
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 52.85 185.49 52.95 186 ;
      END
   END FE_OFN90079_n_40674

   PIN FE_OFN90099_FE_OCPN63313_n_40689
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 35.35 0.51 35.45 ;
      END
   END FE_OFN90099_FE_OCPN63313_n_40689

   PIN FE_OFN92681_n_40584
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 62.75 0.51 62.85 ;
      END
   END FE_OFN92681_n_40584

   PIN FE_OFN92683_n_40586
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 133.35 0.51 133.45 ;
      END
   END FE_OFN92683_n_40586

   PIN FE_OFN92826_n_40562
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 86.95 0.51 87.05 ;
      END
   END FE_OFN92826_n_40562

   PIN FE_OFN92897_n_40742
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 134.95 0.51 135.05 ;
      END
   END FE_OFN92897_n_40742

   PIN FE_OFN93006_n_40725
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 22.35 0.51 22.45 ;
      END
   END FE_OFN93006_n_40725

   PIN FE_OFN93027_n_40885
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 79.35 0.51 79.45 ;
      END
   END FE_OFN93027_n_40885

   PIN FE_OFN93041_n_40615
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 133.15 0.51 133.25 ;
      END
   END FE_OFN93041_n_40615

   PIN FE_OFN93057_n_40326
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 132.15 0.51 132.25 ;
      END
   END FE_OFN93057_n_40326

   PIN FE_OFN93058_n_40380
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 48.95 0.51 49.05 ;
      END
   END FE_OFN93058_n_40380

   PIN FE_OFN93060_n_40468
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 150.95 0.51 151.05 ;
      END
   END FE_OFN93060_n_40468

   PIN FE_OFN93171_n_40656
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 60.35 0.51 60.45 ;
      END
   END FE_OFN93171_n_40656

   PIN FE_OFN93173_n_41200
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 121.35 0.51 121.45 ;
      END
   END FE_OFN93173_n_41200

   PIN FE_OFN93186_n_40422
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 104.95 0.51 105.05 ;
      END
   END FE_OFN93186_n_40422

   PIN FE_OFN93289_n_40441
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 162.95 0.51 163.05 ;
      END
   END FE_OFN93289_n_40441

   PIN FE_OFN93291_n_40578
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 79.15 0.51 79.25 ;
      END
   END FE_OFN93291_n_40578

   PIN FE_OFN93292_n_40587
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 42.15 0.51 42.25 ;
      END
   END FE_OFN93292_n_40587

   PIN FE_OFN93294_n_40680
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 43.35 0.51 43.45 ;
      END
   END FE_OFN93294_n_40680

   PIN FE_OFN93352_n_40623
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 142.35 0.51 142.45 ;
      END
   END FE_OFN93352_n_40623

   PIN FE_OFN93353_n_40382
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 8.15 0.51 8.25 ;
      END
   END FE_OFN93353_n_40382

   PIN FE_OFN94636_n_40702
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 131.95 0.51 132.05 ;
      END
   END FE_OFN94636_n_40702

   PIN FE_OFN94776_n_40849
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 36.75 0.51 36.85 ;
      END
   END FE_OFN94776_n_40849

   PIN FE_OFN94918_n_40413
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 113.55 0.51 113.65 ;
      END
   END FE_OFN94918_n_40413

   PIN FE_OFN95014_n_41213
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 122.35 0.51 122.45 ;
      END
   END FE_OFN95014_n_41213

   PIN FE_OFN95068_n_40835
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 62.55 0.51 62.65 ;
      END
   END FE_OFN95068_n_40835

   PIN FE_OFN95079_n_40444
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 69.35 0.51 69.45 ;
      END
   END FE_OFN95079_n_40444

   PIN FE_OFN95120_n_40529
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 158.95 0.51 159.05 ;
      END
   END FE_OFN95120_n_40529

   PIN FE_OFN95165_n_40353
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 87.55 161.4 87.65 ;
      END
   END FE_OFN95165_n_40353

   PIN FE_OFN95201_n_40714
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 131.75 0.51 131.85 ;
      END
   END FE_OFN95201_n_40714

   PIN FE_OFN96060_FE_OCPN59260_n_40732
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 32.55 0.51 32.65 ;
      END
   END FE_OFN96060_FE_OCPN59260_n_40732

   PIN FE_OFN96766_FE_OCPN60886_n_40646
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 69.15 0.51 69.25 ;
      END
   END FE_OFN96766_FE_OCPN60886_n_40646

   PIN FE_OFN96958_n_40592
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 149.35 0.51 149.45 ;
      END
   END FE_OFN96958_n_40592

   PIN FE_OFN97291_n_40798
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 86.35 0.51 86.45 ;
      END
   END FE_OFN97291_n_40798

   PIN FE_OFN97312_n_40440
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 68.95 0.51 69.05 ;
      END
   END FE_OFN97312_n_40440

   PIN FE_OFN97388_n_40734
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 21.55 0.51 21.65 ;
      END
   END FE_OFN97388_n_40734

   PIN FE_OFN97595_FE_OCPN61185_n_40442
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 70.35 0.51 70.45 ;
      END
   END FE_OFN97595_FE_OCPN61185_n_40442

   PIN FE_RN_2180_0
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 110.25 185.49 110.35 186 ;
      END
   END FE_RN_2180_0

   PIN n_40316
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 86.75 0.51 86.85 ;
      END
   END n_40316

   PIN n_40337
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 121.15 0.51 121.25 ;
      END
   END n_40337

   PIN n_40354
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 134.95 0.51 135.05 ;
      END
   END n_40354

   PIN n_40363
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 6.05 185.49 6.15 186 ;
      END
   END n_40363

   PIN n_40393
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 104.75 0.51 104.85 ;
      END
   END n_40393

   PIN n_40397
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 21.35 0.51 21.45 ;
      END
   END n_40397

   PIN n_40404
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 131.55 0.51 131.65 ;
      END
   END n_40404

   PIN n_40409
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 131.35 0.51 131.45 ;
      END
   END n_40409

   PIN n_40414
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 132.35 0.51 132.45 ;
      END
   END n_40414

   PIN n_40418
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 150.75 0.51 150.85 ;
      END
   END n_40418

   PIN n_40423
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 150.55 0.51 150.65 ;
      END
   END n_40423

   PIN n_40449
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 36.35 0.51 36.45 ;
      END
   END n_40449

   PIN n_40460
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 68.75 0.51 68.85 ;
      END
   END n_40460

   PIN n_40505
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 113.35 0.51 113.45 ;
      END
   END n_40505

   PIN n_40516
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 16.85 185.49 16.95 186 ;
      END
   END n_40516

   PIN n_40526
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 135.35 0.51 135.45 ;
      END
   END n_40526

   PIN n_40556
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 95.45 185.49 95.55 186 ;
      END
   END n_40556

   PIN n_40579
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 36.15 0.51 36.25 ;
      END
   END n_40579

   PIN n_40593
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 122.15 0.51 122.25 ;
      END
   END n_40593

   PIN n_40598
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 120.95 0.51 121.05 ;
      END
   END n_40598

   PIN n_40616
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 149.15 0.51 149.25 ;
      END
   END n_40616

   PIN n_40637
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 142.35 0.51 142.45 ;
      END
   END n_40637

   PIN n_40666
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 115.15 0.51 115.25 ;
      END
   END n_40666

   PIN n_40685
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 115.75 0.51 115.85 ;
      END
   END n_40685

   PIN n_40690
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 164.95 0.51 165.05 ;
      END
   END n_40690

   PIN n_40701
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 70.25 185.49 70.35 186 ;
      END
   END n_40701

   PIN n_40706
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 114.35 0.51 114.45 ;
      END
   END n_40706

   PIN n_40710
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 131.15 0.51 131.25 ;
      END
   END n_40710

   PIN n_40720
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 142.15 0.51 142.25 ;
      END
   END n_40720

   PIN n_40729
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 18.85 185.49 18.95 186 ;
      END
   END n_40729

   PIN n_40741
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 86.05 185.49 86.15 186 ;
      END
   END n_40741

   PIN n_40743
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 104.55 0.51 104.65 ;
      END
   END n_40743

   PIN n_40745
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 107.15 0.51 107.25 ;
      END
   END n_40745

   PIN n_40765
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 113.15 0.51 113.25 ;
      END
   END n_40765

   PIN n_40768
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 132.15 0.51 132.25 ;
      END
   END n_40768

   PIN n_40770
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 119.35 0.51 119.45 ;
      END
   END n_40770

   PIN n_40777
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 5.85 185.49 5.95 186 ;
      END
   END n_40777

   PIN n_40783
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 71.25 185.49 71.35 186 ;
      END
   END n_40783

   PIN n_41024
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 150.35 0.51 150.45 ;
      END
   END n_41024

   PIN n_41051
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 140.75 0.51 140.85 ;
      END
   END n_41051

   PIN n_41057
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 150.15 161.4 150.25 ;
      END
   END n_41057

   PIN n_41085
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 7.95 0.51 8.05 ;
      END
   END n_41085

   PIN n_41094
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 78.95 0.51 79.05 ;
      END
   END n_41094

   PIN n_41111
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 95.35 0.51 95.45 ;
      END
   END n_41111

   PIN n_41129
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 123.45 185.49 123.55 186 ;
      END
   END n_41129

   PIN n_41136
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 123.15 0.51 123.25 ;
      END
   END n_41136

   PIN n_41188
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 140.55 0.51 140.65 ;
      END
   END n_41188

   PIN n_41231
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 78.15 0.51 78.25 ;
      END
   END n_41231

   PIN n_42980
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 160.89 123.35 161.4 123.45 ;
      END
   END n_42980

   PIN n_42981
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 131.25 185.49 131.35 186 ;
      END
   END n_42981

   PIN n_42983
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 131.05 185.49 131.15 186 ;
      END
   END n_42983

   PIN n_45340
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 68.45 185.49 68.55 186 ;
      END
   END n_45340

   PIN n_45516
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 140.25 185.49 140.35 186 ;
      END
   END n_45516

   PIN n_51367
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 152.25 185.49 152.35 186 ;
      END
   END n_51367

   PIN n_51369
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 151.65 185.49 151.75 186 ;
      END
   END n_51369

   PIN n_53993
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 43.15 0.51 43.25 ;
      END
   END n_53993

   PIN n_54048
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 130.95 0.51 131.05 ;
      END
   END n_54048

   PIN n_54049
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 5.65 185.49 5.75 186 ;
      END
   END n_54049

   PIN n_54050
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 59.05 185.49 59.15 186 ;
      END
   END n_54050

   PIN n_54051
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 87.95 0.51 88.05 ;
      END
   END n_54051

   PIN n_54054
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 106.95 0.51 107.05 ;
      END
   END n_54054

   PIN n_54088
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 5.45 185.49 5.55 186 ;
      END
   END n_54088

   PIN n_54101
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 140.35 0.51 140.45 ;
      END
   END n_54101

   PIN n_54219
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 14.45 185.49 14.55 186 ;
      END
   END n_54219

   PIN n_54222
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 177.55 0.51 177.65 ;
      END
   END n_54222

   PIN n_56439
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 131.95 0.51 132.05 ;
      END
   END n_56439

   PIN n_57586
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 68.55 0.51 68.65 ;
      END
   END n_57586

   PIN n_58039
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 59.65 185.49 59.75 186 ;
      END
   END n_58039

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 161.4 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 161.4 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 161.4 8.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 11.745 161.4 12.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 15.745 161.4 16.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 19.745 161.4 20.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 23.745 161.4 24.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 27.745 161.4 28.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 31.745 161.4 32.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 35.745 161.4 36.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 39.745 161.4 40.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 43.745 161.4 44.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 47.745 161.4 48.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 51.745 161.4 52.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 55.745 161.4 56.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 59.745 161.4 60.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 63.745 161.4 64.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 67.745 161.4 68.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 71.745 161.4 72.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 75.745 161.4 76.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 79.745 161.4 80.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 83.745 161.4 84.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 87.745 161.4 88.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 91.745 161.4 92.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 95.745 161.4 96.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 99.745 161.4 100.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 103.745 161.4 104.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 107.745 161.4 108.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 111.745 161.4 112.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 115.745 161.4 116.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 119.745 161.4 120.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 123.745 161.4 124.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 127.745 161.4 128.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 131.745 161.4 132.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 135.745 161.4 136.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 139.745 161.4 140.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 143.745 161.4 144.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 147.745 161.4 148.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 151.745 161.4 152.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 155.745 161.4 156.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 159.745 161.4 160.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 163.745 161.4 164.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 167.745 161.4 168.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 171.745 161.4 172.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 175.745 161.4 176.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 179.745 161.4 180.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 183.745 161.4 184.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 161.4 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 161.4 6.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 9.745 161.4 10.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 13.745 161.4 14.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 17.745 161.4 18.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 21.745 161.4 22.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 25.745 161.4 26.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 29.745 161.4 30.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 33.745 161.4 34.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 37.745 161.4 38.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 41.745 161.4 42.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 45.745 161.4 46.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 49.745 161.4 50.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 53.745 161.4 54.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 57.745 161.4 58.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 61.745 161.4 62.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 65.745 161.4 66.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 69.745 161.4 70.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 73.745 161.4 74.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 77.745 161.4 78.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 81.745 161.4 82.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 85.745 161.4 86.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 89.745 161.4 90.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 93.745 161.4 94.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 97.745 161.4 98.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 101.745 161.4 102.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 105.745 161.4 106.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 109.745 161.4 110.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 113.745 161.4 114.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 117.745 161.4 118.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 121.745 161.4 122.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 125.745 161.4 126.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 129.745 161.4 130.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 133.745 161.4 134.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 137.745 161.4 138.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 141.745 161.4 142.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 145.745 161.4 146.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 149.745 161.4 150.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 153.745 161.4 154.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 157.745 161.4 158.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 161.745 161.4 162.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 165.745 161.4 166.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 169.745 161.4 170.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 173.745 161.4 174.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 177.745 161.4 178.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 181.745 161.4 182.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 185.745 161.4 186.255 ;
      END
   END vdd

   OBS
      LAYER metal1 ;
         RECT 0 0 161.4 186 ;
   END
   OBS
      LAYER metal2 ;
         RECT 0 0 161.4 186 ;
   END
   OBS
      LAYER metal3 ;
         RECT 0 0 161.4 186 ;
   END
   OBS
      LAYER metal4 ;
         RECT 0 0 161.4 186 ;
   END
   OBS
      LAYER metal5 ;
         RECT 0 0 161.4 186 ;
   END
END h6

MACRO h3
   CLASS BLOCK ;
   SIZE 180.2 BY 202 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   PIN FE_OCPN56827_n_23035
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 114.45 201.49 114.55 202 ;
      END
   END FE_OCPN56827_n_23035

   PIN FE_OCPN57195_FE_OFN46384_n_23035
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 191.15 0.51 191.25 ;
      END
   END FE_OCPN57195_FE_OFN46384_n_23035

   PIN FE_OCPN57332_FE_OFN48190_n_22999
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 138.15 180.2 138.25 ;
      END
   END FE_OCPN57332_FE_OFN48190_n_22999

   PIN FE_OCPN58002_FE_OFN46384_n_23035
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 191.35 0.51 191.45 ;
      END
   END FE_OCPN58002_FE_OFN46384_n_23035

   PIN FE_OCPN58799_FE_OFN41801_n_23039
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 75.55 0.51 75.65 ;
      END
   END FE_OCPN58799_FE_OFN41801_n_23039

   PIN FE_OCPN59420_FE_OFN47458_n_22985
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 148.95 0.51 149.05 ;
      END
   END FE_OCPN59420_FE_OFN47458_n_22985

   PIN FE_OCPN59424_FE_OFN47458_n_22985
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 179.69 152.95 180.2 153.05 ;
      END
   END FE_OCPN59424_FE_OFN47458_n_22985

   PIN FE_OCPN59425_FE_OFN47458_n_22985
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 152.95 0.51 153.05 ;
      END
   END FE_OCPN59425_FE_OFN47458_n_22985

   PIN FE_OCPN59960_FE_OFN48190_n_22999
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 91.15 180.2 91.25 ;
      END
   END FE_OCPN59960_FE_OFN48190_n_22999

   PIN FE_OCPN60172_FE_OFN47326_n_67216
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 93.35 0.51 93.45 ;
      END
   END FE_OCPN60172_FE_OFN47326_n_67216

   PIN FE_OCPN60404_FE_OFN48179_n_22997
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 65.75 180.2 65.85 ;
      END
   END FE_OCPN60404_FE_OFN48179_n_22997

   PIN FE_OCPN61220_n_24492
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 179.69 84.55 180.2 84.65 ;
      END
   END FE_OCPN61220_n_24492

   PIN FE_OCPN61492_FE_OFN48190_n_22999
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 126.05 201.49 126.15 202 ;
      END
   END FE_OCPN61492_FE_OFN48190_n_22999

   PIN FE_OCPN63674_n_23815
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 154.95 180.2 155.05 ;
      END
   END FE_OCPN63674_n_23815

   PIN FE_OCPN76133_FE_OFN41801_n_23039
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 75.75 0.51 75.85 ;
      END
   END FE_OCPN76133_FE_OFN41801_n_23039

   PIN FE_OCPN76840_FE_OFN47632_n_22865
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 93.55 0.51 93.65 ;
      END
   END FE_OCPN76840_FE_OFN47632_n_22865

   PIN FE_OCPN76842_FE_OFN47632_n_22865
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 39.65 0 39.75 0.51 ;
      END
   END FE_OCPN76842_FE_OFN47632_n_22865

   PIN FE_OCPN77030_FE_OFN75657_n_22948
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 183.55 0.51 183.65 ;
      END
   END FE_OCPN77030_FE_OFN75657_n_22948

   PIN FE_OCP_RBN77248_FE_OCPN57193_FE_OFN46384_n_23035
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 107.05 0 107.15 0.51 ;
      END
   END FE_OCP_RBN77248_FE_OCPN57193_FE_OFN46384_n_23035

   PIN FE_OCP_RBN77364_FE_OCPN57515_FE_OFN47099_n_23039
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 165.85 0 165.95 0.51 ;
      END
   END FE_OCP_RBN77364_FE_OCPN57515_FE_OFN47099_n_23039

   PIN FE_OFN13351_n_25338
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 51.05 0 51.15 0.51 ;
      END
   END FE_OFN13351_n_25338

   PIN FE_OFN13710_n_23652
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 57.55 0.51 57.65 ;
      END
   END FE_OFN13710_n_23652

   PIN FE_OFN13716_n_24566
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 30.15 180.2 30.25 ;
      END
   END FE_OFN13716_n_24566

   PIN FE_OFN29431_n_522
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 69.45 0 69.55 0.51 ;
      END
   END FE_OFN29431_n_522

   PIN FE_OFN33789_n_3396
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 130.25 0 130.35 0.51 ;
      END
   END FE_OFN33789_n_3396

   PIN FE_OFN34206_n_82
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 69.25 0 69.35 0.51 ;
      END
   END FE_OFN34206_n_82

   PIN FE_OFN34223_n_81
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 102.35 180.2 102.45 ;
      END
   END FE_OFN34223_n_81

   PIN FE_OFN34312_n_77
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 50.95 0.51 51.05 ;
      END
   END FE_OFN34312_n_77

   PIN FE_OFN34580_n_223
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 22.55 180.2 22.65 ;
      END
   END FE_OFN34580_n_223

   PIN FE_OFN34592_n_223
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 39.95 180.2 40.05 ;
      END
   END FE_OFN34592_n_223

   PIN FE_OFN34595_n_223
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 112.95 180.2 113.05 ;
      END
   END FE_OFN34595_n_223

   PIN FE_OFN34606_n_223
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 66.55 180.2 66.65 ;
      END
   END FE_OFN34606_n_223

   PIN FE_OFN41924_n_227
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 57.75 0.51 57.85 ;
      END
   END FE_OFN41924_n_227

   PIN FE_OFN41991_n_228
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 120.35 180.2 120.45 ;
      END
   END FE_OFN41991_n_228

   PIN FE_OFN42299_n_47
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 39.55 180.2 39.65 ;
      END
   END FE_OFN42299_n_47

   PIN FE_OFN42492_n_33
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 153.55 180.2 153.65 ;
      END
   END FE_OFN42492_n_33

   PIN FE_OFN42501_n_33
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 172.85 0 172.95 0.51 ;
      END
   END FE_OFN42501_n_33

   PIN FE_OFN42529_n_32
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 129.35 180.2 129.45 ;
      END
   END FE_OFN42529_n_32

   PIN FE_OFN42808_n_10
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 57.75 180.2 57.85 ;
      END
   END FE_OFN42808_n_10

   PIN FE_OFN42954_n_3289
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 12.95 180.2 13.05 ;
      END
   END FE_OFN42954_n_3289

   PIN FE_OFN42968_n_1990
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 165.15 180.2 165.25 ;
      END
   END FE_OFN42968_n_1990

   PIN FE_OFN43882_n_67219
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 131.15 0.51 131.25 ;
      END
   END FE_OFN43882_n_67219

   PIN FE_OFN43982_mux_g_ln477_q_1311_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 27.05 0 27.15 0.51 ;
      END
   END FE_OFN43982_mux_g_ln477_q_1311_

   PIN FE_OFN47020_n_67217
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 78.85 0 78.95 0.51 ;
      END
   END FE_OFN47020_n_67217

   PIN FE_OFN47329_n_67216
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 102.55 0.51 102.65 ;
      END
   END FE_OFN47329_n_67216

   PIN FE_OFN47630_n_22865
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 146.95 0.51 147.05 ;
      END
   END FE_OFN47630_n_22865

   PIN FE_OFN47632_n_22865
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 179.69 66.55 180.2 66.65 ;
      END
   END FE_OFN47632_n_22865

   PIN FE_OFN48892_n_24195
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 39.35 180.2 39.45 ;
      END
   END FE_OFN48892_n_24195

   PIN FE_OFN51049_n_23652
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 101.95 180.2 102.05 ;
      END
   END FE_OFN51049_n_23652

   PIN FE_OFN51274_n_25014
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 111.35 180.2 111.45 ;
      END
   END FE_OFN51274_n_25014

   PIN FE_OFN51275_n_25016
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 111.55 180.2 111.65 ;
      END
   END FE_OFN51275_n_25016

   PIN FE_OFN51548_n_23656
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 138.95 180.2 139.05 ;
      END
   END FE_OFN51548_n_23656

   PIN FE_OFN51552_n_23702
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 138.35 180.2 138.45 ;
      END
   END FE_OFN51552_n_23702

   PIN FE_OFN51947_n_23990
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 190.95 180.2 191.05 ;
      END
   END FE_OFN51947_n_23990

   PIN FE_OFN52123_n_23549
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 152.95 180.2 153.05 ;
      END
   END FE_OFN52123_n_23549

   PIN FE_OFN53748_n_3398
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 96.65 0 96.75 0.51 ;
      END
   END FE_OFN53748_n_3398

   PIN FE_OFN53753_n_71
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 132.25 201.49 132.35 202 ;
      END
   END FE_OFN53753_n_71

   PIN FE_OFN53899_n_89
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 155.65 0 155.75 0.51 ;
      END
   END FE_OFN53899_n_89

   PIN FE_OFN54457_n_23864
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 51.25 0 51.35 0.51 ;
      END
   END FE_OFN54457_n_23864

   PIN FE_OFN54621_n_23573
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 179.69 111.55 180.2 111.65 ;
      END
   END FE_OFN54621_n_23573

   PIN FE_OFN54630_n_23981
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 179.69 138.35 180.2 138.45 ;
      END
   END FE_OFN54630_n_23981

   PIN FE_OFN54631_n_23986
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 179.69 138.55 180.2 138.65 ;
      END
   END FE_OFN54631_n_23986

   PIN FE_OFN54638_n_24584
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 120.75 180.2 120.85 ;
      END
   END FE_OFN54638_n_24584

   PIN FE_OFN54639_n_24584
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 84.75 0.51 84.85 ;
      END
   END FE_OFN54639_n_24584

   PIN FE_OFN54891_n_23983
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 102.55 180.2 102.65 ;
      END
   END FE_OFN54891_n_23983

   PIN FE_OFN56004_n_5228837_bar
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 192.95 0.51 193.05 ;
      END
   END FE_OFN56004_n_5228837_bar

   PIN FE_OFN71792_eq_15722_64_n_18
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 150.45 0 150.55 0.51 ;
      END
   END FE_OFN71792_eq_15722_64_n_18

   PIN FE_OFN73040_n_23035
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 40.15 180.2 40.25 ;
      END
   END FE_OFN73040_n_23035

   PIN FE_OFN73486_n_11
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 110.05 0 110.15 0.51 ;
      END
   END FE_OFN73486_n_11

   PIN FE_OFN73506_n_10
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 191.95 180.2 192.05 ;
      END
   END FE_OFN73506_n_10

   PIN FE_OFN73546_n_30
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 114.45 0 114.55 0.51 ;
      END
   END FE_OFN73546_n_30

   PIN FE_OFN73612_n_43
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 153.15 180.2 153.25 ;
      END
   END FE_OFN73612_n_43

   PIN FE_OFN73633_n_31
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 34.75 180.2 34.85 ;
      END
   END FE_OFN73633_n_31

   PIN FE_OFN73665_n_33
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 172.65 201.49 172.75 202 ;
      END
   END FE_OFN73665_n_33

   PIN FE_OFN73711_n_222
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 29.45 0 29.55 0.51 ;
      END
   END FE_OFN73711_n_222

   PIN FE_OFN74312_n_61
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 78.45 0 78.55 0.51 ;
      END
   END FE_OFN74312_n_61

   PIN FE_OFN75677_n_22920
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 155.95 0.51 156.05 ;
      END
   END FE_OFN75677_n_22920

   PIN FE_OFN81211_n_24583
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 42.25 0 42.35 0.51 ;
      END
   END FE_OFN81211_n_24583

   PIN FE_OFN85501_n_223
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 71.25 0 71.35 0.51 ;
      END
   END FE_OFN85501_n_223

   PIN FE_OFN86522_n_518
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 21.55 0.51 21.65 ;
      END
   END FE_OFN86522_n_518

   PIN FE_OFN87976_FE_OCPN56158_FE_OFN47027_n_67213
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 150.95 180.2 151.05 ;
      END
   END FE_OFN87976_FE_OCPN56158_FE_OFN47027_n_67213

   PIN FE_OFN88160_n_22979
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 151.35 0.51 151.45 ;
      END
   END FE_OFN88160_n_22979

   PIN FE_OFN88164_n_22979
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 153.15 0.51 153.25 ;
      END
   END FE_OFN88164_n_22979

   PIN FE_OFN89154_n_865
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 23.45 201.49 23.55 202 ;
      END
   END FE_OFN89154_n_865

   PIN FE_OFN90772_FE_OCPN60312_FE_OFN47628_n_22865
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 153.35 0.51 153.45 ;
      END
   END FE_OFN90772_FE_OCPN60312_FE_OFN47628_n_22865

   PIN FE_OFN90794_n_22919
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 158.95 0.51 159.05 ;
      END
   END FE_OFN90794_n_22919

   PIN FE_OFN90904_n_67217
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 39.75 0.51 39.85 ;
      END
   END FE_OFN90904_n_67217

   PIN FE_OFN90954_FE_RN_2244_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 153.35 180.2 153.45 ;
      END
   END FE_OFN90954_FE_RN_2244_0

   PIN FE_OFN91045_n_25028
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 151.15 180.2 151.25 ;
      END
   END FE_OFN91045_n_25028

   PIN FE_OFN93717_n_67217
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 39.05 0 39.15 0.51 ;
      END
   END FE_OFN93717_n_67217

   PIN FE_OFN93911_n_23836
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 137.95 180.2 138.05 ;
      END
   END FE_OFN93911_n_23836

   PIN FE_OFN94059_n_23989
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 174.55 180.2 174.65 ;
      END
   END FE_OFN94059_n_23989

   PIN FE_OFN94140_n_879
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 166.25 201.49 166.35 202 ;
      END
   END FE_OFN94140_n_879

   PIN FE_OFN94180_FE_OCPN77031_FE_OFN75657_n_22948
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 173.55 0.51 173.65 ;
      END
   END FE_OFN94180_FE_OCPN77031_FE_OFN75657_n_22948

   PIN FE_OFN98114_n_50
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 132.65 0 132.75 0.51 ;
      END
   END FE_OFN98114_n_50

   PIN FE_OFN98267_n_71
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 33.45 201.49 33.55 202 ;
      END
   END FE_OFN98267_n_71

   PIN FE_RN_4736_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 159.45 0 159.55 0.51 ;
      END
   END FE_RN_4736_0

   PIN FE_RN_4810_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 84.15 180.2 84.25 ;
      END
   END FE_RN_4810_0

   PIN FE_RN_5927_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 48.95 180.2 49.05 ;
      END
   END FE_RN_5927_0

   PIN mux_g_ln477_q_1304_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 165.05 0 165.15 0.51 ;
      END
   END mux_g_ln477_q_1304_

   PIN mux_g_ln477_q_1307_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 111.75 180.2 111.85 ;
      END
   END mux_g_ln477_q_1307_

   PIN mux_g_ln477_q_1311_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 179.69 176.15 180.2 176.25 ;
      END
   END mux_g_ln477_q_1311_

   PIN mux_g_ln477_q_1347_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 49.95 0.51 50.05 ;
      END
   END mux_g_ln477_q_1347_

   PIN mux_g_ln477_q_1350_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 15.45 0 15.55 0.51 ;
      END
   END mux_g_ln477_q_1350_

   PIN mux_g_ln477_q_1355_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 6.05 0 6.15 0.51 ;
      END
   END mux_g_ln477_q_1355_

   PIN mux_g_ln477_q_1364_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 6.65 0 6.75 0.51 ;
      END
   END mux_g_ln477_q_1364_

   PIN mux_g_ln477_q_1366_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 105.05 0 105.15 0.51 ;
      END
   END mux_g_ln477_q_1366_

   PIN mux_g_ln477_q_1480_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 75.15 0.51 75.25 ;
      END
   END mux_g_ln477_q_1480_

   PIN mux_g_ln477_q_1484_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 138.75 180.2 138.85 ;
      END
   END mux_g_ln477_q_1484_

   PIN mux_g_ln477_q_1488_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 24.65 0 24.75 0.51 ;
      END
   END mux_g_ln477_q_1488_

   PIN mux_g_ln477_q_1496_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 147.15 0.51 147.25 ;
      END
   END mux_g_ln477_q_1496_

   PIN mux_g_ln477_q_1497_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 108.95 0.51 109.05 ;
      END
   END mux_g_ln477_q_1497_

   PIN mux_g_ln477_q_1500_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 91.35 180.2 91.45 ;
      END
   END mux_g_ln477_q_1500_

   PIN mux_g_ln477_q_1503_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 165.55 0.51 165.65 ;
      END
   END mux_g_ln477_q_1503_

   PIN mux_g_ln477_q_1534_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 78.85 201.49 78.95 202 ;
      END
   END mux_g_ln477_q_1534_

   PIN mux_g_ln477_q_578_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 171.45 0 171.55 0.51 ;
      END
   END mux_g_ln477_q_578_

   PIN mux_g_ln477_q_592_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 84.25 0 84.35 0.51 ;
      END
   END mux_g_ln477_q_592_

   PIN mux_g_ln477_q_593_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 51.45 0 51.55 0.51 ;
      END
   END mux_g_ln477_q_593_

   PIN mux_g_ln477_q_597_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 105.45 0 105.55 0.51 ;
      END
   END mux_g_ln477_q_597_

   PIN mux_g_ln477_q_601_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 105.65 0 105.75 0.51 ;
      END
   END mux_g_ln477_q_601_

   PIN mux_g_ln477_q_602_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 69.05 0 69.15 0.51 ;
      END
   END mux_g_ln477_q_602_

   PIN mux_g_ln477_q_604_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 99.65 0 99.75 0.51 ;
      END
   END mux_g_ln477_q_604_

   PIN n_2109
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 168.45 0 168.55 0.51 ;
      END
   END n_2109

   PIN n_2226
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 75.75 180.2 75.85 ;
      END
   END n_2226

   PIN n_23565
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 156.35 0.51 156.45 ;
      END
   END n_23565

   PIN n_23712
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 10.95 180.2 11.05 ;
      END
   END n_23712

   PIN n_23850
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 84.95 180.2 85.05 ;
      END
   END n_23850

   PIN n_23872
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 51.35 180.2 51.45 ;
      END
   END n_23872

   PIN n_23898
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 147.35 180.2 147.45 ;
      END
   END n_23898

   PIN n_23911
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 66.15 180.2 66.25 ;
      END
   END n_23911

   PIN n_24578
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 130.95 180.2 131.05 ;
      END
   END n_24578

   PIN n_24650
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 70.55 180.2 70.65 ;
      END
   END n_24650

   PIN n_24655
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 39.15 180.2 39.25 ;
      END
   END n_24655

   PIN n_24658
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 87.25 0 87.35 0.51 ;
      END
   END n_24658

   PIN n_24848
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 179.69 22.15 180.2 22.25 ;
      END
   END n_24848

   PIN n_25026
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 151.35 180.2 151.45 ;
      END
   END n_25026

   PIN n_25030
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 33.45 0 33.55 0.51 ;
      END
   END n_25030

   PIN n_25035
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 132.45 201.49 132.55 202 ;
      END
   END n_25035

   PIN n_25044
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 156.55 0.51 156.65 ;
      END
   END n_25044

   PIN n_25299
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 92.95 180.2 93.05 ;
      END
   END n_25299

   PIN n_25309
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 102.95 180.2 103.05 ;
      END
   END n_25309

   PIN n_2712
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 22.15 180.2 22.25 ;
      END
   END n_2712

   PIN n_2800
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 78.05 0 78.15 0.51 ;
      END
   END n_2800

   PIN n_2812
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 9.15 180.2 9.25 ;
      END
   END n_2812

   PIN n_3110
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 65.95 180.2 66.05 ;
      END
   END n_3110

   PIN n_3283
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 8.95 180.2 9.05 ;
      END
   END n_3283

   PIN n_3290
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 168.45 0 168.55 0.51 ;
      END
   END n_3290

   PIN n_4733
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 102.75 0.51 102.85 ;
      END
   END n_4733

   PIN n_5562
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 40.85 0 40.95 0.51 ;
      END
   END n_5562

   PIN n_5563
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 13.85 0 13.95 0.51 ;
      END
   END n_5563

   PIN n_5890
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 31.15 0.51 31.25 ;
      END
   END n_5890

   PIN n_6316
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 70.55 0.51 70.65 ;
      END
   END n_6316

   PIN n_6739
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 150.65 0 150.75 0.51 ;
      END
   END n_6739

   PIN FE_OCPN56158_FE_OFN47027_n_67213
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 140.95 180.2 141.05 ;
      END
   END FE_OCPN56158_FE_OFN47027_n_67213

   PIN FE_OCPN56824_n_23035
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 132.95 180.2 133.05 ;
      END
   END FE_OCPN56824_n_23035

   PIN FE_OCPN57568_FE_OFN47196_n_67214
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 77.85 0 77.95 0.51 ;
      END
   END FE_OCPN57568_FE_OFN47196_n_67214

   PIN FE_OCPN58871_FE_OFN43374_n_22937
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 93.35 180.2 93.45 ;
      END
   END FE_OCPN58871_FE_OFN43374_n_22937

   PIN FE_OCPN59418_FE_OFN47458_n_22985
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 22.35 180.2 22.45 ;
      END
   END FE_OCPN59418_FE_OFN47458_n_22985

   PIN FE_OCPN59878_FE_OFN47327_n_67216
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 179.69 57.55 180.2 57.65 ;
      END
   END FE_OCPN59878_FE_OFN47327_n_67216

   PIN FE_OCPN59929_FE_OFN47456_n_22985
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 84.75 180.2 84.85 ;
      END
   END FE_OCPN59929_FE_OFN47456_n_22985

   PIN FE_OCPN59934_n_24570
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 47.95 180.2 48.05 ;
      END
   END FE_OCPN59934_n_24570

   PIN FE_OCPN60169_FE_OFN47326_n_67216
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 21.55 180.2 21.65 ;
      END
   END FE_OCPN60169_FE_OFN47326_n_67216

   PIN FE_OCPN60170_FE_OFN47326_n_67216
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 31.35 180.2 31.45 ;
      END
   END FE_OCPN60170_FE_OFN47326_n_67216

   PIN FE_OCPN60246_FE_OFN47005_n_67217
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 58.15 180.2 58.25 ;
      END
   END FE_OCPN60246_FE_OFN47005_n_67217

   PIN FE_OCPN60333_FE_OFN41824_n_23039
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 122.95 180.2 123.05 ;
      END
   END FE_OCPN60333_FE_OFN41824_n_23039

   PIN FE_OCPN60351_FE_OFN43508_n_22865
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 132.25 0 132.35 0.51 ;
      END
   END FE_OCPN60351_FE_OFN43508_n_22865

   PIN FE_OCPN60402_FE_OFN48179_n_22997
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 60.95 180.2 61.05 ;
      END
   END FE_OCPN60402_FE_OFN48179_n_22997

   PIN FE_OCPN61219_n_24492
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 34.85 201.49 34.95 202 ;
      END
   END FE_OCPN61219_n_24492

   PIN FE_OCPN63510_FE_OFN41801_n_23039
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 39.75 180.2 39.85 ;
      END
   END FE_OCPN63510_FE_OFN41801_n_23039

   PIN FE_OCPN77813_n_23035
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 57.95 180.2 58.05 ;
      END
   END FE_OCPN77813_n_23035

   PIN FE_OCPN77821_FE_OFN47978_n_23035
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 105.25 0 105.35 0.51 ;
      END
   END FE_OCPN77821_FE_OFN47978_n_23035

   PIN FE_OCPN77894_n_23972
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 169.15 180.2 169.25 ;
      END
   END FE_OCPN77894_n_23972

   PIN FE_OCPN78264_FE_OFN47649_n_22866
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 130.85 0 130.95 0.51 ;
      END
   END FE_OCPN78264_FE_OFN47649_n_22866

   PIN FE_OCPN95395_FE_OFN46375_n_23035
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 66.35 180.2 66.45 ;
      END
   END FE_OCPN95395_FE_OFN46375_n_23035

   PIN FE_OCPN95638_FE_OFN48190_n_22999
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 51.15 180.2 51.25 ;
      END
   END FE_OCPN95638_FE_OFN48190_n_22999

   PIN FE_OCPUNCON99093_FE_OCP_RBN77363_FE_OCPN57515_FE_OFN47099_n_23039
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 24.25 201.49 24.35 202 ;
      END
   END FE_OCPUNCON99093_FE_OCP_RBN77363_FE_OCPN57515_FE_OFN47099_n_23039

   PIN FE_OCP_RBN77173_FE_OFN46375_n_23035
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 92.05 0 92.15 0.51 ;
      END
   END FE_OCP_RBN77173_FE_OFN46375_n_23035

   PIN FE_OFN13154_n_25272
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 70.35 180.2 70.45 ;
      END
   END FE_OFN13154_n_25272

   PIN FE_OFN13349_n_25338
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 29.95 180.2 30.05 ;
      END
   END FE_OFN13349_n_25338

   PIN FE_OFN15344_n_24443
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 50.95 180.2 51.05 ;
      END
   END FE_OFN15344_n_24443

   PIN FE_OFN29701_n_518
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 68.25 0 68.35 0.51 ;
      END
   END FE_OFN29701_n_518

   PIN FE_OFN34029_n_89
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 134.05 201.49 134.15 202 ;
      END
   END FE_OFN34029_n_89

   PIN FE_OFN34082_n_87
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 60.45 0 60.55 0.51 ;
      END
   END FE_OFN34082_n_87

   PIN FE_OFN34202_n_82
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 113.35 180.2 113.45 ;
      END
   END FE_OFN34202_n_82

   PIN FE_OFN34291_n_78
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 169.35 180.2 169.45 ;
      END
   END FE_OFN34291_n_78

   PIN FE_OFN34467_n_59
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 145.05 0 145.15 0.51 ;
      END
   END FE_OFN34467_n_59

   PIN FE_OFN34549_n_223
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 91.55 180.2 91.65 ;
      END
   END FE_OFN34549_n_223

   PIN FE_OFN34560_n_223
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 78.25 0 78.35 0.51 ;
      END
   END FE_OFN34560_n_223

   PIN FE_OFN35094_n_5228270_bar
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 127.05 201.49 127.15 202 ;
      END
   END FE_OFN35094_n_5228270_bar

   PIN FE_OFN35482_eq_15722_64_n_18
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 172.45 201.49 172.55 202 ;
      END
   END FE_OFN35482_eq_15722_64_n_18

   PIN FE_OFN42005_n_231
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 57.05 201.49 57.15 202 ;
      END
   END FE_OFN42005_n_231

   PIN FE_OFN42081_n_222
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 101.65 0 101.75 0.51 ;
      END
   END FE_OFN42081_n_222

   PIN FE_OFN42082_n_222
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 42.05 0 42.15 0.51 ;
      END
   END FE_OFN42082_n_222

   PIN FE_OFN42113_n_222
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 151.65 201.49 151.75 202 ;
      END
   END FE_OFN42113_n_222

   PIN FE_OFN42143_n_57
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 69.45 201.49 69.55 202 ;
      END
   END FE_OFN42143_n_57

   PIN FE_OFN42297_n_47
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 111.15 180.2 111.25 ;
      END
   END FE_OFN42297_n_47

   PIN FE_OFN42346_n_45
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 138.55 180.2 138.65 ;
      END
   END FE_OFN42346_n_45

   PIN FE_OFN42388_n_43
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 60.65 201.49 60.75 202 ;
      END
   END FE_OFN42388_n_43

   PIN FE_OFN42435_n_41
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 143.45 201.49 143.55 202 ;
      END
   END FE_OFN42435_n_41

   PIN FE_OFN42544_n_31
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 138.85 201.49 138.95 202 ;
      END
   END FE_OFN42544_n_31

   PIN FE_OFN42570_n_30
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 115.85 201.49 115.95 202 ;
      END
   END FE_OFN42570_n_30

   PIN FE_OFN42595_n_29
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 60.25 201.49 60.35 202 ;
      END
   END FE_OFN42595_n_29

   PIN FE_OFN42596_n_29
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 60.45 201.49 60.55 202 ;
      END
   END FE_OFN42596_n_29

   PIN FE_OFN42629_n_20
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 179.69 150.95 180.2 151.05 ;
      END
   END FE_OFN42629_n_20

   PIN FE_OFN42789_n_11
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 90.95 180.2 91.05 ;
      END
   END FE_OFN42789_n_11

   PIN FE_OFN42953_n_3289
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 39.55 0.51 39.65 ;
      END
   END FE_OFN42953_n_3289

   PIN FE_OFN43845_n_67218
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 45.2 0 45.4 0.255 ;
      END
   END FE_OFN43845_n_67218

   PIN FE_OFN43847_n_67218
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 15 0 15.2 0.255 ;
      END
   END FE_OFN43847_n_67218

   PIN FE_OFN46995_n_67217
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 75.55 180.2 75.65 ;
      END
   END FE_OFN46995_n_67217

   PIN FE_OFN46996_n_67217
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 70.75 180.2 70.85 ;
      END
   END FE_OFN46996_n_67217

   PIN FE_OFN47017_n_67217
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 150.45 0 150.55 0.51 ;
      END
   END FE_OFN47017_n_67217

   PIN FE_OFN47019_n_67217
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 118.85 0 118.95 0.51 ;
      END
   END FE_OFN47019_n_67217

   PIN FE_OFN47328_n_67216
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 68.95 180.2 69.05 ;
      END
   END FE_OFN47328_n_67216

   PIN FE_OFN47628_n_22865
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 151.55 180.2 151.65 ;
      END
   END FE_OFN47628_n_22865

   PIN FE_OFN47808_n_22977
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 55.85 0 55.95 0.51 ;
      END
   END FE_OFN47808_n_22977

   PIN FE_OFN47977_n_23035
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 105.25 0 105.35 0.51 ;
      END
   END FE_OFN47977_n_23035

   PIN FE_OFN48729_n_865
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 183.75 0.51 183.85 ;
      END
   END FE_OFN48729_n_865

   PIN FE_OFN48776_n_879
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 87.45 0 87.55 0.51 ;
      END
   END FE_OFN48776_n_879

   PIN FE_OFN50050_n_71
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 52.2 0 52.4 0.255 ;
      END
   END FE_OFN50050_n_71

   PIN FE_OFN51564_n_23989
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 151.15 0.51 151.25 ;
      END
   END FE_OFN51564_n_23989

   PIN FE_OFN51946_n_23990
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 190.95 0.51 191.05 ;
      END
   END FE_OFN51946_n_23990

   PIN FE_OFN53694_n_91
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 70.35 0.51 70.45 ;
      END
   END FE_OFN53694_n_91

   PIN FE_OFN53750_n_71
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 88.85 201.49 88.95 202 ;
      END
   END FE_OFN53750_n_71

   PIN FE_OFN53910_n_77
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 31.15 180.2 31.25 ;
      END
   END FE_OFN53910_n_77

   PIN FE_OFN53911_n_77
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 170.45 0 170.55 0.51 ;
      END
   END FE_OFN53911_n_77

   PIN FE_OFN72259_n_3398
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 153.05 201.49 153.15 202 ;
      END
   END FE_OFN72259_n_3398

   PIN FE_OFN73407_n_14
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 113.15 180.2 113.25 ;
      END
   END FE_OFN73407_n_14

   PIN FE_OFN73437_n_40
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 84.35 0.51 84.45 ;
      END
   END FE_OFN73437_n_40

   PIN FE_OFN73503_n_10
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 171.65 201.49 171.75 202 ;
      END
   END FE_OFN73503_n_10

   PIN FE_OFN73527_n_42
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 102.75 180.2 102.85 ;
      END
   END FE_OFN73527_n_42

   PIN FE_OFN73542_n_30
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 75.15 180.2 75.25 ;
      END
   END FE_OFN73542_n_30

   PIN FE_OFN73592_n_44
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 114.25 201.49 114.35 202 ;
      END
   END FE_OFN73592_n_44

   PIN FE_OFN73597_n_44
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 131.15 180.2 131.25 ;
      END
   END FE_OFN73597_n_44

   PIN FE_OFN73753_n_227
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 21.95 180.2 22.05 ;
      END
   END FE_OFN73753_n_227

   PIN FE_OFN74310_n_61
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 147.15 180.2 147.25 ;
      END
   END FE_OFN74310_n_61

   PIN FE_OFN74425_n_81
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 57.55 180.2 57.65 ;
      END
   END FE_OFN74425_n_81

   PIN FE_OFN74585_n_79
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 179.69 92.15 180.2 92.25 ;
      END
   END FE_OFN74585_n_79

   PIN FE_OFN74729_n_522
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 75.35 0.51 75.45 ;
      END
   END FE_OFN74729_n_522

   PIN FE_OFN74760_n_528
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 41.45 0 41.55 0.51 ;
      END
   END FE_OFN74760_n_528

   PIN FE_OFN75614_n_67219
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 104.45 201.49 104.55 202 ;
      END
   END FE_OFN75614_n_67219

   PIN FE_OFN79568_n_24853
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 30.95 180.2 31.05 ;
      END
   END FE_OFN79568_n_24853

   PIN FE_OFN81210_n_24583
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 72.95 180.2 73.05 ;
      END
   END FE_OFN81210_n_24583

   PIN FE_OFN85037_n_16
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 101.05 201.49 101.15 202 ;
      END
   END FE_OFN85037_n_16

   PIN FE_OFN85123_n_33
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 87.65 0 87.75 0.51 ;
      END
   END FE_OFN85123_n_33

   PIN FE_OFN85133_n_222
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 102.15 180.2 102.25 ;
      END
   END FE_OFN85133_n_222

   PIN FE_OFN85161_n_228
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 163.65 201.49 163.75 202 ;
      END
   END FE_OFN85161_n_228

   PIN FE_OFN88159_n_22979
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 78.45 201.49 78.55 202 ;
      END
   END FE_OFN88159_n_22979

   PIN FE_OFN88474_n_23035
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 57.35 180.2 57.45 ;
      END
   END FE_OFN88474_n_23035

   PIN FE_OFN90605_n_22920
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 165.55 180.2 165.65 ;
      END
   END FE_OFN90605_n_22920

   PIN FE_OFN90793_n_22919
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 158.95 180.2 159.05 ;
      END
   END FE_OFN90793_n_22919

   PIN FE_OFN91248_n_22948
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 179.69 165.55 180.2 165.65 ;
      END
   END FE_OFN91248_n_22948

   PIN FE_OFN91275_n_24566
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 52.75 180.2 52.85 ;
      END
   END FE_OFN91275_n_24566

   PIN FE_OFN91539_n_24449
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 120.55 180.2 120.65 ;
      END
   END FE_OFN91539_n_24449

   PIN FE_OFN93720_n_22938
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 130.95 0.51 131.05 ;
      END
   END FE_OFN93720_n_22938

   PIN FE_OFN94058_n_23983
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 24.45 0 24.55 0.51 ;
      END
   END FE_OFN94058_n_23983

   PIN FE_OFN98113_n_50
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 90.95 0.51 91.05 ;
      END
   END FE_OFN98113_n_50

   PIN FE_OFN98889_n_67217
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 141.25 0 141.35 0.51 ;
      END
   END FE_OFN98889_n_67217

   PIN FE_RN_2244_0
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 57.15 180.2 57.25 ;
      END
   END FE_RN_2244_0

   PIN FE_RN_4805_0
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 6.45 0 6.55 0.51 ;
      END
   END FE_RN_4805_0

   PIN a_in_203_0
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 129.55 0.51 129.65 ;
      END
   END a_in_203_0

   PIN a_in_208_0
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 94.15 0.51 94.25 ;
      END
   END a_in_208_0

   PIN a_in_208_3
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 48.75 0.51 48.85 ;
      END
   END a_in_208_3

   PIN a_in_209_2
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 129.75 0.51 129.85 ;
      END
   END a_in_209_2

   PIN a_in_20_0
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 60.65 0 60.75 0.51 ;
      END
   END a_in_20_0

   PIN a_in_20_1
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 93.55 0.51 93.65 ;
      END
   END a_in_20_1

   PIN a_in_20_2
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 12.75 0.51 12.85 ;
      END
   END a_in_20_2

   PIN a_in_20_3
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 66.75 0.51 66.85 ;
      END
   END a_in_20_3

   PIN a_in_210_2
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 129.35 0.51 129.45 ;
      END
   END a_in_210_2

   PIN a_in_210_3
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 129.55 0.51 129.65 ;
      END
   END a_in_210_3

   PIN a_in_213_0
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 192.55 0.51 192.65 ;
      END
   END a_in_213_0

   PIN a_in_22_0
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 48.55 0.51 48.65 ;
      END
   END a_in_22_0

   PIN a_in_22_1
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 125.05 0 125.15 0.51 ;
      END
   END a_in_22_1

   PIN a_in_23_0
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 132.45 0 132.55 0.51 ;
      END
   END a_in_23_0

   PIN a_in_242_2
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 148.15 0.51 148.25 ;
      END
   END a_in_242_2

   PIN a_in_243_2
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 147.95 0.51 148.05 ;
      END
   END a_in_243_2

   PIN a_in_246_1
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 111.55 0.51 111.65 ;
      END
   END a_in_246_1

   PIN a_in_247_1
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 93.15 0.51 93.25 ;
      END
   END a_in_247_1

   PIN a_in_251_2
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 174.35 0.51 174.45 ;
      END
   END a_in_251_2

   PIN a_in_253_1
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 123.45 0 123.55 0.51 ;
      END
   END a_in_253_1

   PIN a_in_253_2
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 129.15 0.51 129.25 ;
      END
   END a_in_253_2

   PIN a_in_255_2
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 191.75 0.51 191.85 ;
      END
   END a_in_255_2

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 30.5 0.255 30.7 ;
      END
   END ispd_clk

   PIN memread_edit_dist_g2_ln254_unr113_q_6_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 33.45 0 33.55 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr113_q_6_

   PIN memread_edit_dist_g2_ln254_unr48_q_0_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 96.45 0 96.55 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr48_q_0_

   PIN memread_edit_dist_g2_ln254_unr48_q_4_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 172.65 0 172.75 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr48_q_4_

   PIN memread_edit_dist_g2_ln254_unr49_q_10_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 87.45 0 87.55 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr49_q_10_

   PIN memread_edit_dist_g2_ln254_unr49_q_1_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 111.05 0 111.15 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr49_q_1_

   PIN memread_edit_dist_g2_ln254_unr49_q_2_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 163.65 0 163.75 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr49_q_2_

   PIN memread_edit_dist_g2_ln254_unr49_q_3_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 74.85 0 74.95 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr49_q_3_

   PIN memread_edit_dist_g2_ln254_unr49_q_6_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 24.05 0 24.15 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr49_q_6_

   PIN memread_edit_dist_g2_ln254_unr49_q_7_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 24.25 0 24.35 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr49_q_7_

   PIN memread_edit_dist_g2_ln254_unr49_q_8_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 32.65 0 32.75 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr49_q_8_

   PIN mux_g_ln477_q_1324_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 150.65 0 150.75 0.51 ;
      END
   END mux_g_ln477_q_1324_

   PIN mux_g_ln477_q_1344_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 48.65 0 48.75 0.51 ;
      END
   END mux_g_ln477_q_1344_

   PIN mux_g_ln477_q_1354_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 84.55 0.51 84.65 ;
      END
   END mux_g_ln477_q_1354_

   PIN mux_g_ln477_q_1481_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 110.75 180.2 110.85 ;
      END
   END mux_g_ln477_q_1481_

   PIN mux_g_ln477_q_1482_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 150.95 0.51 151.05 ;
      END
   END mux_g_ln477_q_1482_

   PIN mux_g_ln477_q_1486_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 138.75 0.51 138.85 ;
      END
   END mux_g_ln477_q_1486_

   PIN mux_g_ln477_q_1501_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 156.15 0.51 156.25 ;
      END
   END mux_g_ln477_q_1501_

   PIN mux_g_ln477_q_1518_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 6.85 201.49 6.95 202 ;
      END
   END mux_g_ln477_q_1518_

   PIN mux_g_ln477_q_1525_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 15.45 201.49 15.55 202 ;
      END
   END mux_g_ln477_q_1525_

   PIN mux_g_ln477_q_1526_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 33.25 0 33.35 0.51 ;
      END
   END mux_g_ln477_q_1526_

   PIN mux_g_ln477_q_600_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 65.25 0 65.35 0.51 ;
      END
   END mux_g_ln477_q_600_

   PIN n_1788
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 120.75 0.51 120.85 ;
      END
   END n_1788

   PIN n_1861
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 78.65 0 78.75 0.51 ;
      END
   END n_1861

   PIN n_1990
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 142.05 0 142.15 0.51 ;
      END
   END n_1990

   PIN n_2013
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 157.45 0 157.55 0.51 ;
      END
   END n_2013

   PIN n_2044
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 96.45 0 96.55 0.51 ;
      END
   END n_2044

   PIN n_2050
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 120.55 0.51 120.65 ;
      END
   END n_2050

   PIN n_2070
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 6.45 0 6.55 0.51 ;
      END
   END n_2070

   PIN n_2108
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 64.05 0 64.15 0.51 ;
      END
   END n_2108

   PIN n_2202
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 21.75 180.2 21.85 ;
      END
   END n_2202

   PIN n_2260
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 169.15 0.51 169.25 ;
      END
   END n_2260

   PIN n_23549
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 138.55 0.51 138.65 ;
      END
   END n_23549

   PIN n_23573
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 19.45 0 19.55 0.51 ;
      END
   END n_23573

   PIN n_23650
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 31.35 0.51 31.45 ;
      END
   END n_23650

   PIN n_23702
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 132.95 0.51 133.05 ;
      END
   END n_23702

   PIN n_23746
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 70.75 0.51 70.85 ;
      END
   END n_23746

   PIN n_23815
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 165.35 0.51 165.45 ;
      END
   END n_23815

   PIN n_23843
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 84.55 180.2 84.65 ;
      END
   END n_23843

   PIN n_23864
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 45.65 0 45.75 0.51 ;
      END
   END n_23864

   PIN n_23901
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 168.95 180.2 169.05 ;
      END
   END n_23901

   PIN n_23981
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 111.55 0.51 111.65 ;
      END
   END n_23981

   PIN n_23986
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 128.95 0.51 129.05 ;
      END
   END n_23986

   PIN n_2402
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 51.65 0 51.75 0.51 ;
      END
   END n_2402

   PIN n_2412
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 114.25 0 114.35 0.51 ;
      END
   END n_2412

   PIN n_24195
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 132.05 0 132.15 0.51 ;
      END
   END n_24195

   PIN n_24445
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 93.15 180.2 93.25 ;
      END
   END n_24445

   PIN n_24462
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 75.35 180.2 75.45 ;
      END
   END n_24462

   PIN n_24465
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 56.95 180.2 57.05 ;
      END
   END n_24465

   PIN n_2450
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 155.95 180.2 156.05 ;
      END
   END n_2450

   PIN n_24851
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 96.05 0 96.15 0.51 ;
      END
   END n_24851

   PIN n_24855
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 84.35 180.2 84.45 ;
      END
   END n_24855

   PIN n_25014
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 111.35 0.51 111.45 ;
      END
   END n_25014

   PIN n_25016
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 120.35 0.51 120.45 ;
      END
   END n_25016

   PIN n_2513
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 30.95 0.51 31.05 ;
      END
   END n_2513

   PIN n_25319
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 110.95 180.2 111.05 ;
      END
   END n_25319

   PIN n_2593
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 96.25 0 96.35 0.51 ;
      END
   END n_2593

   PIN n_2628
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 29.25 0 29.35 0.51 ;
      END
   END n_2628

   PIN n_2642
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 145.25 0 145.35 0.51 ;
      END
   END n_2642

   PIN n_2754
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 21.75 0.51 21.85 ;
      END
   END n_2754

   PIN n_2809
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 71.35 0.51 71.45 ;
      END
   END n_2809

   PIN n_2826
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 168.95 0.51 169.05 ;
      END
   END n_2826

   PIN n_2944
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 111.15 0.51 111.25 ;
      END
   END n_2944

   PIN n_2986
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 10.95 0.51 11.05 ;
      END
   END n_2986

   PIN n_3111
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 57.35 0.51 57.45 ;
      END
   END n_3111

   PIN n_3265
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 12.55 0.51 12.65 ;
      END
   END n_3265

   PIN n_3303
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 78.45 0 78.55 0.51 ;
      END
   END n_3303

   PIN n_48
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 110.95 0.51 111.05 ;
      END
   END n_48

   PIN n_5228837_bar
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 26.85 201.49 26.95 202 ;
      END
   END n_5228837_bar

   PIN n_5347
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 48.95 0.51 49.05 ;
      END
   END n_5347

   PIN n_5409
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 134.65 201.49 134.75 202 ;
      END
   END n_5409

   PIN n_6457
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.69 165.35 180.2 165.45 ;
      END
   END n_6457

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 180.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 180.2 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 180.2 8.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 11.745 180.2 12.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 15.745 180.2 16.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 19.745 180.2 20.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 23.745 180.2 24.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 27.745 180.2 28.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 31.745 180.2 32.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 35.745 180.2 36.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 39.745 180.2 40.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 43.745 180.2 44.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 47.745 180.2 48.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 51.745 180.2 52.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 55.745 180.2 56.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 59.745 180.2 60.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 63.745 180.2 64.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 67.745 180.2 68.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 71.745 180.2 72.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 75.745 180.2 76.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 79.745 180.2 80.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 83.745 180.2 84.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 87.745 180.2 88.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 91.745 180.2 92.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 95.745 180.2 96.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 99.745 180.2 100.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 103.745 180.2 104.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 107.745 180.2 108.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 111.745 180.2 112.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 115.745 180.2 116.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 119.745 180.2 120.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 123.745 180.2 124.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 127.745 180.2 128.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 131.745 180.2 132.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 135.745 180.2 136.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 139.745 180.2 140.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 143.745 180.2 144.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 147.745 180.2 148.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 151.745 180.2 152.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 155.745 180.2 156.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 159.745 180.2 160.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 163.745 180.2 164.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 167.745 180.2 168.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 171.745 180.2 172.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 175.745 180.2 176.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 179.745 180.2 180.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 183.745 180.2 184.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 187.745 180.2 188.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 191.745 180.2 192.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 195.745 180.2 196.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 199.745 180.2 200.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 180.2 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 180.2 6.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 9.745 180.2 10.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 13.745 180.2 14.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 17.745 180.2 18.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 21.745 180.2 22.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 25.745 180.2 26.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 29.745 180.2 30.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 33.745 180.2 34.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 37.745 180.2 38.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 41.745 180.2 42.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 45.745 180.2 46.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 49.745 180.2 50.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 53.745 180.2 54.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 57.745 180.2 58.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 61.745 180.2 62.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 65.745 180.2 66.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 69.745 180.2 70.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 73.745 180.2 74.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 77.745 180.2 78.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 81.745 180.2 82.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 85.745 180.2 86.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 89.745 180.2 90.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 93.745 180.2 94.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 97.745 180.2 98.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 101.745 180.2 102.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 105.745 180.2 106.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 109.745 180.2 110.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 113.745 180.2 114.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 117.745 180.2 118.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 121.745 180.2 122.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 125.745 180.2 126.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 129.745 180.2 130.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 133.745 180.2 134.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 137.745 180.2 138.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 141.745 180.2 142.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 145.745 180.2 146.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 149.745 180.2 150.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 153.745 180.2 154.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 157.745 180.2 158.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 161.745 180.2 162.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 165.745 180.2 166.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 169.745 180.2 170.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 173.745 180.2 174.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 177.745 180.2 178.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 181.745 180.2 182.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 185.745 180.2 186.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 189.745 180.2 190.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 193.745 180.2 194.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 197.745 180.2 198.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 201.745 180.2 202.255 ;
      END
   END vdd

   OBS
      LAYER metal1 ;
         RECT 0 0 180.2 202 ;
   END
   OBS
      LAYER metal2 ;
         RECT 0 0 180.2 202 ;
   END
   OBS
      LAYER metal3 ;
         RECT 0 0 180.2 202 ;
   END
   OBS
      LAYER metal4 ;
         RECT 0 0 180.2 202 ;
   END
   OBS
      LAYER metal5 ;
         RECT 0 0 180.2 202 ;
   END
END h3

MACRO h2
   CLASS BLOCK ;
   SIZE 180.4 BY 116 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   PIN FE_OCPN61466_FE_OFN48299_n_31625
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 179.89 32.55 180.4 32.65 ;
      END
   END FE_OCPN61466_FE_OFN48299_n_31625

   PIN FE_OCPN78682_n_32759
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 77.75 0.51 77.85 ;
      END
   END FE_OCPN78682_n_32759

   PIN FE_OCPN99272_FE_OFN46361_n_67216
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 40.85 0 40.95 0.51 ;
      END
   END FE_OCPN99272_FE_OFN46361_n_67216

   PIN FE_OCPUNCON78515_ternarymux_ln49_0_unr82_z_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 41.35 180.4 41.45 ;
      END
   END FE_OCPUNCON78515_ternarymux_ln49_0_unr82_z_3_

   PIN FE_OFN30000_n_35944
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 85.15 0.51 85.25 ;
      END
   END FE_OFN30000_n_35944

   PIN FE_OFN30327_n_36003
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 59.35 0.51 59.45 ;
      END
   END FE_OFN30327_n_36003

   PIN FE_OFN30401_n_35970
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 32.95 0.51 33.05 ;
      END
   END FE_OFN30401_n_35970

   PIN FE_OFN30534_n_36241
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 59.15 0.51 59.25 ;
      END
   END FE_OFN30534_n_36241

   PIN FE_OFN30638_n_36637
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 71.55 0.51 71.65 ;
      END
   END FE_OFN30638_n_36637

   PIN FE_OFN35164_memwrite_edit_dist_g2_ln280_unr61_en_0__4469706
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 19.35 0.51 19.45 ;
      END
   END FE_OFN35164_memwrite_edit_dist_g2_ln280_unr61_en_0__4469706

   PIN FE_OFN42686_n_15
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 7.75 180.4 7.85 ;
      END
   END FE_OFN42686_n_15

   PIN FE_OFN42687_n_15
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 161.85 115.49 161.95 116 ;
      END
   END FE_OFN42687_n_15

   PIN FE_OFN42689_n_15
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 171.65 0 171.75 0.51 ;
      END
   END FE_OFN42689_n_15

   PIN FE_OFN42935_n_2966
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 149.45 0 149.55 0.51 ;
      END
   END FE_OFN42935_n_2966

   PIN FE_OFN46788_n_26948
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 18.35 0.51 18.45 ;
      END
   END FE_OFN46788_n_26948

   PIN FE_OFN49891_n_93
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 171.25 0 171.35 0.51 ;
      END
   END FE_OFN49891_n_93

   PIN FE_OFN53694_n_91
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 7.15 0.51 7.25 ;
      END
   END FE_OFN53694_n_91

   PIN FE_OFN54144_ternarymux_ln49_0_unr61_z_10__4330982
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 77.95 0.51 78.05 ;
      END
   END FE_OFN54144_ternarymux_ln49_0_unr61_z_10__4330982

   PIN FE_OFN54360_memread_edit_dist_a_ln268_unr124_a_33__4330321
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 7.15 180.4 7.25 ;
      END
   END FE_OFN54360_memread_edit_dist_a_ln268_unr124_a_33__4330321

   PIN FE_OFN64405_a_in_3_3
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 111.45 115.49 111.55 116 ;
      END
   END FE_OFN64405_a_in_3_3

   PIN FE_OFN73421_n_32
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 154.25 0 154.35 0.51 ;
      END
   END FE_OFN73421_n_32

   PIN FE_OFN73591_n_44
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 113.45 115.49 113.55 116 ;
      END
   END FE_OFN73591_n_44

   PIN FE_OFN73647_n_15
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 7.35 180.4 7.45 ;
      END
   END FE_OFN73647_n_15

   PIN FE_OFN74017_n_31641
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 179.89 6.95 180.4 7.05 ;
      END
   END FE_OFN74017_n_31641

   PIN FE_OFN74682_n_524
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 19.35 180.4 19.45 ;
      END
   END FE_OFN74682_n_524

   PIN FE_OFN85123_n_33
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 175.45 0 175.55 0.51 ;
      END
   END FE_OFN85123_n_33

   PIN FE_OFN85607_n_82
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 128.25 115.49 128.35 116 ;
      END
   END FE_OFN85607_n_82

   PIN FE_OFN85608_n_82
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 121.45 0 121.55 0.51 ;
      END
   END FE_OFN85608_n_82

   PIN FE_OFN86767_n_36757
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 71.75 0.51 71.85 ;
      END
   END FE_OFN86767_n_36757

   PIN FE_OFN91935_n_31635
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 7.55 180.4 7.65 ;
      END
   END FE_OFN91935_n_31635

   PIN FE_OFN91977_n_857
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 141.05 115.49 141.15 116 ;
      END
   END FE_OFN91977_n_857

   PIN FE_OFN93495_ternarymux_ln49_0_unr61_z_9__4330986
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 82.95 0.51 83.05 ;
      END
   END FE_OFN93495_ternarymux_ln49_0_unr61_z_9__4330986

   PIN FE_OFN98121_n_32
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 178.65 115.49 178.75 116 ;
      END
   END FE_OFN98121_n_32

   PIN FE_RN_1501_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 18.75 180.4 18.85 ;
      END
   END FE_RN_1501_0

   PIN FE_RN_5563_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 59.95 180.4 60.05 ;
      END
   END FE_RN_5563_0

   PIN FE_RN_5983_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 59.35 0.51 59.45 ;
      END
   END FE_RN_5983_0

   PIN add_ln174_1_unr61_z_10__2985680
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 108.35 0.51 108.45 ;
      END
   END add_ln174_1_unr61_z_10__2985680

   PIN add_ln174_1_unr61_z_8__2227506
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 78.15 0.51 78.25 ;
      END
   END add_ln174_1_unr61_z_8__2227506

   PIN g2_m_82__5_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 108.15 180.4 108.25 ;
      END
   END g2_m_82__5_

   PIN g2_q63_10_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 51.55 180.4 51.65 ;
      END
   END g2_q63_10_

   PIN g2_q63_11_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 108.35 180.4 108.45 ;
      END
   END g2_q63_11_

   PIN g2_q63_2__4327386
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 18.55 180.4 18.65 ;
      END
   END g2_q63_2__4327386

   PIN g2_q63_4__4327390
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 7.95 180.4 8.05 ;
      END
   END g2_q63_4__4327390

   PIN g2_q63_6__4327379
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 71.75 180.4 71.85 ;
      END
   END g2_q63_6__4327379

   PIN g2_q63_7__4327380
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 156.65 115.49 156.75 116 ;
      END
   END g2_q63_7__4327380

   PIN g2_q63_9_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 147.65 115.49 147.75 116 ;
      END
   END g2_q63_9_

   PIN memread_edit_dist_g2_ln254_unr61_q_0_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 45.35 180.4 45.45 ;
      END
   END memread_edit_dist_g2_ln254_unr61_q_0_

   PIN memread_edit_dist_g2_ln254_unr61_q_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 14.75 180.4 14.85 ;
      END
   END memread_edit_dist_g2_ln254_unr61_q_1_

   PIN memread_edit_dist_g2_ln254_unr61_q_5_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 86.35 180.4 86.45 ;
      END
   END memread_edit_dist_g2_ln254_unr61_q_5_

   PIN memread_edit_dist_g2_ln254_unr61_q_8_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 58.95 180.4 59.05 ;
      END
   END memread_edit_dist_g2_ln254_unr61_q_8_

   PIN n_24340
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 33.55 180.4 33.65 ;
      END
   END n_24340

   PIN n_26697
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 33.55 0.51 33.65 ;
      END
   END n_26697

   PIN n_27298
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 59.15 180.4 59.25 ;
      END
   END n_27298

   PIN n_27299
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 78.55 180.4 78.65 ;
      END
   END n_27299

   PIN n_27447
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 33.9 0.255 34.1 ;
      END
   END n_27447

   PIN n_31764
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 173.05 0 173.15 0.51 ;
      END
   END n_31764

   PIN n_31953
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 115.45 115.49 115.55 116 ;
      END
   END n_31953

   PIN n_32018
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 51.15 180.4 51.25 ;
      END
   END n_32018

   PIN n_32973
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 111.85 115.49 111.95 116 ;
      END
   END n_32973

   PIN n_33099
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 156.85 115.49 156.95 116 ;
      END
   END n_33099

   PIN n_33228
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 67.95 0.51 68.05 ;
      END
   END n_33228

   PIN n_33242
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 95.55 0.51 95.65 ;
      END
   END n_33242

   PIN n_33306
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 108.15 0.51 108.25 ;
      END
   END n_33306

   PIN n_33604
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 50.75 0.51 50.85 ;
      END
   END n_33604

   PIN n_33628
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 97.15 0.51 97.25 ;
      END
   END n_33628

   PIN n_33629
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 107.95 0.51 108.05 ;
      END
   END n_33629

   PIN n_33671
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 59.55 0.51 59.65 ;
      END
   END n_33671

   PIN n_33727
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 71.95 0.51 72.05 ;
      END
   END n_33727

   PIN n_33944
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 23.55 0.51 23.65 ;
      END
   END n_33944

   PIN n_34407
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 107.75 0.51 107.85 ;
      END
   END n_34407

   PIN n_35212
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 77.1 0.255 77.3 ;
      END
   END n_35212

   PIN n_39172
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 33.15 0.51 33.25 ;
      END
   END n_39172

   PIN n_39327
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 33.35 0.51 33.45 ;
      END
   END n_39327

   PIN n_39343
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 45.75 0.51 45.85 ;
      END
   END n_39343

   PIN n_39370
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 41.15 0.51 41.25 ;
      END
   END n_39370

   PIN n_43334
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 78.05 0 78.15 0.51 ;
      END
   END n_43334

   PIN n_60455
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 102.65 0 102.75 0.51 ;
      END
   END n_60455

   PIN n_60469
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 5.55 180.4 5.65 ;
      END
   END n_60469

   PIN n_60475
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 77.35 180.4 77.45 ;
      END
   END n_60475

   PIN n_60667
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 5.75 180.4 5.85 ;
      END
   END n_60667

   PIN n_64828
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 180.145 77.7 180.4 77.9 ;
      END
   END n_64828

   PIN n_66478
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 51.15 0.51 51.25 ;
      END
   END n_66478

   PIN ternarymux_ln49_0_unr61_z_8__4330990
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 113.65 0 113.75 0.51 ;
      END
   END ternarymux_ln49_0_unr61_z_8__4330990

   PIN ternarymux_ln49_0_unr62_z_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 14.55 0.51 14.65 ;
      END
   END ternarymux_ln49_0_unr62_z_1_

   PIN ternarymux_ln49_0_unr62_z_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 49.95 0.51 50.05 ;
      END
   END ternarymux_ln49_0_unr62_z_3_

   PIN ternarymux_ln49_0_unr62_z_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 50.35 0.51 50.45 ;
      END
   END ternarymux_ln49_0_unr62_z_4_

   PIN ternarymux_ln49_0_unr62_z_5_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 58.95 0.51 59.05 ;
      END
   END ternarymux_ln49_0_unr62_z_5_

   PIN ternarymux_ln49_0_unr62_z_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 50.55 0.51 50.65 ;
      END
   END ternarymux_ln49_0_unr62_z_7_

   PIN ternarymux_ln49_0_unr82_z_10__4331318
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 107.55 0.51 107.65 ;
      END
   END ternarymux_ln49_0_unr82_z_10__4331318

   PIN ternarymux_ln49_0_unr82_z_8__4331326
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 51.35 180.4 51.45 ;
      END
   END ternarymux_ln49_0_unr82_z_8__4331326

   PIN ternarymux_ln49_5_unr62_z_0_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 77.55 0.51 77.65 ;
      END
   END ternarymux_ln49_5_unr62_z_0_

   PIN ternarymux_ln49_6_unr82_z_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 45.55 180.4 45.65 ;
      END
   END ternarymux_ln49_6_unr82_z_12_

   PIN ternarymux_ln49_8_unr82_z_11_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 67.95 180.4 68.05 ;
      END
   END ternarymux_ln49_8_unr82_z_11_

   PIN FE_OCPN57527_FE_OFN47118_n_23039
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 33.35 180.4 33.45 ;
      END
   END FE_OCPN57527_FE_OFN47118_n_23039

   PIN FE_OCPN57867_n_93
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 45.15 180.4 45.25 ;
      END
   END FE_OCPN57867_n_93

   PIN FE_OCPN58733_FE_OFN46361_n_67216
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 151.65 115.49 151.75 116 ;
      END
   END FE_OCPN58733_FE_OFN46361_n_67216

   PIN FE_OCPN60536_FE_OFN48705_n_59125
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 135.85 0 135.95 0.51 ;
      END
   END FE_OCPN60536_FE_OFN48705_n_59125

   PIN FE_OCPN62476_n_65256
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 59.65 115.49 59.75 116 ;
      END
   END FE_OCPN62476_n_65256

   PIN FE_OCPN78686_ternarymux_ln49_0_unr62_z_4_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 71.35 0.51 71.45 ;
      END
   END FE_OCPN78686_ternarymux_ln49_0_unr62_z_4_

   PIN FE_OCPN78960_add_ln174_1_unr81_z_8__2227792
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 83.95 180.4 84.05 ;
      END
   END FE_OCPN78960_add_ln174_1_unr81_z_8__2227792

   PIN FE_OCP_DRV_N76505_n_32047
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 59.35 180.4 59.45 ;
      END
   END FE_OCP_DRV_N76505_n_32047

   PIN FE_OFN29317_n_524
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 12.85 0 12.95 0.51 ;
      END
   END FE_OFN29317_n_524

   PIN FE_OFN30108_n_36239
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 49.95 180.4 50.05 ;
      END
   END FE_OFN30108_n_36239

   PIN FE_OFN30153_n_36584
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 44.95 180.4 45.05 ;
      END
   END FE_OFN30153_n_36584

   PIN FE_OFN30155_n_36438
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 147.85 0 147.95 0.51 ;
      END
   END FE_OFN30155_n_36438

   PIN FE_OFN30163_n_36334
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 20.95 180.4 21.05 ;
      END
   END FE_OFN30163_n_36334

   PIN FE_OFN30326_n_36003
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 23.35 180.4 23.45 ;
      END
   END FE_OFN30326_n_36003

   PIN FE_OFN30400_n_35970
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 33.15 180.4 33.25 ;
      END
   END FE_OFN30400_n_35970

   PIN FE_OFN30637_n_36637
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 50.95 180.4 51.05 ;
      END
   END FE_OFN30637_n_36637

   PIN FE_OFN30801_n_36371
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 6.95 180.4 7.05 ;
      END
   END FE_OFN30801_n_36371

   PIN FE_OFN31996_n_31637
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 84.95 0.51 85.05 ;
      END
   END FE_OFN31996_n_31637

   PIN FE_OFN34194_n_82
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 165.85 115.49 165.95 116 ;
      END
   END FE_OFN34194_n_82

   PIN FE_OFN42374_n_44
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 113.65 0 113.75 0.51 ;
      END
   END FE_OFN42374_n_44

   PIN FE_OFN42487_n_33
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 149.25 115.49 149.35 116 ;
      END
   END FE_OFN42487_n_33

   PIN FE_OFN46247_a_in_6_2
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 45.55 0.51 45.65 ;
      END
   END FE_OFN46247_a_in_6_2

   PIN FE_OFN46272_a_in_3_3
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 111.65 115.49 111.75 116 ;
      END
   END FE_OFN46272_a_in_3_3

   PIN FE_OFN47675_n_22885
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 174.45 0 174.55 0.51 ;
      END
   END FE_OFN47675_n_22885

   PIN FE_OFN47898_n_31635
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 6.95 0.51 7.05 ;
      END
   END FE_OFN47898_n_31635

   PIN FE_OFN48370_n_31641
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 95.75 0.51 95.85 ;
      END
   END FE_OFN48370_n_31641

   PIN FE_OFN50337_n_64841
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 96.95 0.51 97.05 ;
      END
   END FE_OFN50337_n_64841

   PIN FE_OFN50338_n_64841
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 50.55 0.51 50.65 ;
      END
   END FE_OFN50338_n_64841

   PIN FE_OFN50556_lt_ln49_6_unr82_z
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 180.145 33.9 180.4 34.1 ;
      END
   END FE_OFN50556_lt_ln49_6_unr82_z

   PIN FE_OFN50580_lt_ln49_6_unr61_z
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 70.9 0.255 71.1 ;
      END
   END FE_OFN50580_lt_ln49_6_unr61_z

   PIN FE_OFN53691_n_91
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 21.85 0 21.95 0.51 ;
      END
   END FE_OFN53691_n_91

   PIN FE_OFN55966_ternarymux_ln49_0_unr61_z_5_
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 179.89 5.55 180.4 5.65 ;
      END
   END FE_OFN55966_ternarymux_ln49_0_unr61_z_5_

   PIN FE_OFN55978_ternarymux_ln49_0_unr61_z_10__4330982
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 168.05 0 168.15 0.51 ;
      END
   END FE_OFN55978_ternarymux_ln49_0_unr61_z_10__4330982

   PIN FE_OFN70914_memwrite_edit_dist_g2_ln280_unr61_en_0__4469706
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 44.45 115.49 44.55 116 ;
      END
   END FE_OFN70914_memwrite_edit_dist_g2_ln280_unr61_en_0__4469706

   PIN FE_OFN70915_n_21264
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 55.45 115.49 55.55 116 ;
      END
   END FE_OFN70915_n_21264

   PIN FE_OFN85983_FE_OCPN60599_FE_OFN48344_n_31639
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 98.15 0.51 98.25 ;
      END
   END FE_OFN85983_FE_OCPN60599_FE_OFN48344_n_31639

   PIN FE_OFN86656_n_36241
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 41.15 180.4 41.25 ;
      END
   END FE_OFN86656_n_36241

   PIN FE_OFN86766_n_36757
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 50.75 180.4 50.85 ;
      END
   END FE_OFN86766_n_36757

   PIN FE_OFN88247_n_31634
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 14.95 180.4 15.05 ;
      END
   END FE_OFN88247_n_31634

   PIN FE_OFN90783_n_67217
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 32.95 180.4 33.05 ;
      END
   END FE_OFN90783_n_67217

   PIN FE_OFN91976_n_857
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 142.65 0 142.75 0.51 ;
      END
   END FE_OFN91976_n_857

   PIN FE_OFN92515_n_31642
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 48.45 115.49 48.55 116 ;
      END
   END FE_OFN92515_n_31642

   PIN FE_OFN93183_FE_OCPN61464_FE_OFN48299_n_31625
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 129.85 115.49 129.95 116 ;
      END
   END FE_OFN93183_FE_OCPN61464_FE_OFN48299_n_31625

   PIN FE_OFN98340_ternarymux_ln49_0_unr62_z_2_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 57.95 0.51 58.05 ;
      END
   END FE_OFN98340_ternarymux_ln49_0_unr62_z_2_

   PIN FE_RN_1499_0
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 165.45 0 165.55 0.51 ;
      END
   END FE_RN_1499_0

   PIN a_in_3_3
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 86.55 0.51 86.65 ;
      END
   END a_in_3_3

   PIN add_ln174_1_unr60_z_10__2985662
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 175.25 0 175.35 0.51 ;
      END
   END add_ln174_1_unr60_z_10__2985662

   PIN add_ln174_1_unr60_z_8__2227484
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 174.85 0 174.95 0.51 ;
      END
   END add_ln174_1_unr60_z_8__2227484

   PIN add_ln174_1_unr60_z_9__2985661
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 175.05 0 175.15 0.51 ;
      END
   END add_ln174_1_unr60_z_9__2985661

   PIN add_ln174_1_unr81_z_10__2985914
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 154.25 115.49 154.35 116 ;
      END
   END add_ln174_1_unr81_z_10__2985914

   PIN add_ln174_1_unr81_z_9__2985913
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 97.35 180.4 97.45 ;
      END
   END add_ln174_1_unr81_z_9__2985913

   PIN g2_m_81__6_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 95.95 0.51 96.05 ;
      END
   END g2_m_81__6_

   PIN g2_q63_3__4327387
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 149.65 0 149.75 0.51 ;
      END
   END g2_q63_3__4327387

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 131 0 131.2 0.255 ;
      END
   END ispd_clk

   PIN memread_edit_dist_a_ln268_unr124_a_33__4330321
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 12.85 0 12.95 0.51 ;
      END
   END memread_edit_dist_a_ln268_unr124_a_33__4330321

   PIN mux_g_ln477_q_538_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 166.05 115.49 166.15 116 ;
      END
   END mux_g_ln477_q_538_

   PIN n_15
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 57.85 0 57.95 0.51 ;
      END
   END n_15

   PIN n_26724
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 77.15 180.4 77.25 ;
      END
   END n_26724

   PIN n_27093
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 32.95 0.51 33.05 ;
      END
   END n_27093

   PIN n_27289
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 76.95 180.4 77.05 ;
      END
   END n_27289

   PIN n_27691
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 106.65 0 106.75 0.51 ;
      END
   END n_27691

   PIN n_28399
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 180.145 96.9 180.4 97.1 ;
      END
   END n_28399

   PIN n_28421
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 68.35 180.4 68.45 ;
      END
   END n_28421

   PIN n_28422
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 71.55 180.4 71.65 ;
      END
   END n_28422

   PIN n_28515
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 71.35 180.4 71.45 ;
      END
   END n_28515

   PIN n_2966
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 149.65 115.49 149.75 116 ;
      END
   END n_2966

   PIN n_31796
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 140.85 115.49 140.95 116 ;
      END
   END n_31796

   PIN n_32
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 138.85 0 138.95 0.51 ;
      END
   END n_32

   PIN n_33098
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 156.85 115.49 156.95 116 ;
      END
   END n_33098

   PIN n_33248
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 82.45 0 82.55 0.51 ;
      END
   END n_33248

   PIN n_33317
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 59.75 180.4 59.85 ;
      END
   END n_33317

   PIN n_33768
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 112.65 0 112.75 0.51 ;
      END
   END n_33768

   PIN n_34371
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 50.15 0.51 50.25 ;
      END
   END n_34371

   PIN n_35200
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 64.05 0 64.15 0.51 ;
      END
   END n_35200

   PIN n_35944
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 59.55 180.4 59.65 ;
      END
   END n_35944

   PIN n_36245
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 14.55 180.4 14.65 ;
      END
   END n_36245

   PIN n_39238
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 77.55 0.51 77.65 ;
      END
   END n_39238

   PIN n_48546
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 180.145 50.3 180.4 50.5 ;
      END
   END n_48546

   PIN n_51746
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 45.35 0.51 45.45 ;
      END
   END n_51746

   PIN n_59964
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 180.145 70.9 180.4 71.1 ;
      END
   END n_59964

   PIN n_60462
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 18.55 0.51 18.65 ;
      END
   END n_60462

   PIN n_60666
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 84.95 180.4 85.05 ;
      END
   END n_60666

   PIN n_61220
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 78.35 180.4 78.45 ;
      END
   END n_61220

   PIN n_61225
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 67.75 180.4 67.85 ;
      END
   END n_61225

   PIN n_62440
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 45.15 0.51 45.25 ;
      END
   END n_62440

   PIN n_62441
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 44.95 0.51 45.05 ;
      END
   END n_62441

   PIN n_62442
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 18.75 0.51 18.85 ;
      END
   END n_62442

   PIN n_62443
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 75.85 0 75.95 0.51 ;
      END
   END n_62443

   PIN n_64842
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 71.95 180.4 72.05 ;
      END
   END n_64842

   PIN n_66477
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 166.45 0 166.55 0.51 ;
      END
   END n_66477

   PIN ternarymux_ln49_0_unr61_z_0_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 105.25 0 105.35 0.51 ;
      END
   END ternarymux_ln49_0_unr61_z_0_

   PIN ternarymux_ln49_0_unr61_z_1_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 58.65 0 58.75 0.51 ;
      END
   END ternarymux_ln49_0_unr61_z_1_

   PIN ternarymux_ln49_0_unr61_z_2_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 94.45 0 94.55 0.51 ;
      END
   END ternarymux_ln49_0_unr61_z_2_

   PIN ternarymux_ln49_0_unr61_z_3_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 54.45 0 54.55 0.51 ;
      END
   END ternarymux_ln49_0_unr61_z_3_

   PIN ternarymux_ln49_0_unr61_z_4_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 50.95 0.51 51.05 ;
      END
   END ternarymux_ln49_0_unr61_z_4_

   PIN ternarymux_ln49_0_unr61_z_6_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 70.65 0 70.75 0.51 ;
      END
   END ternarymux_ln49_0_unr61_z_6_

   PIN ternarymux_ln49_0_unr61_z_7_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 43.85 0 43.95 0.51 ;
      END
   END ternarymux_ln49_0_unr61_z_7_

   PIN ternarymux_ln49_0_unr61_z_9__4330986
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 127.45 0 127.55 0.51 ;
      END
   END ternarymux_ln49_0_unr61_z_9__4330986

   PIN ternarymux_ln49_0_unr62_z_8__4331006
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 58.95 0.51 59.05 ;
      END
   END ternarymux_ln49_0_unr62_z_8__4331006

   PIN ternarymux_ln49_0_unr62_z_9__4331002
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 83.15 0.51 83.25 ;
      END
   END ternarymux_ln49_0_unr62_z_9__4331002

   PIN ternarymux_ln49_0_unr82_z_3_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 78.15 180.4 78.25 ;
      END
   END ternarymux_ln49_0_unr82_z_3_

   PIN ternarymux_ln49_0_unr82_z_5_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 107.95 180.4 108.05 ;
      END
   END ternarymux_ln49_0_unr82_z_5_

   PIN ternarymux_ln49_8_unr82_z_9_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 179.89 68.15 180.4 68.25 ;
      END
   END ternarymux_ln49_8_unr82_z_9_

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 180.4 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 180.4 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 180.4 8.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 11.745 180.4 12.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 15.745 180.4 16.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 19.745 180.4 20.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 23.745 180.4 24.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 27.745 180.4 28.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 31.745 180.4 32.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 35.745 180.4 36.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 39.745 180.4 40.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 43.745 180.4 44.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 47.745 180.4 48.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 51.745 180.4 52.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 55.745 180.4 56.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 59.745 180.4 60.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 63.745 180.4 64.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 67.745 180.4 68.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 71.745 180.4 72.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 75.745 180.4 76.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 79.745 180.4 80.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 83.745 180.4 84.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 87.745 180.4 88.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 91.745 180.4 92.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 95.745 180.4 96.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 99.745 180.4 100.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 103.745 180.4 104.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 107.745 180.4 108.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 111.745 180.4 112.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 115.745 180.4 116.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 180.4 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 180.4 6.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 9.745 180.4 10.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 13.745 180.4 14.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 17.745 180.4 18.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 21.745 180.4 22.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 25.745 180.4 26.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 29.745 180.4 30.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 33.745 180.4 34.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 37.745 180.4 38.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 41.745 180.4 42.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 45.745 180.4 46.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 49.745 180.4 50.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 53.745 180.4 54.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 57.745 180.4 58.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 61.745 180.4 62.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 65.745 180.4 66.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 69.745 180.4 70.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 73.745 180.4 74.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 77.745 180.4 78.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 81.745 180.4 82.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 85.745 180.4 86.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 89.745 180.4 90.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 93.745 180.4 94.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 97.745 180.4 98.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 101.745 180.4 102.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 105.745 180.4 106.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 109.745 180.4 110.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 113.745 180.4 114.255 ;
      END
   END vdd

   OBS
      LAYER metal1 ;
         RECT 0 0 180.4 116 ;
   END
   OBS
      LAYER metal2 ;
         RECT 0 0 180.4 116 ;
   END
   OBS
      LAYER metal3 ;
         RECT 0 0 180.4 116 ;
   END
   OBS
      LAYER metal4 ;
         RECT 0 0 180.4 116 ;
   END
   OBS
      LAYER metal5 ;
         RECT 0 0 180.4 116 ;
   END
END h2

MACRO h1
   CLASS BLOCK ;
   SIZE 183 BY 250 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   PIN FE_OCPN56133_n_35331
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 169.95 183 170.05 ;
      END
   END FE_OCPN56133_n_35331

   PIN FE_OCPN57867_n_93
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 178.05 0 178.15 0.51 ;
      END
   END FE_OCPN57867_n_93

   PIN FE_OCPN58711_n_33467_bar
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 110.85 0 110.95 0.51 ;
      END
   END FE_OCPN58711_n_33467_bar

   PIN FE_OCPN60456_memread_edit_dist_a_ln268_unr124_a_9__4329837
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 54.95 183 55.05 ;
      END
   END FE_OCPN60456_memread_edit_dist_a_ln268_unr124_a_9__4329837

   PIN FE_OCPN60530_FE_OFN48705_n_59125
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 29.65 0 29.75 0.51 ;
      END
   END FE_OCPN60530_FE_OFN48705_n_59125

   PIN FE_OCPN61465_FE_OFN48299_n_31625
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 144.15 0.51 144.25 ;
      END
   END FE_OCPN61465_FE_OFN48299_n_31625

   PIN FE_OCPN62334_n_58046
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 196.55 0.51 196.65 ;
      END
   END FE_OCPN62334_n_58046

   PIN FE_OCPN62350_n_65199
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 136.05 0 136.15 0.51 ;
      END
   END FE_OCPN62350_n_65199

   PIN FE_OCPN62854_n_33487_bar
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 127.45 0 127.55 0.51 ;
      END
   END FE_OCPN62854_n_33487_bar

   PIN FE_OCPN63056_FE_OFN47982_n_23035
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 62.75 183 62.85 ;
      END
   END FE_OCPN63056_FE_OFN47982_n_23035

   PIN FE_OCPN63788_FE_OFN48830_n_31626
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 56.85 0 56.95 0.51 ;
      END
   END FE_OCPN63788_FE_OFN48830_n_31626

   PIN FE_OCPN63795_FE_OFN48307_n_31634
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 38.85 0 38.95 0.51 ;
      END
   END FE_OCPN63795_FE_OFN48307_n_31634

   PIN FE_OCPN78052_FE_OFN48367_n_31641
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 235.35 0.51 235.45 ;
      END
   END FE_OCPN78052_FE_OFN48367_n_31641

   PIN FE_OCPN95861_n_58050
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 56.85 249.49 56.95 250 ;
      END
   END FE_OCPN95861_n_58050

   PIN FE_OFN28637_n_36328
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 143.35 183 143.45 ;
      END
   END FE_OFN28637_n_36328

   PIN FE_OFN28734_n_40187
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 20.8 0 21 0.255 ;
      END
   END FE_OFN28734_n_40187

   PIN FE_OFN30022_n_36839
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 206.75 0.51 206.85 ;
      END
   END FE_OFN30022_n_36839

   PIN FE_OFN30049_n_36035
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 110.95 0.51 111.05 ;
      END
   END FE_OFN30049_n_36035

   PIN FE_OFN30051_n_36014
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 180.55 0.51 180.65 ;
      END
   END FE_OFN30051_n_36014

   PIN FE_OFN30065_n_37068
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 200.15 0.51 200.25 ;
      END
   END FE_OFN30065_n_37068

   PIN FE_OFN30075_n_36916
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 134.35 0.51 134.45 ;
      END
   END FE_OFN30075_n_36916

   PIN FE_OFN30206_n_36803
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 80.95 0.51 81.05 ;
      END
   END FE_OFN30206_n_36803

   PIN FE_OFN30245_n_37046
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 161.35 0.51 161.45 ;
      END
   END FE_OFN30245_n_37046

   PIN FE_OFN30248_n_37029
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 97.95 0.51 98.05 ;
      END
   END FE_OFN30248_n_37029

   PIN FE_OFN30266_n_36785
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 133.95 0.51 134.05 ;
      END
   END FE_OFN30266_n_36785

   PIN FE_OFN30301_n_36379
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 53.35 0.51 53.45 ;
      END
   END FE_OFN30301_n_36379

   PIN FE_OFN30337_n_36733
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 161.55 0.51 161.65 ;
      END
   END FE_OFN30337_n_36733

   PIN FE_OFN30356_n_35984
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 206.35 0.51 206.45 ;
      END
   END FE_OFN30356_n_35984

   PIN FE_OFN30389_n_34771
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 177.45 0 177.55 0.51 ;
      END
   END FE_OFN30389_n_34771

   PIN FE_OFN30460_n_36563
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 151.95 0.51 152.05 ;
      END
   END FE_OFN30460_n_36563

   PIN FE_OFN30471_n_35975
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 220.95 0.51 221.05 ;
      END
   END FE_OFN30471_n_35975

   PIN FE_OFN30521_n_36965
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 82.95 0.51 83.05 ;
      END
   END FE_OFN30521_n_36965

   PIN FE_OFN30531_n_36390
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 179.35 0.51 179.45 ;
      END
   END FE_OFN30531_n_36390

   PIN FE_OFN30574_n_36953
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 187.95 0.51 188.05 ;
      END
   END FE_OFN30574_n_36953

   PIN FE_OFN30590_n_36899
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 125.15 0.51 125.25 ;
      END
   END FE_OFN30590_n_36899

   PIN FE_OFN30594_n_36874
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 107.55 0.51 107.65 ;
      END
   END FE_OFN30594_n_36874

   PIN FE_OFN30641_n_36622
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 134.55 0.51 134.65 ;
      END
   END FE_OFN30641_n_36622

   PIN FE_OFN30660_n_36401
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 215.35 0.51 215.45 ;
      END
   END FE_OFN30660_n_36401

   PIN FE_OFN30662_n_36399
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 206.55 0.51 206.65 ;
      END
   END FE_OFN30662_n_36399

   PIN FE_OFN30685_n_36201
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 90.95 0.51 91.05 ;
      END
   END FE_OFN30685_n_36201

   PIN FE_OFN30698_n_36086
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 109.55 0.51 109.65 ;
      END
   END FE_OFN30698_n_36086

   PIN FE_OFN30707_n_36073
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 134.15 0.51 134.25 ;
      END
   END FE_OFN30707_n_36073

   PIN FE_OFN30717_n_36030
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 99.15 0.51 99.25 ;
      END
   END FE_OFN30717_n_36030

   PIN FE_OFN30724_n_36015
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 172.15 0.51 172.25 ;
      END
   END FE_OFN30724_n_36015

   PIN FE_OFN30729_n_35986
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 72.95 0.51 73.05 ;
      END
   END FE_OFN30729_n_35986

   PIN FE_OFN30733_n_35978
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 226.95 0.51 227.05 ;
      END
   END FE_OFN30733_n_35978

   PIN FE_OFN30796_n_36565
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 103.35 0.51 103.45 ;
      END
   END FE_OFN30796_n_36565

   PIN FE_OFN30810_n_34732
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 111.25 0 111.35 0.51 ;
      END
   END FE_OFN30810_n_34732

   PIN FE_OFN30812_n_34732
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 107.35 183 107.45 ;
      END
   END FE_OFN30812_n_34732

   PIN FE_OFN30828_n_36787
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 81.65 249.49 81.75 250 ;
      END
   END FE_OFN30828_n_36787

   PIN FE_OFN30862_n_34779
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 102.05 0 102.15 0.51 ;
      END
   END FE_OFN30862_n_34779

   PIN FE_OFN30869_n_36922
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 244.95 0.51 245.05 ;
      END
   END FE_OFN30869_n_36922

   PIN FE_OFN30904_n_35995
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 134.35 0.51 134.45 ;
      END
   END FE_OFN30904_n_35995

   PIN FE_OFN31034_n_34785
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 160.05 0 160.15 0.51 ;
      END
   END FE_OFN31034_n_34785

   PIN FE_OFN32007_n_31638
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 134.75 0.51 134.85 ;
      END
   END FE_OFN32007_n_31638

   PIN FE_OFN32021_n_31639
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 43.95 0.51 44.05 ;
      END
   END FE_OFN32021_n_31639

   PIN FE_OFN32360_n_21259
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 161.35 0.51 161.45 ;
      END
   END FE_OFN32360_n_21259

   PIN FE_OFN33793_n_3370
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 101.85 0 101.95 0.51 ;
      END
   END FE_OFN33793_n_3370

   PIN FE_OFN34105_n_86
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 52.25 0 52.35 0.51 ;
      END
   END FE_OFN34105_n_86

   PIN FE_OFN34914_n_53413
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 152.15 0.51 152.25 ;
      END
   END FE_OFN34914_n_53413

   PIN FE_OFN34942_n_51091
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 161.75 0.51 161.85 ;
      END
   END FE_OFN34942_n_51091

   PIN FE_OFN41931_n_230
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 137.85 0 137.95 0.51 ;
      END
   END FE_OFN41931_n_230

   PIN FE_OFN42169_n_53
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 173.85 249.49 173.95 250 ;
      END
   END FE_OFN42169_n_53

   PIN FE_OFN42913_n_3242
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 174.75 183 174.85 ;
      END
   END FE_OFN42913_n_3242

   PIN FE_OFN43005_n_35325
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 173.65 0 173.75 0.51 ;
      END
   END FE_OFN43005_n_35325

   PIN FE_OFN43958_mux_g_ln477_q_520_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 125.05 249.49 125.15 250 ;
      END
   END FE_OFN43958_mux_g_ln477_q_520_

   PIN FE_OFN47854_n_23045
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 105.25 249.49 105.35 250 ;
      END
   END FE_OFN47854_n_23045

   PIN FE_OFN48299_n_31625
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 84.05 0 84.15 0.51 ;
      END
   END FE_OFN48299_n_31625

   PIN FE_OFN48313_n_31634
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 178.9 0.255 179.1 ;
      END
   END FE_OFN48313_n_31634

   PIN FE_OFN48316_n_31634
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 144.95 0.51 145.05 ;
      END
   END FE_OFN48316_n_31634

   PIN FE_OFN48344_n_31639
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 11.85 0 11.95 0.51 ;
      END
   END FE_OFN48344_n_31639

   PIN FE_OFN48367_n_31641
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 116.75 0.51 116.85 ;
      END
   END FE_OFN48367_n_31641

   PIN FE_OFN48368_n_31641
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 7.65 0 7.75 0.51 ;
      END
   END FE_OFN48368_n_31641

   PIN FE_OFN48708_n_59125
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 115.95 0.51 116.05 ;
      END
   END FE_OFN48708_n_59125

   PIN FE_OFN48845_n_31626
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 116.15 0.51 116.25 ;
      END
   END FE_OFN48845_n_31626

   PIN FE_OFN48846_n_31626
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 233.55 0.51 233.65 ;
      END
   END FE_OFN48846_n_31626

   PIN FE_OFN48848_n_31626
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 146.45 0 146.55 0.51 ;
      END
   END FE_OFN48848_n_31626

   PIN FE_OFN49702_n_87
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 57.05 249.49 57.15 250 ;
      END
   END FE_OFN49702_n_87

   PIN FE_OFN49703_n_87
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 93.05 249.49 93.15 250 ;
      END
   END FE_OFN49703_n_87

   PIN FE_OFN50544_lt_ln49_6_unr75_z
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 180.15 0.51 180.25 ;
      END
   END FE_OFN50544_lt_ln49_6_unr75_z

   PIN FE_OFN50546_lt_ln49_6_unr75_z
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 168.95 0.51 169.05 ;
      END
   END FE_OFN50546_lt_ln49_6_unr75_z

   PIN FE_OFN70357_n_36808
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 217.15 183 217.25 ;
      END
   END FE_OFN70357_n_36808

   PIN FE_OFN71105_memwrite_edit_dist_g2_ln280_unr73_en_0__4469519
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 233.55 0.51 233.65 ;
      END
   END FE_OFN71105_memwrite_edit_dist_g2_ln280_unr73_en_0__4469519

   PIN FE_OFN71827_n_51730
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 205.55 0.51 205.65 ;
      END
   END FE_OFN71827_n_51730

   PIN FE_OFN73372_n_20
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 160.65 249.49 160.75 250 ;
      END
   END FE_OFN73372_n_20

   PIN FE_OFN73646_n_15
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 108.85 249.49 108.95 250 ;
      END
   END FE_OFN73646_n_15

   PIN FE_OFN73661_n_29
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 65.85 249.49 65.95 250 ;
      END
   END FE_OFN73661_n_29

   PIN FE_OFN73975_n_32261
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 166.95 0.51 167.05 ;
      END
   END FE_OFN73975_n_32261

   PIN FE_OFN74037_n_31638
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 83.85 0 83.95 0.51 ;
      END
   END FE_OFN74037_n_31638

   PIN FE_OFN74082_n_59052
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 52.75 0.51 52.85 ;
      END
   END FE_OFN74082_n_59052

   PIN FE_OFN74310_n_61
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 5.15 183 5.25 ;
      END
   END FE_OFN74310_n_61

   PIN FE_OFN74580_n_79
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 57.05 0 57.15 0.51 ;
      END
   END FE_OFN74580_n_79

   PIN FE_OFN74879_n_36980
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 62.55 0.51 62.65 ;
      END
   END FE_OFN74879_n_36980

   PIN FE_OFN74969_n_36218
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 74.95 0.51 75.05 ;
      END
   END FE_OFN74969_n_36218

   PIN FE_OFN75080_n_34770
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 178.05 0 178.15 0.51 ;
      END
   END FE_OFN75080_n_34770

   PIN FE_OFN75216_n_35297
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 146.65 249.49 146.75 250 ;
      END
   END FE_OFN75216_n_35297

   PIN FE_OFN75258_n_35301
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 15.35 183 15.45 ;
      END
   END FE_OFN75258_n_35301

   PIN FE_OFN75313_n_35325
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 143.75 183 143.85 ;
      END
   END FE_OFN75313_n_35325

   PIN FE_OFN75550_FE_OCPN62021_FE_OFN50813_n_67216
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 18.35 183 18.45 ;
      END
   END FE_OFN75550_FE_OCPN62021_FE_OFN50813_n_67216

   PIN FE_OFN75725_n_35331
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 245.15 183 245.25 ;
      END
   END FE_OFN75725_n_35331

   PIN FE_OFN84025_n_21287
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 116.35 0.51 116.45 ;
      END
   END FE_OFN84025_n_21287

   PIN FE_OFN84037_n_7936
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 27.15 183 27.25 ;
      END
   END FE_OFN84037_n_7936

   PIN FE_OFN85021_n_57
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 148.85 249.49 148.95 250 ;
      END
   END FE_OFN85021_n_57

   PIN FE_OFN85096_n_30
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 74.85 249.49 74.95 250 ;
      END
   END FE_OFN85096_n_30

   PIN FE_OFN85107_n_53
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 142.85 249.49 142.95 250 ;
      END
   END FE_OFN85107_n_53

   PIN FE_OFN85118_n_15
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 236.95 183 237.05 ;
      END
   END FE_OFN85118_n_15

   PIN FE_OFN85990_n_31637
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 141.15 0.51 141.25 ;
      END
   END FE_OFN85990_n_31637

   PIN FE_OFN86082_g2_q72_2__4327665
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 89.35 183 89.45 ;
      END
   END FE_OFN86082_g2_q72_2__4327665

   PIN FE_OFN86624_n_36643
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 155.15 0.51 155.25 ;
      END
   END FE_OFN86624_n_36643

   PIN FE_OFN86680_n_36864
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 152.75 0.51 152.85 ;
      END
   END FE_OFN86680_n_36864

   PIN FE_OFN86686_n_35998
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 74.15 0.51 74.25 ;
      END
   END FE_OFN86686_n_35998

   PIN FE_OFN86751_n_36820
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 161.55 0.51 161.65 ;
      END
   END FE_OFN86751_n_36820

   PIN FE_OFN86757_n_36061
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 98.15 0.51 98.25 ;
      END
   END FE_OFN86757_n_36061

   PIN FE_OFN86879_n_36948
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 49.35 0.51 49.45 ;
      END
   END FE_OFN86879_n_36948

   PIN FE_OFN86936_n_36221
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 242.55 0.51 242.65 ;
      END
   END FE_OFN86936_n_36221

   PIN FE_OFN87036_n_35936
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 107.75 0.51 107.85 ;
      END
   END FE_OFN87036_n_35936

   PIN FE_OFN87056_n_36888
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 180.75 0.51 180.85 ;
      END
   END FE_OFN87056_n_36888

   PIN FE_OFN87975_n_35283
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 72.95 183 73.05 ;
      END
   END FE_OFN87975_n_35283

   PIN FE_OFN88306_n_65239
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 170.95 0.51 171.05 ;
      END
   END FE_OFN88306_n_65239

   PIN FE_OFN94568_n_31625
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 62.05 0 62.15 0.51 ;
      END
   END FE_OFN94568_n_31625

   PIN FE_OFN94908_n_31626
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 4.95 183 5.05 ;
      END
   END FE_OFN94908_n_31626

   PIN FE_OFN95909_n_65250
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 125.35 0.51 125.45 ;
      END
   END FE_OFN95909_n_65250

   PIN FE_OFN98159_n_230
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 164.45 249.49 164.55 250 ;
      END
   END FE_OFN98159_n_230

   PIN FE_OFN98509_n_37004
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 161.75 0.51 161.85 ;
      END
   END FE_OFN98509_n_37004

   PIN FE_OFN98531_n_36062
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 85.35 0.51 85.45 ;
      END
   END FE_OFN98531_n_36062

   PIN FE_RN_3498_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 215.35 0.51 215.45 ;
      END
   END FE_RN_3498_0

   PIN add_85532_72_n_4327722
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 216.95 0.51 217.05 ;
      END
   END add_85532_72_n_4327722

   PIN add_85538_72_n_4327812
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 92.45 0 92.55 0.51 ;
      END
   END add_85538_72_n_4327812

   PIN g2_bridge202_rtl_ce_en_3755253_bar
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 216.3 0.255 216.5 ;
      END
   END g2_bridge202_rtl_ce_en_3755253_bar

   PIN g2_bridge208_rtl_ce_en_3756288
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 43.35 0.51 43.45 ;
      END
   END g2_bridge208_rtl_ce_en_3756288

   PIN g2_q72_1__4327663
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 109.15 0.51 109.25 ;
      END
   END g2_q72_1__4327663

   PIN g2_q77_1__4327814
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 62.35 183 62.45 ;
      END
   END g2_q77_1__4327814

   PIN g2_q77_3__4327817
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 72.15 183 72.25 ;
      END
   END g2_q77_3__4327817

   PIN g2_q78_10_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 100.45 0 100.55 0.51 ;
      END
   END g2_q78_10_

   PIN g2_q78_8_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 119.85 0 119.95 0.51 ;
      END
   END g2_q78_8_

   PIN gt_93966_62_n_89
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 53.95 0.51 54.05 ;
      END
   END gt_93966_62_n_89

   PIN memread_edit_dist_a_ln268_unr124_a_21__4330189
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 95.15 183 95.25 ;
      END
   END memread_edit_dist_a_ln268_unr124_a_21__4330189

   PIN memread_edit_dist_g2_ln254_unr67_q_10_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 26.35 183 26.45 ;
      END
   END memread_edit_dist_g2_ln254_unr67_q_10_

   PIN memread_edit_dist_g2_ln254_unr67_q_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 176.65 0 176.75 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr67_q_1_

   PIN memread_edit_dist_g2_ln254_unr67_q_5_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 71.95 183 72.05 ;
      END
   END memread_edit_dist_g2_ln254_unr67_q_5_

   PIN memread_edit_dist_g2_ln254_unr68_q_10_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 92.65 0 92.75 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr68_q_10_

   PIN memread_edit_dist_g2_ln254_unr68_q_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 175.65 0 175.75 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr68_q_3_

   PIN memread_edit_dist_g2_ln254_unr69_q_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 35.75 183 35.85 ;
      END
   END memread_edit_dist_g2_ln254_unr69_q_4_

   PIN memread_edit_dist_g2_ln254_unr70_q_0_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 111.15 183 111.25 ;
      END
   END memread_edit_dist_g2_ln254_unr70_q_0_

   PIN memread_edit_dist_g2_ln254_unr70_q_10_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 126.65 0 126.75 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr70_q_10_

   PIN memread_edit_dist_g2_ln254_unr70_q_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 15.55 183 15.65 ;
      END
   END memread_edit_dist_g2_ln254_unr70_q_1_

   PIN memread_edit_dist_g2_ln254_unr70_q_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 8.75 183 8.85 ;
      END
   END memread_edit_dist_g2_ln254_unr70_q_3_

   PIN memread_edit_dist_g2_ln254_unr70_q_5_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 35.95 183 36.05 ;
      END
   END memread_edit_dist_g2_ln254_unr70_q_5_

   PIN memread_edit_dist_g2_ln254_unr70_q_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 93.15 183 93.25 ;
      END
   END memread_edit_dist_g2_ln254_unr70_q_7_

   PIN memread_edit_dist_g2_ln254_unr71_q_0_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 134.35 183 134.45 ;
      END
   END memread_edit_dist_g2_ln254_unr71_q_0_

   PIN memread_edit_dist_g2_ln254_unr71_q_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 8.95 183 9.05 ;
      END
   END memread_edit_dist_g2_ln254_unr71_q_1_

   PIN memread_edit_dist_g2_ln254_unr71_q_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 80.55 183 80.65 ;
      END
   END memread_edit_dist_g2_ln254_unr71_q_2_

   PIN memread_edit_dist_g2_ln254_unr71_q_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 170.55 183 170.65 ;
      END
   END memread_edit_dist_g2_ln254_unr71_q_3_

   PIN memread_edit_dist_g2_ln254_unr71_q_5_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 126.95 183 127.05 ;
      END
   END memread_edit_dist_g2_ln254_unr71_q_5_

   PIN memread_edit_dist_g2_ln254_unr71_q_6_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 44.15 183 44.25 ;
      END
   END memread_edit_dist_g2_ln254_unr71_q_6_

   PIN memread_edit_dist_g2_ln254_unr71_q_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 53.55 183 53.65 ;
      END
   END memread_edit_dist_g2_ln254_unr71_q_7_

   PIN memread_edit_dist_g2_ln254_unr72_q_0_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 125.15 183 125.25 ;
      END
   END memread_edit_dist_g2_ln254_unr72_q_0_

   PIN memread_edit_dist_g2_ln254_unr72_q_11_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 53.75 183 53.85 ;
      END
   END memread_edit_dist_g2_ln254_unr72_q_11_

   PIN memread_edit_dist_g2_ln254_unr72_q_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 165.05 0 165.15 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr72_q_1_

   PIN memread_edit_dist_g2_ln254_unr72_q_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 53.95 183 54.05 ;
      END
   END memread_edit_dist_g2_ln254_unr72_q_2_

   PIN memread_edit_dist_g2_ln254_unr72_q_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 170.75 183 170.85 ;
      END
   END memread_edit_dist_g2_ln254_unr72_q_3_

   PIN memread_edit_dist_g2_ln254_unr72_q_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 143.95 183 144.05 ;
      END
   END memread_edit_dist_g2_ln254_unr72_q_4_

   PIN memread_edit_dist_g2_ln254_unr72_q_5_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 179.55 183 179.65 ;
      END
   END memread_edit_dist_g2_ln254_unr72_q_5_

   PIN memread_edit_dist_g2_ln254_unr76_q_0_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 125.25 0 125.35 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr76_q_0_

   PIN memread_edit_dist_g2_ln254_unr76_q_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 136.65 0 136.75 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr76_q_1_

   PIN memread_edit_dist_g2_ln254_unr76_q_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 141.65 0 141.75 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr76_q_2_

   PIN memread_edit_dist_g2_ln254_unr76_q_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 155.45 0 155.55 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr76_q_3_

   PIN memread_edit_dist_g2_ln254_unr76_q_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 44.35 183 44.45 ;
      END
   END memread_edit_dist_g2_ln254_unr76_q_4_

   PIN memread_edit_dist_g2_ln254_unr76_q_5_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 178.95 183 179.05 ;
      END
   END memread_edit_dist_g2_ln254_unr76_q_5_

   PIN memread_edit_dist_g2_ln254_unr76_q_6_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 152.65 0 152.75 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr76_q_6_

   PIN memread_edit_dist_g2_ln254_unr76_q_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 9.15 183 9.25 ;
      END
   END memread_edit_dist_g2_ln254_unr76_q_7_

   PIN memread_edit_dist_g2_ln254_unr76_q_9_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 182.49 35.55 183 35.65 ;
      END
   END memread_edit_dist_g2_ln254_unr76_q_9_

   PIN memread_edit_dist_g2_ln254_unr77_q_0_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 123.05 0 123.15 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr77_q_0_

   PIN memread_edit_dist_g2_ln254_unr77_q_10_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 164.85 0 164.95 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr77_q_10_

   PIN memread_edit_dist_g2_ln254_unr77_q_11_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 135.45 0 135.55 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr77_q_11_

   PIN memread_edit_dist_g2_ln254_unr77_q_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 92.85 0 92.95 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr77_q_1_

   PIN memread_edit_dist_g2_ln254_unr77_q_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 128.85 0 128.95 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr77_q_2_

   PIN memread_edit_dist_g2_ln254_unr77_q_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 135.65 0 135.75 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr77_q_3_

   PIN memread_edit_dist_g2_ln254_unr77_q_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 119.85 0 119.95 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr77_q_4_

   PIN memread_edit_dist_g2_ln254_unr77_q_5_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 93.05 0 93.15 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr77_q_5_

   PIN memread_edit_dist_g2_ln254_unr77_q_6_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 111.05 0 111.15 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr77_q_6_

   PIN memread_edit_dist_g2_ln254_unr77_q_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 137.25 0 137.35 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr77_q_7_

   PIN memread_edit_dist_g2_ln254_unr77_q_8_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 144.65 0 144.75 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr77_q_8_

   PIN memread_edit_dist_g2_ln254_unr77_q_9_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 34.95 183 35.05 ;
      END
   END memread_edit_dist_g2_ln254_unr77_q_9_

   PIN mux_g_ln251_z_911__4472811
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 129.35 0.51 129.45 ;
      END
   END mux_g_ln251_z_911__4472811

   PIN mux_g_ln251_z_923__4472819
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 83.75 0.51 83.85 ;
      END
   END mux_g_ln251_z_923__4472819

   PIN mux_g_ln251_z_935__4472827
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 35.15 0.51 35.25 ;
      END
   END mux_g_ln251_z_935__4472827

   PIN mux_g_ln477_q_823_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 123.15 183 123.25 ;
      END
   END mux_g_ln477_q_823_

   PIN mux_g_ln477_q_931_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 137.85 0 137.95 0.51 ;
      END
   END mux_g_ln477_q_931_

   PIN n_1796
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 133.55 183 133.65 ;
      END
   END n_1796

   PIN n_1809
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 18.15 183 18.25 ;
      END
   END n_1809

   PIN n_2052
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 89.55 183 89.65 ;
      END
   END n_2052

   PIN n_2059
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 44.55 183 44.65 ;
      END
   END n_2059

   PIN n_2093
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 177.25 0 177.35 0.51 ;
      END
   END n_2093

   PIN n_2122
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 62.15 183 62.25 ;
      END
   END n_2122

   PIN n_21658
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 35.95 0.51 36.05 ;
      END
   END n_21658

   PIN n_23468
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 102.55 183 102.65 ;
      END
   END n_23468

   PIN n_23568
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 16.95 183 17.05 ;
      END
   END n_23568

   PIN n_23738
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 24.95 183 25.05 ;
      END
   END n_23738

   PIN n_2401
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 9.35 183 9.45 ;
      END
   END n_2401

   PIN n_2442
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 177.85 0 177.95 0.51 ;
      END
   END n_2442

   PIN n_24712
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 54.15 183 54.25 ;
      END
   END n_24712

   PIN n_25142
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 6.95 183 7.05 ;
      END
   END n_25142

   PIN n_25200
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 98.15 183 98.25 ;
      END
   END n_25200

   PIN n_2559
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 113.35 183 113.45 ;
      END
   END n_2559

   PIN n_2653
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 36.15 183 36.25 ;
      END
   END n_2653

   PIN n_27360
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 42.95 0.51 43.05 ;
      END
   END n_27360

   PIN n_29502
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 89.9 0.255 90.1 ;
      END
   END n_29502

   PIN n_29627
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 132.95 0.51 133.05 ;
      END
   END n_29627

   PIN n_29628
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 129.15 0.51 129.25 ;
      END
   END n_29628

   PIN n_29630
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 129.55 0.51 129.65 ;
      END
   END n_29630

   PIN n_29802
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 78.95 0.51 79.05 ;
      END
   END n_29802

   PIN n_29893
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 80.95 0.51 81.05 ;
      END
   END n_29893

   PIN n_29895
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 83.15 0.51 83.25 ;
      END
   END n_29895

   PIN n_30118
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 79.75 0.51 79.85 ;
      END
   END n_30118

   PIN n_30120
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 83.35 0.51 83.45 ;
      END
   END n_30120

   PIN n_30316
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 142.55 0.51 142.65 ;
      END
   END n_30316

   PIN n_30339
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 125.55 0.51 125.65 ;
      END
   END n_30339

   PIN n_30590
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 88.95 0.51 89.05 ;
      END
   END n_30590

   PIN n_30594
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 88.75 0.51 88.85 ;
      END
   END n_30594

   PIN n_30671
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 70.95 0.51 71.05 ;
      END
   END n_30671

   PIN n_30672
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 83.55 0.51 83.65 ;
      END
   END n_30672

   PIN n_30693
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 75.35 0.51 75.45 ;
      END
   END n_30693

   PIN n_30772
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 75.15 0.51 75.25 ;
      END
   END n_30772

   PIN n_30898
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 70.75 0.51 70.85 ;
      END
   END n_30898

   PIN n_3116
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 44.75 183 44.85 ;
      END
   END n_3116

   PIN n_31197
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 235.15 0.51 235.25 ;
      END
   END n_31197

   PIN n_31199
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 152.35 0.51 152.45 ;
      END
   END n_31199

   PIN n_31664
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 102.75 0.51 102.85 ;
      END
   END n_31664

   PIN n_31908
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 73.15 0.51 73.25 ;
      END
   END n_31908

   PIN n_3216
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 177.65 0 177.75 0.51 ;
      END
   END n_3216

   PIN n_32226
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 225.55 0.51 225.65 ;
      END
   END n_32226

   PIN n_32312
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 188.75 0.51 188.85 ;
      END
   END n_32312

   PIN n_32314
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 171.15 0.51 171.25 ;
      END
   END n_32314

   PIN n_32320
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 217.75 0.51 217.85 ;
      END
   END n_32320

   PIN n_32321
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 217.55 0.51 217.65 ;
      END
   END n_32321

   PIN n_32383
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 245.15 0.51 245.25 ;
      END
   END n_32383

   PIN n_32385
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 134.55 0.51 134.65 ;
      END
   END n_32385

   PIN n_33478
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 52.95 0.51 53.05 ;
      END
   END n_33478

   PIN n_33638
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 179.95 0.51 180.05 ;
      END
   END n_33638

   PIN n_34651
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 8.55 0.51 8.65 ;
      END
   END n_34651

   PIN n_34723
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 188.5 0.255 188.7 ;
      END
   END n_34723

   PIN n_35137
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 62.15 0.51 62.25 ;
      END
   END n_35137

   PIN n_35948
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 161.95 0.51 162.05 ;
      END
   END n_35948

   PIN n_35972
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 233.75 0.51 233.85 ;
      END
   END n_35972

   PIN n_35982
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 152.35 0.51 152.45 ;
      END
   END n_35982

   PIN n_36120
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 233.75 0.51 233.85 ;
      END
   END n_36120

   PIN n_36223
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 214.95 183 215.05 ;
      END
   END n_36223

   PIN n_36620
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 179.75 0.51 179.85 ;
      END
   END n_36620

   PIN n_36773
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 233.95 0.51 234.05 ;
      END
   END n_36773

   PIN n_36798
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 111.15 0.51 111.25 ;
      END
   END n_36798

   PIN n_36805
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 152.55 0.51 152.65 ;
      END
   END n_36805

   PIN n_36870
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 98.35 0.51 98.45 ;
      END
   END n_36870

   PIN n_39212
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 47.25 249.49 47.35 250 ;
      END
   END n_39212

   PIN n_39292
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 225.75 0.51 225.85 ;
      END
   END n_39292

   PIN n_39330
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 206.15 0.51 206.25 ;
      END
   END n_39330

   PIN n_46010
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 25.15 0.51 25.25 ;
      END
   END n_46010

   PIN n_46011
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 17.55 0.51 17.65 ;
      END
   END n_46011

   PIN n_49326
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 34.75 0.51 34.85 ;
      END
   END n_49326

   PIN n_51070
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 206.95 0.51 207.05 ;
      END
   END n_51070

   PIN n_51313
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 120.75 0.51 120.85 ;
      END
   END n_51313

   PIN n_51468
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 207.15 0.51 207.25 ;
      END
   END n_51468

   PIN n_52148
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 44.15 0.51 44.25 ;
      END
   END n_52148

   PIN n_57659
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 189.15 0.51 189.25 ;
      END
   END n_57659

   PIN n_57660
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 199.15 0.51 199.25 ;
      END
   END n_57660

   PIN n_58140
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 188.95 0.51 189.05 ;
      END
   END n_58140

   PIN n_58801
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 44.35 0.51 44.45 ;
      END
   END n_58801

   PIN n_60533
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 17.75 0.51 17.85 ;
      END
   END n_60533

   PIN n_61491
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 206.55 0.51 206.65 ;
      END
   END n_61491

   PIN n_61495
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 124.95 0.51 125.05 ;
      END
   END n_61495

   PIN n_61496
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 135.15 0.51 135.25 ;
      END
   END n_61496

   PIN n_62362
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 189.35 0.51 189.45 ;
      END
   END n_62362

   PIN n_62363
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 196.75 0.51 196.85 ;
      END
   END n_62363

   PIN n_64805
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 53.15 0.51 53.25 ;
      END
   END n_64805

   PIN n_65187
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 120.05 0 120.15 0.51 ;
      END
   END n_65187

   PIN n_65196
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 8.55 0.51 8.65 ;
      END
   END n_65196

   PIN n_67247
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 44.95 0.51 45.05 ;
      END
   END n_67247

   PIN n_8305
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 43.15 0.51 43.25 ;
      END
   END n_8305

   PIN n_8307
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 34.95 0.51 35.05 ;
      END
   END n_8307

   PIN ternarymux_ln49_0_unr72_z_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 225.95 0.51 226.05 ;
      END
   END ternarymux_ln49_0_unr72_z_2_

   PIN ternarymux_ln49_0_unr72_z_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 226.15 0.51 226.25 ;
      END
   END ternarymux_ln49_0_unr72_z_3_

   PIN ternarymux_ln49_0_unr76_z_10__4331222
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 187.75 0.51 187.85 ;
      END
   END ternarymux_ln49_0_unr76_z_10__4331222

   PIN ternarymux_ln49_0_unr76_z_8__4331230
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 180.35 0.51 180.45 ;
      END
   END ternarymux_ln49_0_unr76_z_8__4331230

   PIN ternarymux_ln49_0_unr78_z_0_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 8.75 0.51 8.85 ;
      END
   END ternarymux_ln49_0_unr78_z_0_

   PIN ternarymux_ln49_0_unr78_z_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 17.95 0.51 18.05 ;
      END
   END ternarymux_ln49_0_unr78_z_1_

   PIN ternarymux_ln49_0_unr78_z_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 14.95 0.51 15.05 ;
      END
   END ternarymux_ln49_0_unr78_z_2_

   PIN ternarymux_ln49_0_unr78_z_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 25.35 0.51 25.45 ;
      END
   END ternarymux_ln49_0_unr78_z_3_

   PIN ternarymux_ln49_0_unr78_z_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 26.35 0.51 26.45 ;
      END
   END ternarymux_ln49_0_unr78_z_4_

   PIN ternarymux_ln49_0_unr78_z_5_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 26.15 0.51 26.25 ;
      END
   END ternarymux_ln49_0_unr78_z_5_

   PIN ternarymux_ln49_0_unr78_z_6_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 63.35 0.51 63.45 ;
      END
   END ternarymux_ln49_0_unr78_z_6_

   PIN ternarymux_ln49_0_unr78_z_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 36.15 0.51 36.25 ;
      END
   END ternarymux_ln49_0_unr78_z_7_

   PIN ternarymux_ln49_0_unr78_z_8__4331262
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 36.35 0.51 36.45 ;
      END
   END ternarymux_ln49_0_unr78_z_8__4331262

   PIN ternarymux_ln49_0_unr78_z_9__4331258
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 53.35 0.51 53.45 ;
      END
   END ternarymux_ln49_0_unr78_z_9__4331258

   PIN ternarymux_ln49_5_unr72_z_0_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 197.15 0.51 197.25 ;
      END
   END ternarymux_ln49_5_unr72_z_0_

   PIN ternarymux_ln49_6_unr75_z_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 205.35 0.51 205.45 ;
      END
   END ternarymux_ln49_6_unr75_z_2_

   PIN ternarymux_ln49_6_unr78_z_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 35.35 0.51 35.45 ;
      END
   END ternarymux_ln49_6_unr78_z_12_

   PIN ternarymux_ln49_unr77_z_8_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 71.15 0.51 71.25 ;
      END
   END ternarymux_ln49_unr77_z_8_

   PIN FE_OCPN56260_ctrlor_ln251_z_0__4471604_bar
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 25.15 183 25.25 ;
      END
   END FE_OCPN56260_ctrlor_ln251_z_0__4471604_bar

   PIN FE_OCPN57864_n_93
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 242.55 183 242.65 ;
      END
   END FE_OCPN57864_n_93

   PIN FE_OCPN62021_FE_OFN50813_n_67216
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 83.15 183 83.25 ;
      END
   END FE_OCPN62021_FE_OFN50813_n_67216

   PIN FE_OCPN62025_FE_OFN50813_n_67216
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 45.35 183 45.45 ;
      END
   END FE_OCPN62025_FE_OFN50813_n_67216

   PIN FE_OCPN62349_n_65199
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 133.95 183 134.05 ;
      END
   END FE_OCPN62349_n_65199

   PIN FE_OCPN62379_FE_OFN47982_n_23035
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 45.15 183 45.25 ;
      END
   END FE_OCPN62379_FE_OFN47982_n_23035

   PIN FE_OCPN62552_FE_OFN47982_n_23035
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 110.85 0 110.95 0.51 ;
      END
   END FE_OCPN62552_FE_OFN47982_n_23035

   PIN FE_OCPN62858_n_33487_bar
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 182.49 26.35 183 26.45 ;
      END
   END FE_OCPN62858_n_33487_bar

   PIN FE_OCPN76859_FE_OFN48337_n_31639
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 92.85 249.49 92.95 250 ;
      END
   END FE_OCPN76859_FE_OFN48337_n_31639

   PIN FE_OCPN76904_n_58046
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 143.15 183 143.25 ;
      END
   END FE_OCPN76904_n_58046

   PIN FE_OCPN77874_FE_OFN48363_n_31641
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 8.85 249.49 8.95 250 ;
      END
   END FE_OCPN77874_FE_OFN48363_n_31641

   PIN FE_OFN28531_n_36394
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 119.85 249.49 119.95 250 ;
      END
   END FE_OFN28531_n_36394

   PIN FE_OFN28589_n_36353
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 138.65 249.49 138.75 250 ;
      END
   END FE_OFN28589_n_36353

   PIN FE_OFN28736_n_59342
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 43.55 183 43.65 ;
      END
   END FE_OFN28736_n_59342

   PIN FE_OFN30021_n_36839
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 227.15 183 227.25 ;
      END
   END FE_OFN30021_n_36839

   PIN FE_OFN30124_n_36029
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 116.55 0.51 116.65 ;
      END
   END FE_OFN30124_n_36029

   PIN FE_OFN30126_n_36012
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 115.75 0.51 115.85 ;
      END
   END FE_OFN30126_n_36012

   PIN FE_OFN30134_n_35994
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 118.95 0.51 119.05 ;
      END
   END FE_OFN30134_n_35994

   PIN FE_OFN30141_n_34781
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.745 63.5 183 63.7 ;
      END
   END FE_OFN30141_n_34781

   PIN FE_OFN30157_n_36428
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 23.45 0 23.55 0.51 ;
      END
   END FE_OFN30157_n_36428

   PIN FE_OFN30217_n_36501
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 24.35 183 24.45 ;
      END
   END FE_OFN30217_n_36501

   PIN FE_OFN30294_n_36448
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 129.05 0 129.15 0.51 ;
      END
   END FE_OFN30294_n_36448

   PIN FE_OFN30298_n_36432
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 162.05 0 162.15 0.51 ;
      END
   END FE_OFN30298_n_36432

   PIN FE_OFN30300_n_36379
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 155.25 0 155.35 0.51 ;
      END
   END FE_OFN30300_n_36379

   PIN FE_OFN30384_n_34771
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 152.35 183 152.45 ;
      END
   END FE_OFN30384_n_34771

   PIN FE_OFN30485_n_34770
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 160.95 183 161.05 ;
      END
   END FE_OFN30485_n_34770

   PIN FE_OFN30528_n_36408
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 35.55 183 35.65 ;
      END
   END FE_OFN30528_n_36408

   PIN FE_OFN30575_n_36929
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 101.85 0 101.95 0.51 ;
      END
   END FE_OFN30575_n_36929

   PIN FE_OFN30593_n_36874
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 43.95 183 44.05 ;
      END
   END FE_OFN30593_n_36874

   PIN FE_OFN30767_n_34754
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.745 64.9 183 65.1 ;
      END
   END FE_OFN30767_n_34754

   PIN FE_OFN30784_n_34754
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 119.65 249.49 119.75 250 ;
      END
   END FE_OFN30784_n_34754

   PIN FE_OFN30785_n_34754
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.745 14.9 183 15.1 ;
      END
   END FE_OFN30785_n_34754

   PIN FE_OFN30819_n_36961
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 83.85 0 83.95 0.51 ;
      END
   END FE_OFN30819_n_36961

   PIN FE_OFN30851_n_36114
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 49.65 0 49.75 0.51 ;
      END
   END FE_OFN30851_n_36114

   PIN FE_OFN30860_n_34779
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 53.15 183 53.25 ;
      END
   END FE_OFN30860_n_34779

   PIN FE_OFN32392_n_51426
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 55.35 183 55.45 ;
      END
   END FE_OFN32392_n_51426

   PIN FE_OFN32394_n_46215
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 70.95 183 71.05 ;
      END
   END FE_OFN32394_n_46215

   PIN FE_OFN32422_n_62230
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 128.5 0.255 128.7 ;
      END
   END FE_OFN32422_n_62230

   PIN FE_OFN32426_g2_bridge200_rtl_ce_en_3754908
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 133.75 0.51 133.85 ;
      END
   END FE_OFN32426_g2_bridge200_rtl_ce_en_3754908

   PIN FE_OFN34918_n_51730
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 182.49 172.15 183 172.25 ;
      END
   END FE_OFN34918_n_51730

   PIN FE_OFN34931_n_51721
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 118.95 183 119.05 ;
      END
   END FE_OFN34931_n_51721

   PIN FE_OFN34933_memwrite_edit_dist_g2_ln280_unr78_en_0__4469092
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 63.15 0.51 63.25 ;
      END
   END FE_OFN34933_memwrite_edit_dist_g2_ln280_unr78_en_0__4469092

   PIN FE_OFN35565_n_48865
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 122.95 183 123.05 ;
      END
   END FE_OFN35565_n_48865

   PIN FE_OFN41927_n_230
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 174.25 249.49 174.35 250 ;
      END
   END FE_OFN41927_n_230

   PIN FE_OFN42046_n_232
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 17.95 183 18.05 ;
      END
   END FE_OFN42046_n_232

   PIN FE_OFN42135_n_222
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 168.85 0 168.95 0.51 ;
      END
   END FE_OFN42135_n_222

   PIN FE_OFN42586_n_29
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 152.65 0 152.75 0.51 ;
      END
   END FE_OFN42586_n_29

   PIN FE_OFN42590_n_29
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 66.05 0 66.15 0.51 ;
      END
   END FE_OFN42590_n_29

   PIN FE_OFN42976_n_35330
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 169.75 183 169.85 ;
      END
   END FE_OFN42976_n_35330

   PIN FE_OFN43000_n_35325
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 164.95 183 165.05 ;
      END
   END FE_OFN43000_n_35325

   PIN FE_OFN43003_n_35325
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 172.95 183 173.05 ;
      END
   END FE_OFN43003_n_35325

   PIN FE_OFN43167_n_35301
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 104.95 183 105.05 ;
      END
   END FE_OFN43167_n_35301

   PIN FE_OFN43216_n_35283
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 176.45 0 176.55 0.51 ;
      END
   END FE_OFN43216_n_35283

   PIN FE_OFN43225_n_35284
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 62.55 183 62.65 ;
      END
   END FE_OFN43225_n_35284

   PIN FE_OFN43271_n_35276
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.745 63.1 183 63.3 ;
      END
   END FE_OFN43271_n_35276

   PIN FE_OFN43925_mux_g_ln477_q_821_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 173.15 183 173.25 ;
      END
   END FE_OFN43925_mux_g_ln477_q_821_

   PIN FE_OFN43998_n_35331
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 55.15 183 55.25 ;
      END
   END FE_OFN43998_n_35331

   PIN FE_OFN46306_n_35331
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 224.95 183 225.05 ;
      END
   END FE_OFN46306_n_35331

   PIN FE_OFN47138_n_23039
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 151.05 0 151.15 0.51 ;
      END
   END FE_OFN47138_n_23039

   PIN FE_OFN47317_n_35285
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 133.35 183 133.45 ;
      END
   END FE_OFN47317_n_35285

   PIN FE_OFN47849_n_23045
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 233.55 183 233.65 ;
      END
   END FE_OFN47849_n_23045

   PIN FE_OFN48291_n_31625
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 161.45 249.49 161.55 250 ;
      END
   END FE_OFN48291_n_31625

   PIN FE_OFN48300_n_31625
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 101.85 249.49 101.95 250 ;
      END
   END FE_OFN48300_n_31625

   PIN FE_OFN48307_n_31634
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 223.75 0.51 223.85 ;
      END
   END FE_OFN48307_n_31634

   PIN FE_OFN48343_n_31639
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 10.45 249.49 10.55 250 ;
      END
   END FE_OFN48343_n_31639

   PIN FE_OFN48353_n_31638
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 83.85 249.49 83.95 250 ;
      END
   END FE_OFN48353_n_31638

   PIN FE_OFN48358_n_31637
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 140.95 0.51 141.05 ;
      END
   END FE_OFN48358_n_31637

   PIN FE_OFN48629_n_31308
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 122.85 249.49 122.95 250 ;
      END
   END FE_OFN48629_n_31308

   PIN FE_OFN48687_n_59052
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 178.25 249.49 178.35 250 ;
      END
   END FE_OFN48687_n_59052

   PIN FE_OFN49699_n_87
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 226.95 183 227.05 ;
      END
   END FE_OFN49699_n_87

   PIN FE_OFN49700_n_87
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 143.55 183 143.65 ;
      END
   END FE_OFN49700_n_87

   PIN FE_OFN50548_lt_ln49_6_unr78_z
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 55.3 0.255 55.5 ;
      END
   END FE_OFN50548_lt_ln49_6_unr78_z

   PIN FE_OFN50882_n_35300
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 130.45 0 130.55 0.51 ;
      END
   END FE_OFN50882_n_35300

   PIN FE_OFN51004_n_23330
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 43.75 183 43.85 ;
      END
   END FE_OFN51004_n_23330

   PIN FE_OFN53892_n_71
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 165.4 0 165.6 0.255 ;
      END
   END FE_OFN53892_n_71

   PIN FE_OFN55363_n_59053
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 92.65 249.49 92.75 250 ;
      END
   END FE_OFN55363_n_59053

   PIN FE_OFN64277_n_57747
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 245.35 183 245.45 ;
      END
   END FE_OFN64277_n_57747

   PIN FE_OFN70360_n_36808
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 155.45 249.49 155.55 250 ;
      END
   END FE_OFN70360_n_36808

   PIN FE_OFN70362_n_36328
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 188.55 0.51 188.65 ;
      END
   END FE_OFN70362_n_36328

   PIN FE_OFN71104_memwrite_edit_dist_g2_ln280_unr73_en_0__4469519
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 170.35 183 170.45 ;
      END
   END FE_OFN71104_memwrite_edit_dist_g2_ln280_unr73_en_0__4469519

   PIN FE_OFN71829_n_53368
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 182.49 233.55 183 233.65 ;
      END
   END FE_OFN71829_n_53368

   PIN FE_OFN73300_n_57
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 165.65 0 165.75 0.51 ;
      END
   END FE_OFN73300_n_57

   PIN FE_OFN73345_n_41
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 215.15 183 215.25 ;
      END
   END FE_OFN73345_n_41

   PIN FE_OFN74070_n_59125
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 101.65 249.49 101.75 250 ;
      END
   END FE_OFN74070_n_59125

   PIN FE_OFN74248_n_223
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 102.75 183 102.85 ;
      END
   END FE_OFN74248_n_223

   PIN FE_OFN74309_n_61
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 155.85 0 155.95 0.51 ;
      END
   END FE_OFN74309_n_61

   PIN FE_OFN74356_n_86
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 83.65 249.49 83.75 250 ;
      END
   END FE_OFN74356_n_86

   PIN FE_OFN74575_n_93
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 178.25 249.49 178.35 250 ;
      END
   END FE_OFN74575_n_93

   PIN FE_OFN74579_n_79
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 176.25 249.49 176.35 250 ;
      END
   END FE_OFN74579_n_79

   PIN FE_OFN74596_n_856
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 143.65 0 143.75 0.51 ;
      END
   END FE_OFN74596_n_856

   PIN FE_OFN74836_n_34785
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 230.95 183 231.05 ;
      END
   END FE_OFN74836_n_34785

   PIN FE_OFN75116_n_34732
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 132.95 183 133.05 ;
      END
   END FE_OFN75116_n_34732

   PIN FE_OFN75232_n_35287
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 142.95 183 143.05 ;
      END
   END FE_OFN75232_n_35287

   PIN FE_OFN75274_n_35301
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 154.45 249.49 154.55 250 ;
      END
   END FE_OFN75274_n_35301

   PIN FE_OFN83829_n_36361
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 122.05 249.49 122.15 250 ;
      END
   END FE_OFN83829_n_36361

   PIN FE_OFN84036_n_7936
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 26.95 183 27.05 ;
      END
   END FE_OFN84036_n_7936

   PIN FE_OFN85095_n_30
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 110.85 249.49 110.95 250 ;
      END
   END FE_OFN85095_n_30

   PIN FE_OFN85116_n_15
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 177.05 0 177.15 0.51 ;
      END
   END FE_OFN85116_n_15

   PIN FE_OFN85912_ternarymux_ln49_0_unr75_z_1_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 198.95 0.51 199.05 ;
      END
   END FE_OFN85912_ternarymux_ln49_0_unr75_z_1_

   PIN FE_OFN86076_n_59125
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 38.25 249.49 38.35 250 ;
      END
   END FE_OFN86076_n_59125

   PIN FE_OFN86112_mux_g_ln251_z_933__4472823
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 32.95 183 33.05 ;
      END
   END FE_OFN86112_mux_g_ln251_z_933__4472823

   PIN FE_OFN86557_n_36439
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 101.65 0 101.75 0.51 ;
      END
   END FE_OFN86557_n_36439

   PIN FE_OFN86620_n_35995
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 137.65 0 137.75 0.51 ;
      END
   END FE_OFN86620_n_35995

   PIN FE_OFN86638_n_36832
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 110.65 0 110.75 0.51 ;
      END
   END FE_OFN86638_n_36832

   PIN FE_OFN86665_n_36390
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 71.75 183 71.85 ;
      END
   END FE_OFN86665_n_36390

   PIN FE_OFN86720_n_36698
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 148.95 183 149.05 ;
      END
   END FE_OFN86720_n_36698

   PIN FE_OFN86741_n_37010
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 80.35 183 80.45 ;
      END
   END FE_OFN86741_n_37010

   PIN FE_OFN86745_n_36401
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 134.15 183 134.25 ;
      END
   END FE_OFN86745_n_36401

   PIN FE_OFN86746_n_36399
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 150.65 0 150.75 0.51 ;
      END
   END FE_OFN86746_n_36399

   PIN FE_OFN86876_n_37029
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 182.49 8.55 183 8.65 ;
      END
   END FE_OFN86876_n_37029

   PIN FE_OFN86890_n_37046
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 131.15 183 131.25 ;
      END
   END FE_OFN86890_n_37046

   PIN FE_OFN86897_n_36447
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 71.55 183 71.65 ;
      END
   END FE_OFN86897_n_36447

   PIN FE_OFN87024_n_34784
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 110.95 183 111.05 ;
      END
   END FE_OFN87024_n_34784

   PIN FE_OFN88035_mux_g_ln477_q_848_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 53.35 183 53.45 ;
      END
   END FE_OFN88035_mux_g_ln477_q_848_

   PIN FE_OFN88305_n_65239
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 216.95 183 217.05 ;
      END
   END FE_OFN88305_n_65239

   PIN FE_OFN88312_n_65240
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 133.75 183 133.85 ;
      END
   END FE_OFN88312_n_65240

   PIN FE_OFN88350_n_26962
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 215.75 0.51 215.85 ;
      END
   END FE_OFN88350_n_26962

   PIN FE_OFN89020_n_31626
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 205.75 0.51 205.85 ;
      END
   END FE_OFN89020_n_31626

   PIN FE_OFN89196_FE_OCPN63783_FE_OFN48830_n_31626
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 56.65 249.49 56.75 250 ;
      END
   END FE_OFN89196_FE_OCPN63783_FE_OFN48830_n_31626

   PIN FE_OFN90979_n_22947
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 44.95 183 45.05 ;
      END
   END FE_OFN90979_n_22947

   PIN FE_OFN95872_n_58716
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 71.35 183 71.45 ;
      END
   END FE_OFN95872_n_58716

   PIN FE_OFN98488_n_35997
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 107.55 183 107.65 ;
      END
   END FE_OFN98488_n_35997

   PIN FE_OFN98505_n_36246
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 165.85 0 165.95 0.51 ;
      END
   END FE_OFN98505_n_36246

   PIN FE_OFN98507_n_36073
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 68.95 183 69.05 ;
      END
   END FE_OFN98507_n_36073

   PIN FE_OFN98899_n_35297
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 169.05 249.49 169.15 250 ;
      END
   END FE_OFN98899_n_35297

   PIN FE_RN_2506_0
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 157.35 0.51 157.45 ;
      END
   END FE_RN_2506_0

   PIN FE_RN_3497_0
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 205.95 0.51 206.05 ;
      END
   END FE_RN_3497_0

   PIN FE_RN_4443_0
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 179.55 0.51 179.65 ;
      END
   END FE_RN_4443_0

   PIN FE_RN_4457_0
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 134.75 0.51 134.85 ;
      END
   END FE_RN_4457_0

   PIN a_in_104_3
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 44.55 0.51 44.65 ;
      END
   END a_in_104_3

   PIN a_in_71_3
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 89.55 0.51 89.65 ;
      END
   END a_in_71_3

   PIN a_in_73_3
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 98.55 0.51 98.65 ;
      END
   END a_in_73_3

   PIN a_in_78_0
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 46.15 0.51 46.25 ;
      END
   END a_in_78_0

   PIN a_in_81_2
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 102.15 0.51 102.25 ;
      END
   END a_in_81_2

   PIN a_in_87_3
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 80.55 0.51 80.65 ;
      END
   END a_in_87_3

   PIN add_85528_72_n_1794471
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 113.15 0.51 113.25 ;
      END
   END add_85528_72_n_1794471

   PIN add_85528_72_n_4327661
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 116.35 0.51 116.45 ;
      END
   END add_85528_72_n_4327661

   PIN add_ln174_1_unr75_z_8__2227682
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 151.75 0.51 151.85 ;
      END
   END add_ln174_1_unr75_z_8__2227682

   PIN b_in_2_3
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 155.65 249.49 155.75 250 ;
      END
   END b_in_2_3

   PIN g2_q69_10_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 98.95 0.51 99.05 ;
      END
   END g2_q69_10_

   PIN g2_q69_1__4327571
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 97.75 0.51 97.85 ;
      END
   END g2_q69_1__4327571

   PIN g2_q69_2__4327573
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 62.35 0.51 62.45 ;
      END
   END g2_q69_2__4327573

   PIN g2_q69_3__4327574
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 106.95 0.51 107.05 ;
      END
   END g2_q69_3__4327574

   PIN g2_q69_5__4327578
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 98.75 0.51 98.85 ;
      END
   END g2_q69_5__4327578

   PIN g2_q69_7__4327567
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 116.55 0.51 116.65 ;
      END
   END g2_q69_7__4327567

   PIN g2_q70_10_
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 24.95 0.51 25.05 ;
      END
   END g2_q70_10_

   PIN g2_q70_11_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 161.15 0.51 161.25 ;
      END
   END g2_q70_11_

   PIN g2_q70_3__4327605
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 115.35 0.51 115.45 ;
      END
   END g2_q70_3__4327605

   PIN g2_q70_5__4327609
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 124.75 0.51 124.85 ;
      END
   END g2_q70_5__4327609

   PIN g2_q70_8_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 124.55 0.51 124.65 ;
      END
   END g2_q70_8_

   PIN g2_q71_4__4327638
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 152.55 0.51 152.65 ;
      END
   END g2_q71_4__4327638

   PIN g2_q71_8_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 142.75 0.51 142.85 ;
      END
   END g2_q71_8_

   PIN g2_q72_10_
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 32.95 0.51 33.05 ;
      END
   END g2_q72_10_

   PIN g2_q72_2__4327665
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 112.95 0.51 113.05 ;
      END
   END g2_q72_2__4327665

   PIN g2_q72_3__4327666
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 114.95 0.51 115.05 ;
      END
   END g2_q72_3__4327666

   PIN g2_q72_5__4327670
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 93.15 0.51 93.25 ;
      END
   END g2_q72_5__4327670

   PIN g2_q72_6__4327658
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 125.55 0.51 125.65 ;
      END
   END g2_q72_6__4327658

   PIN g2_q72_7__4327659
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 92.95 0.51 93.05 ;
      END
   END g2_q72_7__4327659

   PIN g2_q73_11_
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 134.15 0.51 134.25 ;
      END
   END g2_q73_11_

   PIN g2_q73_3__4327696
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 245.35 0.51 245.45 ;
      END
   END g2_q73_3__4327696

   PIN g2_q73_5__4327700
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 160.75 0.51 160.85 ;
      END
   END g2_q73_5__4327700

   PIN g2_q73_6__4327688
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 125.35 0.51 125.45 ;
      END
   END g2_q73_6__4327688

   PIN g2_q73_7__4327689
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 188.35 0.51 188.45 ;
      END
   END g2_q73_7__4327689

   PIN g2_q74_11_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 234.95 0.51 235.05 ;
      END
   END g2_q74_11_

   PIN g2_q74_4__4327730
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 234.95 0.51 235.05 ;
      END
   END g2_q74_4__4327730

   PIN g2_q74_5__4327731
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 228.15 0.51 228.25 ;
      END
   END g2_q74_5__4327731

   PIN g2_q77_2__4327816
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 102.65 249.49 102.75 250 ;
      END
   END g2_q77_2__4327816

   PIN gt_93958_62_n_148_bar
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 179.55 0.51 179.65 ;
      END
   END gt_93958_62_n_148_bar

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 154.8 0 155 0.255 ;
      END
   END ispd_clk

   PIN memread_edit_dist_a_ln268_unr124_a_9__4329837
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 97.95 183 98.05 ;
      END
   END memread_edit_dist_a_ln268_unr124_a_9__4329837

   PIN memread_edit_dist_g2_ln254_unr66_q_11_
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 107.35 0.51 107.45 ;
      END
   END memread_edit_dist_g2_ln254_unr66_q_11_

   PIN memread_edit_dist_g2_ln254_unr67_q_6_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 137.45 0 137.55 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr67_q_6_

   PIN memread_edit_dist_g2_ln254_unr68_q_0_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 143.15 0.51 143.25 ;
      END
   END memread_edit_dist_g2_ln254_unr68_q_0_

   PIN memread_edit_dist_g2_ln254_unr68_q_4_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 134.95 0.51 135.05 ;
      END
   END memread_edit_dist_g2_ln254_unr68_q_4_

   PIN memread_edit_dist_g2_ln254_unr68_q_7_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 152.95 0.51 153.05 ;
      END
   END memread_edit_dist_g2_ln254_unr68_q_7_

   PIN memread_edit_dist_g2_ln254_unr69_q_10_
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 110.95 0.51 111.05 ;
      END
   END memread_edit_dist_g2_ln254_unr69_q_10_

   PIN memread_edit_dist_g2_ln254_unr69_q_3_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 150.85 0 150.95 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr69_q_3_

   PIN memread_edit_dist_g2_ln254_unr69_q_6_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 146.65 0 146.75 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr69_q_6_

   PIN memread_edit_dist_g2_ln254_unr69_q_7_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 164.85 0 164.95 0.51 ;
      END
   END memread_edit_dist_g2_ln254_unr69_q_7_

   PIN memread_edit_dist_g2_ln254_unr70_q_11_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 61.15 183 61.25 ;
      END
   END memread_edit_dist_g2_ln254_unr70_q_11_

   PIN memread_edit_dist_g2_ln254_unr70_q_8_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 62.95 0.51 63.05 ;
      END
   END memread_edit_dist_g2_ln254_unr70_q_8_

   PIN memwrite_edit_dist_g2_ln280_unr75_en_0__4469773
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 215.55 0.51 215.65 ;
      END
   END memwrite_edit_dist_g2_ln280_unr75_en_0__4469773

   PIN memwrite_edit_dist_g2_ln280_unr76_en_0__4469257
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 138.75 0.51 138.85 ;
      END
   END memwrite_edit_dist_g2_ln280_unr76_en_0__4469257

   PIN mux_g_ln477_q_11_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 155.05 249.49 155.15 250 ;
      END
   END mux_g_ln477_q_11_

   PIN mux_g_ln477_q_520_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 120.75 183 120.85 ;
      END
   END mux_g_ln477_q_520_

   PIN mux_g_ln477_q_799_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 107.15 183 107.25 ;
      END
   END mux_g_ln477_q_799_

   PIN mux_g_ln477_q_803_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 61.95 183 62.05 ;
      END
   END mux_g_ln477_q_803_

   PIN mux_g_ln477_q_806_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 166.05 0 166.15 0.51 ;
      END
   END mux_g_ln477_q_806_

   PIN mux_g_ln477_q_810_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 35.35 183 35.45 ;
      END
   END mux_g_ln477_q_810_

   PIN mux_g_ln477_q_811_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 61.75 183 61.85 ;
      END
   END mux_g_ln477_q_811_

   PIN mux_g_ln477_q_814_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 26.15 183 26.25 ;
      END
   END mux_g_ln477_q_814_

   PIN mux_g_ln477_q_815_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 61.55 183 61.65 ;
      END
   END mux_g_ln477_q_815_

   PIN mux_g_ln477_q_816_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 174.65 0 174.75 0.51 ;
      END
   END mux_g_ln477_q_816_

   PIN mux_g_ln477_q_818_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 161.15 183 161.25 ;
      END
   END mux_g_ln477_q_818_

   PIN mux_g_ln477_q_820_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 165.45 0 165.55 0.51 ;
      END
   END mux_g_ln477_q_820_

   PIN mux_g_ln477_q_827_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 25.95 183 26.05 ;
      END
   END mux_g_ln477_q_827_

   PIN mux_g_ln477_q_831_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 155.65 0 155.75 0.51 ;
      END
   END mux_g_ln477_q_831_

   PIN mux_g_ln477_q_834_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 25.75 183 25.85 ;
      END
   END mux_g_ln477_q_834_

   PIN mux_g_ln477_q_835_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 113.15 183 113.25 ;
      END
   END mux_g_ln477_q_835_

   PIN mux_g_ln477_q_836_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 82.95 183 83.05 ;
      END
   END mux_g_ln477_q_836_

   PIN mux_g_ln477_q_841_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 177.65 0 177.75 0.51 ;
      END
   END mux_g_ln477_q_841_

   PIN mux_g_ln477_q_846_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 92.95 183 93.05 ;
      END
   END mux_g_ln477_q_846_

   PIN mux_g_ln477_q_851_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 17.75 183 17.85 ;
      END
   END mux_g_ln477_q_851_

   PIN n_21259
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 130.95 183 131.05 ;
      END
   END n_21259

   PIN n_21278
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 121.35 183 121.45 ;
      END
   END n_21278

   PIN n_21287
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 208.95 183 209.05 ;
      END
   END n_21287

   PIN n_23142
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 94.95 183 95.05 ;
      END
   END n_23142

   PIN n_23298
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 108.95 0.51 109.05 ;
      END
   END n_23298

   PIN n_23337
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 100.95 0.51 101.05 ;
      END
   END n_23337

   PIN n_23348
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 94.65 0 94.75 0.51 ;
      END
   END n_23348

   PIN n_26820
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 215.95 0.51 216.05 ;
      END
   END n_26820

   PIN n_27167
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 217.35 0.51 217.45 ;
      END
   END n_27167

   PIN n_27169
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 197.35 0.51 197.45 ;
      END
   END n_27169

   PIN n_27172
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 244.95 0.51 245.05 ;
      END
   END n_27172

   PIN n_27478
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 214.9 0.255 215.1 ;
      END
   END n_27478

   PIN n_28223
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 206.35 0.51 206.45 ;
      END
   END n_28223

   PIN n_28405
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 204.9 0.255 205.1 ;
      END
   END n_28405

   PIN n_28469
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 217.15 0.51 217.25 ;
      END
   END n_28469

   PIN n_28821
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 155.25 0 155.35 0.51 ;
      END
   END n_28821

   PIN n_28879
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 153.25 0 153.35 0.51 ;
      END
   END n_28879

   PIN n_29799
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 128.95 0.51 129.05 ;
      END
   END n_29799

   PIN n_30353
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 141.5 0.255 141.7 ;
      END
   END n_30353

   PIN n_3063
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 43.75 0.51 43.85 ;
      END
   END n_3063

   PIN n_30960
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 92.95 0.51 93.05 ;
      END
   END n_30960

   PIN n_30965
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 91.15 0.51 91.25 ;
      END
   END n_30965

   PIN n_31888
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 157.55 0.51 157.65 ;
      END
   END n_31888

   PIN n_32070
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 109.35 0.51 109.45 ;
      END
   END n_32070

   PIN n_32511
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 179.35 0.51 179.45 ;
      END
   END n_32511

   PIN n_33240
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 156.75 0.51 156.85 ;
      END
   END n_33240

   PIN n_33245
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 55.75 0.51 55.85 ;
      END
   END n_33245

   PIN n_33384
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 160.95 0.51 161.05 ;
      END
   END n_33384

   PIN n_33386
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 169.95 0.51 170.05 ;
      END
   END n_33386

   PIN n_33467_bar
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 25.55 183 25.65 ;
      END
   END n_33467_bar

   PIN n_33556
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 186.95 0.51 187.05 ;
      END
   END n_33556

   PIN n_33599
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 187.15 0.51 187.25 ;
      END
   END n_33599

   PIN n_33639
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 154.95 0.51 155.05 ;
      END
   END n_33639

   PIN n_3370
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 114.95 183 115.05 ;
      END
   END n_3370

   PIN n_34235
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 169.75 0.51 169.85 ;
      END
   END n_34235

   PIN n_34404
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 54.9 0.255 55.1 ;
      END
   END n_34404

   PIN n_34535
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 195.75 0.51 195.85 ;
      END
   END n_34535

   PIN n_35331
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 52.95 183 53.05 ;
      END
   END n_35331

   PIN n_35936
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 165.25 0 165.35 0.51 ;
      END
   END n_35936

   PIN n_35978
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 71.15 183 71.25 ;
      END
   END n_35978

   PIN n_35984
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 172.45 0 172.55 0.51 ;
      END
   END n_35984

   PIN n_36005
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 170.15 183 170.25 ;
      END
   END n_36005

   PIN n_36014
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 17.55 183 17.65 ;
      END
   END n_36014

   PIN n_36015
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 100.95 183 101.05 ;
      END
   END n_36015

   PIN n_36035
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 52.75 183 52.85 ;
      END
   END n_36035

   PIN n_36060
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 80.15 183 80.25 ;
      END
   END n_36060

   PIN n_36062
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 35.15 183 35.25 ;
      END
   END n_36062

   PIN n_36086
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 70.75 183 70.85 ;
      END
   END n_36086

   PIN n_36113
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 72.05 0 72.15 0.51 ;
      END
   END n_36113

   PIN n_36221
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 155.65 0 155.75 0.51 ;
      END
   END n_36221

   PIN n_36250
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 182.49 52.95 183 53.05 ;
      END
   END n_36250

   PIN n_36339
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 182.49 26.55 183 26.65 ;
      END
   END n_36339

   PIN n_36355
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 96.45 249.49 96.55 250 ;
      END
   END n_36355

   PIN n_36486
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 155.45 0 155.55 0.51 ;
      END
   END n_36486

   PIN n_36520
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 182.49 18.15 183 18.25 ;
      END
   END n_36520

   PIN n_36547
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 10.25 0 10.35 0.51 ;
      END
   END n_36547

   PIN n_36563
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 115.95 183 116.05 ;
      END
   END n_36563

   PIN n_36622
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 34.75 183 34.85 ;
      END
   END n_36622

   PIN n_36733
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 8.55 183 8.65 ;
      END
   END n_36733

   PIN n_36748
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 42.95 183 43.05 ;
      END
   END n_36748

   PIN n_36785
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 112.95 183 113.05 ;
      END
   END n_36785

   PIN n_36787
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 61.35 183 61.45 ;
      END
   END n_36787

   PIN n_36803
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 158.45 0 158.55 0.51 ;
      END
   END n_36803

   PIN n_36899
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 70.55 183 70.65 ;
      END
   END n_36899

   PIN n_36922
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 52.55 183 52.65 ;
      END
   END n_36922

   PIN n_36928
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 133.15 183 133.25 ;
      END
   END n_36928

   PIN n_36944
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 173.85 0 173.95 0.51 ;
      END
   END n_36944

   PIN n_36948
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 171.85 0 171.95 0.51 ;
      END
   END n_36948

   PIN n_36953
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 52.35 183 52.45 ;
      END
   END n_36953

   PIN n_36965
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 52.15 183 52.25 ;
      END
   END n_36965

   PIN n_36980
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 119.65 0 119.75 0.51 ;
      END
   END n_36980

   PIN n_39130
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 52.55 0.51 52.65 ;
      END
   END n_39130

   PIN n_39362
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 24.95 0.51 25.05 ;
      END
   END n_39362

   PIN n_42401
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 115.55 0.51 115.65 ;
      END
   END n_42401

   PIN n_43309
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 195.3 0.255 195.5 ;
      END
   END n_43309

   PIN n_45751
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 196.95 0.51 197.05 ;
      END
   END n_45751

   PIN n_45752
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 76.85 249.49 76.95 250 ;
      END
   END n_45752

   PIN n_46296
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 38.45 249.49 38.55 250 ;
      END
   END n_46296

   PIN n_51091
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 204.95 183 205.05 ;
      END
   END n_51091

   PIN n_53413
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 146.95 183 147.05 ;
      END
   END n_53413

   PIN n_56864
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 194.95 0.51 195.05 ;
      END
   END n_56864

   PIN n_56944
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 163.85 249.49 163.95 250 ;
      END
   END n_56944

   PIN n_57
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 56.85 0 56.95 0.51 ;
      END
   END n_57

   PIN n_57749
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 161.35 183 161.45 ;
      END
   END n_57749

   PIN n_57753
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 152.75 183 152.85 ;
      END
   END n_57753

   PIN n_58050
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 152.55 183 152.65 ;
      END
   END n_58050

   PIN n_58450
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 137.85 249.49 137.95 250 ;
      END
   END n_58450

   PIN n_58539
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 174.05 249.49 174.15 250 ;
      END
   END n_58539

   PIN n_58771
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 182.49 132.95 183 133.05 ;
      END
   END n_58771

   PIN n_58784
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 60.95 0.51 61.05 ;
      END
   END n_58784

   PIN n_6033
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 89.15 183 89.25 ;
      END
   END n_6033

   PIN n_60540
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 35.55 0.51 35.65 ;
      END
   END n_60540

   PIN n_60542
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 67.35 0.51 67.45 ;
      END
   END n_60542

   PIN n_60548
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 81.95 0.51 82.05 ;
      END
   END n_60548

   PIN n_60638
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 188.15 0.51 188.25 ;
      END
   END n_60638

   PIN n_64833
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 143.5 0.255 143.7 ;
      END
   END n_64833

   PIN n_64835
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 170.5 0.255 170.7 ;
      END
   END n_64835

   PIN n_65250
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 182.49 244.95 183 245.05 ;
      END
   END n_65250

   PIN n_66515
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 35.75 0.51 35.85 ;
      END
   END n_66515

   PIN n_67153
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 139.35 0.51 139.45 ;
      END
   END n_67153

   PIN ternarymux_ln49_0_unr72_z_1_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 170.15 0.51 170.25 ;
      END
   END ternarymux_ln49_0_unr72_z_1_

   PIN ternarymux_ln49_0_unr75_z_0_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 225.35 0.51 225.45 ;
      END
   END ternarymux_ln49_0_unr75_z_0_

   PIN ternarymux_ln49_0_unr75_z_2_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 214.35 0.51 214.45 ;
      END
   END ternarymux_ln49_0_unr75_z_2_

   PIN ternarymux_ln49_0_unr75_z_3_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 224.95 0.51 225.05 ;
      END
   END ternarymux_ln49_0_unr75_z_3_

   PIN ternarymux_ln49_0_unr75_z_4_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 225.15 0.51 225.25 ;
      END
   END ternarymux_ln49_0_unr75_z_4_

   PIN ternarymux_ln49_0_unr75_z_5_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 179.75 0.51 179.85 ;
      END
   END ternarymux_ln49_0_unr75_z_5_

   PIN ternarymux_ln49_0_unr75_z_6_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 169.55 0.51 169.65 ;
      END
   END ternarymux_ln49_0_unr75_z_6_

   PIN ternarymux_ln49_0_unr75_z_7_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 169.35 0.51 169.45 ;
      END
   END ternarymux_ln49_0_unr75_z_7_

   PIN ternarymux_ln49_0_unr76_z_5_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 167.95 0.51 168.05 ;
      END
   END ternarymux_ln49_0_unr76_z_5_

   PIN ternarymux_ln49_0_unr76_z_6_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 171.35 0.51 171.45 ;
      END
   END ternarymux_ln49_0_unr76_z_6_

   PIN ternarymux_ln49_0_unr76_z_7_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 162.95 0.51 163.05 ;
      END
   END ternarymux_ln49_0_unr76_z_7_

   PIN ternarymux_ln49_0_unr76_z_9__4331226
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 142.95 0.51 143.05 ;
      END
   END ternarymux_ln49_0_unr76_z_9__4331226

   PIN ternarymux_ln49_6_unr77_z_8_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 90.95 0.51 91.05 ;
      END
   END ternarymux_ln49_6_unr77_z_8_

   PIN ternarymux_ln49_8_unr72_z_0_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 214.15 0.51 214.25 ;
      END
   END ternarymux_ln49_8_unr72_z_0_

   PIN ternarymux_ln49_8_unr72_z_1_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 214.55 0.51 214.65 ;
      END
   END ternarymux_ln49_8_unr72_z_1_

   PIN ternarymux_ln49_8_unr78_z_10_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 23.95 0.51 24.05 ;
      END
   END ternarymux_ln49_8_unr78_z_10_

   PIN ternarymux_ln49_unr75_z_0_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 216.95 0.51 217.05 ;
      END
   END ternarymux_ln49_unr75_z_0_

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 183 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 183 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 183 8.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 11.745 183 12.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 15.745 183 16.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 19.745 183 20.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 23.745 183 24.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 27.745 183 28.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 31.745 183 32.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 35.745 183 36.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 39.745 183 40.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 43.745 183 44.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 47.745 183 48.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 51.745 183 52.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 55.745 183 56.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 59.745 183 60.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 63.745 183 64.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 67.745 183 68.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 71.745 183 72.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 75.745 183 76.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 79.745 183 80.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 83.745 183 84.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 87.745 183 88.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 91.745 183 92.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 95.745 183 96.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 99.745 183 100.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 103.745 183 104.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 107.745 183 108.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 111.745 183 112.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 115.745 183 116.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 119.745 183 120.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 123.745 183 124.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 127.745 183 128.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 131.745 183 132.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 135.745 183 136.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 139.745 183 140.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 143.745 183 144.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 147.745 183 148.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 151.745 183 152.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 155.745 183 156.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 159.745 183 160.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 163.745 183 164.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 167.745 183 168.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 171.745 183 172.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 175.745 183 176.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 179.745 183 180.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 183.745 183 184.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 187.745 183 188.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 191.745 183 192.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 195.745 183 196.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 199.745 183 200.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 203.745 183 204.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 207.745 183 208.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 211.745 183 212.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 215.745 183 216.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 219.745 183 220.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 223.745 183 224.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 227.745 183 228.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 231.745 183 232.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 235.745 183 236.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 239.745 183 240.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 243.745 183 244.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 247.745 183 248.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 183 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 183 6.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 9.745 183 10.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 13.745 183 14.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 17.745 183 18.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 21.745 183 22.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 25.745 183 26.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 29.745 183 30.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 33.745 183 34.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 37.745 183 38.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 41.745 183 42.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 45.745 183 46.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 49.745 183 50.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 53.745 183 54.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 57.745 183 58.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 61.745 183 62.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 65.745 183 66.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 69.745 183 70.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 73.745 183 74.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 77.745 183 78.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 81.745 183 82.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 85.745 183 86.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 89.745 183 90.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 93.745 183 94.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 97.745 183 98.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 101.745 183 102.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 105.745 183 106.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 109.745 183 110.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 113.745 183 114.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 117.745 183 118.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 121.745 183 122.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 125.745 183 126.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 129.745 183 130.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 133.745 183 134.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 137.745 183 138.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 141.745 183 142.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 145.745 183 146.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 149.745 183 150.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 153.745 183 154.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 157.745 183 158.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 161.745 183 162.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 165.745 183 166.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 169.745 183 170.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 173.745 183 174.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 177.745 183 178.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 181.745 183 182.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 185.745 183 186.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 189.745 183 190.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 193.745 183 194.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 197.745 183 198.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 201.745 183 202.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 205.745 183 206.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 209.745 183 210.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 213.745 183 214.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 217.745 183 218.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 221.745 183 222.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 225.745 183 226.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 229.745 183 230.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 233.745 183 234.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 237.745 183 238.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 241.745 183 242.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 245.745 183 246.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 249.745 183 250.255 ;
      END
   END vdd

   OBS
      LAYER metal1 ;
         RECT 0 0 183 250 ;
   END
   OBS
      LAYER metal2 ;
         RECT 0 0 183 250 ;
   END
   OBS
      LAYER metal3 ;
         RECT 0 0 183 250 ;
   END
   OBS
      LAYER metal4 ;
         RECT 0 0 183 250 ;
   END
   OBS
      LAYER metal5 ;
         RECT 0 0 183 250 ;
   END
END h1

MACRO ms00f80
   CLASS CORE ;
   SIZE 1.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN ck
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END ck

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.05 0.5 1.15 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.6 2.255 ;
      END
   END vdd

END ms00f80

MACRO in01f01
   CLASS CORE ;
   SIZE 0.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 0.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 0.4 2.255 ;
      END
   END vdd

END in01f01

MACRO oa12f01
   CLASS CORE ;
   SIZE 1.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
   END vdd

END oa12f01

MACRO na03f01
   CLASS CORE ;
   SIZE 1.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
   END vdd

END na03f01

MACRO na04m01
   CLASS CORE ;
   SIZE 1.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.6 2.255 ;
      END
   END vdd

END na04m01

MACRO na02f01
   CLASS CORE ;
   SIZE 0.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 0.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 0.8 2.255 ;
      END
   END vdd

END na02f01

MACRO no02f01
   CLASS CORE ;
   SIZE 0.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 0.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 0.8 2.255 ;
      END
   END vdd

END no02f01

MACRO ao12f01
   CLASS CORE ;
   SIZE 1.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
   END vdd

END ao12f01

MACRO ao22s01
   CLASS CORE ;
   SIZE 1.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.6 2.255 ;
      END
   END vdd

END ao22s01

MACRO oa22f01
   CLASS CORE ;
   SIZE 1.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 1.35 0.95 1.55 1.05 ;
         LAYER metal2 ;
             RECT 1.25 0.5 1.35 1.05 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.6 2.255 ;
      END
   END vdd

END oa22f01

MACRO no03m01
   CLASS CORE ;
   SIZE 1.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
   END vdd

END no03m01

MACRO oa22m01
   CLASS CORE ;
   SIZE 1.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.6 2.255 ;
      END
   END vdd

END oa22m01

MACRO no04s01
   CLASS CORE ;
   SIZE 1.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.6 2.255 ;
      END
   END vdd

END no04s01

MACRO in01s80
   CLASS CORE ;
   SIZE 51.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.2 2.255 ;
      END
   END vdd

END in01s80

MACRO in01f01X2HE
   CLASS CORE ;
   SIZE 1.2 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 1.2 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
   END vdd

END in01f01X2HE

MACRO in01f01X2HO
   CLASS CORE ;
   SIZE 0.8 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 0.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 0.8 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 0.8 2.255 ;
      END
   END vss

END in01f01X2HO

MACRO in01f01X3H
   CLASS CORE ;
   SIZE 1.2 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 4.5 0.55 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 1.2 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 1.2 6.255 ;
      END
   END vdd

END in01f01X3H

MACRO in01f01X4HE
   CLASS CORE ;
   SIZE 1.2 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 4.5 0.75 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 1.2 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 1.2 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 1.2 6.255 ;
      END
   END vdd

END in01f01X4HE

MACRO in01f01X4HO
   CLASS CORE ;
   SIZE 1.6 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 4.5 0.95 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 1.6 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 1.6 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.6 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 1.6 6.255 ;
      END
   END vss

END in01f01X4HO

MACRO in01s80X2HE
   CLASS CORE ;
   SIZE 51.2 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 51.2 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.2 2.255 ;
      END
   END vdd

END in01s80X2HE

MACRO in01s80X2HO
   CLASS CORE ;
   SIZE 51.2 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 51.2 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.2 2.255 ;
      END
   END vss

END in01s80X2HO

MACRO in01s80X3H
   CLASS CORE ;
   SIZE 51.2 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 4.5 0.15 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 51.2 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.2 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 51.2 6.255 ;
      END
   END vdd

END in01s80X3H

MACRO in01s80X4HE
   CLASS CORE ;
   SIZE 51.2 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 4.5 25.75 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 51.2 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 51.2 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.2 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 51.2 6.255 ;
      END
   END vdd

END in01s80X4HE

MACRO in01s80X4HO
   CLASS CORE ;
   SIZE 51.2 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 4.5 25.75 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 51.2 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 51.2 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.2 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 51.2 6.255 ;
      END
   END vss

END in01s80X4HO

END LIBRARY
