module top ();
 LOGIC1_X1 t1 (.Z(n1));
 BUF_X1 u0 (.A(n1));
 BUF_X1 u1 (.A(n1));
 BUF_X1 u2 (.A(n1));
 BUF_X1 u3 (.A(n1));
 BUF_X1 u4 (.A(n1));
 BUF_X1 u5 (.A(n1));
 BUF_X1 u6 (.A(n1));
 BUF_X1 u7 (.A(n1));
 BUF_X1 u8 (.A(n1));
 BUF_X1 u9 (.A(n1));
 BUF_X1 u10 (.A(n1));
 BUF_X1 u11 (.A(n1));
 BUF_X1 u12 (.A(n1));
 BUF_X1 u13 (.A(n1));
 BUF_X1 u14 (.A(n1));
 BUF_X1 u15 (.A(n1));
 BUF_X1 u16 (.A(n1));
 BUF_X1 u17 (.A(n1));
 BUF_X1 u18 (.A(n1));
 BUF_X1 u19 (.A(n1));
 BUF_X1 u20 (.A(n1));
 BUF_X1 u21 (.A(n1));
 BUF_X1 u22 (.A(n1));
 BUF_X1 u23 (.A(n1));
 BUF_X1 u24 (.A(n1));
 BUF_X1 u25 (.A(n1));
 BUF_X1 u26 (.A(n1));
 BUF_X1 u27 (.A(n1));
 BUF_X1 u28 (.A(n1));
 BUF_X1 u29 (.A(n1));
 BUF_X1 u30 (.A(n1));
 BUF_X1 u31 (.A(n1));
 BUF_X1 u32 (.A(n1));
 BUF_X1 u33 (.A(n1));
 BUF_X1 u34 (.A(n1));
 BUF_X1 u35 (.A(n1));
 BUF_X1 u36 (.A(n1));
 BUF_X1 u37 (.A(n1));
 BUF_X1 u38 (.A(n1));
 BUF_X1 u39 (.A(n1));
 BUF_X1 u40 (.A(n1));
 BUF_X1 u41 (.A(n1));
 BUF_X1 u42 (.A(n1));
 BUF_X1 u43 (.A(n1));
 BUF_X1 u44 (.A(n1));
 BUF_X1 u45 (.A(n1));
 BUF_X1 u46 (.A(n1));
 BUF_X1 u47 (.A(n1));
 BUF_X1 u48 (.A(n1));
 BUF_X1 u49 (.A(n1));
 BUF_X1 u50 (.A(n1));
 BUF_X1 u51 (.A(n1));
 BUF_X1 u52 (.A(n1));
 BUF_X1 u53 (.A(n1));
 BUF_X1 u54 (.A(n1));
 BUF_X1 u55 (.A(n1));
 BUF_X1 u56 (.A(n1));
 BUF_X1 u57 (.A(n1));
 BUF_X1 u58 (.A(n1));
 BUF_X1 u59 (.A(n1));
 BUF_X1 u60 (.A(n1));
 BUF_X1 u61 (.A(n1));
 BUF_X1 u62 (.A(n1));
 BUF_X1 u63 (.A(n1));
 BUF_X1 u64 (.A(n1));
 BUF_X1 u65 (.A(n1));
 BUF_X1 u66 (.A(n1));
 BUF_X1 u67 (.A(n1));
 BUF_X1 u68 (.A(n1));
 BUF_X1 u69 (.A(n1));
 BUF_X1 u70 (.A(n1));
 BUF_X1 u71 (.A(n1));
 BUF_X1 u72 (.A(n1));
 BUF_X1 u73 (.A(n1));
 BUF_X1 u74 (.A(n1));
 BUF_X1 u75 (.A(n1));
 BUF_X1 u76 (.A(n1));
 BUF_X1 u77 (.A(n1));
 BUF_X1 u78 (.A(n1));
 BUF_X1 u79 (.A(n1));
 BUF_X1 u80 (.A(n1));
 BUF_X1 u81 (.A(n1));
 BUF_X1 u82 (.A(n1));
 BUF_X1 u83 (.A(n1));
 BUF_X1 u84 (.A(n1));
 BUF_X1 u85 (.A(n1));
 BUF_X1 u86 (.A(n1));
 BUF_X1 u87 (.A(n1));
 BUF_X1 u88 (.A(n1));
 BUF_X1 u89 (.A(n1));
 BUF_X1 u90 (.A(n1));
 BUF_X1 u91 (.A(n1));
 PAD pad1 (.IN(n1));
 PAD pad2 (.IN(n1));
 PAD pad3 (.IN(n1));
 PAD pad4 (.IN(n1));
 PAD pad5 (.IN(n1));
 PAD pad6 (.IN(n1));
 PAD pad7 (.IN(n1));
 PAD pad8 (.IN(n1));
 PAD pad9 (.IN(n1));
 PAD pad10 (.IN(n1));
 PAD pad11 (.IN(n1));
endmodule
