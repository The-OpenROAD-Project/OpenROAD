VERSION 5.5 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO ms00f80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN ck
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END ck

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.05 0.5 1.15 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.6 2.255 ;
      END
   END vdd

END ms00f80

MACRO oa22f80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 204.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 40.85 0.5 40.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 81.85 0.5 81.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 122.8 0.5 122.9 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 163.9 0.5 164 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 204.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 204.8 2.255 ;
      END
   END vdd

END oa22f80

MACRO oa22f40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 102.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 20.45 0.5 20.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 40.85 0.5 40.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 61.45 0.5 61.55 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 81.85 0.5 81.95 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 102.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 102.4 2.255 ;
      END
   END vdd

END oa22f40

MACRO oa22f20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 51.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 10.25 0.5 10.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 20.45 0.5 20.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 30.65 0.5 30.75 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 40.85 0.5 40.95 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.2 2.255 ;
      END
   END vdd

END oa22f20

MACRO oa22f10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.05 0.5 5.15 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 10.25 0.5 10.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 15.25 0.5 15.35 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 20.45 0.5 20.55 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.6 2.255 ;
      END
   END vdd

END oa22f10

MACRO oa22f08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.05 0.5 5.15 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 7.65 0.5 7.75 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 10.25 0.5 10.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
   END vdd

END oa22f08

MACRO oa22f06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 9.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.85 0.5 3.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.65 0.5 5.75 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 7.65 0.5 7.75 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 9.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 9.6 2.255 ;
      END
   END vdd

END oa22f06

MACRO oa22f04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.85 0.5 3.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.05 0.5 5.15 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6.4 2.255 ;
      END
   END vdd

END oa22f04

MACRO oa22f03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.85 0.5 2.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.85 0.5 3.95 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4.8 2.255 ;
      END
   END vdd

END oa22f03

MACRO oa22f02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.2 2.255 ;
      END
   END vdd

END oa22f02

MACRO oa22f01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 1 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 0 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.6 2.255 ;
      END
   END vdd

END oa22f01

MACRO oa22m80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 204.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 40.85 0.5 40.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 81.85 0.5 81.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 122.8 0.5 122.9 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 163.9 0.5 164 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 204.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 204.8 2.255 ;
      END
   END vdd

END oa22m80

MACRO oa22m40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 102.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 20.45 0.5 20.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 40.85 0.5 40.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 61.45 0.5 61.55 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 81.85 0.5 81.95 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 102.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 102.4 2.255 ;
      END
   END vdd

END oa22m40

MACRO oa22m20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 51.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 10.25 0.5 10.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 20.45 0.5 20.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 30.65 0.5 30.75 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 40.85 0.5 40.95 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.2 2.255 ;
      END
   END vdd

END oa22m20

MACRO oa22m10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.05 0.5 5.15 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 10.25 0.5 10.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 15.25 0.5 15.35 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 20.45 0.5 20.55 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.6 2.255 ;
      END
   END vdd

END oa22m10

MACRO oa22m08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.05 0.5 5.15 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 7.65 0.5 7.75 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 10.25 0.5 10.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
   END vdd

END oa22m08

MACRO oa22m06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 9.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.85 0.5 3.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.65 0.5 5.75 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 7.65 0.5 7.75 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 9.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 9.6 2.255 ;
      END
   END vdd

END oa22m06

MACRO oa22m04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.85 0.5 3.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.05 0.5 5.15 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6.4 2.255 ;
      END
   END vdd

END oa22m04

MACRO oa22m03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.85 0.5 2.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.85 0.5 3.95 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4.8 2.255 ;
      END
   END vdd

END oa22m03

MACRO oa22m02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.2 2.255 ;
      END
   END vdd

END oa22m02

MACRO oa22m01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.6 2.255 ;
      END
   END vdd

END oa22m01

MACRO oa22s80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 204.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 40.85 0.5 40.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 81.85 0.5 81.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 122.8 0.5 122.9 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 163.9 0.5 164 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 204.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 204.8 2.255 ;
      END
   END vdd

END oa22s80

MACRO oa22s40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 102.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 20.45 0.5 20.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 40.85 0.5 40.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 61.45 0.5 61.55 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 81.85 0.5 81.95 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 102.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 102.4 2.255 ;
      END
   END vdd

END oa22s40

MACRO oa22s20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 51.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 10.25 0.5 10.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 20.45 0.5 20.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 30.65 0.5 30.75 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 40.85 0.5 40.95 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.2 2.255 ;
      END
   END vdd

END oa22s20

MACRO oa22s10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.05 0.5 5.15 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 10.25 0.5 10.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 15.25 0.5 15.35 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 20.45 0.5 20.55 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.6 2.255 ;
      END
   END vdd

END oa22s10

MACRO oa22s08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.05 0.5 5.15 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 7.65 0.5 7.75 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 10.25 0.5 10.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
   END vdd

END oa22s08

MACRO oa22s06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 9.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.85 0.5 3.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.65 0.5 5.75 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 7.65 0.5 7.75 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 9.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 9.6 2.255 ;
      END
   END vdd

END oa22s06

MACRO oa22s04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.85 0.5 3.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.05 0.5 5.15 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6.4 2.255 ;
      END
   END vdd

END oa22s04

MACRO oa22s03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.85 0.5 2.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.85 0.5 3.95 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4.8 2.255 ;
      END
   END vdd

END oa22s03

MACRO oa22s02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.2 2.255 ;
      END
   END vdd

END oa22s02

MACRO oa22s01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.6 2.255 ;
      END
   END vdd

END oa22s01

MACRO oa12f80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 153.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 38.45 0.5 38.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 76.85 0.5 76.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 115.2 0.5 115.3 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 153.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 153.6 2.255 ;
      END
   END vdd

END oa12f80

MACRO oa12f40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 76.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 19.25 0.5 19.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 38.45 0.5 38.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 57.65 0.5 57.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 76.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 76.8 2.255 ;
      END
   END vdd

END oa12f40

MACRO oa12f20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 38.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 9.65 0.5 9.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 19.25 0.5 19.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 28.85 0.5 28.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 38.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 38.4 2.255 ;
      END
   END vdd

END oa12f20

MACRO oa12f10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 19.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 9.65 0.5 9.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 14.45 0.5 14.55 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 19.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 19.2 2.255 ;
      END
   END vdd

END oa12f10

MACRO oa12f08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 9.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 7.25 0.5 7.35 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 9.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 9.6 2.255 ;
      END
   END vdd

END oa12f08

MACRO oa12f06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 7.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.65 0.5 3.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.45 0.5 5.55 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 7.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 7.2 2.255 ;
      END
   END vdd

END oa12f06

MACRO oa12f04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.65 0.5 3.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4.8 2.255 ;
      END
   END vdd

END oa12f04

MACRO oa12f03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.65 0.5 2.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.6 2.255 ;
      END
   END vdd

END oa12f03

MACRO oa12f02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
   END vdd

END oa12f02

MACRO oa12f01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
   END vdd

END oa12f01

MACRO oa12m80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 153.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 38.45 0.5 38.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 76.85 0.5 76.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 115.2 0.5 115.3 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 153.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 153.6 2.255 ;
      END
   END vdd

END oa12m80

MACRO oa12m40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 76.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 19.25 0.5 19.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 38.45 0.5 38.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 57.65 0.5 57.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 76.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 76.8 2.255 ;
      END
   END vdd

END oa12m40

MACRO oa12m20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 38.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 9.65 0.5 9.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 19.25 0.5 19.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 28.85 0.5 28.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 38.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 38.4 2.255 ;
      END
   END vdd

END oa12m20

MACRO oa12m10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 19.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 9.65 0.5 9.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 14.45 0.5 14.55 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 19.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 19.2 2.255 ;
      END
   END vdd

END oa12m10

MACRO oa12m08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 9.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 7.25 0.5 7.35 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 9.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 9.6 2.255 ;
      END
   END vdd

END oa12m08

MACRO oa12m06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 7.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.65 0.5 3.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.45 0.5 5.55 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 7.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 7.2 2.255 ;
      END
   END vdd

END oa12m06

MACRO oa12m04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.65 0.5 3.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4.8 2.255 ;
      END
   END vdd

END oa12m04

MACRO oa12m03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.65 0.5 2.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.6 2.255 ;
      END
   END vdd

END oa12m03

MACRO oa12m02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
   END vdd

END oa12m02

MACRO oa12m01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
   END vdd

END oa12m01

MACRO oa12s80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 153.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 38.45 0.5 38.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 76.85 0.5 76.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 115.2 0.5 115.3 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 153.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 153.6 2.255 ;
      END
   END vdd

END oa12s80

MACRO oa12s40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 76.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 19.25 0.5 19.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 38.45 0.5 38.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 57.65 0.5 57.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 76.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 76.8 2.255 ;
      END
   END vdd

END oa12s40

MACRO oa12s20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 38.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 9.65 0.5 9.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 19.25 0.5 19.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 28.85 0.5 28.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 38.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 38.4 2.255 ;
      END
   END vdd

END oa12s20

MACRO oa12s10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 19.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 9.65 0.5 9.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 14.45 0.5 14.55 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 19.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 19.2 2.255 ;
      END
   END vdd

END oa12s10

MACRO oa12s08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 9.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 7.25 0.5 7.35 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 9.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 9.6 2.255 ;
      END
   END vdd

END oa12s08

MACRO oa12s06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 7.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.65 0.5 3.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.45 0.5 5.55 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 7.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 7.2 2.255 ;
      END
   END vdd

END oa12s06

MACRO oa12s04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.65 0.5 3.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4.8 2.255 ;
      END
   END vdd

END oa12s04

MACRO oa12s03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.65 0.5 2.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.6 2.255 ;
      END
   END vdd

END oa12s03

MACRO oa12s02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
   END vdd

END oa12s02

MACRO oa12s01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
   END vdd

END oa12s01

MACRO ao22f80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 204.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 40.85 0.5 40.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 81.85 0.5 81.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 122.8 0.5 122.9 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 163.9 0.5 164 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 204.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 204.8 2.255 ;
      END
   END vdd

END ao22f80

MACRO ao22f40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 102.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 20.45 0.5 20.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 40.85 0.5 40.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 61.45 0.5 61.55 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 81.85 0.5 81.95 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 102.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 102.4 2.255 ;
      END
   END vdd

END ao22f40

MACRO ao22f20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 51.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 10.25 0.5 10.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 20.45 0.5 20.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 30.65 0.5 30.75 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 40.85 0.5 40.95 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.2 2.255 ;
      END
   END vdd

END ao22f20

MACRO ao22f10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.05 0.5 5.15 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 10.25 0.5 10.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 15.25 0.5 15.35 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 20.45 0.5 20.55 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.6 2.255 ;
      END
   END vdd

END ao22f10

MACRO ao22f08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.05 0.5 5.15 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 7.65 0.5 7.75 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 10.25 0.5 10.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
   END vdd

END ao22f08

MACRO ao22f06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 9.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.85 0.5 3.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.65 0.5 5.75 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 7.65 0.5 7.75 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 9.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 9.6 2.255 ;
      END
   END vdd

END ao22f06

MACRO ao22f04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.85 0.5 3.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.05 0.5 5.15 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6.4 2.255 ;
      END
   END vdd

END ao22f04

MACRO ao22f03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.85 0.5 2.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.85 0.5 3.95 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4.8 2.255 ;
      END
   END vdd

END ao22f03

MACRO ao22f02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.2 2.255 ;
      END
   END vdd

END ao22f02

MACRO ao22f01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.6 2.255 ;
      END
   END vdd

END ao22f01

MACRO ao22m80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 204.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 40.85 0.5 40.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 81.85 0.5 81.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 122.8 0.5 122.9 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 163.9 0.5 164 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 204.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 204.8 2.255 ;
      END
   END vdd

END ao22m80

MACRO ao22m40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 102.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 20.45 0.5 20.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 40.85 0.5 40.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 61.45 0.5 61.55 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 81.85 0.5 81.95 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 102.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 102.4 2.255 ;
      END
   END vdd

END ao22m40

MACRO ao22m20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 51.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 10.25 0.5 10.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 20.45 0.5 20.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 30.65 0.5 30.75 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 40.85 0.5 40.95 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.2 2.255 ;
      END
   END vdd

END ao22m20

MACRO ao22m10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.05 0.5 5.15 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 10.25 0.5 10.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 15.25 0.5 15.35 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 20.45 0.5 20.55 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.6 2.255 ;
      END
   END vdd

END ao22m10

MACRO ao22m08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.05 0.5 5.15 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 7.65 0.5 7.75 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 10.25 0.5 10.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
   END vdd

END ao22m08

MACRO ao22m06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 9.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.85 0.5 3.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.65 0.5 5.75 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 7.65 0.5 7.75 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 9.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 9.6 2.255 ;
      END
   END vdd

END ao22m06

MACRO ao22m04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.85 0.5 3.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.05 0.5 5.15 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6.4 2.255 ;
      END
   END vdd

END ao22m04

MACRO ao22m03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.85 0.5 2.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.85 0.5 3.95 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4.8 2.255 ;
      END
   END vdd

END ao22m03

MACRO ao22m02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.2 2.255 ;
      END
   END vdd

END ao22m02

MACRO ao22m01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.6 2.255 ;
      END
   END vdd

END ao22m01

MACRO ao22s80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 204.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 40.85 0.5 40.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 81.85 0.5 81.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 122.8 0.5 122.9 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 163.9 0.5 164 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 204.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 204.8 2.255 ;
      END
   END vdd

END ao22s80

MACRO ao22s40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 102.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 20.45 0.5 20.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 40.85 0.5 40.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 61.45 0.5 61.55 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 81.85 0.5 81.95 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 102.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 102.4 2.255 ;
      END
   END vdd

END ao22s40

MACRO ao22s20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 51.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 10.25 0.5 10.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 20.45 0.5 20.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 30.65 0.5 30.75 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 40.85 0.5 40.95 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.2 2.255 ;
      END
   END vdd

END ao22s20

MACRO ao22s10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.05 0.5 5.15 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 10.25 0.5 10.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 15.25 0.5 15.35 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 20.45 0.5 20.55 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.6 2.255 ;
      END
   END vdd

END ao22s10

MACRO ao22s08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.05 0.5 5.15 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 7.65 0.5 7.75 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 10.25 0.5 10.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
   END vdd

END ao22s08

MACRO ao22s06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 9.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.85 0.5 3.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.65 0.5 5.75 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 7.65 0.5 7.75 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 9.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 9.6 2.255 ;
      END
   END vdd

END ao22s06

MACRO ao22s04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.85 0.5 3.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.05 0.5 5.15 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6.4 2.255 ;
      END
   END vdd

END ao22s04

MACRO ao22s03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.85 0.5 2.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.85 0.5 3.95 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4.8 2.255 ;
      END
   END vdd

END ao22s03

MACRO ao22s02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.2 2.255 ;
      END
   END vdd

END ao22s02

MACRO ao22s01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 1 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.6 2.255 ;
      END
   END vdd

END ao22s01

MACRO ao12f80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 153.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 38.45 0.5 38.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 76.85 0.5 76.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 115.2 0.5 115.3 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 153.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 153.6 2.255 ;
      END
   END vdd

END ao12f80

MACRO ao12f40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 76.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 19.25 0.5 19.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 38.45 0.5 38.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 57.65 0.5 57.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 76.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 76.8 2.255 ;
      END
   END vdd

END ao12f40

MACRO ao12f20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 38.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 9.65 0.5 9.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 19.25 0.5 19.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 28.85 0.5 28.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 38.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 38.4 2.255 ;
      END
   END vdd

END ao12f20

MACRO ao12f10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 19.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 9.65 0.5 9.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 14.45 0.5 14.55 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 19.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 19.2 2.255 ;
      END
   END vdd

END ao12f10

MACRO ao12f08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 9.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 7.25 0.5 7.35 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 9.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 9.6 2.255 ;
      END
   END vdd

END ao12f08

MACRO ao12f06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 7.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.65 0.5 3.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.45 0.5 5.55 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 7.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 7.2 2.255 ;
      END
   END vdd

END ao12f06

MACRO ao12f04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.65 0.5 3.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4.8 2.255 ;
      END
   END vdd

END ao12f04

MACRO ao12f03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.65 0.5 2.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.6 2.255 ;
      END
   END vdd

END ao12f03

MACRO ao12f02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
   END vdd

END ao12f02

MACRO ao12f01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
   END vdd

END ao12f01

MACRO ao12m80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 153.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 38.45 0.5 38.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 76.85 0.5 76.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 115.2 0.5 115.3 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 153.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 153.6 2.255 ;
      END
   END vdd

END ao12m80

MACRO ao12m40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 76.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 19.25 0.5 19.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 38.45 0.5 38.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 57.65 0.5 57.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 76.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 76.8 2.255 ;
      END
   END vdd

END ao12m40

MACRO ao12m20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 38.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 9.65 0.5 9.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 19.25 0.5 19.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 28.85 0.5 28.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 38.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 38.4 2.255 ;
      END
   END vdd

END ao12m20

MACRO ao12m10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 19.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 9.65 0.5 9.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 14.45 0.5 14.55 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 19.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 19.2 2.255 ;
      END
   END vdd

END ao12m10

MACRO ao12m08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 9.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 7.25 0.5 7.35 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 9.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 9.6 2.255 ;
      END
   END vdd

END ao12m08

MACRO ao12m06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 7.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.65 0.5 3.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.45 0.5 5.55 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 7.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 7.2 2.255 ;
      END
   END vdd

END ao12m06

MACRO ao12m04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.65 0.5 3.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4.8 2.255 ;
      END
   END vdd

END ao12m04

MACRO ao12m03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.65 0.5 2.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.6 2.255 ;
      END
   END vdd

END ao12m03

MACRO ao12m02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
   END vdd

END ao12m02

MACRO ao12m01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
   END vdd

END ao12m01

MACRO ao12s80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 153.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 38.45 0.5 38.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 76.85 0.5 76.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 115.2 0.5 115.3 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 153.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 153.6 2.255 ;
      END
   END vdd

END ao12s80

MACRO ao12s40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 76.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 19.25 0.5 19.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 38.45 0.5 38.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 57.65 0.5 57.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 76.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 76.8 2.255 ;
      END
   END vdd

END ao12s40

MACRO ao12s20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 38.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 9.65 0.5 9.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 19.25 0.5 19.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 28.85 0.5 28.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 38.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 38.4 2.255 ;
      END
   END vdd

END ao12s20

MACRO ao12s10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 19.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 9.65 0.5 9.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 14.45 0.5 14.55 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 19.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 19.2 2.255 ;
      END
   END vdd

END ao12s10

MACRO ao12s08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 9.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 7.25 0.5 7.35 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 9.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 9.6 2.255 ;
      END
   END vdd

END ao12s08

MACRO ao12s06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 7.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.65 0.5 3.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.45 0.5 5.55 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 7.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 7.2 2.255 ;
      END
   END vdd

END ao12s06

MACRO ao12s04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.65 0.5 3.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4.8 2.255 ;
      END
   END vdd

END ao12s04

MACRO ao12s03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.65 0.5 2.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.6 2.255 ;
      END
   END vdd

END ao12s03

MACRO ao12s02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
   END vdd

END ao12s02

MACRO ao12s01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
   END vdd

END ao12s01

MACRO no04f80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 128 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 51.25 0.5 51.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 76.85 0.5 76.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 102.5 0.5 102.6 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 128 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 128 2.255 ;
      END
   END vdd

END no04f80

MACRO no04f40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 64 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 38.45 0.5 38.55 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 51.25 0.5 51.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 64 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 64 2.255 ;
      END
   END vdd

END no04f40

MACRO no04f20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 32 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 19.25 0.5 19.35 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 32 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 32 2.255 ;
      END
   END vdd

END no04f20

MACRO no04f10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 16 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 9.65 0.5 9.75 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 16 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 16 2.255 ;
      END
   END vdd

END no04f10

MACRO no04f08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 8 2.255 ;
      END
   END vdd

END no04f08

MACRO no04f06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.85 0.5 3.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.05 0.5 5.15 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6.4 2.255 ;
      END
   END vdd

END no04f06

MACRO no04f04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4 2.255 ;
      END
   END vdd

END no04f04

MACRO no04f03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.2 2.255 ;
      END
   END vdd

END no04f03

MACRO no04f02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.45 0.5 1.55 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
   END vdd

END no04f02

MACRO no04f01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.6 2.255 ;
      END
   END vdd

END no04f01

MACRO no04m80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 128 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 51.25 0.5 51.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 76.85 0.5 76.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 102.5 0.5 102.6 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 128 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 128 2.255 ;
      END
   END vdd

END no04m80

MACRO no04m40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 64 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 38.45 0.5 38.55 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 51.25 0.5 51.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 64 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 64 2.255 ;
      END
   END vdd

END no04m40

MACRO no04m20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 32 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 19.25 0.5 19.35 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 32 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 32 2.255 ;
      END
   END vdd

END no04m20

MACRO no04m10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 16 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 9.65 0.5 9.75 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 16 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 16 2.255 ;
      END
   END vdd

END no04m10

MACRO no04m08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 8 2.255 ;
      END
   END vdd

END no04m08

MACRO no04m06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.85 0.5 3.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.05 0.5 5.15 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6.4 2.255 ;
      END
   END vdd

END no04m06

MACRO no04m04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4 2.255 ;
      END
   END vdd

END no04m04

MACRO no04m03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.2 2.255 ;
      END
   END vdd

END no04m03

MACRO no04m02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.45 0.5 1.55 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
   END vdd

END no04m02

MACRO no04m01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.6 2.255 ;
      END
   END vdd

END no04m01

MACRO no04s80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 128 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 51.25 0.5 51.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 76.85 0.5 76.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 102.5 0.5 102.6 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 128 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 128 2.255 ;
      END
   END vdd

END no04s80

MACRO no04s40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 64 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 38.45 0.5 38.55 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 51.25 0.5 51.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 64 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 64 2.255 ;
      END
   END vdd

END no04s40

MACRO no04s20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 32 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 19.25 0.5 19.35 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 32 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 32 2.255 ;
      END
   END vdd

END no04s20

MACRO no04s10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 16 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 9.65 0.5 9.75 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 16 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 16 2.255 ;
      END
   END vdd

END no04s10

MACRO no04s08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 8 2.255 ;
      END
   END vdd

END no04s08

MACRO no04s06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.85 0.5 3.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.05 0.5 5.15 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6.4 2.255 ;
      END
   END vdd

END no04s06

MACRO no04s04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4 2.255 ;
      END
   END vdd

END no04s04

MACRO no04s03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.2 2.255 ;
      END
   END vdd

END no04s03

MACRO no04s02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.45 0.5 1.55 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
   END vdd

END no04s02

MACRO no04s01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.6 2.255 ;
      END
   END vdd

END no04s01

MACRO no03f80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 102.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 51.25 0.5 51.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 76.85 0.5 76.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 102.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 102.6 2.255 ;
      END
   END vdd

END no03f80

MACRO no03f40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 51.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.85 0.5 25.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 38.65 0.5 38.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.6 2.255 ;
      END
   END vdd

END no03f40

MACRO no03f20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 19.25 0.5 19.35 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.8 2.255 ;
      END
   END vdd

END no03f20

MACRO no03f10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 13.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.65 0.5 6.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 9.85 0.5 9.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 13.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 13.2 2.255 ;
      END
   END vdd

END no03f10

MACRO no03f08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6.6 2.255 ;
      END
   END vdd

END no03f08

MACRO no03f06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.65 0.5 3.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4.8 2.255 ;
      END
   END vdd

END no03f06

MACRO no03f04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.65 0.5 2.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.6 2.255 ;
      END
   END vdd

END no03f04

MACRO no03f03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
   END vdd

END no03f03

MACRO no03f02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.8 2.255 ;
      END
   END vdd

END no03f02

MACRO no03f01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
   END vdd

END no03f01

MACRO no03m80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 102.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 51.25 0.5 51.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 76.85 0.5 76.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 102.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 102.6 2.255 ;
      END
   END vdd

END no03m80

MACRO no03m40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 51.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.85 0.5 25.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 38.65 0.5 38.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.6 2.255 ;
      END
   END vdd

END no03m40

MACRO no03m20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 19.25 0.5 19.35 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.8 2.255 ;
      END
   END vdd

END no03m20

MACRO no03m10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 13.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.65 0.5 6.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 9.85 0.5 9.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 13.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 13.2 2.255 ;
      END
   END vdd

END no03m10

MACRO no03m08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6.6 2.255 ;
      END
   END vdd

END no03m08

MACRO no03m06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.65 0.5 3.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4.8 2.255 ;
      END
   END vdd

END no03m06

MACRO no03m04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.65 0.5 2.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.6 2.255 ;
      END
   END vdd

END no03m04

MACRO no03m03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
   END vdd

END no03m03

MACRO no03m02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.8 2.255 ;
      END
   END vdd

END no03m02

MACRO no03m01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
   END vdd

END no03m01

MACRO no03s80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 102.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 51.25 0.5 51.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 76.85 0.5 76.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 102.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 102.6 2.255 ;
      END
   END vdd

END no03s80

MACRO no03s40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 51.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.85 0.5 25.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 38.65 0.5 38.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.6 2.255 ;
      END
   END vdd

END no03s40

MACRO no03s20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 19.25 0.5 19.35 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.8 2.255 ;
      END
   END vdd

END no03s20

MACRO no03s10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 13.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.65 0.5 6.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 9.85 0.5 9.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 13.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 13.2 2.255 ;
      END
   END vdd

END no03s10

MACRO no03s08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6.6 2.255 ;
      END
   END vdd

END no03s08

MACRO no03s06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.65 0.5 3.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4.8 2.255 ;
      END
   END vdd

END no03s06

MACRO no03s04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.65 0.5 2.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.6 2.255 ;
      END
   END vdd

END no03s04

MACRO no03s03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
   END vdd

END no03s03

MACRO no03s02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.8 2.255 ;
      END
   END vdd

END no03s02

MACRO no03s01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
   END vdd

END no03s01

MACRO no02f80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 76.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 51.25 0.5 51.35 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 76.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 76.8 2.255 ;
      END
   END vdd

END no02f80

MACRO no02f40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 38.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 38.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 38.4 2.255 ;
      END
   END vdd

END no02f40

MACRO no02f20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 19.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 19.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 19.2 2.255 ;
      END
   END vdd

END no02f20

MACRO no02f10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 9.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 9.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 9.6 2.255 ;
      END
   END vdd

END no02f10

MACRO no02f08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4.8 2.255 ;
      END
   END vdd

END no02f08

MACRO no02f06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.6 2.255 ;
      END
   END vdd

END no02f06

MACRO no02f04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
   END vdd

END no02f04

MACRO no02f03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2 2.255 ;
      END
   END vdd

END no02f03

MACRO no02f02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
   END vdd

END no02f02

MACRO no02f01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 0.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 0.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 0.8 2.255 ;
      END
   END vdd

END no02f01

MACRO no02m80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 76.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 51.25 0.5 51.35 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 76.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 76.8 2.255 ;
      END
   END vdd

END no02m80

MACRO no02m40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 38.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 38.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 38.4 2.255 ;
      END
   END vdd

END no02m40

MACRO no02m20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 19.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 19.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 19.2 2.255 ;
      END
   END vdd

END no02m20

MACRO no02m10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 9.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 9.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 9.6 2.255 ;
      END
   END vdd

END no02m10

MACRO no02m08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4.8 2.255 ;
      END
   END vdd

END no02m08

MACRO no02m06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.6 2.255 ;
      END
   END vdd

END no02m06

MACRO no02m04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
   END vdd

END no02m04

MACRO no02m03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2 2.255 ;
      END
   END vdd

END no02m03

MACRO no02m02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
   END vdd

END no02m02

MACRO no02m01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 0.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 0.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 0.8 2.255 ;
      END
   END vdd

END no02m01

MACRO no02s80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 76.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 51.25 0.5 51.35 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 76.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 76.8 2.255 ;
      END
   END vdd

END no02s80

MACRO no02s40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 38.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 38.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 38.4 2.255 ;
      END
   END vdd

END no02s40

MACRO no02s20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 19.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 19.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 19.2 2.255 ;
      END
   END vdd

END no02s20

MACRO no02s10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 9.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 9.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 9.6 2.255 ;
      END
   END vdd

END no02s10

MACRO no02s08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4.8 2.255 ;
      END
   END vdd

END no02s08

MACRO no02s06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.6 2.255 ;
      END
   END vdd

END no02s06

MACRO no02s04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
   END vdd

END no02s04

MACRO no02s03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2 2.255 ;
      END
   END vdd

END no02s03

MACRO no02s02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
   END vdd

END no02s02

MACRO no02s01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 0.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 0.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 0.8 2.255 ;
      END
   END vdd

END no02s01

MACRO na04f80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 128 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 51.25 0.5 51.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 76.85 0.5 76.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 102.5 0.5 102.6 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 128 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 128 2.255 ;
      END
   END vdd

END na04f80

MACRO na04f40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 64 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 38.45 0.5 38.55 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 51.25 0.5 51.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 64 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 64 2.255 ;
      END
   END vdd

END na04f40

MACRO na04f20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 32 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 19.25 0.5 19.35 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 32 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 32 2.255 ;
      END
   END vdd

END na04f20

MACRO na04f10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 16 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 9.65 0.5 9.75 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 16 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 16 2.255 ;
      END
   END vdd

END na04f10

MACRO na04f08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 8 2.255 ;
      END
   END vdd

END na04f08

MACRO na04f06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.85 0.5 3.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.05 0.5 5.15 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6.4 2.255 ;
      END
   END vdd

END na04f06

MACRO na04f04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4 2.255 ;
      END
   END vdd

END na04f04

MACRO na04f03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.2 2.255 ;
      END
   END vdd

END na04f03

MACRO na04f02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.45 0.5 1.55 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
   END vdd

END na04f02

MACRO na04f01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.6 2.255 ;
      END
   END vdd

END na04f01

MACRO na04m80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 128 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 51.25 0.5 51.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 76.85 0.5 76.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 102.5 0.5 102.6 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 128 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 128 2.255 ;
      END
   END vdd

END na04m80

MACRO na04m40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 64 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 38.45 0.5 38.55 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 51.25 0.5 51.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 64 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 64 2.255 ;
      END
   END vdd

END na04m40

MACRO na04m20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 32 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 19.25 0.5 19.35 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 32 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 32 2.255 ;
      END
   END vdd

END na04m20

MACRO na04m10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 16 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 9.65 0.5 9.75 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 16 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 16 2.255 ;
      END
   END vdd

END na04m10

MACRO na04m08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 8 2.255 ;
      END
   END vdd

END na04m08

MACRO na04m06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.85 0.5 3.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.05 0.5 5.15 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6.4 2.255 ;
      END
   END vdd

END na04m06

MACRO na04m04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4 2.255 ;
      END
   END vdd

END na04m04

MACRO na04m03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.2 2.255 ;
      END
   END vdd

END na04m03

MACRO na04m02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.45 0.5 1.55 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
   END vdd

END na04m02

MACRO na04m01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.6 2.255 ;
      END
   END vdd

END na04m01

MACRO na04s80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 128 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 51.25 0.5 51.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 76.85 0.5 76.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 102.5 0.5 102.6 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 128 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 128 2.255 ;
      END
   END vdd

END na04s80

MACRO na04s40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 64 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 38.45 0.5 38.55 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 51.25 0.5 51.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 64 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 64 2.255 ;
      END
   END vdd

END na04s40

MACRO na04s20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 32 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 19.25 0.5 19.35 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 32 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 32 2.255 ;
      END
   END vdd

END na04s20

MACRO na04s10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 16 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 9.65 0.5 9.75 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 16 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 16 2.255 ;
      END
   END vdd

END na04s10

MACRO na04s08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 8 2.255 ;
      END
   END vdd

END na04s08

MACRO na04s06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.85 0.5 3.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.05 0.5 5.15 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6.4 2.255 ;
      END
   END vdd

END na04s06

MACRO na04s04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4 2.255 ;
      END
   END vdd

END na04s04

MACRO na04s03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.2 2.255 ;
      END
   END vdd

END na04s03

MACRO na04s02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.45 0.5 1.55 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
   END vdd

END na04s02

MACRO na04s01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.6 2.255 ;
      END
   END vdd

END na04s01

MACRO na03f80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 102.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 51.25 0.5 51.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 76.85 0.5 76.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 102.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 102.6 2.255 ;
      END
   END vdd

END na03f80

MACRO na03f40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 51.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.85 0.5 25.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 38.65 0.5 38.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.6 2.255 ;
      END
   END vdd

END na03f40

MACRO na03f20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 19.25 0.5 19.35 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.8 2.255 ;
      END
   END vdd

END na03f20

MACRO na03f10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 13.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.65 0.5 6.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 9.85 0.5 9.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 13.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 13.2 2.255 ;
      END
   END vdd

END na03f10

MACRO na03f08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6.6 2.255 ;
      END
   END vdd

END na03f08

MACRO na03f06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.65 0.5 3.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4.8 2.255 ;
      END
   END vdd

END na03f06

MACRO na03f04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.65 0.5 2.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.6 2.255 ;
      END
   END vdd

END na03f04

MACRO na03f03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
   END vdd

END na03f03

MACRO na03f02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.8 2.255 ;
      END
   END vdd

END na03f02

MACRO na03f01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
   END vdd

END na03f01

MACRO na03m80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 102.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 51.25 0.5 51.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 76.85 0.5 76.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 102.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 102.6 2.255 ;
      END
   END vdd

END na03m80

MACRO na03m40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 51.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.85 0.5 25.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 38.65 0.5 38.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.6 2.255 ;
      END
   END vdd

END na03m40

MACRO na03m20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 19.25 0.5 19.35 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.8 2.255 ;
      END
   END vdd

END na03m20

MACRO na03m10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 13.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.65 0.5 6.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 9.85 0.5 9.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 13.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 13.2 2.255 ;
      END
   END vdd

END na03m10

MACRO na03m08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6.6 2.255 ;
      END
   END vdd

END na03m08

MACRO na03m06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.65 0.5 3.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4.8 2.255 ;
      END
   END vdd

END na03m06

MACRO na03m04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.65 0.5 2.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.6 2.255 ;
      END
   END vdd

END na03m04

MACRO na03m03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
   END vdd

END na03m03

MACRO na03m02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.8 2.255 ;
      END
   END vdd

END na03m02

MACRO na03m01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
   END vdd

END na03m01

MACRO na03s80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 102.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 51.25 0.5 51.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 76.85 0.5 76.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 102.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 102.6 2.255 ;
      END
   END vdd

END na03s80

MACRO na03s40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 51.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.85 0.5 25.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 38.65 0.5 38.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.6 2.255 ;
      END
   END vdd

END na03s40

MACRO na03s20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 19.25 0.5 19.35 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.8 2.255 ;
      END
   END vdd

END na03s20

MACRO na03s10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 13.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.65 0.5 6.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 9.85 0.5 9.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 13.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 13.2 2.255 ;
      END
   END vdd

END na03s10

MACRO na03s08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6.6 2.255 ;
      END
   END vdd

END na03s08

MACRO na03s06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.65 0.5 3.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4.8 2.255 ;
      END
   END vdd

END na03s06

MACRO na03s04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.65 0.5 2.75 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.6 2.255 ;
      END
   END vdd

END na03s04

MACRO na03s03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
   END vdd

END na03s03

MACRO na03s02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.8 2.255 ;
      END
   END vdd

END na03s02

MACRO na03s01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
   END vdd

END na03s01

MACRO na02f80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 76.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 51.25 0.5 51.35 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 76.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 76.8 2.255 ;
      END
   END vdd

END na02f80

MACRO na02f40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 38.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 38.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 38.4 2.255 ;
      END
   END vdd

END na02f40

MACRO na02f20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 19.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 19.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 19.2 2.255 ;
      END
   END vdd

END na02f20

MACRO na02f10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 9.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 9.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 9.6 2.255 ;
      END
   END vdd

END na02f10

MACRO na02f08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4.8 2.255 ;
      END
   END vdd

END na02f08

MACRO na02f06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.6 2.255 ;
      END
   END vdd

END na02f06

MACRO na02f04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
   END vdd

END na02f04

MACRO na02f03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2 2.255 ;
      END
   END vdd

END na02f03

MACRO na02f02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
   END vdd

END na02f02

MACRO na02f01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 0.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 0.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 0.8 2.255 ;
      END
   END vdd

END na02f01

MACRO na02m80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 76.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 51.25 0.5 51.35 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 76.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 76.8 2.255 ;
      END
   END vdd

END na02m80

MACRO na02m40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 38.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 38.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 38.4 2.255 ;
      END
   END vdd

END na02m40

MACRO na02m20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 19.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 19.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 19.2 2.255 ;
      END
   END vdd

END na02m20

MACRO na02m10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 9.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 9.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 9.6 2.255 ;
      END
   END vdd

END na02m10

MACRO na02m08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4.8 2.255 ;
      END
   END vdd

END na02m08

MACRO na02m06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.6 2.255 ;
      END
   END vdd

END na02m06

MACRO na02m04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
   END vdd

END na02m04

MACRO na02m03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2 2.255 ;
      END
   END vdd

END na02m03

MACRO na02m02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
   END vdd

END na02m02

MACRO na02m01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 0.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 0.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 0.8 2.255 ;
      END
   END vdd

END na02m01

MACRO na02s80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 76.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 51.25 0.5 51.35 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 76.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 76.8 2.255 ;
      END
   END vdd

END na02s80

MACRO na02s40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 38.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 38.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 38.4 2.255 ;
      END
   END vdd

END na02s40

MACRO na02s20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 19.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 19.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 19.2 2.255 ;
      END
   END vdd

END na02s20

MACRO na02s10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 9.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 9.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 9.6 2.255 ;
      END
   END vdd

END na02s10

MACRO na02s08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4.8 2.255 ;
      END
   END vdd

END na02s08

MACRO na02s06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.6 2.255 ;
      END
   END vdd

END na02s06

MACRO na02s04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
   END vdd

END na02s04

MACRO na02s03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2 2.255 ;
      END
   END vdd

END na02s03

MACRO na02s02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
   END vdd

END na02s02

MACRO na02s01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 0.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 0.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 0.8 2.255 ;
      END
   END vdd

END na02s01

MACRO in01f80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 51.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.2 2.255 ;
      END
   END vdd

END in01f80

MACRO in01f40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.6 2.255 ;
      END
   END vdd

END in01f40

MACRO in01f20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
   END vdd

END in01f20

MACRO in01f10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6.4 2.255 ;
      END
   END vdd

END in01f10

MACRO in01f08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.2 2.255 ;
      END
   END vdd

END in01f08

MACRO in01f06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
   END vdd

END in01f06

MACRO in01f04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.6 2.255 ;
      END
   END vdd

END in01f04

MACRO in01f03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
   END vdd

END in01f03

MACRO in01f02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 0.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 0.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 0.8 2.255 ;
      END
   END vdd

END in01f02

MACRO in01f01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 0.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 0.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 0.4 2.255 ;
      END
   END vdd

END in01f01

MACRO in01m80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 51.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.2 2.255 ;
      END
   END vdd

END in01m80

MACRO in01m40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.6 2.255 ;
      END
   END vdd

END in01m40

MACRO in01m20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
   END vdd

END in01m20

MACRO in01m10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6.4 2.255 ;
      END
   END vdd

END in01m10

MACRO in01m08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.2 2.255 ;
      END
   END vdd

END in01m08

MACRO in01m06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
   END vdd

END in01m06

MACRO in01m04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.6 2.255 ;
      END
   END vdd

END in01m04

MACRO in01m03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
   END vdd

END in01m03

MACRO in01m02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 0.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 0.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 0.8 2.255 ;
      END
   END vdd

END in01m02

MACRO in01m01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 0.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 0.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 0.4 2.255 ;
      END
   END vdd

END in01m01

MACRO in01s80
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 51.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.2 2.255 ;
      END
   END vdd

END in01s80

MACRO in01s40
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.6 2.255 ;
      END
   END vdd

END in01s40

MACRO in01s20
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
   END vdd

END in01s20

MACRO in01s10
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6.4 2.255 ;
      END
   END vdd

END in01s10

MACRO in01s08
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.2 2.255 ;
      END
   END vdd

END in01s08

MACRO in01s06
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
   END vdd

END in01s06

MACRO in01s04
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.6 2.255 ;
      END
   END vdd

END in01s04

MACRO in01s03
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
   END vdd

END in01s03

MACRO in01s02
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 0.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 0.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 0.8 2.255 ;
      END
   END vdd

END in01s02

MACRO in01s01
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 0.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 0.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 0.4 2.255 ;
      END
   END vdd

END in01s01

MACRO in01f80X2HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 51.2 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 51.2 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.2 2.255 ;
      END
   END vdd

END in01f80X2HE

MACRO in01f80X2HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 51.2 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 51.2 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.2 2.255 ;
      END
   END vss

END in01f80X2HO

MACRO in01f80X3H
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 51.2 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 4.5 0.15 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 51.2 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.2 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 51.2 6.255 ;
      END
   END vdd

END in01f80X3H

MACRO in01f80X4HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 51.2 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 4.5 25.75 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 51.2 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 51.2 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.2 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 51.2 6.255 ;
      END
   END vdd

END in01f80X4HE

MACRO in01f80X4HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 51.2 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 4.5 25.75 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 51.2 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 51.2 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.2 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 51.2 6.255 ;
      END
   END vss

END in01f80X4HO

MACRO in01f40X2HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.6 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 25.6 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.6 2.255 ;
      END
   END vdd

END in01f40X2HE

MACRO in01f40X2HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.6 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 25.6 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.6 2.255 ;
      END
   END vss

END in01f40X2HO

MACRO in01f40X3H
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.6 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 4.5 0.15 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 25.6 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.6 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 25.6 6.255 ;
      END
   END vdd

END in01f40X3H

MACRO in01f40X4HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.6 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 4.5 12.95 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 25.6 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 25.6 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.6 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 25.6 6.255 ;
      END
   END vdd

END in01f40X4HE

MACRO in01f40X4HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.6 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 4.5 12.95 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 25.6 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 25.6 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.6 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 25.6 6.255 ;
      END
   END vss

END in01f40X4HO

MACRO in01f20X2HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 12.8 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
   END vdd

END in01f20X2HE

MACRO in01f20X2HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 12.8 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
   END vss

END in01f20X2HO

MACRO in01f20X3H
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 4.5 0.15 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 12.8 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 12.8 6.255 ;
      END
   END vdd

END in01f20X3H

MACRO in01f20X4HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 4.5 6.55 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 12.8 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 12.8 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 12.8 6.255 ;
      END
   END vdd

END in01f20X4HE

MACRO in01f20X4HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 4.5 6.55 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 12.8 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 12.8 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 12.8 6.255 ;
      END
   END vss

END in01f20X4HO

MACRO in01f10X2HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6.4 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6.4 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 6.4 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6.4 2.255 ;
      END
   END vdd

END in01f10X2HE

MACRO in01f10X2HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6.4 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6.4 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 6.4 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6.4 2.255 ;
      END
   END vss

END in01f10X2HO

MACRO in01f10X3H
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6.4 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 4.5 0.15 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6.4 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 6.4 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6.4 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 6.4 6.255 ;
      END
   END vdd

END in01f10X3H

MACRO in01f10X4HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 19.2 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 9.65 4.5 9.75 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 19.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 19.2 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 19.2 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 19.2 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 19.2 6.255 ;
      END
   END vdd

END in01f10X4HE

MACRO in01f10X4HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 4.5 6.55 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 12.8 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 12.8 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 12.8 6.255 ;
      END
   END vss

END in01f10X4HO

MACRO in01f08X2HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 9.6 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 9.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 9.6 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 9.6 2.255 ;
      END
   END vdd

END in01f08X2HE

MACRO in01f08X2HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 9.6 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 9.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 9.6 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 9.6 2.255 ;
      END
   END vss

END in01f08X2HO

MACRO in01f08X3H
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 4.5 4.95 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 12.8 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 12.8 6.255 ;
      END
   END vdd

END in01f08X3H

MACRO in01f08X4HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.6 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 11.25 0.5 11.35 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 4.5 12.95 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 25.6 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 25.6 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.6 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 25.6 6.255 ;
      END
   END vdd

END in01f08X4HE

MACRO in01f08X4HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 4.5 6.55 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 12.8 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 12.8 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 12.8 6.255 ;
      END
   END vss

END in01f08X4HO

MACRO in01f06X2HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 16.8 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 7.25 0.5 7.35 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 8.45 0.5 8.55 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 16.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 16.8 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 16.8 2.255 ;
      END
   END vdd

END in01f06X2HE

MACRO in01f06X2HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4.8 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 4.8 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4.8 2.255 ;
      END
   END vss

END in01f06X2HO

MACRO in01f06X3H
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 14.4 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.05 4.5 6.15 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 7.25 0.5 7.35 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 14.4 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 14.4 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 14.4 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 14.4 6.255 ;
      END
   END vdd

END in01f06X3H

MACRO in01f06X4HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 19.2 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 8.45 0.5 8.55 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 9.65 4.5 9.75 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 19.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 19.2 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 19.2 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 19.2 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 19.2 6.255 ;
      END
   END vdd

END in01f06X4HE

MACRO in01f06X4HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.05 4.5 6.15 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 12 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 12 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 12 6.255 ;
      END
   END vss

END in01f06X4HO

MACRO in01f04X2HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 9.6 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.05 0.5 4.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 9.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 9.6 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 9.6 2.255 ;
      END
   END vdd

END in01f04X2HE

MACRO in01f04X2HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.2 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 3.2 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.2 2.255 ;
      END
   END vss

END in01f04X2HO

MACRO in01f04X3H
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.65 4.5 5.75 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 12.8 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 12.8 6.255 ;
      END
   END vdd

END in01f04X3H

MACRO in01f04X4HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.2 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 4.5 1.75 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 3.2 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 3.2 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.2 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 3.2 6.255 ;
      END
   END vdd

END in01f04X4HE

MACRO in01f04X4HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.65 0.5 5.75 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 4.5 6.55 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 12.8 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 12.8 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 12.8 6.255 ;
      END
   END vss

END in01f04X4HO

MACRO in01f03X2HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.05 0.5 3.15 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 6 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6 2.255 ;
      END
   END vdd

END in01f03X2HE

MACRO in01f03X2HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.6 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 3.6 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.6 2.255 ;
      END
   END vss

END in01f03X2HO

MACRO in01f03X3H
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 8.4 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.65 4.5 3.75 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.25 0.5 4.35 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 8.4 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 8.4 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 8.4 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 8.4 6.255 ;
      END
   END vdd

END in01f03X3H

MACRO in01f03X4HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.6 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 4.5 1.95 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 3.6 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 3.6 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.6 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 3.6 6.255 ;
      END
   END vdd

END in01f03X4HE

MACRO in01f03X4HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.05 4.5 3.15 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 6 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 6 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 6 6.255 ;
      END
   END vss

END in01f03X4HO

MACRO in01f02X2HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.2 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 3.2 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.2 2.255 ;
      END
   END vdd

END in01f02X2HE

MACRO in01f02X2HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.2 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 3.2 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.2 2.255 ;
      END
   END vss

END in01f02X2HO

MACRO in01f02X3H
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6.4 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.85 4.5 2.95 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6.4 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 6.4 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6.4 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 6.4 6.255 ;
      END
   END vdd

END in01f02X3H

MACRO in01f02X4HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.6 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 4.5 0.95 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 1.6 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 1.6 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.6 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 1.6 6.255 ;
      END
   END vdd

END in01f02X4HE

MACRO in01f02X4HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.2 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 4.5 1.75 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 3.2 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 3.2 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.2 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 3.2 6.255 ;
      END
   END vss

END in01f02X4HO

MACRO in01f01X2HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.2 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.45 0.5 1.55 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 3.2 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.2 2.255 ;
      END
   END vdd

END in01f01X2HE

MACRO in01f01X2HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.6 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 1.6 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.6 2.255 ;
      END
   END vss

END in01f01X2HO

MACRO in01f01X3H
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.2 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.45 4.5 1.55 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 3.2 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.2 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 3.2 6.255 ;
      END
   END vdd

END in01f01X3H

MACRO in01f01X4HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.05 0.5 1.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 4.5 1.35 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 2.4 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 2.4 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 2.4 6.255 ;
      END
   END vdd

END in01f01X4HE

MACRO in01f01X4HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 0.8 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 4.5 0.55 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 0.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 0.8 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 0.8 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 0.8 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 0.8 6.255 ;
      END
   END vss

END in01f01X4HO

MACRO in01m80X2HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 51.2 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 51.2 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.2 2.255 ;
      END
   END vdd

END in01m80X2HE

MACRO in01m80X2HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 51.2 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 51.2 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.2 2.255 ;
      END
   END vss

END in01m80X2HO

MACRO in01m80X3H
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 51.2 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 4.5 0.15 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 51.2 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.2 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 51.2 6.255 ;
      END
   END vdd

END in01m80X3H

MACRO in01m80X4HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 51.2 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 4.5 25.75 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 51.2 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 51.2 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.2 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 51.2 6.255 ;
      END
   END vdd

END in01m80X4HE

MACRO in01m80X4HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 51.2 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 4.5 25.75 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 51.2 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 51.2 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.2 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 51.2 6.255 ;
      END
   END vss

END in01m80X4HO

MACRO in01m40X2HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.6 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 25.6 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.6 2.255 ;
      END
   END vdd

END in01m40X2HE

MACRO in01m40X2HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.6 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 25.6 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.6 2.255 ;
      END
   END vss

END in01m40X2HO

MACRO in01m40X3H
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.6 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 4.5 0.15 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 25.6 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.6 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 25.6 6.255 ;
      END
   END vdd

END in01m40X3H

MACRO in01m40X4HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.6 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 4.5 12.95 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 25.6 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 25.6 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.6 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 25.6 6.255 ;
      END
   END vdd

END in01m40X4HE

MACRO in01m40X4HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.6 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 4.5 12.95 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 25.6 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 25.6 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.6 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 25.6 6.255 ;
      END
   END vss

END in01m40X4HO

MACRO in01m20X2HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 12.8 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
   END vdd

END in01m20X2HE

MACRO in01m20X2HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 12.8 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
   END vss

END in01m20X2HO

MACRO in01m20X3H
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 4.5 0.15 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 12.8 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 12.8 6.255 ;
      END
   END vdd

END in01m20X3H

MACRO in01m20X4HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 4.5 6.55 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 12.8 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 12.8 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 12.8 6.255 ;
      END
   END vdd

END in01m20X4HE

MACRO in01m20X4HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 4.5 6.55 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 12.8 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 12.8 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 12.8 6.255 ;
      END
   END vss

END in01m20X4HO

MACRO in01m10X2HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6.4 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6.4 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 6.4 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6.4 2.255 ;
      END
   END vdd

END in01m10X2HE

MACRO in01m10X2HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6.4 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6.4 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 6.4 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6.4 2.255 ;
      END
   END vss

END in01m10X2HO

MACRO in01m10X3H
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6.4 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 4.5 0.15 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6.4 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 6.4 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6.4 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 6.4 6.255 ;
      END
   END vdd

END in01m10X3H

MACRO in01m10X4HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 19.2 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 9.65 4.5 9.75 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 19.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 19.2 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 19.2 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 19.2 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 19.2 6.255 ;
      END
   END vdd

END in01m10X4HE

MACRO in01m10X4HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.6 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 9.65 0.5 9.75 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 4.5 12.95 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 25.6 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 25.6 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.6 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 25.6 6.255 ;
      END
   END vss

END in01m10X4HO

MACRO in01m08X2HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 9.6 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 9.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 9.6 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 9.6 2.255 ;
      END
   END vdd

END in01m08X2HE

MACRO in01m08X2HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.6 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 11.25 0.5 11.35 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 25.6 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.6 2.255 ;
      END
   END vss

END in01m08X2HO

MACRO in01m08X3H
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6.4 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 4.5 1.75 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6.4 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 6.4 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6.4 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 6.4 6.255 ;
      END
   END vdd

END in01m08X3H

MACRO in01m08X4HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.6 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 11.25 0.5 11.35 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 4.5 12.95 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 25.6 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 25.6 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.6 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 25.6 6.255 ;
      END
   END vdd

END in01m08X4HE

MACRO in01m08X4HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 4.5 6.55 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 12.8 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 12.8 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 12.8 6.255 ;
      END
   END vss

END in01m08X4HO

MACRO in01m06X2HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.05 0.5 6.15 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 12 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12 2.255 ;
      END
   END vdd

END in01m06X2HE

MACRO in01m06X2HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4.8 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 4.8 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4.8 2.255 ;
      END
   END vss

END in01m06X2HO

MACRO in01m06X3H
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 9.6 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.65 4.5 3.75 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 9.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 9.6 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 9.6 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 9.6 6.255 ;
      END
   END vdd

END in01m06X3H

MACRO in01m06X4HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 9.6 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.65 0.5 3.75 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 4.5 4.95 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 9.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 9.6 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 9.6 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 9.6 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 9.6 6.255 ;
      END
   END vdd

END in01m06X4HE

MACRO in01m06X4HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 14.4 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.05 0.5 6.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 7.25 4.5 7.35 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 14.4 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 14.4 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 14.4 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 14.4 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 14.4 6.255 ;
      END
   END vss

END in01m06X4HO

MACRO in01m04X2HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.65 0.5 5.75 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 12.8 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
   END vdd

END in01m04X2HE

MACRO in01m04X2HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4.8 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 4.8 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4.8 2.255 ;
      END
   END vss

END in01m04X2HO

MACRO in01m04X3H
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 8 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 4.5 3.35 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.05 0.5 4.15 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 8 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 8 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 8 6.255 ;
      END
   END vdd

END in01m04X3H

MACRO in01m04X4HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.2 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 4.5 1.75 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 3.2 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 3.2 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.2 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 3.2 6.255 ;
      END
   END vdd

END in01m04X4HE

MACRO in01m04X4HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 9.6 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.05 0.5 4.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 4.5 4.95 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 9.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 9.6 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 9.6 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 9.6 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 9.6 6.255 ;
      END
   END vss

END in01m04X4HO

MACRO in01m03X2HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4.8 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 4.8 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4.8 2.255 ;
      END
   END vdd

END in01m03X2HE

MACRO in01m03X2HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.6 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 3.6 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.6 2.255 ;
      END
   END vss

END in01m03X2HO

MACRO in01m03X3H
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 7.2 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.05 4.5 3.15 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.65 0.5 3.75 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 7.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 7.2 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 7.2 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 7.2 6.255 ;
      END
   END vdd

END in01m03X3H

MACRO in01m03X4HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 4.5 1.35 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 2.4 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 2.4 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 2.4 6.255 ;
      END
   END vdd

END in01m03X4HE

MACRO in01m03X4HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 8.4 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.65 0.5 3.75 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.25 4.5 4.35 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 8.4 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 8.4 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 8.4 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 8.4 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 8.4 6.255 ;
      END
   END vss

END in01m03X4HO

MACRO in01m02X2HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.2 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 3.2 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.2 2.255 ;
      END
   END vdd

END in01m02X2HE

MACRO in01m02X2HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.05 0.5 2.15 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 4 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4 2.255 ;
      END
   END vss

END in01m02X2HO

MACRO in01m02X3H
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 4.5 0.95 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 2.4 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 2.4 6.255 ;
      END
   END vdd

END in01m02X3H

MACRO in01m02X4HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4.8 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.05 0.5 2.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 4.5 2.55 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 4.8 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 4.8 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4.8 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 4.8 6.255 ;
      END
   END vdd

END in01m02X4HE

MACRO in01m02X4HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.6 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 4.5 0.95 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 1.6 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 1.6 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.6 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 1.6 6.255 ;
      END
   END vss

END in01m02X4HO

MACRO in01m01X2HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 0.8 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 0.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 0.8 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 0.8 2.255 ;
      END
   END vdd

END in01m01X2HE

MACRO in01m01X2HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.05 0.5 1.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 2.4 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
   END vss

END in01m01X2HO

MACRO in01m01X3H
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.05 4.5 1.15 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 2.4 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 2.4 6.255 ;
      END
   END vdd

END in01m01X3H

MACRO in01m01X4HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.2 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 4.5 0.75 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 1.2 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 1.2 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 1.2 6.255 ;
      END
   END vdd

END in01m01X4HE

MACRO in01m01X4HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.8 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.45 4.5 1.55 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 2.8 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 2.8 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.8 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 2.8 6.255 ;
      END
   END vss

END in01m01X4HO

MACRO in01s80X2HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 51.2 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 51.2 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.2 2.255 ;
      END
   END vdd

END in01s80X2HE

MACRO in01s80X2HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 51.2 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 51.2 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.2 2.255 ;
      END
   END vss

END in01s80X2HO

MACRO in01s80X3H
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 51.2 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 4.5 0.15 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 0.5 25.75 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 51.2 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.2 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 51.2 6.255 ;
      END
   END vdd

END in01s80X3H

MACRO in01s80X4HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 51.2 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 4.5 25.75 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 51.2 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 51.2 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.2 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 51.2 6.255 ;
      END
   END vdd

END in01s80X4HE

MACRO in01s80X4HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 51.2 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 25.65 4.5 25.75 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 51.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 51.2 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 51.2 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 51.2 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 51.2 6.255 ;
      END
   END vss

END in01s80X4HO

MACRO in01s40X2HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.6 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 25.6 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.6 2.255 ;
      END
   END vdd

END in01s40X2HE

MACRO in01s40X2HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.6 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 25.6 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.6 2.255 ;
      END
   END vss

END in01s40X2HO

MACRO in01s40X3H
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.6 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 4.5 0.15 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 25.6 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.6 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 25.6 6.255 ;
      END
   END vdd

END in01s40X3H

MACRO in01s40X4HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.6 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 4.5 12.95 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 25.6 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 25.6 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.6 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 25.6 6.255 ;
      END
   END vdd

END in01s40X4HE

MACRO in01s40X4HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.6 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 4.5 12.95 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 25.6 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 25.6 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.6 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 25.6 6.255 ;
      END
   END vss

END in01s40X4HO

MACRO in01s20X2HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 12.8 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
   END vdd

END in01s20X2HE

MACRO in01s20X2HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 12.8 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
   END vss

END in01s20X2HO

MACRO in01s20X3H
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 4.5 0.15 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 12.8 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 12.8 6.255 ;
      END
   END vdd

END in01s20X3H

MACRO in01s20X4HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 4.5 6.55 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 12.8 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 12.8 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 12.8 6.255 ;
      END
   END vdd

END in01s20X4HE

MACRO in01s20X4HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 4.5 6.55 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 12.8 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 12.8 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 12.8 6.255 ;
      END
   END vss

END in01s20X4HO

MACRO in01s10X2HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6.4 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6.4 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 6.4 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6.4 2.255 ;
      END
   END vdd

END in01s10X2HE

MACRO in01s10X2HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6.4 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6.4 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 6.4 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6.4 2.255 ;
      END
   END vss

END in01s10X2HO

MACRO in01s10X3H
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 6.4 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 4.5 0.15 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 6.4 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 6.4 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 6.4 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 6.4 6.255 ;
      END
   END vdd

END in01s10X3H

MACRO in01s10X4HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 4.5 6.55 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 12.8 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 12.8 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 12.8 6.255 ;
      END
   END vdd

END in01s10X4HE

MACRO in01s10X4HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 32 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 16.05 4.5 16.15 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 32 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 32 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 32 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 32 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 32 6.255 ;
      END
   END vss

END in01s10X4HO

MACRO in01s08X2HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 12.8 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
   END vdd

END in01s08X2HE

MACRO in01s08X2HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.6 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 11.25 0.5 11.35 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 0.5 12.95 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 25.6 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.6 2.255 ;
      END
   END vss

END in01s08X2HO

MACRO in01s08X3H
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 22.4 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 9.65 4.5 9.75 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 11.25 0.5 11.35 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 22.4 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 22.4 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 22.4 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 22.4 6.255 ;
      END
   END vdd

END in01s08X3H

MACRO in01s08X4HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 25.6 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 11.25 0.5 11.35 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 12.85 4.5 12.95 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 25.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 25.6 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 25.6 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 25.6 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 25.6 6.255 ;
      END
   END vdd

END in01s08X4HE

MACRO in01s08X4HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 16 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 0.5 6.55 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 8.05 4.5 8.15 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 16 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 16 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 16 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 16 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 16 6.255 ;
      END
   END vss

END in01s08X4HO

MACRO in01s06X2HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 9.6 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.65 0.5 3.75 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 9.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 9.6 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 9.6 2.255 ;
      END
   END vdd

END in01s06X2HE

MACRO in01s06X2HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 7.2 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.65 0.5 3.75 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 7.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 7.2 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 7.2 2.255 ;
      END
   END vss

END in01s06X2HO

MACRO in01s06X3H
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 16.8 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 7.25 4.5 7.35 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 8.45 0.5 8.55 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 16.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 16.8 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 16.8 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 16.8 6.255 ;
      END
   END vdd

END in01s06X3H

MACRO in01s06X4HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 16.8 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 7.25 0.5 7.35 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 8.45 4.5 8.55 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 16.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 16.8 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 16.8 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 16.8 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 16.8 6.255 ;
      END
   END vdd

END in01s06X4HE

MACRO in01s06X4HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4.8 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 4.5 2.55 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 4.8 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 4.8 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4.8 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 4.8 6.255 ;
      END
   END vss

END in01s06X4HO

MACRO in01s04X2HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 8 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.25 0.5 3.35 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.05 0.5 4.15 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 8 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 8 2.255 ;
      END
   END vdd

END in01s04X2HE

MACRO in01s04X2HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 11.2 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 0.5 4.95 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.65 0.5 5.75 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 11.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 11.2 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 11.2 2.255 ;
      END
   END vss

END in01s04X2HO

MACRO in01s04X3H
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 11.2 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 4.85 4.5 4.95 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.65 0.5 5.75 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 11.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 11.2 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 11.2 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 11.2 6.255 ;
      END
   END vdd

END in01s04X3H

MACRO in01s04X4HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 12.8 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 5.65 0.5 5.75 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 6.45 4.5 6.55 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 12.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 12.8 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 12.8 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 12.8 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 12.8 6.255 ;
      END
   END vdd

END in01s04X4HE

MACRO in01s04X4HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.2 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 4.5 1.75 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 3.2 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 3.2 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.2 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 3.2 6.255 ;
      END
   END vss

END in01s04X4HO

MACRO in01s03X2HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 2.4 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
   END vdd

END in01s03X2HE

MACRO in01s03X2HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 7.2 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.05 0.5 3.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 3.65 0.5 3.75 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 7.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 7.2 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 7.2 2.255 ;
      END
   END vss

END in01s03X2HO

MACRO in01s03X3H
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 4.5 0.75 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 2.4 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 2.4 6.255 ;
      END
   END vdd

END in01s03X3H

MACRO in01s03X4HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.6 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 4.5 1.95 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 3.6 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 3.6 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.6 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 3.6 6.255 ;
      END
   END vdd

END in01s03X4HE

MACRO in01s03X4HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.6 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 4.5 1.95 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 3.6 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 3.6 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.6 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 3.6 6.255 ;
      END
   END vss

END in01s03X4HO

MACRO in01s02X2HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.6 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 1.6 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.6 2.255 ;
      END
   END vdd

END in01s02X2HE

MACRO in01s02X2HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 4 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.05 0.5 2.15 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 4 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 4 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 4 2.255 ;
      END
   END vss

END in01s02X2HO

MACRO in01s02X3H
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 4.5 0.95 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 2.4 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 2.4 6.255 ;
      END
   END vdd

END in01s02X3H

MACRO in01s02X4HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 5.6 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.45 0.5 2.55 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 2.85 4.5 2.95 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 5.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 5.6 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 5.6 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 5.6 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 5.6 6.255 ;
      END
   END vdd

END in01s02X4HE

MACRO in01s02X4HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 3.2 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 4.5 1.75 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 3.2 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 3.2 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.2 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 3.2 6.255 ;
      END
   END vss

END in01s02X4HO

MACRO in01s01X2HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 2.4 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.05 0.5 1.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 2.4 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 2.4 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 2.4 2.255 ;
      END
   END vdd

END in01s01X2HE

MACRO in01s01X2HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.2 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 1.2 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
   END vss

END in01s01X2HO

MACRO in01s01X3H
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 0.8 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 4.5 0.35 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 0.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 0.8 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 0.8 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 0.8 6.255 ;
      END
   END vdd

END in01s01X3H

MACRO in01s01X4HE
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 1.2 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 4.5 0.75 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 1.2 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 1.2 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 1.2 6.255 ;
      END
   END vdd

END in01s01X4HE

MACRO in01s01X4HO
   PROPERTY LEF58_EDGETYPE "
    EDGETYPE LEFT 2 ;
    EDGETYPE RIGHT 2 ;
  " ;
   CLASS CORE ;
   SIZE 0.8 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 4.5 0.55 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 0.8 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 0.8 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 0.8 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 0.8 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 0.8 6.255 ;
      END
   END vss

END in01s01X4HO

END LIBRARY
