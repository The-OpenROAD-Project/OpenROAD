module gcd (clk,
    req_rdy,
    req_val,
    reset,
    resp_rdy,
    resp_val,
    req_msg,
    resp_msg);
 input clk;
 output req_rdy;
 input req_val;
 input reset;
 input resp_rdy;
 output resp_val;
 input [31:0] req_msg;
 output [15:0] resp_msg;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _127_;
 wire _128_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _142_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire \ctrl.state.out[1] ;
 wire \ctrl.state.out[2] ;
 wire \dpath.a_lt_b$in0[0] ;
 wire \dpath.a_lt_b$in0[10] ;
 wire \dpath.a_lt_b$in0[11] ;
 wire \dpath.a_lt_b$in0[12] ;
 wire \dpath.a_lt_b$in0[13] ;
 wire \dpath.a_lt_b$in0[14] ;
 wire \dpath.a_lt_b$in0[15] ;
 wire \dpath.a_lt_b$in0[1] ;
 wire \dpath.a_lt_b$in0[2] ;
 wire \dpath.a_lt_b$in0[3] ;
 wire \dpath.a_lt_b$in0[4] ;
 wire \dpath.a_lt_b$in0[5] ;
 wire \dpath.a_lt_b$in0[6] ;
 wire \dpath.a_lt_b$in0[7] ;
 wire \dpath.a_lt_b$in0[8] ;
 wire \dpath.a_lt_b$in0[9] ;
 wire \dpath.a_lt_b$in1[0] ;
 wire \dpath.a_lt_b$in1[10] ;
 wire \dpath.a_lt_b$in1[11] ;
 wire \dpath.a_lt_b$in1[12] ;
 wire \dpath.a_lt_b$in1[13] ;
 wire \dpath.a_lt_b$in1[14] ;
 wire \dpath.a_lt_b$in1[15] ;
 wire \dpath.a_lt_b$in1[1] ;
 wire \dpath.a_lt_b$in1[2] ;
 wire \dpath.a_lt_b$in1[3] ;
 wire \dpath.a_lt_b$in1[4] ;
 wire \dpath.a_lt_b$in1[5] ;
 wire \dpath.a_lt_b$in1[6] ;
 wire \dpath.a_lt_b$in1[7] ;
 wire \dpath.a_lt_b$in1[8] ;
 wire \dpath.a_lt_b$in1[9] ;
 wire nPWRUP;

 sky130_fd_sc_hd__xnor2_1 _247_ (.A(\dpath.a_lt_b$in1[8] ),
    .B(\dpath.a_lt_b$in0[8] ),
    .Y(_035_));
 sky130_fd_sc_hd__and2b_1 _248_ (.A_N(\dpath.a_lt_b$in0[10] ),
    .B(\dpath.a_lt_b$in1[10] ),
    .X(_036_));
 sky130_fd_sc_hd__nand2b_1 _249_ (.A_N(\dpath.a_lt_b$in1[10] ),
    .B(\dpath.a_lt_b$in0[10] ),
    .Y(_037_));
 sky130_fd_sc_hd__nor2b_1 _250_ (.A(_036_),
    .B_N(_037_),
    .Y(_038_));
 sky130_fd_sc_hd__nor2b_1 _251_ (.A(\dpath.a_lt_b$in1[11] ),
    .B_N(\dpath.a_lt_b$in0[11] ),
    .Y(_039_));
 sky130_fd_sc_hd__nand2b_1 _252_ (.A_N(\dpath.a_lt_b$in0[11] ),
    .B(\dpath.a_lt_b$in1[11] ),
    .Y(_040_));
 sky130_fd_sc_hd__nor2b_1 _253_ (.A(_039_),
    .B_N(_040_),
    .Y(_041_));
 sky130_fd_sc_hd__nand2b_1 _254_ (.A_N(\dpath.a_lt_b$in1[9] ),
    .B(\dpath.a_lt_b$in0[9] ),
    .Y(_042_));
 sky130_fd_sc_hd__nand2b_1 _255_ (.A_N(\dpath.a_lt_b$in0[9] ),
    .B(\dpath.a_lt_b$in1[9] ),
    .Y(_043_));
 sky130_fd_sc_hd__and2_1 _256_ (.A(_042_),
    .B(_043_),
    .X(_044_));
 sky130_fd_sc_hd__and4_1 _257_ (.A(_035_),
    .B(_038_),
    .C(_041_),
    .D(_044_),
    .X(_045_));
 sky130_fd_sc_hd__xor2_1 _258_ (.A(\dpath.a_lt_b$in1[4] ),
    .B(\dpath.a_lt_b$in0[4] ),
    .X(_046_));
 sky130_fd_sc_hd__xor2_1 _259_ (.A(\dpath.a_lt_b$in1[5] ),
    .B(\dpath.a_lt_b$in0[5] ),
    .X(_047_));
 sky130_fd_sc_hd__xor2_1 _261_ (.A(\dpath.a_lt_b$in1[6] ),
    .B(\dpath.a_lt_b$in0[6] ),
    .X(_049_));
 sky130_fd_sc_hd__xor2_1 _262_ (.A(\dpath.a_lt_b$in1[7] ),
    .B(\dpath.a_lt_b$in0[7] ),
    .X(_050_));
 sky130_fd_sc_hd__nor4_2 _263_ (.A(_046_),
    .B(_047_),
    .C(_049_),
    .D(_050_),
    .Y(_051_));
 sky130_fd_sc_hd__inv_1 _264_ (.A(\dpath.a_lt_b$in0[0] ),
    .Y(_052_));
 sky130_fd_sc_hd__nand2b_1 _266_ (.A_N(\dpath.a_lt_b$in1[1] ),
    .B(\dpath.a_lt_b$in0[1] ),
    .Y(_054_));
 sky130_fd_sc_hd__nor2b_1 _267_ (.A(\dpath.a_lt_b$in0[1] ),
    .B_N(\dpath.a_lt_b$in1[1] ),
    .Y(_055_));
 sky130_fd_sc_hd__a31oi_1 _268_ (.A1(_052_),
    .A2(\dpath.a_lt_b$in1[0] ),
    .A3(_054_),
    .B1(_055_),
    .Y(_056_));
 sky130_fd_sc_hd__nor2b_1 _269_ (.A(\dpath.a_lt_b$in1[2] ),
    .B_N(\dpath.a_lt_b$in0[2] ),
    .Y(_057_));
 sky130_fd_sc_hd__nor2b_1 _270_ (.A(\dpath.a_lt_b$in0[2] ),
    .B_N(\dpath.a_lt_b$in1[2] ),
    .Y(_058_));
 sky130_fd_sc_hd__nand2b_1 _271_ (.A_N(\dpath.a_lt_b$in0[3] ),
    .B(_058_),
    .Y(_059_));
 sky130_fd_sc_hd__inv_1 _272_ (.A(\dpath.a_lt_b$in1[3] ),
    .Y(_060_));
 sky130_fd_sc_hd__o311ai_2 _273_ (.A1(\dpath.a_lt_b$in0[3] ),
    .A2(_056_),
    .A3(_057_),
    .B1(_059_),
    .C1(_060_),
    .Y(_061_));
 sky130_fd_sc_hd__a311oi_2 _274_ (.A1(_052_),
    .A2(\dpath.a_lt_b$in1[0] ),
    .A3(_054_),
    .B1(_055_),
    .C1(_058_),
    .Y(_062_));
 sky130_fd_sc_hd__o21ai_1 _275_ (.A1(_057_),
    .A2(_062_),
    .B1(\dpath.a_lt_b$in0[3] ),
    .Y(_063_));
 sky130_fd_sc_hd__nand2_4 _276_ (.A(_061_),
    .B(_063_),
    .Y(_064_));
 sky130_fd_sc_hd__inv_1 _277_ (.A(\dpath.a_lt_b$in1[8] ),
    .Y(_065_));
 sky130_fd_sc_hd__inv_1 _278_ (.A(\dpath.a_lt_b$in0[9] ),
    .Y(_066_));
 sky130_fd_sc_hd__a21oi_1 _279_ (.A1(\dpath.a_lt_b$in1[9] ),
    .A2(_066_),
    .B1(_036_),
    .Y(_067_));
 sky130_fd_sc_hd__o21ai_0 _280_ (.A1(_042_),
    .A2(_036_),
    .B1(_037_),
    .Y(_068_));
 sky130_fd_sc_hd__a31o_2 _281_ (.A1(_065_),
    .A2(\dpath.a_lt_b$in0[8] ),
    .A3(_067_),
    .B1(_068_),
    .X(_069_));
 sky130_fd_sc_hd__nor2b_1 _282_ (.A(\dpath.a_lt_b$in1[7] ),
    .B_N(\dpath.a_lt_b$in0[7] ),
    .Y(_070_));
 sky130_fd_sc_hd__inv_1 _283_ (.A(\dpath.a_lt_b$in0[7] ),
    .Y(_071_));
 sky130_fd_sc_hd__inv_1 _284_ (.A(\dpath.a_lt_b$in0[6] ),
    .Y(_072_));
 sky130_fd_sc_hd__a22oi_1 _285_ (.A1(\dpath.a_lt_b$in1[7] ),
    .A2(_071_),
    .B1(_072_),
    .B2(\dpath.a_lt_b$in1[6] ),
    .Y(_073_));
 sky130_fd_sc_hd__nand2b_1 _286_ (.A_N(\dpath.a_lt_b$in1[6] ),
    .B(\dpath.a_lt_b$in0[6] ),
    .Y(_074_));
 sky130_fd_sc_hd__nand2b_1 _287_ (.A_N(\dpath.a_lt_b$in0[5] ),
    .B(\dpath.a_lt_b$in1[5] ),
    .Y(_075_));
 sky130_fd_sc_hd__nor2b_1 _288_ (.A(\dpath.a_lt_b$in1[4] ),
    .B_N(\dpath.a_lt_b$in0[4] ),
    .Y(_076_));
 sky130_fd_sc_hd__nor2b_1 _289_ (.A(\dpath.a_lt_b$in1[5] ),
    .B_N(\dpath.a_lt_b$in0[5] ),
    .Y(_077_));
 sky130_fd_sc_hd__a211oi_1 _290_ (.A1(_075_),
    .A2(_076_),
    .B1(_077_),
    .C1(_070_),
    .Y(_078_));
 sky130_fd_sc_hd__a2bb2oi_1 _291_ (.A1_N(_070_),
    .A2_N(_073_),
    .B1(_074_),
    .B2(_078_),
    .Y(_079_));
 sky130_fd_sc_hd__a221o_1 _292_ (.A1(_040_),
    .A2(_069_),
    .B1(_045_),
    .B2(_079_),
    .C1(_039_),
    .X(_080_));
 sky130_fd_sc_hd__a31oi_4 _293_ (.A1(_045_),
    .A2(_051_),
    .A3(_064_),
    .B1(_080_),
    .Y(_081_));
 sky130_fd_sc_hd__xor2_1 _294_ (.A(\dpath.a_lt_b$in1[13] ),
    .B(\dpath.a_lt_b$in0[13] ),
    .X(_082_));
 sky130_fd_sc_hd__xnor2_1 _295_ (.A(\dpath.a_lt_b$in1[14] ),
    .B(\dpath.a_lt_b$in0[14] ),
    .Y(_083_));
 sky130_fd_sc_hd__xnor2_1 _296_ (.A(\dpath.a_lt_b$in1[12] ),
    .B(\dpath.a_lt_b$in0[12] ),
    .Y(_084_));
 sky130_fd_sc_hd__nand2_1 _297_ (.A(_083_),
    .B(_084_),
    .Y(_085_));
 sky130_fd_sc_hd__inv_1 _298_ (.A(\dpath.a_lt_b$in0[14] ),
    .Y(_086_));
 sky130_fd_sc_hd__inv_1 _299_ (.A(\dpath.a_lt_b$in0[12] ),
    .Y(_087_));
 sky130_fd_sc_hd__nor2b_1 _300_ (.A(\dpath.a_lt_b$in0[13] ),
    .B_N(\dpath.a_lt_b$in1[13] ),
    .Y(_088_));
 sky130_fd_sc_hd__nand2b_1 _301_ (.A_N(\dpath.a_lt_b$in1[13] ),
    .B(\dpath.a_lt_b$in0[13] ),
    .Y(_089_));
 sky130_fd_sc_hd__o31a_1 _302_ (.A1(\dpath.a_lt_b$in1[12] ),
    .A2(_087_),
    .A3(_088_),
    .B1(_089_),
    .X(_090_));
 sky130_fd_sc_hd__maj3_1 _303_ (.A(\dpath.a_lt_b$in1[14] ),
    .B(_086_),
    .C(_090_),
    .X(_091_));
 sky130_fd_sc_hd__o31ai_1 _304_ (.A1(_081_),
    .A2(_082_),
    .A3(_085_),
    .B1(_091_),
    .Y(_092_));
 sky130_fd_sc_hd__xor2_1 _305_ (.A(\dpath.a_lt_b$in1[15] ),
    .B(\dpath.a_lt_b$in0[15] ),
    .X(_093_));
 sky130_fd_sc_hd__xnor2_1 _306_ (.A(_092_),
    .B(_093_),
    .Y(resp_msg[15]));
 sky130_fd_sc_hd__nand2_1 _307_ (.A(_052_),
    .B(\dpath.a_lt_b$in1[0] ),
    .Y(_094_));
 sky130_fd_sc_hd__xor2_1 _308_ (.A(\dpath.a_lt_b$in1[1] ),
    .B(\dpath.a_lt_b$in0[1] ),
    .X(_095_));
 sky130_fd_sc_hd__xnor2_1 _309_ (.A(_094_),
    .B(_095_),
    .Y(resp_msg[1]));
 sky130_fd_sc_hd__nor2_1 _310_ (.A(_057_),
    .B(_058_),
    .Y(_096_));
 sky130_fd_sc_hd__xor2_1 _311_ (.A(_056_),
    .B(_096_),
    .X(resp_msg[2]));
 sky130_fd_sc_hd__xor2_1 _312_ (.A(\dpath.a_lt_b$in1[3] ),
    .B(\dpath.a_lt_b$in0[3] ),
    .X(_097_));
 sky130_fd_sc_hd__o21ai_0 _313_ (.A1(_057_),
    .A2(_062_),
    .B1(_097_),
    .Y(_098_));
 sky130_fd_sc_hd__or3_1 _314_ (.A(_057_),
    .B(_062_),
    .C(_097_),
    .X(_099_));
 sky130_fd_sc_hd__nand2_1 _315_ (.A(_098_),
    .B(_099_),
    .Y(resp_msg[3]));
 sky130_fd_sc_hd__xnor2_1 _316_ (.A(_046_),
    .B(_064_),
    .Y(resp_msg[4]));
 sky130_fd_sc_hd__inv_1 _317_ (.A(\dpath.a_lt_b$in1[4] ),
    .Y(_100_));
 sky130_fd_sc_hd__maj3_1 _318_ (.A(_100_),
    .B(\dpath.a_lt_b$in0[4] ),
    .C(_064_),
    .X(_101_));
 sky130_fd_sc_hd__xnor2_1 _319_ (.A(_047_),
    .B(_101_),
    .Y(resp_msg[5]));
 sky130_fd_sc_hd__nand2_1 _320_ (.A(\dpath.a_lt_b$in0[4] ),
    .B(_075_),
    .Y(_102_));
 sky130_fd_sc_hd__a21oi_1 _321_ (.A1(_061_),
    .A2(_063_),
    .B1(_102_),
    .Y(_103_));
 sky130_fd_sc_hd__a21o_1 _322_ (.A1(_075_),
    .A2(_076_),
    .B1(_077_),
    .X(_104_));
 sky130_fd_sc_hd__a311oi_2 _323_ (.A1(_100_),
    .A2(_075_),
    .A3(_064_),
    .B1(_103_),
    .C1(_104_),
    .Y(_105_));
 sky130_fd_sc_hd__xor2_1 _324_ (.A(_049_),
    .B(_105_),
    .X(resp_msg[6]));
 sky130_fd_sc_hd__maj3_1 _325_ (.A(\dpath.a_lt_b$in1[6] ),
    .B(_072_),
    .C(_105_),
    .X(_106_));
 sky130_fd_sc_hd__xor2_1 _326_ (.A(_050_),
    .B(_106_),
    .X(resp_msg[7]));
 sky130_fd_sc_hd__a21oi_1 _327_ (.A1(_051_),
    .A2(_064_),
    .B1(_079_),
    .Y(_107_));
 sky130_fd_sc_hd__xnor2_1 _328_ (.A(_035_),
    .B(_107_),
    .Y(resp_msg[8]));
 sky130_fd_sc_hd__nand2_1 _329_ (.A(\dpath.a_lt_b$in0[8] ),
    .B(_051_),
    .Y(_108_));
 sky130_fd_sc_hd__a21oi_1 _330_ (.A1(_061_),
    .A2(_063_),
    .B1(_108_),
    .Y(_109_));
 sky130_fd_sc_hd__nand2_1 _331_ (.A(_065_),
    .B(_051_),
    .Y(_110_));
 sky130_fd_sc_hd__a21oi_1 _332_ (.A1(_061_),
    .A2(_063_),
    .B1(_110_),
    .Y(_111_));
 sky130_fd_sc_hd__maj3_1 _333_ (.A(_065_),
    .B(\dpath.a_lt_b$in0[8] ),
    .C(_079_),
    .X(_112_));
 sky130_fd_sc_hd__nor3_2 _334_ (.A(_109_),
    .B(_111_),
    .C(_112_),
    .Y(_113_));
 sky130_fd_sc_hd__xnor2_1 _335_ (.A(_044_),
    .B(_113_),
    .Y(resp_msg[9]));
 sky130_fd_sc_hd__o31ai_1 _336_ (.A1(_109_),
    .A2(_111_),
    .A3(_112_),
    .B1(_043_),
    .Y(_114_));
 sky130_fd_sc_hd__and2_1 _337_ (.A(_042_),
    .B(_114_),
    .X(_115_));
 sky130_fd_sc_hd__xnor2_1 _338_ (.A(_038_),
    .B(_115_),
    .Y(resp_msg[10]));
 sky130_fd_sc_hd__o21ai_0 _339_ (.A1(_036_),
    .A2(_115_),
    .B1(_037_),
    .Y(_116_));
 sky130_fd_sc_hd__xor2_1 _340_ (.A(_041_),
    .B(_116_),
    .X(resp_msg[11]));
 sky130_fd_sc_hd__xnor2_1 _341_ (.A(_081_),
    .B(_084_),
    .Y(resp_msg[12]));
 sky130_fd_sc_hd__maj3_1 _342_ (.A(\dpath.a_lt_b$in1[12] ),
    .B(_087_),
    .C(_081_),
    .X(_117_));
 sky130_fd_sc_hd__xor2_1 _343_ (.A(_082_),
    .B(_117_),
    .X(resp_msg[13]));
 sky130_fd_sc_hd__a21oi_1 _344_ (.A1(_089_),
    .A2(_117_),
    .B1(_088_),
    .Y(_118_));
 sky130_fd_sc_hd__xor2_1 _345_ (.A(_083_),
    .B(_118_),
    .X(resp_msg[14]));
 sky130_fd_sc_hd__xor2_1 _346_ (.A(\dpath.a_lt_b$in0[0] ),
    .B(\dpath.a_lt_b$in1[0] ),
    .X(resp_msg[0]));
 sky130_fd_sc_hd__nor4_1 _349_ (.A(\dpath.a_lt_b$in1[10] ),
    .B(\dpath.a_lt_b$in1[11] ),
    .C(\dpath.a_lt_b$in1[12] ),
    .D(\dpath.a_lt_b$in1[1] ),
    .Y(_121_));
 sky130_fd_sc_hd__nor4_1 _350_ (.A(\dpath.a_lt_b$in1[13] ),
    .B(\dpath.a_lt_b$in1[14] ),
    .C(\dpath.a_lt_b$in1[15] ),
    .D(\dpath.a_lt_b$in1[0] ),
    .Y(_122_));
 sky130_fd_sc_hd__nor4_1 _351_ (.A(\dpath.a_lt_b$in1[2] ),
    .B(\dpath.a_lt_b$in1[3] ),
    .C(\dpath.a_lt_b$in1[4] ),
    .D(\dpath.a_lt_b$in1[9] ),
    .Y(_123_));
 sky130_fd_sc_hd__nor4_1 _352_ (.A(\dpath.a_lt_b$in1[5] ),
    .B(\dpath.a_lt_b$in1[6] ),
    .C(\dpath.a_lt_b$in1[7] ),
    .D(\dpath.a_lt_b$in1[8] ),
    .Y(_124_));
 sky130_fd_sc_hd__nand4_1 _353_ (.A(_121_),
    .B(_122_),
    .C(_123_),
    .D(_124_),
    .Y(_125_));
 sky130_fd_sc_hd__a22oi_1 _355_ (.A1(req_rdy),
    .A2(req_val),
    .B1(_125_),
    .B2(\ctrl.state.out[2] ),
    .Y(_127_));
 sky130_fd_sc_hd__nor2_1 _356_ (.A(reset),
    .B(_127_),
    .Y(_002_));
 sky130_fd_sc_hd__inv_1 _357_ (.A(\ctrl.state.out[1] ),
    .Y(_128_));
 sky130_fd_sc_hd__nor3_1 _358_ (.A(\ctrl.state.out[2] ),
    .B(req_rdy),
    .C(_128_),
    .Y(resp_val));
 sky130_fd_sc_hd__inv_1 _360_ (.A(req_val),
    .Y(_130_));
 sky130_fd_sc_hd__a221o_1 _361_ (.A1(req_rdy),
    .A2(_130_),
    .B1(resp_rdy),
    .B2(resp_val),
    .C1(reset),
    .X(_000_));
 sky130_fd_sc_hd__inv_1 _362_ (.A(req_rdy),
    .Y(_131_));
 sky130_fd_sc_hd__a21o_1 _363_ (.A1(_131_),
    .A2(resp_rdy),
    .B1(_128_),
    .X(_132_));
 sky130_fd_sc_hd__inv_1 _364_ (.A(\ctrl.state.out[2] ),
    .Y(_133_));
 sky130_fd_sc_hd__a21o_1 _365_ (.A1(_128_),
    .A2(_125_),
    .B1(_133_),
    .X(_134_));
 sky130_fd_sc_hd__a21oi_1 _366_ (.A1(_132_),
    .A2(_134_),
    .B1(reset),
    .Y(_001_));
 sky130_fd_sc_hd__inv_1 _368_ (.A(\dpath.a_lt_b$in0[15] ),
    .Y(_136_));
 sky130_fd_sc_hd__or3_1 _369_ (.A(_136_),
    .B(_082_),
    .C(_085_),
    .X(_137_));
 sky130_fd_sc_hd__o221ai_2 _370_ (.A1(_136_),
    .A2(_091_),
    .B1(_137_),
    .B2(_081_),
    .C1(\dpath.a_lt_b$in1[15] ),
    .Y(_138_));
 sky130_fd_sc_hd__o311ai_4 _371_ (.A1(_081_),
    .A2(_082_),
    .A3(_085_),
    .B1(_091_),
    .C1(_136_),
    .Y(_139_));
 sky130_fd_sc_hd__a21oi_4 _372_ (.A1(_138_),
    .A2(_139_),
    .B1(_133_),
    .Y(_140_));
 sky130_fd_sc_hd__mux2i_1 _374_ (.A0(\dpath.a_lt_b$in1[0] ),
    .A1(\dpath.a_lt_b$in0[0] ),
    .S(_140_),
    .Y(_142_));
 sky130_fd_sc_hd__nand2_1 _376_ (.A(req_rdy),
    .B(req_msg[0]),
    .Y(_144_));
 sky130_fd_sc_hd__o21ai_1 _377_ (.A1(req_rdy),
    .A2(_142_),
    .B1(_144_),
    .Y(_003_));
 sky130_fd_sc_hd__mux2i_1 _378_ (.A0(\dpath.a_lt_b$in1[1] ),
    .A1(\dpath.a_lt_b$in0[1] ),
    .S(_140_),
    .Y(_145_));
 sky130_fd_sc_hd__nand2_1 _379_ (.A(req_rdy),
    .B(req_msg[1]),
    .Y(_146_));
 sky130_fd_sc_hd__o21ai_1 _380_ (.A1(req_rdy),
    .A2(_145_),
    .B1(_146_),
    .Y(_004_));
 sky130_fd_sc_hd__mux2i_1 _382_ (.A0(\dpath.a_lt_b$in1[2] ),
    .A1(\dpath.a_lt_b$in0[2] ),
    .S(_140_),
    .Y(_148_));
 sky130_fd_sc_hd__nand2_1 _383_ (.A(req_rdy),
    .B(req_msg[2]),
    .Y(_149_));
 sky130_fd_sc_hd__o21ai_1 _384_ (.A1(req_rdy),
    .A2(_148_),
    .B1(_149_),
    .Y(_005_));
 sky130_fd_sc_hd__mux2i_1 _385_ (.A0(\dpath.a_lt_b$in1[3] ),
    .A1(\dpath.a_lt_b$in0[3] ),
    .S(_140_),
    .Y(_150_));
 sky130_fd_sc_hd__nand2_1 _386_ (.A(req_rdy),
    .B(req_msg[3]),
    .Y(_151_));
 sky130_fd_sc_hd__o21ai_1 _387_ (.A1(req_rdy),
    .A2(_150_),
    .B1(_151_),
    .Y(_006_));
 sky130_fd_sc_hd__mux2i_1 _388_ (.A0(\dpath.a_lt_b$in1[4] ),
    .A1(\dpath.a_lt_b$in0[4] ),
    .S(_140_),
    .Y(_152_));
 sky130_fd_sc_hd__nand2_1 _389_ (.A(req_rdy),
    .B(req_msg[4]),
    .Y(_153_));
 sky130_fd_sc_hd__o21ai_1 _390_ (.A1(req_rdy),
    .A2(_152_),
    .B1(_153_),
    .Y(_007_));
 sky130_fd_sc_hd__mux2i_1 _391_ (.A0(\dpath.a_lt_b$in1[5] ),
    .A1(\dpath.a_lt_b$in0[5] ),
    .S(_140_),
    .Y(_154_));
 sky130_fd_sc_hd__nand2_1 _392_ (.A(req_rdy),
    .B(req_msg[5]),
    .Y(_155_));
 sky130_fd_sc_hd__o21ai_1 _393_ (.A1(req_rdy),
    .A2(_154_),
    .B1(_155_),
    .Y(_008_));
 sky130_fd_sc_hd__mux2i_1 _394_ (.A0(\dpath.a_lt_b$in1[6] ),
    .A1(\dpath.a_lt_b$in0[6] ),
    .S(_140_),
    .Y(_156_));
 sky130_fd_sc_hd__nand2_1 _395_ (.A(req_rdy),
    .B(req_msg[6]),
    .Y(_157_));
 sky130_fd_sc_hd__o21ai_1 _396_ (.A1(req_rdy),
    .A2(_156_),
    .B1(_157_),
    .Y(_009_));
 sky130_fd_sc_hd__mux2i_1 _397_ (.A0(\dpath.a_lt_b$in1[7] ),
    .A1(\dpath.a_lt_b$in0[7] ),
    .S(_140_),
    .Y(_158_));
 sky130_fd_sc_hd__nand2_1 _398_ (.A(req_rdy),
    .B(req_msg[7]),
    .Y(_159_));
 sky130_fd_sc_hd__o21ai_1 _399_ (.A1(req_rdy),
    .A2(_158_),
    .B1(_159_),
    .Y(_010_));
 sky130_fd_sc_hd__mux2i_1 _400_ (.A0(\dpath.a_lt_b$in1[8] ),
    .A1(\dpath.a_lt_b$in0[8] ),
    .S(_140_),
    .Y(_160_));
 sky130_fd_sc_hd__nand2_1 _401_ (.A(req_rdy),
    .B(req_msg[8]),
    .Y(_161_));
 sky130_fd_sc_hd__o21ai_1 _402_ (.A1(req_rdy),
    .A2(_160_),
    .B1(_161_),
    .Y(_011_));
 sky130_fd_sc_hd__mux2i_1 _403_ (.A0(\dpath.a_lt_b$in1[9] ),
    .A1(\dpath.a_lt_b$in0[9] ),
    .S(_140_),
    .Y(_162_));
 sky130_fd_sc_hd__nand2_1 _404_ (.A(req_rdy),
    .B(req_msg[9]),
    .Y(_163_));
 sky130_fd_sc_hd__o21ai_1 _405_ (.A1(req_rdy),
    .A2(_162_),
    .B1(_163_),
    .Y(_012_));
 sky130_fd_sc_hd__mux2i_1 _406_ (.A0(\dpath.a_lt_b$in1[10] ),
    .A1(\dpath.a_lt_b$in0[10] ),
    .S(_140_),
    .Y(_164_));
 sky130_fd_sc_hd__nand2_1 _407_ (.A(req_rdy),
    .B(req_msg[10]),
    .Y(_165_));
 sky130_fd_sc_hd__o21ai_1 _408_ (.A1(req_rdy),
    .A2(_164_),
    .B1(_165_),
    .Y(_013_));
 sky130_fd_sc_hd__mux2i_1 _409_ (.A0(\dpath.a_lt_b$in1[11] ),
    .A1(\dpath.a_lt_b$in0[11] ),
    .S(_140_),
    .Y(_166_));
 sky130_fd_sc_hd__nand2_1 _410_ (.A(req_rdy),
    .B(req_msg[11]),
    .Y(_167_));
 sky130_fd_sc_hd__o21ai_1 _411_ (.A1(req_rdy),
    .A2(_166_),
    .B1(_167_),
    .Y(_014_));
 sky130_fd_sc_hd__mux2i_1 _412_ (.A0(\dpath.a_lt_b$in1[12] ),
    .A1(\dpath.a_lt_b$in0[12] ),
    .S(_140_),
    .Y(_168_));
 sky130_fd_sc_hd__nand2_1 _413_ (.A(req_rdy),
    .B(req_msg[12]),
    .Y(_169_));
 sky130_fd_sc_hd__o21ai_1 _414_ (.A1(req_rdy),
    .A2(_168_),
    .B1(_169_),
    .Y(_015_));
 sky130_fd_sc_hd__mux2i_1 _415_ (.A0(\dpath.a_lt_b$in1[13] ),
    .A1(\dpath.a_lt_b$in0[13] ),
    .S(_140_),
    .Y(_170_));
 sky130_fd_sc_hd__nand2_1 _416_ (.A(req_rdy),
    .B(req_msg[13]),
    .Y(_171_));
 sky130_fd_sc_hd__o21ai_1 _417_ (.A1(req_rdy),
    .A2(_170_),
    .B1(_171_),
    .Y(_016_));
 sky130_fd_sc_hd__mux2i_1 _418_ (.A0(\dpath.a_lt_b$in1[14] ),
    .A1(\dpath.a_lt_b$in0[14] ),
    .S(_140_),
    .Y(_172_));
 sky130_fd_sc_hd__nand2_1 _419_ (.A(req_rdy),
    .B(req_msg[14]),
    .Y(_173_));
 sky130_fd_sc_hd__o21ai_1 _420_ (.A1(req_rdy),
    .A2(_172_),
    .B1(_173_),
    .Y(_017_));
 sky130_fd_sc_hd__o21ai_0 _421_ (.A1(_133_),
    .A2(\dpath.a_lt_b$in0[15] ),
    .B1(\dpath.a_lt_b$in1[15] ),
    .Y(_174_));
 sky130_fd_sc_hd__nand2_1 _422_ (.A(req_rdy),
    .B(req_msg[15]),
    .Y(_175_));
 sky130_fd_sc_hd__o21ai_0 _423_ (.A1(req_rdy),
    .A2(_174_),
    .B1(_175_),
    .Y(_018_));
 sky130_fd_sc_hd__inv_1 _424_ (.A(req_msg[16]),
    .Y(_176_));
 sky130_fd_sc_hd__nand2_1 _425_ (.A(\dpath.a_lt_b$in0[0] ),
    .B(\dpath.a_lt_b$in1[0] ),
    .Y(_177_));
 sky130_fd_sc_hd__and2_1 _426_ (.A(_138_),
    .B(_139_),
    .X(_178_));
 sky130_fd_sc_hd__mux2i_1 _428_ (.A0(\dpath.a_lt_b$in1[0] ),
    .A1(_177_),
    .S(_178_),
    .Y(_180_));
 sky130_fd_sc_hd__nor2_1 _429_ (.A(_133_),
    .B(req_rdy),
    .Y(_181_));
 sky130_fd_sc_hd__a211oi_1 _430_ (.A1(\ctrl.state.out[2] ),
    .A2(\dpath.a_lt_b$in1[0] ),
    .B1(\dpath.a_lt_b$in0[0] ),
    .C1(req_rdy),
    .Y(_182_));
 sky130_fd_sc_hd__a221oi_1 _431_ (.A1(req_rdy),
    .A2(_176_),
    .B1(_180_),
    .B2(_181_),
    .C1(_182_),
    .Y(_019_));
 sky130_fd_sc_hd__nand2_1 _432_ (.A(\ctrl.state.out[2] ),
    .B(_131_),
    .Y(_183_));
 sky130_fd_sc_hd__mux2i_1 _434_ (.A0(\dpath.a_lt_b$in1[1] ),
    .A1(resp_msg[1]),
    .S(_178_),
    .Y(_185_));
 sky130_fd_sc_hd__nor2_1 _435_ (.A(\ctrl.state.out[2] ),
    .B(req_rdy),
    .Y(_186_));
 sky130_fd_sc_hd__a22oi_1 _436_ (.A1(req_msg[17]),
    .A2(req_rdy),
    .B1(\dpath.a_lt_b$in0[1] ),
    .B2(_186_),
    .Y(_187_));
 sky130_fd_sc_hd__o21ai_1 _437_ (.A1(_183_),
    .A2(_185_),
    .B1(_187_),
    .Y(_020_));
 sky130_fd_sc_hd__mux2i_1 _438_ (.A0(\dpath.a_lt_b$in1[2] ),
    .A1(resp_msg[2]),
    .S(_178_),
    .Y(_188_));
 sky130_fd_sc_hd__a22oi_1 _439_ (.A1(req_msg[18]),
    .A2(req_rdy),
    .B1(\dpath.a_lt_b$in0[2] ),
    .B2(_186_),
    .Y(_189_));
 sky130_fd_sc_hd__o21ai_1 _440_ (.A1(_183_),
    .A2(_188_),
    .B1(_189_),
    .Y(_021_));
 sky130_fd_sc_hd__a21oi_1 _441_ (.A1(_138_),
    .A2(_139_),
    .B1(_060_),
    .Y(_190_));
 sky130_fd_sc_hd__a21oi_1 _442_ (.A1(resp_msg[3]),
    .A2(_178_),
    .B1(_190_),
    .Y(_191_));
 sky130_fd_sc_hd__a22oi_1 _443_ (.A1(req_msg[19]),
    .A2(req_rdy),
    .B1(\dpath.a_lt_b$in0[3] ),
    .B2(_186_),
    .Y(_192_));
 sky130_fd_sc_hd__o21ai_1 _444_ (.A1(_183_),
    .A2(_191_),
    .B1(_192_),
    .Y(_022_));
 sky130_fd_sc_hd__a21oi_1 _445_ (.A1(_138_),
    .A2(_139_),
    .B1(_100_),
    .Y(_193_));
 sky130_fd_sc_hd__a21oi_1 _446_ (.A1(resp_msg[4]),
    .A2(_178_),
    .B1(_193_),
    .Y(_194_));
 sky130_fd_sc_hd__a22oi_1 _447_ (.A1(req_msg[20]),
    .A2(req_rdy),
    .B1(\dpath.a_lt_b$in0[4] ),
    .B2(_186_),
    .Y(_195_));
 sky130_fd_sc_hd__o21ai_1 _448_ (.A1(_183_),
    .A2(_194_),
    .B1(_195_),
    .Y(_023_));
 sky130_fd_sc_hd__mux2i_1 _449_ (.A0(\dpath.a_lt_b$in1[5] ),
    .A1(resp_msg[5]),
    .S(_178_),
    .Y(_196_));
 sky130_fd_sc_hd__a22oi_1 _450_ (.A1(req_msg[21]),
    .A2(req_rdy),
    .B1(\dpath.a_lt_b$in0[5] ),
    .B2(_186_),
    .Y(_197_));
 sky130_fd_sc_hd__o21ai_0 _451_ (.A1(_183_),
    .A2(_196_),
    .B1(_197_),
    .Y(_024_));
 sky130_fd_sc_hd__nand2_1 _452_ (.A(\ctrl.state.out[2] ),
    .B(\dpath.a_lt_b$in0[6] ),
    .Y(_198_));
 sky130_fd_sc_hd__mux2i_1 _453_ (.A0(\dpath.a_lt_b$in0[6] ),
    .A1(_198_),
    .S(_105_),
    .Y(_199_));
 sky130_fd_sc_hd__o21bai_1 _454_ (.A1(_140_),
    .A2(_199_),
    .B1_N(\dpath.a_lt_b$in1[6] ),
    .Y(_200_));
 sky130_fd_sc_hd__and2_1 _455_ (.A(_072_),
    .B(_105_),
    .X(_201_));
 sky130_fd_sc_hd__nor3_1 _456_ (.A(_133_),
    .B(_072_),
    .C(_105_),
    .Y(_202_));
 sky130_fd_sc_hd__o211ai_1 _457_ (.A1(_201_),
    .A2(_202_),
    .B1(_178_),
    .C1(\dpath.a_lt_b$in1[6] ),
    .Y(_203_));
 sky130_fd_sc_hd__a21oi_1 _458_ (.A1(_133_),
    .A2(_072_),
    .B1(req_rdy),
    .Y(_204_));
 sky130_fd_sc_hd__a32o_1 _459_ (.A1(_200_),
    .A2(_203_),
    .A3(_204_),
    .B1(req_rdy),
    .B2(req_msg[22]),
    .X(_025_));
 sky130_fd_sc_hd__mux2i_1 _460_ (.A0(\dpath.a_lt_b$in1[7] ),
    .A1(resp_msg[7]),
    .S(_178_),
    .Y(_205_));
 sky130_fd_sc_hd__o2bb2ai_1 _461_ (.A1_N(_186_),
    .A2_N(_071_),
    .B1(_131_),
    .B2(req_msg[23]),
    .Y(_206_));
 sky130_fd_sc_hd__a21oi_1 _462_ (.A1(_181_),
    .A2(_205_),
    .B1(_206_),
    .Y(_026_));
 sky130_fd_sc_hd__a21oi_1 _463_ (.A1(_138_),
    .A2(_139_),
    .B1(_065_),
    .Y(_207_));
 sky130_fd_sc_hd__a21oi_1 _464_ (.A1(resp_msg[8]),
    .A2(_178_),
    .B1(_207_),
    .Y(_208_));
 sky130_fd_sc_hd__a22oi_1 _465_ (.A1(req_msg[24]),
    .A2(req_rdy),
    .B1(\dpath.a_lt_b$in0[8] ),
    .B2(_186_),
    .Y(_209_));
 sky130_fd_sc_hd__o21ai_1 _466_ (.A1(_183_),
    .A2(_208_),
    .B1(_209_),
    .Y(_027_));
 sky130_fd_sc_hd__xnor2_1 _467_ (.A(_066_),
    .B(_113_),
    .Y(_210_));
 sky130_fd_sc_hd__nor2_1 _468_ (.A(\dpath.a_lt_b$in0[9] ),
    .B(_113_),
    .Y(_211_));
 sky130_fd_sc_hd__nor2_1 _469_ (.A(\ctrl.state.out[2] ),
    .B(_211_),
    .Y(_212_));
 sky130_fd_sc_hd__a211oi_1 _470_ (.A1(_178_),
    .A2(_210_),
    .B1(_212_),
    .C1(\dpath.a_lt_b$in1[9] ),
    .Y(_213_));
 sky130_fd_sc_hd__nand2_1 _471_ (.A(\ctrl.state.out[2] ),
    .B(\dpath.a_lt_b$in0[9] ),
    .Y(_214_));
 sky130_fd_sc_hd__nand2_1 _472_ (.A(_066_),
    .B(_113_),
    .Y(_215_));
 sky130_fd_sc_hd__o21ai_0 _473_ (.A1(_113_),
    .A2(_214_),
    .B1(_215_),
    .Y(_216_));
 sky130_fd_sc_hd__nor2_1 _474_ (.A(\ctrl.state.out[2] ),
    .B(\dpath.a_lt_b$in0[9] ),
    .Y(_217_));
 sky130_fd_sc_hd__a311o_1 _475_ (.A1(\dpath.a_lt_b$in1[9] ),
    .A2(_178_),
    .A3(_216_),
    .B1(_217_),
    .C1(req_rdy),
    .X(_218_));
 sky130_fd_sc_hd__nand2_1 _476_ (.A(req_msg[25]),
    .B(req_rdy),
    .Y(_219_));
 sky130_fd_sc_hd__o21ai_1 _477_ (.A1(_213_),
    .A2(_218_),
    .B1(_219_),
    .Y(_028_));
 sky130_fd_sc_hd__inv_1 _478_ (.A(\dpath.a_lt_b$in1[10] ),
    .Y(_220_));
 sky130_fd_sc_hd__a22oi_1 _479_ (.A1(req_msg[26]),
    .A2(req_rdy),
    .B1(\dpath.a_lt_b$in0[10] ),
    .B2(_186_),
    .Y(_221_));
 sky130_fd_sc_hd__nand3_1 _480_ (.A(resp_msg[10]),
    .B(_178_),
    .C(_181_),
    .Y(_222_));
 sky130_fd_sc_hd__o311ai_2 _481_ (.A1(_220_),
    .A2(_178_),
    .A3(_183_),
    .B1(_221_),
    .C1(_222_),
    .Y(_029_));
 sky130_fd_sc_hd__inv_1 _482_ (.A(\dpath.a_lt_b$in0[11] ),
    .Y(_223_));
 sky130_fd_sc_hd__a311oi_1 _483_ (.A1(_042_),
    .A2(_037_),
    .A3(_114_),
    .B1(_036_),
    .C1(_223_),
    .Y(_224_));
 sky130_fd_sc_hd__and4_1 _484_ (.A(_223_),
    .B(_066_),
    .C(_037_),
    .D(_113_),
    .X(_225_));
 sky130_fd_sc_hd__nand2_1 _485_ (.A(\dpath.a_lt_b$in1[9] ),
    .B(_037_),
    .Y(_226_));
 sky130_fd_sc_hd__nor2_1 _486_ (.A(\dpath.a_lt_b$in0[11] ),
    .B(_226_),
    .Y(_227_));
 sky130_fd_sc_hd__nor3_1 _487_ (.A(\dpath.a_lt_b$in0[11] ),
    .B(\dpath.a_lt_b$in0[9] ),
    .C(_226_),
    .Y(_228_));
 sky130_fd_sc_hd__a221o_1 _488_ (.A1(_223_),
    .A2(_036_),
    .B1(_113_),
    .B2(_227_),
    .C1(_228_),
    .X(_229_));
 sky130_fd_sc_hd__o311ai_1 _489_ (.A1(_224_),
    .A2(_225_),
    .A3(_229_),
    .B1(_139_),
    .C1(_138_),
    .Y(_230_));
 sky130_fd_sc_hd__xor2_1 _490_ (.A(\dpath.a_lt_b$in1[11] ),
    .B(_230_),
    .X(_231_));
 sky130_fd_sc_hd__a22oi_1 _491_ (.A1(req_msg[27]),
    .A2(req_rdy),
    .B1(\dpath.a_lt_b$in0[11] ),
    .B2(_186_),
    .Y(_232_));
 sky130_fd_sc_hd__o21ai_1 _492_ (.A1(_183_),
    .A2(_231_),
    .B1(_232_),
    .Y(_030_));
 sky130_fd_sc_hd__mux2i_1 _493_ (.A0(\dpath.a_lt_b$in1[12] ),
    .A1(resp_msg[12]),
    .S(_178_),
    .Y(_233_));
 sky130_fd_sc_hd__a22oi_1 _494_ (.A1(req_msg[28]),
    .A2(req_rdy),
    .B1(\dpath.a_lt_b$in0[12] ),
    .B2(_186_),
    .Y(_234_));
 sky130_fd_sc_hd__o21ai_0 _495_ (.A1(_183_),
    .A2(_233_),
    .B1(_234_),
    .Y(_031_));
 sky130_fd_sc_hd__mux2i_1 _496_ (.A0(\dpath.a_lt_b$in1[13] ),
    .A1(resp_msg[13]),
    .S(_178_),
    .Y(_235_));
 sky130_fd_sc_hd__or3_1 _497_ (.A(\ctrl.state.out[2] ),
    .B(req_rdy),
    .C(\dpath.a_lt_b$in0[13] ),
    .X(_236_));
 sky130_fd_sc_hd__o21ai_0 _498_ (.A1(req_msg[29]),
    .A2(_131_),
    .B1(_236_),
    .Y(_237_));
 sky130_fd_sc_hd__a21oi_1 _499_ (.A1(_181_),
    .A2(_235_),
    .B1(_237_),
    .Y(_032_));
 sky130_fd_sc_hd__and3_1 _500_ (.A(_138_),
    .B(_139_),
    .C(_181_),
    .X(_238_));
 sky130_fd_sc_hd__nand2_1 _501_ (.A(\dpath.a_lt_b$in1[14] ),
    .B(\ctrl.state.out[2] ),
    .Y(_239_));
 sky130_fd_sc_hd__o22ai_1 _502_ (.A1(\ctrl.state.out[2] ),
    .A2(_086_),
    .B1(_178_),
    .B2(_239_),
    .Y(_240_));
 sky130_fd_sc_hd__and2_1 _503_ (.A(req_msg[30]),
    .B(req_rdy),
    .X(_241_));
 sky130_fd_sc_hd__a221o_1 _504_ (.A1(resp_msg[14]),
    .A2(_238_),
    .B1(_240_),
    .B2(_131_),
    .C1(_241_),
    .X(_033_));
 sky130_fd_sc_hd__nor2_1 _505_ (.A(\dpath.a_lt_b$in1[15] ),
    .B(_136_),
    .Y(_242_));
 sky130_fd_sc_hd__nand2_1 _506_ (.A(\dpath.a_lt_b$in1[15] ),
    .B(\ctrl.state.out[2] ),
    .Y(_243_));
 sky130_fd_sc_hd__a21oi_1 _507_ (.A1(\dpath.a_lt_b$in0[15] ),
    .A2(_092_),
    .B1(_243_),
    .Y(_244_));
 sky130_fd_sc_hd__a221oi_1 _508_ (.A1(_133_),
    .A2(\dpath.a_lt_b$in0[15] ),
    .B1(_092_),
    .B2(_242_),
    .C1(_244_),
    .Y(_245_));
 sky130_fd_sc_hd__nand2_1 _509_ (.A(req_msg[31]),
    .B(req_rdy),
    .Y(_246_));
 sky130_fd_sc_hd__o21ai_0 _510_ (.A1(req_rdy),
    .A2(_245_),
    .B1(_246_),
    .Y(_034_));
 sky130_fd_sc_hd__dfxtp_1 _511_ (.D(_000_),
    .Q(req_rdy),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _512_ (.D(_001_),
    .Q(\ctrl.state.out[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _513_ (.D(_002_),
    .Q(\ctrl.state.out[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _514_ (.D(_003_),
    .Q(\dpath.a_lt_b$in1[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _515_ (.D(_004_),
    .Q(\dpath.a_lt_b$in1[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _516_ (.D(_005_),
    .Q(\dpath.a_lt_b$in1[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _517_ (.D(_006_),
    .Q(\dpath.a_lt_b$in1[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _518_ (.D(_007_),
    .Q(\dpath.a_lt_b$in1[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _519_ (.D(_008_),
    .Q(\dpath.a_lt_b$in1[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _520_ (.D(_009_),
    .Q(\dpath.a_lt_b$in1[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _521_ (.D(_010_),
    .Q(\dpath.a_lt_b$in1[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _522_ (.D(_011_),
    .Q(\dpath.a_lt_b$in1[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _523_ (.D(_012_),
    .Q(\dpath.a_lt_b$in1[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _524_ (.D(_013_),
    .Q(\dpath.a_lt_b$in1[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _525_ (.D(_014_),
    .Q(\dpath.a_lt_b$in1[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _526_ (.D(_015_),
    .Q(\dpath.a_lt_b$in1[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _527_ (.D(_016_),
    .Q(\dpath.a_lt_b$in1[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _528_ (.D(_017_),
    .Q(\dpath.a_lt_b$in1[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _529_ (.D(_018_),
    .Q(\dpath.a_lt_b$in1[15] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _530_ (.D(_019_),
    .Q(\dpath.a_lt_b$in0[0] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _531_ (.D(_020_),
    .Q(\dpath.a_lt_b$in0[1] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _532_ (.D(_021_),
    .Q(\dpath.a_lt_b$in0[2] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _533_ (.D(_022_),
    .Q(\dpath.a_lt_b$in0[3] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _534_ (.D(_023_),
    .Q(\dpath.a_lt_b$in0[4] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _535_ (.D(_024_),
    .Q(\dpath.a_lt_b$in0[5] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _536_ (.D(_025_),
    .Q(\dpath.a_lt_b$in0[6] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _537_ (.D(_026_),
    .Q(\dpath.a_lt_b$in0[7] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _538_ (.D(_027_),
    .Q(\dpath.a_lt_b$in0[8] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _539_ (.D(_028_),
    .Q(\dpath.a_lt_b$in0[9] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _540_ (.D(_029_),
    .Q(\dpath.a_lt_b$in0[10] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _541_ (.D(_030_),
    .Q(\dpath.a_lt_b$in0[11] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _542_ (.D(_031_),
    .Q(\dpath.a_lt_b$in0[12] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _543_ (.D(_032_),
    .Q(\dpath.a_lt_b$in0[13] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _544_ (.D(_033_),
    .Q(\dpath.a_lt_b$in0[14] ),
    .CLK(clk));
 sky130_fd_sc_hd__dfxtp_1 _545_ (.D(_034_),
    .Q(\dpath.a_lt_b$in0[15] ),
    .CLK(clk));
endmodule
