VERSION 5.6 ;
  BUSBITCHARS "[]" ;
  DIVIDERCHAR "/" ;

MACRO capacitor_test_nf
  CLASS CORE ;
  ORIGIN 0.000 0.000 ;
  FOREIGN capacitor_test_nf 0 0 ;
  SIZE 30.720 BY 36.630 ;
  PIN pin0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 7.860 25.990 29.860 ;
        RECT 3.990 6.670 5.750 7.860 ;
    END
  END pin0
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 8.395 30.720 8.765 ;
      LAYER via ;
        RECT 3.300 8.420 3.560 8.680 ;
        RECT 26.305 8.420 26.565 8.680 ;
      LAYER met2 ;
        RECT 3.200 7.720 3.850 11.315 ;
        RECT 26.130 7.720 26.780 11.315 ;
      LAYER via2 ;
        RECT 3.395 10.515 3.675 10.795 ;
        RECT 3.395 9.685 3.675 9.965 ;
        RECT 3.395 8.830 3.675 9.110 ;
        RECT 3.395 7.945 3.675 8.225 ;
        RECT 26.320 10.515 26.600 10.795 ;
        RECT 26.320 9.685 26.600 9.965 ;
        RECT 26.320 8.830 26.600 9.110 ;
        RECT 26.320 7.945 26.600 8.225 ;
      LAYER met3 ;
        RECT 3.200 7.720 26.780 30.000 ;
    END
  END vgnd
  OBS
#      LAYER nwell ;
#        RECT -0.330 34.445 31.050 37.045 ;
#      LAYER pwell ;
#        RECT -0.130 32.345 30.850 32.775 ;
#      LAYER nwell ;
#        RECT -0.330 26.305 0.810 30.675 ;
#        RECT 29.910 26.305 31.050 30.675 ;
#      LAYER pwell ;
#        RECT -0.130 24.205 0.610 24.635 ;
#        RECT 30.110 24.205 30.850 24.635 ;
#      LAYER nwell ;
#        RECT -0.330 18.165 0.810 22.535 ;
#        RECT 29.910 18.165 31.050 22.535 ;
#      LAYER pwell ;
#        RECT -0.130 16.065 0.610 16.495 ;
#        RECT 30.110 16.065 30.850 16.495 ;
#      LAYER nwell ;
#        RECT -0.330 10.025 0.810 14.395 ;
#        RECT 29.910 10.025 31.050 14.395 ;
#      LAYER pwell ;
#        RECT -0.130 7.925 0.610 8.355 ;
#        RECT 30.110 7.925 30.850 8.355 ;
#      LAYER nwell ;
#        RECT -0.330 4.485 0.810 6.255 ;
#        RECT 29.910 4.485 31.050 6.255 ;
#        RECT -0.330 1.885 31.050 4.485 ;
#      LAYER pwell ;
#        RECT -0.130 -0.215 30.850 0.215 ;
      LAYER li1 ;
        RECT 0.000 36.545 30.720 36.715 ;
        RECT 0.000 32.475 30.720 32.645 ;
        RECT 0.000 28.405 0.480 28.575 ;
        RECT 30.240 28.405 30.720 28.575 ;
        RECT 0.000 24.335 0.480 24.505 ;
        RECT 30.240 24.335 30.720 24.505 ;
        RECT 0.000 20.265 0.480 20.435 ;
        RECT 30.240 20.265 30.720 20.435 ;
        RECT 0.000 16.195 0.480 16.365 ;
        RECT 30.240 16.195 30.720 16.365 ;
        RECT 0.000 12.125 0.480 12.295 ;
        RECT 30.240 12.125 30.720 12.295 ;
        RECT 0.000 8.055 0.480 8.225 ;
        RECT 30.240 8.055 30.720 8.225 ;
        RECT 0.000 3.985 30.720 4.155 ;
        RECT 0.000 -0.085 30.720 0.085 ;
      LAYER mcon ;
        RECT 0.155 36.545 0.325 36.715 ;
        RECT 0.635 36.545 0.805 36.715 ;
        RECT 1.115 36.545 1.285 36.715 ;
        RECT 1.595 36.545 1.765 36.715 ;
        RECT 2.075 36.545 2.245 36.715 ;
        RECT 2.555 36.545 2.725 36.715 ;
        RECT 3.035 36.545 3.205 36.715 ;
        RECT 3.515 36.545 3.685 36.715 ;
        RECT 3.995 36.545 4.165 36.715 ;
        RECT 4.475 36.545 4.645 36.715 ;
        RECT 4.955 36.545 5.125 36.715 ;
        RECT 5.435 36.545 5.605 36.715 ;
        RECT 5.915 36.545 6.085 36.715 ;
        RECT 6.395 36.545 6.565 36.715 ;
        RECT 6.875 36.545 7.045 36.715 ;
        RECT 7.355 36.545 7.525 36.715 ;
        RECT 7.835 36.545 8.005 36.715 ;
        RECT 8.315 36.545 8.485 36.715 ;
        RECT 8.795 36.545 8.965 36.715 ;
        RECT 9.275 36.545 9.445 36.715 ;
        RECT 9.755 36.545 9.925 36.715 ;
        RECT 10.235 36.545 10.405 36.715 ;
        RECT 10.715 36.545 10.885 36.715 ;
        RECT 11.195 36.545 11.365 36.715 ;
        RECT 11.675 36.545 11.845 36.715 ;
        RECT 12.155 36.545 12.325 36.715 ;
        RECT 12.635 36.545 12.805 36.715 ;
        RECT 13.115 36.545 13.285 36.715 ;
        RECT 13.595 36.545 13.765 36.715 ;
        RECT 14.075 36.545 14.245 36.715 ;
        RECT 14.555 36.545 14.725 36.715 ;
        RECT 15.035 36.545 15.205 36.715 ;
        RECT 15.515 36.545 15.685 36.715 ;
        RECT 15.995 36.545 16.165 36.715 ;
        RECT 16.475 36.545 16.645 36.715 ;
        RECT 16.955 36.545 17.125 36.715 ;
        RECT 17.435 36.545 17.605 36.715 ;
        RECT 17.915 36.545 18.085 36.715 ;
        RECT 18.395 36.545 18.565 36.715 ;
        RECT 18.875 36.545 19.045 36.715 ;
        RECT 19.355 36.545 19.525 36.715 ;
        RECT 19.835 36.545 20.005 36.715 ;
        RECT 20.315 36.545 20.485 36.715 ;
        RECT 20.795 36.545 20.965 36.715 ;
        RECT 21.275 36.545 21.445 36.715 ;
        RECT 21.755 36.545 21.925 36.715 ;
        RECT 22.235 36.545 22.405 36.715 ;
        RECT 22.715 36.545 22.885 36.715 ;
        RECT 23.195 36.545 23.365 36.715 ;
        RECT 23.675 36.545 23.845 36.715 ;
        RECT 24.155 36.545 24.325 36.715 ;
        RECT 24.635 36.545 24.805 36.715 ;
        RECT 25.115 36.545 25.285 36.715 ;
        RECT 25.595 36.545 25.765 36.715 ;
        RECT 26.075 36.545 26.245 36.715 ;
        RECT 26.555 36.545 26.725 36.715 ;
        RECT 27.035 36.545 27.205 36.715 ;
        RECT 27.515 36.545 27.685 36.715 ;
        RECT 27.995 36.545 28.165 36.715 ;
        RECT 28.475 36.545 28.645 36.715 ;
        RECT 28.955 36.545 29.125 36.715 ;
        RECT 29.435 36.545 29.605 36.715 ;
        RECT 29.915 36.545 30.085 36.715 ;
        RECT 30.395 36.545 30.565 36.715 ;
        RECT 0.155 32.475 0.325 32.645 ;
        RECT 0.635 32.475 0.805 32.645 ;
        RECT 1.115 32.475 1.285 32.645 ;
        RECT 1.595 32.475 1.765 32.645 ;
        RECT 2.075 32.475 2.245 32.645 ;
        RECT 2.555 32.475 2.725 32.645 ;
        RECT 3.035 32.475 3.205 32.645 ;
        RECT 3.515 32.475 3.685 32.645 ;
        RECT 3.995 32.475 4.165 32.645 ;
        RECT 4.475 32.475 4.645 32.645 ;
        RECT 4.955 32.475 5.125 32.645 ;
        RECT 5.435 32.475 5.605 32.645 ;
        RECT 5.915 32.475 6.085 32.645 ;
        RECT 6.395 32.475 6.565 32.645 ;
        RECT 6.875 32.475 7.045 32.645 ;
        RECT 7.355 32.475 7.525 32.645 ;
        RECT 7.835 32.475 8.005 32.645 ;
        RECT 8.315 32.475 8.485 32.645 ;
        RECT 8.795 32.475 8.965 32.645 ;
        RECT 9.275 32.475 9.445 32.645 ;
        RECT 9.755 32.475 9.925 32.645 ;
        RECT 10.235 32.475 10.405 32.645 ;
        RECT 10.715 32.475 10.885 32.645 ;
        RECT 11.195 32.475 11.365 32.645 ;
        RECT 11.675 32.475 11.845 32.645 ;
        RECT 12.155 32.475 12.325 32.645 ;
        RECT 12.635 32.475 12.805 32.645 ;
        RECT 13.115 32.475 13.285 32.645 ;
        RECT 13.595 32.475 13.765 32.645 ;
        RECT 14.075 32.475 14.245 32.645 ;
        RECT 14.555 32.475 14.725 32.645 ;
        RECT 15.035 32.475 15.205 32.645 ;
        RECT 15.515 32.475 15.685 32.645 ;
        RECT 15.995 32.475 16.165 32.645 ;
        RECT 16.475 32.475 16.645 32.645 ;
        RECT 16.955 32.475 17.125 32.645 ;
        RECT 17.435 32.475 17.605 32.645 ;
        RECT 17.915 32.475 18.085 32.645 ;
        RECT 18.395 32.475 18.565 32.645 ;
        RECT 18.875 32.475 19.045 32.645 ;
        RECT 19.355 32.475 19.525 32.645 ;
        RECT 19.835 32.475 20.005 32.645 ;
        RECT 20.315 32.475 20.485 32.645 ;
        RECT 20.795 32.475 20.965 32.645 ;
        RECT 21.275 32.475 21.445 32.645 ;
        RECT 21.755 32.475 21.925 32.645 ;
        RECT 22.235 32.475 22.405 32.645 ;
        RECT 22.715 32.475 22.885 32.645 ;
        RECT 23.195 32.475 23.365 32.645 ;
        RECT 23.675 32.475 23.845 32.645 ;
        RECT 24.155 32.475 24.325 32.645 ;
        RECT 24.635 32.475 24.805 32.645 ;
        RECT 25.115 32.475 25.285 32.645 ;
        RECT 25.595 32.475 25.765 32.645 ;
        RECT 26.075 32.475 26.245 32.645 ;
        RECT 26.555 32.475 26.725 32.645 ;
        RECT 27.035 32.475 27.205 32.645 ;
        RECT 27.515 32.475 27.685 32.645 ;
        RECT 27.995 32.475 28.165 32.645 ;
        RECT 28.475 32.475 28.645 32.645 ;
        RECT 28.955 32.475 29.125 32.645 ;
        RECT 29.435 32.475 29.605 32.645 ;
        RECT 29.915 32.475 30.085 32.645 ;
        RECT 30.395 32.475 30.565 32.645 ;
        RECT 0.155 28.405 0.325 28.575 ;
        RECT 30.395 28.405 30.565 28.575 ;
        RECT 0.155 24.335 0.325 24.505 ;
        RECT 30.395 24.335 30.565 24.505 ;
        RECT 0.155 20.265 0.325 20.435 ;
        RECT 30.395 20.265 30.565 20.435 ;
        RECT 0.155 16.195 0.325 16.365 ;
        RECT 30.395 16.195 30.565 16.365 ;
        RECT 0.155 12.125 0.325 12.295 ;
        RECT 30.395 12.125 30.565 12.295 ;
        RECT 0.155 8.055 0.325 8.225 ;
        RECT 30.395 8.055 30.565 8.225 ;
        RECT 0.155 3.985 0.325 4.155 ;
        RECT 0.635 3.985 0.805 4.155 ;
        RECT 1.115 3.985 1.285 4.155 ;
        RECT 1.595 3.985 1.765 4.155 ;
        RECT 2.075 3.985 2.245 4.155 ;
        RECT 2.555 3.985 2.725 4.155 ;
        RECT 3.035 3.985 3.205 4.155 ;
        RECT 3.515 3.985 3.685 4.155 ;
        RECT 3.995 3.985 4.165 4.155 ;
        RECT 4.475 3.985 4.645 4.155 ;
        RECT 4.955 3.985 5.125 4.155 ;
        RECT 5.435 3.985 5.605 4.155 ;
        RECT 5.915 3.985 6.085 4.155 ;
        RECT 6.395 3.985 6.565 4.155 ;
        RECT 6.875 3.985 7.045 4.155 ;
        RECT 7.355 3.985 7.525 4.155 ;
        RECT 7.835 3.985 8.005 4.155 ;
        RECT 8.315 3.985 8.485 4.155 ;
        RECT 8.795 3.985 8.965 4.155 ;
        RECT 9.275 3.985 9.445 4.155 ;
        RECT 9.755 3.985 9.925 4.155 ;
        RECT 10.235 3.985 10.405 4.155 ;
        RECT 10.715 3.985 10.885 4.155 ;
        RECT 11.195 3.985 11.365 4.155 ;
        RECT 11.675 3.985 11.845 4.155 ;
        RECT 12.155 3.985 12.325 4.155 ;
        RECT 12.635 3.985 12.805 4.155 ;
        RECT 13.115 3.985 13.285 4.155 ;
        RECT 13.595 3.985 13.765 4.155 ;
        RECT 14.075 3.985 14.245 4.155 ;
        RECT 14.555 3.985 14.725 4.155 ;
        RECT 15.035 3.985 15.205 4.155 ;
        RECT 15.515 3.985 15.685 4.155 ;
        RECT 15.995 3.985 16.165 4.155 ;
        RECT 16.475 3.985 16.645 4.155 ;
        RECT 16.955 3.985 17.125 4.155 ;
        RECT 17.435 3.985 17.605 4.155 ;
        RECT 17.915 3.985 18.085 4.155 ;
        RECT 18.395 3.985 18.565 4.155 ;
        RECT 18.875 3.985 19.045 4.155 ;
        RECT 19.355 3.985 19.525 4.155 ;
        RECT 19.835 3.985 20.005 4.155 ;
        RECT 20.315 3.985 20.485 4.155 ;
        RECT 20.795 3.985 20.965 4.155 ;
        RECT 21.275 3.985 21.445 4.155 ;
        RECT 21.755 3.985 21.925 4.155 ;
        RECT 22.235 3.985 22.405 4.155 ;
        RECT 22.715 3.985 22.885 4.155 ;
        RECT 23.195 3.985 23.365 4.155 ;
        RECT 23.675 3.985 23.845 4.155 ;
        RECT 24.155 3.985 24.325 4.155 ;
        RECT 24.635 3.985 24.805 4.155 ;
        RECT 25.115 3.985 25.285 4.155 ;
        RECT 25.595 3.985 25.765 4.155 ;
        RECT 26.075 3.985 26.245 4.155 ;
        RECT 26.555 3.985 26.725 4.155 ;
        RECT 27.035 3.985 27.205 4.155 ;
        RECT 27.515 3.985 27.685 4.155 ;
        RECT 27.995 3.985 28.165 4.155 ;
        RECT 28.475 3.985 28.645 4.155 ;
        RECT 28.955 3.985 29.125 4.155 ;
        RECT 29.435 3.985 29.605 4.155 ;
        RECT 29.915 3.985 30.085 4.155 ;
        RECT 30.395 3.985 30.565 4.155 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
        RECT 13.595 -0.085 13.765 0.085 ;
        RECT 14.075 -0.085 14.245 0.085 ;
        RECT 14.555 -0.085 14.725 0.085 ;
        RECT 15.035 -0.085 15.205 0.085 ;
        RECT 15.515 -0.085 15.685 0.085 ;
        RECT 15.995 -0.085 16.165 0.085 ;
        RECT 16.475 -0.085 16.645 0.085 ;
        RECT 16.955 -0.085 17.125 0.085 ;
        RECT 17.435 -0.085 17.605 0.085 ;
        RECT 17.915 -0.085 18.085 0.085 ;
        RECT 18.395 -0.085 18.565 0.085 ;
        RECT 18.875 -0.085 19.045 0.085 ;
        RECT 19.355 -0.085 19.525 0.085 ;
        RECT 19.835 -0.085 20.005 0.085 ;
        RECT 20.315 -0.085 20.485 0.085 ;
        RECT 20.795 -0.085 20.965 0.085 ;
        RECT 21.275 -0.085 21.445 0.085 ;
        RECT 21.755 -0.085 21.925 0.085 ;
        RECT 22.235 -0.085 22.405 0.085 ;
        RECT 22.715 -0.085 22.885 0.085 ;
        RECT 23.195 -0.085 23.365 0.085 ;
        RECT 23.675 -0.085 23.845 0.085 ;
        RECT 24.155 -0.085 24.325 0.085 ;
        RECT 24.635 -0.085 24.805 0.085 ;
        RECT 25.115 -0.085 25.285 0.085 ;
        RECT 25.595 -0.085 25.765 0.085 ;
        RECT 26.075 -0.085 26.245 0.085 ;
        RECT 26.555 -0.085 26.725 0.085 ;
        RECT 27.035 -0.085 27.205 0.085 ;
        RECT 27.515 -0.085 27.685 0.085 ;
        RECT 27.995 -0.085 28.165 0.085 ;
        RECT 28.475 -0.085 28.645 0.085 ;
        RECT 28.955 -0.085 29.125 0.085 ;
        RECT 29.435 -0.085 29.605 0.085 ;
        RECT 29.915 -0.085 30.085 0.085 ;
        RECT 30.395 -0.085 30.565 0.085 ;
      LAYER met1 ;
        RECT 0.000 36.515 30.720 36.745 ;
        RECT 0.000 36.005 30.720 36.375 ;
        RECT 0.000 32.815 30.720 33.185 ;
        RECT 0.000 32.445 30.720 32.675 ;
        RECT 0.000 31.935 0.480 32.305 ;
        RECT 30.240 31.935 30.720 32.305 ;
        RECT 0.000 28.745 0.480 29.115 ;
        RECT 30.240 28.745 30.720 29.115 ;
        RECT 0.000 28.375 0.480 28.605 ;
        RECT 30.240 28.375 30.720 28.605 ;
        RECT 0.000 27.865 0.480 28.235 ;
        RECT 30.240 27.865 30.720 28.235 ;
        RECT 0.000 24.675 0.480 25.045 ;
        RECT 30.240 24.675 30.720 25.045 ;
        RECT 0.000 24.305 0.480 24.535 ;
        RECT 30.240 24.305 30.720 24.535 ;
        RECT 0.000 23.795 0.480 24.165 ;
        RECT 30.240 23.795 30.720 24.165 ;
        RECT 0.000 20.605 0.480 20.975 ;
        RECT 30.240 20.605 30.720 20.975 ;
        RECT 0.000 20.235 0.480 20.465 ;
        RECT 30.240 20.235 30.720 20.465 ;
        RECT 0.000 19.725 0.480 20.095 ;
        RECT 30.240 19.725 30.720 20.095 ;
        RECT 0.000 16.535 0.480 16.905 ;
        RECT 30.240 16.535 30.720 16.905 ;
        RECT 0.000 16.165 0.480 16.395 ;
        RECT 30.240 16.165 30.720 16.395 ;
        RECT 0.000 15.655 0.480 16.025 ;
        RECT 30.240 15.655 30.720 16.025 ;
        RECT 0.000 12.465 0.480 12.835 ;
        RECT 30.240 12.465 30.720 12.835 ;
        RECT 0.000 12.095 0.480 12.325 ;
        RECT 30.240 12.095 30.720 12.325 ;
        RECT 0.000 11.585 0.480 11.955 ;
        RECT 30.240 11.585 30.720 11.955 ;
        RECT 0.000 8.025 0.480 8.255 ;
        RECT 30.240 8.025 30.720 8.255 ;
        RECT 0.000 7.515 0.480 7.885 ;
        RECT 30.240 7.515 30.720 7.885 ;
        RECT 0.000 4.325 0.480 4.695 ;
        RECT 30.240 4.325 30.720 4.695 ;
        RECT 0.000 3.955 30.720 4.185 ;
        RECT 0.000 3.445 30.720 3.815 ;
        RECT 0.000 0.255 30.720 0.625 ;
        RECT 0.000 -0.115 30.720 0.115 ;
  END
END capacitor_test_nf
END LIBRARY

