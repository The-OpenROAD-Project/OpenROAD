VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.1 ;

LAYER M1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 ;
  WIDTH 0.1 ;
  OFFSET 0.1 ;
  AREA 0.042 ;
END M1

LAYER M2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 ;
  WIDTH 0.1 ;
  OFFSET 0.1 ;
  AREA 0.052 ;
END M2

SITE site1
  CLASS CORE ;
  SIZE 50 BY 20 ;
END site1

MACRO snl_bufx1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_bufx1

MACRO snl_bufx2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_bufx2

MACRO snl_invx1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_invx1

MACRO snl_and02x1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_and02x1

MACRO snl_nor02x1
 SIZE 50 BY 20 ;
 PIN ZN DIRECTION OUTPUT ; END ZN
 PIN A DIRECTION INPUT ; END A
 PIN B DIRECTION INPUT ; END B
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_nor02x1

MACRO snl_ffqx1
 SIZE 50 BY 20 ;
 PIN Q DIRECTION OUTPUT ; END Q
 PIN D DIRECTION INPUT ; END D
 PIN CP DIRECTION INPUT ; END CP
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_ffqx1

END LIBRARY
