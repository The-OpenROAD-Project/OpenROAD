module top ();
 LOGIC1_X1 t1 (.Z(n1));
 BUF_X1 u0 (.A(n1));
 BUF_X1 u1 (.A(n1));
 BUF_X1 u2 (.A(n1));
 BUF_X1 u3 (.A(n1));
 BUF_X1 u4 (.A(n1));
 BUF_X1 u5 (.A(n1));
 PAD pad1 (.IN(n1));
 PAD pad2 (.IN(n1));
endmodule
