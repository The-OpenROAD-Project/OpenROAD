VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO COVER_MACRO
  CLASS COVER BUMP ;
  ORIGIN 0.0 0.0 ;
  SIZE 100.0 BY 100.0 ;
END COVER_MACRO

END LIBRARY
