module wb_dma_top (
	clk, 
	rst_i, 
	wb0s_data_i, 
	wb0s_data_o, 
	wb0_addr_i, 
	wb0_sel_i, 
	wb0_we_i, 
	wb0_cyc_i, 
	wb0_stb_i, 
	wb0_ack_o, 
	wb0_err_o, 
	wb0_rty_o, 
	wb0m_data_i, 
	wb0m_data_o, 
	wb0_addr_o, 
	wb0_sel_o, 
	wb0_we_o, 
	wb0_cyc_o, 
	wb0_stb_o, 
	wb0_ack_i, 
	wb0_err_i, 
	wb0_rty_i, 
	wb1s_data_i, 
	wb1s_data_o, 
	wb1_addr_i, 
	wb1_sel_i, 
	wb1_we_i, 
	wb1_cyc_i, 
	wb1_stb_i, 
	wb1_ack_o, 
	wb1_err_o, 
	wb1_rty_o, 
	wb1m_data_i, 
	wb1m_data_o, 
	wb1_addr_o, 
	wb1_sel_o, 
	wb1_we_o, 
	wb1_cyc_o, 
	wb1_stb_o, 
	wb1_ack_i, 
	wb1_err_i, 
	wb1_rty_i, 
	dma_req_i, 
	dma_ack_o, 
	dma_nd_i, 
	dma_rest_i, 
	inta_o, 
	intb_o);
   input clk;
   input rst_i;
   input [31:0] wb0s_data_i;
   output [31:0] wb0s_data_o;
   input [31:0] wb0_addr_i;
   input [3:0] wb0_sel_i;
   input wb0_we_i;
   input wb0_cyc_i;
   input wb0_stb_i;
   output wb0_ack_o;
   output wb0_err_o;
   output wb0_rty_o;
   input [31:0] wb0m_data_i;
   output [31:0] wb0m_data_o;
   output [31:0] wb0_addr_o;
   output [3:0] wb0_sel_o;
   output wb0_we_o;
   output wb0_cyc_o;
   output wb0_stb_o;
   input wb0_ack_i;
   input wb0_err_i;
   input wb0_rty_i;
   input [31:0] wb1s_data_i;
   output [31:0] wb1s_data_o;
   input [31:0] wb1_addr_i;
   input [3:0] wb1_sel_i;
   input wb1_we_i;
   input wb1_cyc_i;
   input wb1_stb_i;
   output wb1_ack_o;
   output wb1_err_o;
   output wb1_rty_o;
   input [31:0] wb1m_data_i;
   output [31:0] wb1m_data_o;
   output [31:0] wb1_addr_o;
   output [3:0] wb1_sel_o;
   output wb1_we_o;
   output wb1_cyc_o;
   output wb1_stb_o;
   input wb1_ack_i;
   input wb1_err_i;
   input wb1_rty_i;
   input [0:0] dma_req_i;
   output [0:0] dma_ack_o;
   input [0:0] dma_nd_i;
   input [0:0] dma_rest_i;
   output inta_o;
   output intb_o;

   // Internal wires
   wire FE_OCPN676_n1580;
   wire FE_OCPN675_n1580;
   wire FE_OCPN674_n2186;
   wire FE_OCPN673_n1577;
   wire FE_OCPN672_n1577;
   wire FE_OCPN671_n2356;
   wire FE_OCPN670_n2356;
   wire FE_OCPN669_slv0_adr_4_;
   wire FE_OCPN668_wb1_cyc_o;
   wire FE_OCPN667_wb1_cyc_o;
   wire FE_OCPN666_wb1_cyc_o;
   wire FE_OCPN665_wb1_cyc_o;
   wire FE_OCPN664_FE_RN_16;
   wire FE_OCPN663_n1428;
   wire FE_UNCONNECTED_37;
   wire FE_UNCONNECTED_36;
   wire FE_UNCONNECTED_35;
   wire FE_OCPN659_wb1_cyc_o;
   wire FE_OCPN661_wb1_cyc_o;
   wire FE_OCPN660_wb1_cyc_o;
   wire FE_OCPN658_wb1_cyc_o;
   wire FE_OCPN657_wb1_cyc_o;
   wire FE_OCPN656_wb1_cyc_o;
   wire FE_OCPN655_wb1_cyc_o;
   wire FE_OCPN651_wb1_cyc_o;
   wire FE_OCPN643_wb1_cyc_o;
   wire FE_OCPN642_wb1_cyc_o;
   wire FE_OCPN636_wb1_cyc_o;
   wire FE_OCPN634_wb1_cyc_o;
   wire FE_OCPN633_wb1_cyc_o;
   wire FE_OCPN632_wb1_cyc_o;
   wire FE_OCPN631_wb1_cyc_o;
   wire FE_OCPN630_wb1_cyc_o;
   wire FE_OCPN629_wb1_cyc_o;
   wire FE_OCPN628_wb1_cyc_o;
   wire FE_OCPN627_wb1_cyc_o;
   wire FE_OCPN626_wb1_cyc_o;
   wire FE_OCPN625_wb1_cyc_o;
   wire FE_OCPN624_wb1_cyc_o;
   wire FE_OCPN622_n1516;
   wire FE_OCPN620_n1516;
   wire FE_OCPN619_n1513;
   wire FE_OCPN618_n1591;
   wire FE_OCPN617_slv0_adr_5_;
   wire FE_OCPN615_n1516;
   wire FE_OCPN614_n1516;
   wire FE_OCPN613_n1516;
   wire FE_OCPN612_n1516;
   wire FE_OCPN611_slv0_adr_3_;
   wire FE_OCPN610_slv0_adr_3_;
   wire FE_OCPN609_slv0_adr_3_;
   wire FE_UNCONNECTED_34;
   wire FE_UNCONNECTED_33;
   wire FE_UNCONNECTED_32;
   wire FE_RN_61_0;
   wire FE_RN_60_0;
   wire FE_RN_59_0;
   wire FE_OCPN566_n2357;
   wire FE_OCPN565_n2357;
   wire FE_OCPN562_n2357;
   wire FE_OCPN561_n2357;
   wire FE_OCPN560_n2357;
   wire FE_OCPN559_n2357;
   wire FE_OCPN558_n2357;
   wire FE_RN_18;
   wire FE_RN_58_0;
   wire FE_RN_57_0;
   wire FE_RN_56_0;
   wire FE_OCPN554_n1529;
   wire FE_OCPN553_n1529;
   wire FE_RN_55_0;
   wire FE_RN_54_0;
   wire FE_RN_53_0;
   wire FE_OCPN552_n1424;
   wire FE_OCPN549_n1529;
   wire FE_OCPN547_n1529;
   wire FE_OCPN545_n2159;
   wire FE_OCPN544_n2159;
   wire FE_UNCONNECTED_31;
   wire FE_OCPN540_n1595;
   wire FE_OCPN539_n1595;
   wire FE_OCPN538_n1595;
   wire FE_OCPN537_n1595;
   wire FE_UNCONNECTED_30;
   wire FE_UNCONNECTED_29;
   wire FE_UNCONNECTED_28;
   wire FE_OCPN528_n1597;
   wire FE_RN_17;
   wire FE_RN_16;
   wire FE_OCPN514_slv0_adr_3_;
   wire FE_OCPN513_slv0_adr_3_;
   wire FE_OCPN512_slv0_adr_3_;
   wire FE_OCPN511_slv0_adr_3_;
   wire FE_OCPN510_slv0_adr_3_;
   wire FE_RN_15;
   wire FE_RN_14;
   wire FE_RN_13;
   wire FE_OCPN505_n2304;
   wire FE_UNCONNECTED_27;
   wire FE_UNCONNECTED_26;
   wire FE_UNCONNECTED_25;
   wire FE_UNCONNECTED_24;
   wire FE_UNCONNECTED_23;
   wire FE_UNCONNECTED_22;
   wire FE_RN_12;
   wire FE_RN_11;
   wire FE_RN_5;
   wire FE_OCPN481_n2343;
   wire FE_OCPN480_n1573;
   wire FE_OCPN479_n1573;
   wire FE_OCPN478_n1573;
   wire FE_RN_9;
   wire FE_OCPN464_n1521;
   wire FE_OCPN463_n1521;
   wire FE_OCPN462_n1521;
   wire FE_RN_52_0;
   wire FE_RN_51_0;
   wire FE_RN_50_0;
   wire FE_RN_8;
   wire FE_RN_7;
   wire FE_RN_49_0;
   wire FE_RN_47_0;
   wire FE_RN_46_0;
   wire FE_RN_44_0;
   wire FE_OCPN444_slv0_adr_8_;
   wire FE_OCPN443_slv0_adr_8_;
   wire FE_OCPN442_slv0_adr_8_;
   wire FE_RN_43_0;
   wire FE_RN_42_0;
   wire FE_RN_41_0;
   wire FE_UNCONNECTED_21;
   wire FE_UNCONNECTED_20;
   wire FE_UNCONNECTED_19;
   wire FE_UNCONNECTED_18;
   wire FE_OFN427_wb0_ack_i;
   wire FE_OFN426_wb0_ack_i;
   wire FE_UNCONNECTED_17;
   wire FE_UNCONNECTED_16;
   wire FE_UNCONNECTED_15;
   wire FE_UNCONNECTED_14;
   wire FE_UNCONNECTED_13;
   wire FE_UNCONNECTED_12;
   wire FE_RN_40_0;
   wire FE_RN_39_0;
   wire FE_RN_38_0;
   wire FE_RN_37_0;
   wire FE_RN_36_0;
   wire FE_RN_35_0;
   wire FE_RN_34_0;
   wire FE_OCPN403_n2346;
   wire FE_OCPN402_n2346;
   wire FE_UNCONNECTED_11;
   wire FE_UNCONNECTED_10;
   wire FE_UNCONNECTED_9;
   wire FE_UNCONNECTED_8;
   wire FE_UNCONNECTED_7;
   wire FE_OCPN385_n1579;
   wire FE_OCPN384_n1579;
   wire FE_OCPN383_n1512;
   wire FE_RN_33_0;
   wire FE_RN_31_0;
   wire FE_RN_4;
   wire FE_RN_30_0;
   wire FE_RN_29_0;
   wire FE_RN_28_0;
   wire FE_RN_27_0;
   wire FE_RN_26_0;
   wire FE_RN_25_0;
   wire FE_RN_24_0;
   wire FE_RN_23_0;
   wire FE_RN_22_0;
   wire FE_OCPN370_n2194;
   wire FE_OCPN368_n2194;
   wire FE_OCPN367_n2194;
   wire FE_OCPN366_n2194;
   wire FE_OCPN365_n2194;
   wire FE_OCPN363_n2194;
   wire FE_UNCONNECTED_6;
   wire FE_UNCONNECTED_5;
   wire FE_UNCONNECTED_4;
   wire FE_UNCONNECTED_3;
   wire FE_UNCONNECTED_2;
   wire FE_UNCONNECTED_1;
   wire FE_RN_21_0;
   wire FE_RN_1;
   wire FE_RN_20_0;
   wire FE_RN_19_0;
   wire FE_OCPN277_wb0_cyc_o;
   wire FE_OCPN284_wb0_cyc_o;
   wire FE_OCPN280_wb0_cyc_o;
   wire FE_RN_15_0;
   wire FE_RN_13_0;
   wire FE_OCPN200_n2156;
   wire FE_OCPN192_slv0_adr_9_;
   wire FE_RN_12_0;
   wire FE_RN_11_0;
   wire FE_RN_9_0;
   wire FE_RN_7_0;
   wire FE_OCPN186_n1893;
   wire FE_OCPN180_n1521;
   wire FE_OCPN179_n1521;
   wire FE_OCPN178_n1521;
   wire FE_OCPN176_n1521;
   wire FE_RN_2;
   wire FE_OCPN171_n2346;
   wire FE_OCPN170_n2346;
   wire FE_OCPN169_n2346;
   wire FE_OCPN167_n2346;
   wire FE_OCPN166_n2346;
   wire FE_OCPN165_n2346;
   wire FE_OCPN163_n2346;
   wire FE_OCPN139_slv0_adr_2_;
   wire FE_OCPN138_slv0_adr_2_;
   wire FE_OCPN137_slv0_adr_2_;
   wire FE_OCPN129_n2007;
   wire FE_OCPN126_FE_RN_;
   wire FE_OCPN124_FE_RN_;
   wire FE_OCPN122_FE_RN_;
   wire FE_OCPN120_FE_RN_;
   wire FE_OCPN106_slv0_adr_2_;
   wire FE_RN_;
   wire FE_OCPN80_n1919;
   wire FE_OCPN79_n2056;
   wire FE_OCPN78_n2056;
   wire FE_RN_5_0;
   wire FE_RN_2_0;
   wire FE_RN_0_0;
   wire FE_UNCONNECTED_0;
   wire slv0_re;
   wire slv0_we;
   wire ndnr_0_;
   wire slv1_re;
   wire slv1_we;
   wire u0_N3074;
   wire u0_int_maskb_0_;
   wire u0_int_maskb_1_;
   wire u0_int_maskb_2_;
   wire u0_int_maskb_3_;
   wire u0_int_maskb_4_;
   wire u0_int_maskb_5_;
   wire u0_int_maskb_6_;
   wire u0_int_maskb_7_;
   wire u0_int_maskb_8_;
   wire u0_int_maskb_9_;
   wire u0_int_maskb_10_;
   wire u0_int_maskb_11_;
   wire u0_int_maskb_12_;
   wire u0_int_maskb_13_;
   wire u0_int_maskb_14_;
   wire u0_int_maskb_15_;
   wire u0_int_maskb_16_;
   wire u0_int_maskb_17_;
   wire u0_int_maskb_18_;
   wire u0_int_maskb_19_;
   wire u0_int_maskb_20_;
   wire u0_int_maskb_21_;
   wire u0_int_maskb_22_;
   wire u0_int_maskb_23_;
   wire u0_int_maskb_24_;
   wire u0_int_maskb_25_;
   wire u0_int_maskb_26_;
   wire u0_int_maskb_27_;
   wire u0_int_maskb_28_;
   wire u0_int_maskb_29_;
   wire u0_int_maskb_30_;
   wire u0_int_maska_0_;
   wire u0_int_maska_1_;
   wire u0_int_maska_2_;
   wire u0_int_maska_3_;
   wire u0_int_maska_4_;
   wire u0_int_maska_5_;
   wire u0_int_maska_6_;
   wire u0_int_maska_7_;
   wire u0_int_maska_8_;
   wire u0_int_maska_9_;
   wire u0_int_maska_10_;
   wire u0_int_maska_11_;
   wire u0_int_maska_12_;
   wire u0_int_maska_13_;
   wire u0_int_maska_14_;
   wire u0_int_maska_15_;
   wire u0_int_maska_16_;
   wire u0_int_maska_17_;
   wire u0_int_maska_18_;
   wire u0_int_maska_19_;
   wire u0_int_maska_20_;
   wire u0_int_maska_21_;
   wire u0_int_maska_22_;
   wire u0_int_maska_23_;
   wire u0_int_maska_24_;
   wire u0_int_maska_25_;
   wire u0_int_maska_26_;
   wire u0_int_maska_27_;
   wire u0_int_maska_28_;
   wire u0_int_maska_29_;
   wire u0_int_maska_30_;
   wire u1_N1032;
   wire u3_u1_N5;
   wire u3_u1_N4;
   wire u3_u1_N3;
   wire u3_u1_rf_ack;
   wire u4_u1_N4;
   wire u4_u1_N3;
   wire u4_u1_rf_ack;
   wire n498;
   wire n499;
   wire n500;
   wire n501;
   wire n502;
   wire n503;
   wire n504;
   wire n505;
   wire n506;
   wire n507;
   wire n508;
   wire n509;
   wire n510;
   wire n511;
   wire n512;
   wire n513;
   wire n514;
   wire n515;
   wire n516;
   wire n517;
   wire n518;
   wire n519;
   wire n520;
   wire n521;
   wire n522;
   wire n523;
   wire n524;
   wire n525;
   wire n526;
   wire n527;
   wire n528;
   wire n529;
   wire n530;
   wire n531;
   wire n532;
   wire n533;
   wire n534;
   wire n535;
   wire n536;
   wire n537;
   wire n538;
   wire n539;
   wire n540;
   wire n541;
   wire n542;
   wire n543;
   wire n544;
   wire n545;
   wire n546;
   wire n547;
   wire n548;
   wire n549;
   wire n550;
   wire n551;
   wire n552;
   wire n553;
   wire n554;
   wire n555;
   wire n556;
   wire n557;
   wire n558;
   wire n559;
   wire n560;
   wire n570;
   wire n571;
   wire n581;
   wire n583;
   wire n585;
   wire n587;
   wire n589;
   wire n591;
   wire n593;
   wire n595;
   wire n597;
   wire n599;
   wire n601;
   wire n603;
   wire n605;
   wire n607;
   wire n609;
   wire n611;
   wire n613;
   wire n615;
   wire n617;
   wire n619;
   wire n621;
   wire n623;
   wire n625;
   wire n627;
   wire n629;
   wire n631;
   wire n633;
   wire n635;
   wire n637;
   wire n639;
   wire n641;
   wire n643;
   wire n645;
   wire n647;
   wire n649;
   wire n651;
   wire n653;
   wire n655;
   wire n657;
   wire n659;
   wire n661;
   wire n663;
   wire n665;
   wire n667;
   wire n669;
   wire n671;
   wire n673;
   wire n675;
   wire n677;
   wire n679;
   wire n681;
   wire n683;
   wire n685;
   wire n687;
   wire n689;
   wire n691;
   wire n693;
   wire n695;
   wire n697;
   wire n699;
   wire n701;
   wire n703;
   wire n705;
   wire n707;
   wire n709;
   wire n711;
   wire n713;
   wire n715;
   wire n717;
   wire n719;
   wire n721;
   wire n731;
   wire n732;
   wire n733;
   wire n734;
   wire n742;
   wire n745;
   wire n746;
   wire n747;
   wire n748;
   wire n749;
   wire n750;
   wire n751;
   wire n752;
   wire n753;
   wire n754;
   wire n755;
   wire n756;
   wire n757;
   wire n758;
   wire n759;
   wire n760;
   wire n761;
   wire n762;
   wire n763;
   wire n764;
   wire n765;
   wire n766;
   wire n767;
   wire n800;
   wire n801;
   wire n802;
   wire n803;
   wire n804;
   wire n805;
   wire n806;
   wire n807;
   wire n808;
   wire n809;
   wire n810;
   wire n811;
   wire n812;
   wire n813;
   wire n814;
   wire n815;
   wire n816;
   wire n817;
   wire n818;
   wire n819;
   wire n820;
   wire n821;
   wire n822;
   wire n823;
   wire n824;
   wire n825;
   wire n826;
   wire n827;
   wire n828;
   wire n829;
   wire n830;
   wire n831;
   wire n893;
   wire n1414;
   wire n1416;
   wire n1417;
   wire n1418;
   wire n1419;
   wire n1424;
   wire n1425;
   wire n1426;
   wire n1428;
   wire n1438;
   wire n1442;
   wire n1467;
   wire n1468;
   wire n1469;
   wire n1470;
   wire n1471;
   wire n1472;
   wire n1473;
   wire n1474;
   wire n1476;
   wire n1477;
   wire n1478;
   wire n1479;
   wire n1480;
   wire n1481;
   wire n1484;
   wire n1488;
   wire n1489;
   wire n1490;
   wire n1491;
   wire n1492;
   wire n1493;
   wire n1494;
   wire n1495;
   wire n1496;
   wire n1497;
   wire n1498;
   wire n1499;
   wire n1500;
   wire n1501;
   wire n1502;
   wire n1503;
   wire n1504;
   wire n1505;
   wire n1506;
   wire n1507;
   wire n1510;
   wire n1512;
   wire n1513;
   wire n1515;
   wire n1516;
   wire n1517;
   wire n1521;
   wire n1522;
   wire n1523;
   wire n1524;
   wire n1525;
   wire n1526;
   wire n1527;
   wire n1528;
   wire n1529;
   wire n1530;
   wire n1531;
   wire n1532;
   wire n1533;
   wire n1534;
   wire n1535;
   wire n1536;
   wire n1537;
   wire n1541;
   wire n1542;
   wire n1543;
   wire n1544;
   wire n1545;
   wire n1546;
   wire n1547;
   wire n1548;
   wire n1549;
   wire n1550;
   wire n1551;
   wire n1552;
   wire n1553;
   wire n1554;
   wire n1555;
   wire n1556;
   wire n1557;
   wire n1558;
   wire n1559;
   wire n1560;
   wire n1561;
   wire n1562;
   wire n1563;
   wire n1564;
   wire n1566;
   wire n1573;
   wire n1574;
   wire n1575;
   wire n1576;
   wire n1577;
   wire n1579;
   wire n1580;
   wire n1581;
   wire n1582;
   wire n1583;
   wire n1584;
   wire n1585;
   wire n1591;
   wire n1595;
   wire n1597;
   wire n1605;
   wire n1607;
   wire n1608;
   wire n1609;
   wire n1610;
   wire n1611;
   wire n1612;
   wire n1613;
   wire n1614;
   wire n1615;
   wire n1616;
   wire n1617;
   wire n1618;
   wire n1619;
   wire n1620;
   wire n1621;
   wire n1622;
   wire n1623;
   wire n1624;
   wire n1625;
   wire n1626;
   wire n1628;
   wire n1629;
   wire n1630;
   wire n1631;
   wire n1632;
   wire n1633;
   wire n1634;
   wire n1635;
   wire n1636;
   wire n1637;
   wire n1638;
   wire n1639;
   wire n1641;
   wire n1642;
   wire n1643;
   wire n1644;
   wire n1645;
   wire n1646;
   wire n1647;
   wire n1648;
   wire n1649;
   wire n1650;
   wire n1651;
   wire n1652;
   wire n1653;
   wire n1654;
   wire n1655;
   wire n1656;
   wire n1657;
   wire n1658;
   wire n1659;
   wire n1660;
   wire n1661;
   wire n1662;
   wire n1663;
   wire n1664;
   wire n1665;
   wire n1666;
   wire n1667;
   wire n1668;
   wire n1669;
   wire n1670;
   wire n1671;
   wire n1672;
   wire n1673;
   wire n1674;
   wire n1675;
   wire n1676;
   wire n1677;
   wire n1678;
   wire n1679;
   wire n1681;
   wire n1682;
   wire n1683;
   wire n1684;
   wire n1685;
   wire n1686;
   wire n1687;
   wire n1688;
   wire n1689;
   wire n1690;
   wire n1691;
   wire n1692;
   wire n1693;
   wire n1694;
   wire n1695;
   wire n1696;
   wire n1697;
   wire n1698;
   wire n1699;
   wire n1700;
   wire n1701;
   wire n1702;
   wire n1703;
   wire n1704;
   wire n1705;
   wire n1706;
   wire n1707;
   wire n1708;
   wire n1709;
   wire n1710;
   wire n1711;
   wire n1712;
   wire n1713;
   wire n1714;
   wire n1715;
   wire n1716;
   wire n1717;
   wire n1718;
   wire n1719;
   wire n1720;
   wire n1721;
   wire n1722;
   wire n1723;
   wire n1724;
   wire n1725;
   wire n1726;
   wire n1727;
   wire n1728;
   wire n1729;
   wire n1730;
   wire n1731;
   wire n1732;
   wire n1733;
   wire n1734;
   wire n1735;
   wire n1736;
   wire n1737;
   wire n1738;
   wire n1739;
   wire n1740;
   wire n1741;
   wire n1742;
   wire n1743;
   wire n1744;
   wire n1745;
   wire n1746;
   wire n1747;
   wire n1750;
   wire n1751;
   wire n1752;
   wire n1753;
   wire n1754;
   wire n1755;
   wire n1756;
   wire n1757;
   wire n1758;
   wire n1759;
   wire n1760;
   wire n1761;
   wire n1762;
   wire n1763;
   wire n1764;
   wire n1765;
   wire n1766;
   wire n1767;
   wire n1768;
   wire n1769;
   wire n1770;
   wire n1771;
   wire n1772;
   wire n1773;
   wire n1774;
   wire n1775;
   wire n1776;
   wire n1777;
   wire n1778;
   wire n1779;
   wire n1780;
   wire n1781;
   wire n1782;
   wire n1783;
   wire n1784;
   wire n1785;
   wire n1786;
   wire n1787;
   wire n1788;
   wire n1789;
   wire n1790;
   wire n1791;
   wire n1792;
   wire n1793;
   wire n1794;
   wire n1795;
   wire n1796;
   wire n1797;
   wire n1798;
   wire n1799;
   wire n1800;
   wire n1801;
   wire n1802;
   wire n1803;
   wire n1804;
   wire n1805;
   wire n1806;
   wire n1807;
   wire n1808;
   wire n1809;
   wire n1810;
   wire n1811;
   wire n1812;
   wire n1813;
   wire n1814;
   wire n1815;
   wire n1816;
   wire n1817;
   wire n1818;
   wire n1819;
   wire n1820;
   wire n1821;
   wire n1822;
   wire n1823;
   wire n1824;
   wire n1825;
   wire n1826;
   wire n1827;
   wire n1828;
   wire n1829;
   wire n1830;
   wire n1831;
   wire n1832;
   wire n1833;
   wire n1834;
   wire n1835;
   wire n1836;
   wire n1837;
   wire n1838;
   wire n1839;
   wire n1840;
   wire n1841;
   wire n1842;
   wire n1843;
   wire n1844;
   wire n1845;
   wire n1846;
   wire n1847;
   wire n1848;
   wire n1849;
   wire n1850;
   wire n1851;
   wire n1852;
   wire n1853;
   wire n1854;
   wire n1855;
   wire n1856;
   wire n1857;
   wire n1858;
   wire n1859;
   wire n1860;
   wire n1861;
   wire n1862;
   wire n1863;
   wire n1864;
   wire n1865;
   wire n1866;
   wire n1867;
   wire n1868;
   wire n1870;
   wire n1871;
   wire n1872;
   wire n1873;
   wire n1874;
   wire n1875;
   wire n1876;
   wire n1877;
   wire n1878;
   wire n1879;
   wire n1880;
   wire n1881;
   wire n1882;
   wire n1883;
   wire n1884;
   wire n1885;
   wire n1886;
   wire n1887;
   wire n1888;
   wire n1889;
   wire n1890;
   wire n1891;
   wire n1892;
   wire n1894;
   wire n1895;
   wire n1896;
   wire n1897;
   wire n1898;
   wire n1899;
   wire n1900;
   wire n1901;
   wire n1904;
   wire n1905;
   wire n1906;
   wire n1907;
   wire n1908;
   wire n1909;
   wire n1910;
   wire n1911;
   wire n1912;
   wire n1913;
   wire n1914;
   wire n1915;
   wire n1916;
   wire n1917;
   wire n1918;
   wire n1919;
   wire n1920;
   wire n1921;
   wire n1923;
   wire n1924;
   wire n1925;
   wire n1926;
   wire n1927;
   wire n1928;
   wire n1929;
   wire n1930;
   wire n1931;
   wire n1932;
   wire n1933;
   wire n1934;
   wire n1935;
   wire n1936;
   wire n1937;
   wire n1938;
   wire n1939;
   wire n1940;
   wire n1941;
   wire n1942;
   wire n1943;
   wire n1944;
   wire n1945;
   wire n1946;
   wire n1947;
   wire n1948;
   wire n1949;
   wire n1950;
   wire n1951;
   wire n1952;
   wire n1953;
   wire n1954;
   wire n1955;
   wire n1956;
   wire n1957;
   wire n1958;
   wire n1959;
   wire n1960;
   wire n1961;
   wire n1962;
   wire n1963;
   wire n1964;
   wire n1965;
   wire n1966;
   wire n1967;
   wire n1968;
   wire n1969;
   wire n1970;
   wire n1971;
   wire n1972;
   wire n1973;
   wire n1974;
   wire n1975;
   wire n1976;
   wire n1977;
   wire n1978;
   wire n1979;
   wire n1980;
   wire n1981;
   wire n1982;
   wire n1983;
   wire n1984;
   wire n1985;
   wire n1986;
   wire n1987;
   wire n1988;
   wire n1989;
   wire n1990;
   wire n1991;
   wire n1992;
   wire n1993;
   wire n1994;
   wire n1995;
   wire n1996;
   wire n1997;
   wire n1998;
   wire n1999;
   wire n2000;
   wire n2001;
   wire n2002;
   wire n2003;
   wire n2004;
   wire n2005;
   wire n2006;
   wire n2007;
   wire n2008;
   wire n2009;
   wire n2010;
   wire n2011;
   wire n2012;
   wire n2013;
   wire n2014;
   wire n2015;
   wire n2016;
   wire n2017;
   wire n2018;
   wire n2019;
   wire n2020;
   wire n2021;
   wire n2022;
   wire n2023;
   wire n2024;
   wire n2025;
   wire n2026;
   wire n2027;
   wire n2028;
   wire n2029;
   wire n2030;
   wire n2031;
   wire n2032;
   wire n2033;
   wire n2034;
   wire n2035;
   wire n2036;
   wire n2037;
   wire n2038;
   wire n2039;
   wire n2040;
   wire n2041;
   wire n2042;
   wire n2043;
   wire n2044;
   wire n2045;
   wire n2046;
   wire n2047;
   wire n2048;
   wire n2049;
   wire n2050;
   wire n2051;
   wire n2052;
   wire n2053;
   wire n2054;
   wire n2055;
   wire n2056;
   wire n2060;
   wire n2063;
   wire n2068;
   wire n2069;
   wire n2070;
   wire n2071;
   wire n2072;
   wire n2073;
   wire n2074;
   wire n2075;
   wire n2076;
   wire n2077;
   wire n2078;
   wire n2079;
   wire n2080;
   wire n2081;
   wire n2082;
   wire n2083;
   wire n2084;
   wire n2085;
   wire n2086;
   wire n2087;
   wire n2088;
   wire n2089;
   wire n2090;
   wire n2091;
   wire n2092;
   wire n2093;
   wire n2094;
   wire n2095;
   wire n2096;
   wire n2097;
   wire n2098;
   wire n2099;
   wire n2100;
   wire n2101;
   wire n2102;
   wire n2103;
   wire n2104;
   wire n2105;
   wire n2106;
   wire n2107;
   wire n2108;
   wire n2109;
   wire n2110;
   wire n2111;
   wire n2112;
   wire n2113;
   wire n2114;
   wire n2115;
   wire n2116;
   wire n2117;
   wire n2118;
   wire n2119;
   wire n2120;
   wire n2121;
   wire n2122;
   wire n2123;
   wire n2124;
   wire n2125;
   wire n2126;
   wire n2127;
   wire n2128;
   wire n2129;
   wire n2130;
   wire n2131;
   wire n2132;
   wire n2133;
   wire n2134;
   wire n2135;
   wire n2136;
   wire n2137;
   wire n2138;
   wire n2139;
   wire n2140;
   wire n2141;
   wire n2142;
   wire n2143;
   wire n2144;
   wire n2145;
   wire n2146;
   wire n2147;
   wire n2148;
   wire n2149;
   wire n2150;
   wire n2151;
   wire n2152;
   wire n2153;
   wire n2154;
   wire n2155;
   wire n2156;
   wire n2157;
   wire n2158;
   wire n2159;
   wire n2160;
   wire n2161;
   wire n2162;
   wire n2163;
   wire n2164;
   wire n2165;
   wire n2166;
   wire n2167;
   wire n2168;
   wire n2169;
   wire n2170;
   wire n2171;
   wire n2172;
   wire n2173;
   wire n2174;
   wire n2175;
   wire n2176;
   wire n2177;
   wire n2178;
   wire n2179;
   wire n2180;
   wire n2181;
   wire n2182;
   wire n2183;
   wire n2184;
   wire n2185;
   wire n2186;
   wire n2187;
   wire n2188;
   wire n2189;
   wire n2190;
   wire n2191;
   wire n2192;
   wire n2193;
   wire n2194;
   wire n2195;
   wire n2196;
   wire n2197;
   wire n2198;
   wire n2199;
   wire n2200;
   wire n2201;
   wire n2202;
   wire n2203;
   wire n2204;
   wire n2205;
   wire n2206;
   wire n2207;
   wire n2208;
   wire n2209;
   wire n2210;
   wire n2211;
   wire n2212;
   wire n2213;
   wire n2214;
   wire n2215;
   wire n2216;
   wire n2217;
   wire n2218;
   wire n2219;
   wire n2220;
   wire n2221;
   wire n2222;
   wire n2223;
   wire n2224;
   wire n2225;
   wire n2226;
   wire n2227;
   wire n2228;
   wire n2230;
   wire n2231;
   wire n2232;
   wire n2233;
   wire n2234;
   wire n2235;
   wire n2236;
   wire n2237;
   wire n2238;
   wire n2239;
   wire n2240;
   wire n2241;
   wire n2242;
   wire n2243;
   wire n2244;
   wire n2245;
   wire n2246;
   wire n2247;
   wire n2248;
   wire n2249;
   wire n2250;
   wire n2251;
   wire n2252;
   wire n2253;
   wire n2254;
   wire n2255;
   wire n2256;
   wire n2257;
   wire n2258;
   wire n2259;
   wire n2260;
   wire n2261;
   wire n2262;
   wire n2263;
   wire n2264;
   wire n2265;
   wire n2266;
   wire n2267;
   wire n2268;
   wire n2269;
   wire n2270;
   wire n2271;
   wire n2272;
   wire n2273;
   wire n2274;
   wire n2275;
   wire n2276;
   wire n2277;
   wire n2278;
   wire n2279;
   wire n2280;
   wire n2281;
   wire n2282;
   wire n2284;
   wire n2285;
   wire n2286;
   wire n2287;
   wire n2288;
   wire n2289;
   wire n2292;
   wire n2293;
   wire n2294;
   wire n2295;
   wire n2296;
   wire n2297;
   wire n2299;
   wire n2300;
   wire n2301;
   wire n2302;
   wire n2303;
   wire n2304;
   wire n2305;
   wire n2306;
   wire n2307;
   wire n2308;
   wire n2309;
   wire n2310;
   wire n2311;
   wire n2312;
   wire n2313;
   wire n2314;
   wire n2315;
   wire n2316;
   wire n2317;
   wire n2318;
   wire n2319;
   wire n2320;
   wire n2321;
   wire n2322;
   wire n2323;
   wire n2324;
   wire n2325;
   wire n2326;
   wire n2327;
   wire n2328;
   wire n2329;
   wire n2330;
   wire n2331;
   wire n2332;
   wire n2333;
   wire n2334;
   wire n2335;
   wire n2336;
   wire n2337;
   wire n2338;
   wire n2339;
   wire n2340;
   wire n2341;
   wire n2342;
   wire n2343;
   wire n2345;
   wire n2346;
   wire n2347;
   wire n2349;
   wire n2350;
   wire n2351;
   wire n2352;
   wire n2353;
   wire n2355;
   wire n2356;
   wire n2357;
   wire n2358;
   wire n2359;
   wire n2360;
   wire n2361;
   wire n2362;
   wire n2363;
   wire n2364;
   wire n2365;
   wire n2366;
   wire n2367;
   wire n2368;
   wire n2369;
   wire n2370;
   wire n2371;
   wire n2372;
   wire n2373;
   wire n2374;
   wire n2375;
   wire n2376;
   wire n2377;
   wire n2378;
   wire n2379;
   wire n2380;
   wire n2381;
   wire n2382;
   wire n2383;
   wire n2384;
   wire n2385;
   wire n2386;
   wire n2387;
   wire n2388;
   wire n2389;
   wire n2390;
   wire n2391;
   wire n2392;
   wire n2393;
   wire n2394;
   wire n2395;
   wire n2396;
   wire n2397;
   wire n2398;
   wire n2399;
   wire n2400;
   wire n2401;
   wire n2402;
   wire n2403;
   wire n2404;
   wire n2405;
   wire n2406;
   wire n2407;
   wire n2408;
   wire n2409;
   wire n2410;
   wire n2411;
   wire n2412;
   wire n2413;
   wire n2414;
   wire n2415;
   wire n2416;
   wire n2417;
   wire n2418;
   wire n2419;
   wire n2420;
   wire n2421;
   wire n2422;
   wire n2423;
   wire n2424;
   wire n2425;
   wire n2426;
   wire n2427;
   wire n2428;
   wire n2429;
   wire n2430;
   wire n2431;
   wire n2432;
   wire n2433;
   wire n2434;
   wire n2435;
   wire n2436;
   wire n2437;
   wire n2438;
   wire n2439;
   wire n2440;
   wire n2441;
   wire n2442;
   wire n2443;
   wire n2444;
   wire n2445;
   wire n2446;
   wire n2448;
   wire n2449;
   wire n2450;
   wire n2451;
   wire n2452;
   wire n2453;
   wire n2454;
   wire n2455;
   wire n2456;
   wire n2457;
   wire n2458;
   wire n2459;
   wire n2460;
   wire n2461;
   wire n2462;
   wire n2463;
   wire n2464;
   wire n2465;
   wire n2466;
   wire n2469;
   wire n2470;
   wire n2471;
   wire n2472;
   wire n2473;
   wire n2474;
   wire n2475;
   wire n2476;
   wire n2477;
   wire n2478;
   wire n2479;
   wire n2480;
   wire n2481;
   wire n2482;
   wire n2483;
   wire n2484;
   wire n2485;
   wire n2486;
   wire n2487;
   wire n2488;
   wire n2489;
   wire n2490;
   wire n2491;
   wire n2492;
   wire n2493;
   wire n2494;
   wire n2495;
   wire n2496;
   wire n2497;
   wire n2498;
   wire n2499;
   wire n2500;
   wire n2501;
   wire [9:2] slv0_adr;
   wire [31:0] slv0_dout;
   wire [31:0] slv0_din;
   wire [21:0] ch0_csr;
   wire [26:0] ch0_txsz;
   wire [31:2] ch0_adr0;
   wire [31:2] ch0_adr1;
   wire [31:0] de_csr;

   assign dma_ack_o[0] = 1'b0 ;

   in01f20 FE_OCPC676_n1580 (.o(FE_OCPN676_n1580),
	.a(n1580));
   in01s08 FE_OCPC675_n1580 (.o(FE_OCPN675_n1580),
	.a(n1580));
   in01f02 FE_OCPC674_n2186 (.o(FE_OCPN674_n2186),
	.a(n2186));
   in01f20 FE_OCPC673_n1577 (.o(FE_OCPN673_n1577),
	.a(n1577));
   in01f08 FE_OCPC672_n1577 (.o(FE_OCPN672_n1577),
	.a(n1577));
   in01f20 FE_OCPC671_n2356 (.o(FE_OCPN671_n2356),
	.a(n2356));
   in01f20 FE_OCPC670_n2356 (.o(FE_OCPN670_n2356),
	.a(n2356));
   in01f80 FE_OCPC669_slv0_adr_4_ (.o(FE_OCPN669_slv0_adr_4_),
	.a(slv0_adr[4]));
   in01s02 FE_OCPC668_wb1_cyc_o (.o(FE_OCPN668_wb1_cyc_o),
	.a(FE_OCPN666_wb1_cyc_o));
   in01s06 FE_OCPC667_wb1_cyc_o (.o(FE_OCPN667_wb1_cyc_o),
	.a(FE_OCPN665_wb1_cyc_o));
   in01s10 FE_OCPC666_wb1_cyc_o (.o(FE_OCPN666_wb1_cyc_o),
	.a(FE_OCPN636_wb1_cyc_o));
   in01m04 FE_OCPC665_wb1_cyc_o (.o(FE_OCPN665_wb1_cyc_o),
	.a(FE_OCPN636_wb1_cyc_o));
   in01f20 FE_OCPC664_FE_RN_16 (.o(FE_OCPN664_FE_RN_16),
	.a(FE_RN_16));
   in01f04 FE_OCPC663_n1428 (.o(FE_OCPN663_n1428),
	.a(n1428));
   in01s10 FE_OCPC662_wb1_cyc_o (.o(wb1_cyc_o),
	.a(FE_OCPN660_wb1_cyc_o));
   in01s03 FE_OCPC661_wb1_cyc_o (.o(FE_OCPN661_wb1_cyc_o),
	.a(FE_OCPN660_wb1_cyc_o));
   in01s06 FE_OCPC660_wb1_cyc_o (.o(FE_OCPN660_wb1_cyc_o),
	.a(FE_OCPN659_wb1_cyc_o));
   in01s20 FE_OCPC658_wb1_cyc_o (.o(FE_OCPN658_wb1_cyc_o),
	.a(FE_OCPN655_wb1_cyc_o));
   in01s20 FE_OCPC657_wb1_cyc_o (.o(FE_OCPN657_wb1_cyc_o),
	.a(FE_OCPN655_wb1_cyc_o));
   in01s20 FE_OCPC656_wb1_cyc_o (.o(FE_OCPN656_wb1_cyc_o),
	.a(FE_OCPN655_wb1_cyc_o));
   in01s20 FE_OCPC655_wb1_cyc_o (.o(FE_OCPN655_wb1_cyc_o),
	.a(FE_OCPN625_wb1_cyc_o));
   in01s10 FE_OCPC651_wb1_cyc_o (.o(FE_OCPN651_wb1_cyc_o),
	.a(FE_OCPN634_wb1_cyc_o));
   in01m06 FE_OCPC643_wb1_cyc_o (.o(FE_OCPN643_wb1_cyc_o),
	.a(FE_OCPN632_wb1_cyc_o));
   in01s10 FE_OCPC642_wb1_cyc_o (.o(FE_OCPN642_wb1_cyc_o),
	.a(FE_OCPN632_wb1_cyc_o));
   in01m08 FE_OCPC636_wb1_cyc_o (.o(FE_OCPN636_wb1_cyc_o),
	.a(FE_OCPN659_wb1_cyc_o));
   in01s08 FE_OCPC634_wb1_cyc_o (.o(FE_OCPN634_wb1_cyc_o),
	.a(FE_OCPN659_wb1_cyc_o));
   in01s06 FE_OCPC633_wb1_cyc_o (.o(FE_OCPN633_wb1_cyc_o),
	.a(FE_OCPN659_wb1_cyc_o));
   in01s08 FE_OCPC632_wb1_cyc_o (.o(FE_OCPN632_wb1_cyc_o),
	.a(FE_OCPN659_wb1_cyc_o));
   in01s02 FE_OCPC631_wb1_cyc_o (.o(FE_OCPN631_wb1_cyc_o),
	.a(FE_OCPN659_wb1_cyc_o));
   in01s03 FE_OCPC630_wb1_cyc_o (.o(FE_OCPN630_wb1_cyc_o),
	.a(FE_OCPN659_wb1_cyc_o));
   in01s06 FE_OCPC629_wb1_cyc_o (.o(FE_OCPN629_wb1_cyc_o),
	.a(FE_OCPN659_wb1_cyc_o));
   in01s01 FE_OCPC628_wb1_cyc_o (.o(FE_OCPN628_wb1_cyc_o),
	.a(FE_OCPN659_wb1_cyc_o));
   in01s06 FE_OCPC627_wb1_cyc_o (.o(FE_OCPN627_wb1_cyc_o),
	.a(FE_OCPN659_wb1_cyc_o));
   in01m08 FE_OCPC626_wb1_cyc_o (.o(FE_OCPN626_wb1_cyc_o),
	.a(FE_OCPN659_wb1_cyc_o));
   in01s10 FE_OCPC625_wb1_cyc_o (.o(FE_OCPN625_wb1_cyc_o),
	.a(FE_OCPN659_wb1_cyc_o));
   in01s03 FE_OCPC624_wb1_cyc_o (.o(FE_OCPN624_wb1_cyc_o),
	.a(FE_OCPN659_wb1_cyc_o));
   in01m10 FE_OCPC622_n1516 (.o(FE_OCPN622_n1516),
	.a(FE_OCPN612_n1516));
   in01m04 FE_OCPC620_n1516 (.o(FE_OCPN620_n1516),
	.a(FE_OCPN612_n1516));
   in01m20 FE_OCPC619_n1513 (.o(FE_OCPN619_n1513),
	.a(n1513));
   in01m08 FE_OCPC618_n1591 (.o(FE_OCPN618_n1591),
	.a(n1591));
   in01f80 FE_OCPC617_slv0_adr_5_ (.o(FE_OCPN617_slv0_adr_5_),
	.a(slv0_adr[5]));
   na04m04 FE_RC_129_0 (.o(n2445),
	.d(n1560),
	.c(n1561),
	.b(n2215),
	.a(n2241));
   in01f04 FE_OCPC615_n1516 (.o(FE_OCPN615_n1516),
	.a(n1516));
   in01m06 FE_OCPC614_n1516 (.o(FE_OCPN614_n1516),
	.a(n1516));
   in01m10 FE_OCPC613_n1516 (.o(FE_OCPN613_n1516),
	.a(n1516));
   in01f20 FE_OCPC612_n1516 (.o(FE_OCPN612_n1516),
	.a(n1516));
   no03f08 FE_RC_128_0 (.o(n1965),
	.c(n1962),
	.b(n1963),
	.a(FE_OCPN673_n1577));
   ao22s04 FE_RC_127_0 (.o(n1561),
	.d(n2356),
	.c(ch0_adr1[20]),
	.b(FE_OCPN560_n2357),
	.a(ch0_adr0[20]));
   in01f20 FE_OCPC611_slv0_adr_3_ (.o(FE_OCPN611_slv0_adr_3_),
	.a(FE_OCPN609_slv0_adr_3_));
   in01f20 FE_OCPC610_slv0_adr_3_ (.o(FE_OCPN610_slv0_adr_3_),
	.a(FE_OCPN609_slv0_adr_3_));
   in01f20 FE_OCPC609_slv0_adr_3_ (.o(FE_OCPN609_slv0_adr_3_),
	.a(slv0_adr[3]));
   in01s01 FE_RC_126_0 (.o(FE_RN_59_0),
	.a(slv1_re));
   in01s01 FE_RC_125_0 (.o(FE_RN_60_0),
	.a(slv1_we));
   na02s01 FE_RC_124_0 (.o(FE_RN_61_0),
	.b(FE_RN_60_0),
	.a(FE_RN_59_0));
   na02s01 FE_RC_123_0 (.o(n1728),
	.b(n1727),
	.a(FE_RN_61_0));
   na04s10 FE_RC_122_0 (.o(n1597),
	.d(n2366),
	.c(n2367),
	.b(n2365),
	.a(n2368));
   oa22m02 FE_RC_121_0 (.o(n538),
	.d(FE_OCPN383_n1512),
	.c(n2020),
	.b(n1591),
	.a(n2023));
   in01f10 FE_OCPC566_n2357 (.o(FE_OCPN566_n2357),
	.a(FE_OCPN559_n2357));
   in01m08 FE_OCPC565_n2357 (.o(FE_OCPN565_n2357),
	.a(FE_OCPN559_n2357));
   in01f08 FE_OCPC562_n2357 (.o(FE_OCPN562_n2357),
	.a(FE_OCPN558_n2357));
   in01m06 FE_OCPC561_n2357 (.o(FE_OCPN561_n2357),
	.a(FE_OCPN558_n2357));
   in01s08 FE_OCPC560_n2357 (.o(FE_OCPN560_n2357),
	.a(n2357));
   in01f10 FE_OCPC559_n2357 (.o(FE_OCPN559_n2357),
	.a(n2357));
   in01m08 FE_OCPC558_n2357 (.o(FE_OCPN558_n2357),
	.a(n2357));
   na02f20 U1882_dup (.o(FE_RN_18),
	.b(n1484),
	.a(FE_OCPN163_n2346));
   na03f06 FE_RC_120_0 (.o(n2461),
	.c(n1947),
	.b(n1948),
	.a(n1946));
   na04m80 FE_RC_119_0 (.o(n1626),
	.d(FE_OCPN511_slv0_adr_3_),
	.c(FE_OCPN139_slv0_adr_2_),
	.b(FE_OCPN669_slv0_adr_4_),
	.a(slv0_we));
   in01s01 FE_RC_118_0 (.o(FE_RN_56_0),
	.a(u0_int_maska_13_));
   in01m10 FE_RC_117_0 (.o(FE_RN_57_0),
	.a(n2343));
   no02m08 FE_RC_116_0 (.o(FE_RN_58_0),
	.b(FE_RN_57_0),
	.a(FE_RN_56_0));
   no02f08 FE_RC_115_0 (.o(n2091),
	.b(FE_RN_58_0),
	.a(n2090));
   ao22f08 FE_RC_114_0 (.o(n2269),
	.d(FE_OCPN124_FE_RN_),
	.c(u0_int_maska_24_),
	.b(FE_OCPN552_n1424),
	.a(u0_int_maskb_24_));
   in01m10 FE_OCPC554_n1529 (.o(FE_OCPN554_n1529),
	.a(FE_OCPN553_n1529));
   in01f08 FE_OCPC553_n1529 (.o(FE_OCPN553_n1529),
	.a(n1529));
   in01s01 FE_RC_113_0 (.o(FE_RN_53_0),
	.a(u0_int_maska_26_));
   in01f10 FE_RC_112_0 (.o(FE_RN_54_0),
	.a(FE_OCPN124_FE_RN_));
   no02f08 FE_RC_111_0 (.o(FE_RN_55_0),
	.b(FE_RN_54_0),
	.a(FE_RN_53_0));
   no02f06 FE_RC_110_0 (.o(n2299),
	.b(FE_RN_55_0),
	.a(n2297));
   in01f20 FE_OCPC552_n1424 (.o(FE_OCPN552_n1424),
	.a(n1424));
   in01s04 FE_OCPC549_n1529 (.o(FE_OCPN549_n1529),
	.a(n1529));
   in01s06 FE_OCPC547_n1529 (.o(FE_OCPN547_n1529),
	.a(FE_OCPN549_n1529));
   oa22f08 FE_RC_109_0 (.o(n1979),
	.d(FE_RN_14),
	.c(n1977),
	.b(FE_OCPN670_n2356),
	.a(n1978));
   in01m10 FE_OCPC545_n2159 (.o(FE_OCPN545_n2159),
	.a(n2159));
   in01f20 FE_OCPC544_n2159 (.o(FE_OCPN544_n2159),
	.a(n2159));
   oa22m06 FE_RC_108_0 (.o(n2349),
	.d(n2345),
	.c(FE_OCPN169_n2346),
	.b(FE_OCPN670_n2356),
	.a(n2347));
   oa22f08 FE_RC_107_0 (.o(n2093),
	.d(n2091),
	.c(FE_OCPN170_n2346),
	.b(FE_OCPN671_n2356),
	.a(n2092));
   in01s10 FE_OCPC540_n1595 (.o(FE_OCPN540_n1595),
	.a(n1595));
   in01m08 FE_OCPC539_n1595 (.o(FE_OCPN539_n1595),
	.a(n1595));
   in01m10 FE_OCPC538_n1595 (.o(FE_OCPN538_n1595),
	.a(n1595));
   in01s04 FE_OCPC537_n1595 (.o(FE_OCPN537_n1595),
	.a(n1595));
   in01s10 FE_OCPC528_n1597 (.o(FE_OCPN528_n1597),
	.a(n1597));
   no02s20 U2188_dup (.o(FE_RN_17),
	.b(n1725),
	.a(n2364));
   no02f80 U2938_dup_dup (.o(FE_RN_16),
	.b(slv0_adr[6]),
	.a(slv0_adr[7]));
   in01f20 FE_OCPC514_slv0_adr_3_ (.o(FE_OCPN514_slv0_adr_3_),
	.a(FE_OCPN510_slv0_adr_3_));
   in01f20 FE_OCPC513_slv0_adr_3_ (.o(FE_OCPN513_slv0_adr_3_),
	.a(FE_OCPN510_slv0_adr_3_));
   in01f20 FE_OCPC512_slv0_adr_3_ (.o(FE_OCPN512_slv0_adr_3_),
	.a(slv0_adr[3]));
   in01f80 FE_OCPC511_slv0_adr_3_ (.o(FE_OCPN511_slv0_adr_3_),
	.a(slv0_adr[3]));
   in01f20 FE_OCPC510_slv0_adr_3_ (.o(FE_OCPN510_slv0_adr_3_),
	.a(slv0_adr[3]));
   in01s10 FE_OCPC170_n2346_dup (.o(FE_RN_15),
	.a(FE_OCPN166_n2346));
   in01s20 FE_OCPC169_n2346_dup (.o(FE_RN_14),
	.a(FE_OCPN165_n2346));
   in01m10 FE_OCPC383_n1512_dup (.o(FE_RN_13),
	.a(n1512));
   in01m10 FE_OCPC505_n2304 (.o(FE_OCPN505_n2304),
	.a(n2304));
   no02s10 U2953_dup2 (.o(FE_RN_12),
	.b(n1737),
	.a(n1738));
   no02s10 U2953_dup1 (.o(FE_RN_11),
	.b(n1737),
	.a(n1738));
   na02s08 U2952_dup (.o(FE_RN_5),
	.b(n1733),
	.a(n1734));
   in01s10 FE_OCPC481_n2343 (.o(FE_OCPN481_n2343),
	.a(n2343));
   in01m02 FE_OCPC480_n1573 (.o(FE_OCPN480_n1573),
	.a(n1573));
   in01m10 FE_OCPC479_n1573 (.o(FE_OCPN479_n1573),
	.a(n1573));
   in01s04 FE_OCPC478_n1573 (.o(FE_OCPN478_n1573),
	.a(n1573));
   na02f40 U2945_dup (.o(FE_RN_9),
	.b(FE_RN_8),
	.a(n2343));
   in01s06 FE_OCPC464_n1521 (.o(FE_OCPN464_n1521),
	.a(FE_OCPN176_n1521));
   in01m10 FE_OCPC463_n1521 (.o(FE_OCPN463_n1521),
	.a(FE_OCPN176_n1521));
   in01f20 FE_OCPC462_n1521 (.o(FE_OCPN462_n1521),
	.a(FE_OCPN176_n1521));
   no02s04 FE_RC_105_0 (.o(FE_RN_50_0),
	.b(n1595),
	.a(n1875));
   in01m02 FE_RC_104_0 (.o(FE_RN_51_0),
	.a(n1628));
   in01s02 FE_RC_103_0 (.o(n528),
	.a(FE_RN_52_0));
   no02s04 FE_RC_102_0 (.o(FE_RN_52_0),
	.b(FE_RN_51_0),
	.a(FE_RN_50_0));
   no02f20 U1922_dup (.o(FE_RN_8),
	.b(n1890),
	.a(n1546));
   na03f80 U2300_dup (.o(FE_RN_7),
	.c(FE_OCPN511_slv0_adr_3_),
	.b(FE_OCPN669_slv0_adr_4_),
	.a(FE_OCPN139_slv0_adr_2_));
   in01s01 FE_RC_101_0 (.o(FE_RN_47_0),
	.a(n1894));
   na02s04 FE_RC_99_0 (.o(FE_RN_49_0),
	.b(FE_OCPN540_n1595),
	.a(FE_RN_47_0));
   na02s02 FE_RC_98_0 (.o(n526),
	.b(FE_RN_49_0),
	.a(n1888));
   no03f08 FE_RC_97_0 (.o(n1947),
	.c(n1944),
	.b(n1945),
	.a(FE_OCPN673_n1577));
   oa22f06 FE_RC_96_0 (.o(n509),
	.d(FE_OCPN676_n1580),
	.c(n2191),
	.b(FE_OCPN538_n1595),
	.a(n2192));
   in01s02 FE_RC_95_0 (.o(FE_RN_44_0),
	.a(ch0_txsz[22]));
   no02m10 FE_RC_93_0 (.o(FE_RN_46_0),
	.b(FE_OCPN505_n2304),
	.a(FE_RN_44_0));
   no02m08 FE_RC_92_0 (.o(n2245),
	.b(FE_RN_46_0),
	.a(n2244));
   in01s40 FE_OCPC444_slv0_adr_8_ (.o(FE_OCPN444_slv0_adr_8_),
	.a(slv0_adr[8]));
   in01m06 FE_OCPC443_slv0_adr_8_ (.o(FE_OCPN443_slv0_adr_8_),
	.a(FE_OCPN444_slv0_adr_8_));
   in01s40 FE_OCPC442_slv0_adr_8_ (.o(FE_OCPN442_slv0_adr_8_),
	.a(FE_OCPN444_slv0_adr_8_));
   in01s02 FE_RC_91_0 (.o(FE_RN_41_0),
	.a(n1556));
   in01m03 FE_RC_90_0 (.o(FE_RN_42_0),
	.a(n1559));
   na02f04 FE_RC_89_0 (.o(FE_RN_43_0),
	.b(FE_RN_42_0),
	.a(FE_RN_41_0));
   no02m04 FE_RC_88_0 (.o(n1481),
	.b(n1554),
	.a(FE_RN_43_0));
   in01s04 FE_OFC427_wb0_ack_i (.o(FE_OFN427_wb0_ack_i),
	.a(FE_OFN426_wb0_ack_i));
   in01s02 FE_OFC426_wb0_ack_i (.o(FE_OFN426_wb0_ack_i),
	.a(wb0_ack_i));
   in01s01 FE_RC_86_0 (.o(FE_RN_38_0),
	.a(ch0_txsz[2]));
   in01m04 FE_RC_85_0 (.o(FE_RN_39_0),
	.a(n1924));
   no02m08 FE_RC_84_0 (.o(FE_RN_40_0),
	.b(FE_RN_39_0),
	.a(FE_RN_38_0));
   no02m08 FE_RC_83_0 (.o(n1906),
	.b(FE_RN_40_0),
	.a(n1905));
   ao22f08 FE_RC_82_0 (.o(n2239),
	.d(FE_OCPN124_FE_RN_),
	.c(u0_int_maska_22_),
	.b(FE_OCPN552_n1424),
	.a(u0_int_maskb_22_));
   oa22m04 FE_RC_81_0 (.o(n521),
	.d(FE_OCPN676_n1580),
	.c(n1985),
	.b(FE_OCPN539_n1595),
	.a(n1989));
   na03f06 FE_RC_80_0 (.o(n2456),
	.c(n2031),
	.b(n2029),
	.a(n2030));
   no02s02 FE_RC_79_0 (.o(FE_RN_35_0),
	.b(FE_OCPN657_wb1_cyc_o),
	.a(n1652));
   in01s01 FE_RC_78_0 (.o(FE_RN_36_0),
	.a(FE_OCPN661_wb1_cyc_o));
   in01s01 FE_RC_77_0 (.o(wb1_addr_o[8]),
	.a(FE_RN_37_0));
   no02s02 FE_RC_76_0 (.o(FE_RN_37_0),
	.b(FE_RN_36_0),
	.a(FE_RN_35_0));
   na02s02 FE_RC_75_0 (.o(FE_RN_34_0),
	.b(FE_OCPN651_wb1_cyc_o),
	.a(wb0_addr_i[25]));
   na02s02 FE_RC_74_0 (.o(wb1_addr_o[25]),
	.b(FE_RN_34_0),
	.a(wb1_cyc_o));
   no04s80 FE_RC_73_0 (.o(n1725),
	.d(wb1_addr_i[31]),
	.c(wb1_addr_i[29]),
	.b(wb1_addr_i[30]),
	.a(wb1_addr_i[28]));
   na03f06 FE_RC_70_0 (.o(n2459),
	.c(n1981),
	.b(n1982),
	.a(n1980));
   oa22s04 FE_RC_69_0 (.o(n551),
	.d(FE_OCPN383_n1512),
	.c(n2238),
	.b(n1591),
	.a(n2237));
   na03f80 FE_RC_68_0 (.o(FE_RN_),
	.c(FE_OCPN669_slv0_adr_4_),
	.b(FE_OCPN139_slv0_adr_2_),
	.a(FE_OCPN512_slv0_adr_3_));
   in01m02 FE_OCPC403_n2346 (.o(FE_OCPN403_n2346),
	.a(FE_OCPN402_n2346));
   in01m06 FE_OCPC402_n2346 (.o(FE_OCPN402_n2346),
	.a(n2346));
   oa22f08 FE_RC_66_0 (.o(n2325),
	.d(n2323),
	.c(FE_OCPN167_n2346),
	.b(FE_OCPN670_n2356),
	.a(n2324));
   in01s06 FE_OCPC385_n1579 (.o(FE_OCPN385_n1579),
	.a(FE_RN_18));
   in01s06 FE_OCPC384_n1579 (.o(FE_OCPN384_n1579),
	.a(FE_RN_18));
   in01s20 FE_OCPC383_n1512 (.o(FE_OCPN383_n1512),
	.a(n1512));
   in01s01 FE_RC_64_0 (.o(FE_RN_31_0),
	.a(n1488));
   na02s04 FE_RC_62_0 (.o(FE_RN_33_0),
	.b(FE_OCPN619_n1513),
	.a(FE_RN_31_0));
   na02s02 FE_RC_61_0 (.o(n643),
	.b(FE_RN_33_0),
	.a(n1889));
   no02f80 U2302_dup2 (.o(FE_RN_4),
	.b(slv0_adr[8]),
	.a(slv0_adr[9]));
   no03f08 FE_RC_60_0 (.o(FE_RN_27_0),
	.c(FE_RN_26_0),
	.b(FE_RN_23_0),
	.a(FE_OCPN672_n1577));
   na02m04 FE_RC_59_0 (.o(FE_RN_22_0),
	.b(n2165),
	.a(ch0_adr0[11]));
   no02f08 FE_RC_58_0 (.o(FE_RN_23_0),
	.b(FE_OCPN671_n2356),
	.a(n2063));
   no02f08 FE_RC_57_0 (.o(FE_RN_24_0),
	.b(n1424),
	.a(n2060));
   ao12f06 FE_RC_56_0 (.o(FE_RN_25_0),
	.c(n2343),
	.b(u0_int_maska_11_),
	.a(FE_RN_24_0));
   no02f06 FE_RC_55_0 (.o(FE_RN_26_0),
	.b(FE_RN_25_0),
	.a(FE_OCPN403_n2346));
   in01s01 FE_RC_53_0 (.o(FE_RN_28_0),
	.a(ch0_csr[11]));
   no02m08 FE_RC_52_0 (.o(FE_RN_29_0),
	.b(n2156),
	.a(FE_RN_28_0));
   ao12f06 FE_RC_51_0 (.o(FE_RN_30_0),
	.c(n2225),
	.b(ch0_txsz[11]),
	.a(FE_RN_29_0));
   na03f06 FE_RC_50_0 (.o(n2454),
	.c(FE_RN_30_0),
	.b(FE_RN_27_0),
	.a(FE_RN_22_0));
   in01f20 FE_OCPC370_n2194 (.o(FE_OCPN370_n2194),
	.a(FE_OCPN366_n2194));
   in01s10 FE_OCPC368_n2194 (.o(FE_OCPN368_n2194),
	.a(FE_OCPN365_n2194));
   in01m10 FE_OCPC367_n2194 (.o(FE_OCPN367_n2194),
	.a(FE_OCPN365_n2194));
   in01f10 FE_OCPC366_n2194 (.o(FE_OCPN366_n2194),
	.a(n2194));
   in01f10 FE_OCPC365_n2194 (.o(FE_OCPN365_n2194),
	.a(n2194));
   in01s06 FE_OCPC363_n2194 (.o(FE_OCPN363_n2194),
	.a(n2194));
   oa22f02 FE_RC_48_0 (.o(n593),
	.d(FE_OCPN180_n1521),
	.c(n2013),
	.b(FE_OCPN463_n1521),
	.a(n2005));
   in01s01 FE_RC_47_0 (.o(wb1s_data_o[3]),
	.a(FE_RN_21_0));
   ao22s02 FE_RC_46_0 (.o(FE_RN_21_0),
	.d(FE_OCPN643_wb1_cyc_o),
	.c(wb0m_data_i[3]),
	.b(FE_RN_1),
	.a(de_csr[3]));
   no02s20 U2953_dup (.o(FE_RN_1),
	.b(n1737),
	.a(FE_RN_5));
   na02s02 FE_RC_45_0 (.o(FE_RN_19_0),
	.b(FE_OCPN627_wb1_cyc_o),
	.a(slv0_din[25]));
   in01s01 FE_RC_44_0 (.o(FE_RN_20_0),
	.a(wb1s_data_i[25]));
   oa12s02 FE_RC_43_0 (.o(wb0m_data_o[25]),
	.c(FE_OCPN633_wb1_cyc_o),
	.b(FE_RN_20_0),
	.a(FE_RN_19_0));
   in01s10 FE_OCPC284_wb0_cyc_o (.o(FE_OCPN284_wb0_cyc_o),
	.a(FE_OCPN280_wb0_cyc_o));
   in01s10 FE_OCPC283_wb0_cyc_o (.o(wb0_cyc_o),
	.a(FE_OCPN280_wb0_cyc_o));
   in01f06 FE_OCPC280_wb0_cyc_o (.o(FE_OCPN280_wb0_cyc_o),
	.a(FE_RN_17));
   no04s80 FE_RC_38_0 (.o(n1629),
	.d(wb0_addr_i[29]),
	.c(wb0_addr_i[30]),
	.b(wb0_addr_i[28]),
	.a(wb0_addr_i[31]));
   in01s01 FE_RC_37_0 (.o(FE_RN_13_0),
	.a(n2001));
   na02s02 FE_RC_35_0 (.o(FE_RN_15_0),
	.b(FE_OCPN651_wb1_cyc_o),
	.a(FE_RN_13_0));
   na02s02 FE_RC_34_0 (.o(wb0m_data_o[7]),
	.b(n2000),
	.a(FE_RN_15_0));
   in01s04 FE_OCPC200_n2156 (.o(FE_OCPN200_n2156),
	.a(n2156));
   in01s10 FE_OCPC192_slv0_adr_9_ (.o(FE_OCPN192_slv0_adr_9_),
	.a(n1547));
   in01m06 FE_RC_32_0 (.o(FE_RN_11_0),
	.a(n1416));
   no02f06 FE_RC_31_0 (.o(FE_RN_12_0),
	.b(FE_RN_11_0),
	.a(n1916));
   no02f04 FE_RC_30_0 (.o(n1927),
	.b(FE_RN_12_0),
	.a(n1926));
   in01s01 FE_RC_29_0 (.o(FE_RN_7_0),
	.a(ch0_csr[3]));
   no02s06 FE_RC_27_0 (.o(FE_RN_9_0),
	.b(n2156),
	.a(FE_RN_7_0));
   no02f04 FE_RC_26_0 (.o(n1928),
	.b(FE_RN_9_0),
	.a(n1921));
   in01s20 FE_OCPC186_n1893 (.o(FE_OCPN186_n1893),
	.a(FE_RN_4));
   in01f08 FE_OCPC180_n1521 (.o(FE_OCPN180_n1521),
	.a(n1521));
   in01f08 FE_OCPC179_n1521 (.o(FE_OCPN179_n1521),
	.a(n1521));
   in01f10 FE_OCPC178_n1521 (.o(FE_OCPN178_n1521),
	.a(n1521));
   in01f40 FE_OCPC176_n1521 (.o(FE_OCPN176_n1521),
	.a(n1521));
   no02f20 U2302_dup (.o(FE_RN_2),
	.b(FE_OCPN443_slv0_adr_8_),
	.a(FE_OCPN192_slv0_adr_9_));
   in01s04 FE_OCPC171_n2346 (.o(FE_OCPN171_n2346),
	.a(FE_OCPN166_n2346));
   in01s10 FE_OCPC170_n2346 (.o(FE_OCPN170_n2346),
	.a(FE_OCPN166_n2346));
   in01s20 FE_OCPC169_n2346 (.o(FE_OCPN169_n2346),
	.a(FE_OCPN165_n2346));
   in01s06 FE_OCPC167_n2346 (.o(FE_OCPN167_n2346),
	.a(FE_OCPN402_n2346));
   in01m10 FE_OCPC166_n2346 (.o(FE_OCPN166_n2346),
	.a(n2346));
   in01m20 FE_OCPC165_n2346 (.o(FE_OCPN165_n2346),
	.a(n2346));
   in01s40 FE_OCPC163_n2346 (.o(FE_OCPN163_n2346),
	.a(n2346));
   na03f06 FE_RC_25_0 (.o(n2448),
	.c(n2167),
	.b(n2168),
	.a(n2166));
   in01f80 FE_OCPC139_slv0_adr_2_ (.o(FE_OCPN139_slv0_adr_2_),
	.a(FE_OCPN137_slv0_adr_2_));
   in01s10 FE_OCPC138_slv0_adr_2_ (.o(FE_OCPN138_slv0_adr_2_),
	.a(slv0_adr[2]));
   in01f80 FE_OCPC137_slv0_adr_2_ (.o(FE_OCPN137_slv0_adr_2_),
	.a(slv0_adr[2]));
   in01f10 FE_OCPC129_n2007 (.o(FE_OCPN129_n2007),
	.a(n2007));
   no04f40 FE_RC_24_0 (.o(n1530),
	.d(n1529),
	.c(FE_OCPN617_slv0_adr_5_),
	.b(FE_OCPN442_slv0_adr_8_),
	.a(slv0_adr[9]));
   in01f10 FE_OCPC126_FE_RN_ (.o(FE_OCPN126_FE_RN_),
	.a(FE_OCPN120_FE_RN_));
   in01f20 FE_OCPC124_FE_RN_ (.o(FE_OCPN124_FE_RN_),
	.a(FE_RN_));
   in01f10 FE_OCPC122_FE_RN_ (.o(FE_OCPN122_FE_RN_),
	.a(FE_RN_));
   in01f10 FE_OCPC120_FE_RN_ (.o(FE_OCPN120_FE_RN_),
	.a(FE_RN_));
   in01f20 FE_OCPC106_slv0_adr_2_ (.o(FE_OCPN106_slv0_adr_2_),
	.a(FE_OCPN139_slv0_adr_2_));
   na02f20 FE_RC_22_0 (.o(n1512),
	.b(FE_OCPN552_n1424),
	.a(n1522));
   na03f06 FE_RC_21_0 (.o(n2449),
	.c(n2149),
	.b(n2148),
	.a(n2147));
   in01f06 FE_OCPC80_n1919 (.o(FE_OCPN80_n1919),
	.a(n1919));
   in01s04 FE_OCPC79_n2056 (.o(FE_OCPN79_n2056),
	.a(FE_OCPN78_n2056));
   in01s03 FE_OCPC78_n2056 (.o(FE_OCPN78_n2056),
	.a(n2056));
   no02s08 FE_RC_17_0 (.o(FE_RN_5_0),
	.b(n2156),
	.a(n2369));
   no02f04 FE_RC_16_0 (.o(n1907),
	.b(n1899),
	.a(FE_RN_5_0));
   na03f06 FE_RC_15_0 (.o(n2455),
	.c(n2046),
	.b(n2045),
	.a(n2047));
   in01s01 FE_RC_13_0 (.o(FE_RN_0_0),
	.a(n1884));
   na02s04 FE_RC_11_0 (.o(FE_RN_2_0),
	.b(FE_OCPN200_n2156),
	.a(FE_RN_0_0));
   na02f02 FE_RC_10_0 (.o(n2464),
	.b(n1549),
	.a(FE_RN_2_0));
   oa22m04 FE_RC_9_0 (.o(n518),
	.d(FE_OCPN676_n1580),
	.c(n2034),
	.b(FE_OCPN540_n1595),
	.a(n2037));
   na03f06 FE_RC_7_0 (.o(n2460),
	.c(n1966),
	.b(n1964),
	.a(n1965));
   na03f06 FE_RC_4_0 (.o(n2185),
	.c(n2180),
	.b(n2181),
	.a(n2241));
   na03f06 FE_RC_3_0 (.o(n2450),
	.c(n2130),
	.b(n2131),
	.a(n2129));
   na04f40 FE_RC_2_0 (.o(n1546),
	.d(n1547),
	.c(n1548),
	.b(slv0_adr[5]),
	.a(slv0_we));
   oa22f08 FE_RC_0_0 (.o(n2128),
	.d(n2126),
	.c(FE_RN_15),
	.b(FE_OCPN671_n2356),
	.a(n2127));
   ms00f80 u1_ndnr_reg_0_ (.o(ndnr_0_),
	.d(u1_N1032),
	.ck(clk));
   ms00f80 u3_u1_slv_dout_reg_0_ (.o(slv0_dout[0]),
	.d(wb0m_data_i[0]),
	.ck(clk));
   ms00f80 u3_u1_slv_dout_reg_1_ (.o(slv0_dout[1]),
	.d(wb0m_data_i[1]),
	.ck(clk));
   ms00f80 u3_u1_slv_dout_reg_2_ (.o(slv0_dout[2]),
	.d(wb0m_data_i[2]),
	.ck(clk));
   ms00f80 u3_u1_slv_dout_reg_3_ (.o(slv0_dout[3]),
	.d(wb0m_data_i[3]),
	.ck(clk));
   ms00f80 u3_u1_slv_dout_reg_4_ (.o(slv0_dout[4]),
	.d(wb0m_data_i[4]),
	.ck(clk));
   ms00f80 u3_u1_slv_dout_reg_5_ (.o(slv0_dout[5]),
	.d(wb0m_data_i[5]),
	.ck(clk));
   ms00f80 u3_u1_slv_dout_reg_6_ (.o(slv0_dout[6]),
	.d(wb0m_data_i[6]),
	.ck(clk));
   ms00f80 u3_u1_slv_dout_reg_7_ (.o(slv0_dout[7]),
	.d(wb0m_data_i[7]),
	.ck(clk));
   ms00f80 u3_u1_slv_dout_reg_8_ (.o(slv0_dout[8]),
	.d(wb0m_data_i[8]),
	.ck(clk));
   ms00f80 u3_u1_slv_dout_reg_9_ (.o(slv0_dout[9]),
	.d(wb0m_data_i[9]),
	.ck(clk));
   ms00f80 u3_u1_slv_dout_reg_10_ (.o(slv0_dout[10]),
	.d(wb0m_data_i[10]),
	.ck(clk));
   ms00f80 u3_u1_slv_dout_reg_11_ (.o(slv0_dout[11]),
	.d(wb0m_data_i[11]),
	.ck(clk));
   ms00f80 u3_u1_slv_dout_reg_12_ (.o(slv0_dout[12]),
	.d(wb0m_data_i[12]),
	.ck(clk));
   ms00f80 u3_u1_slv_dout_reg_13_ (.o(slv0_dout[13]),
	.d(wb0m_data_i[13]),
	.ck(clk));
   ms00f80 u3_u1_slv_dout_reg_14_ (.o(slv0_dout[14]),
	.d(wb0m_data_i[14]),
	.ck(clk));
   ms00f80 u3_u1_slv_dout_reg_15_ (.o(slv0_dout[15]),
	.d(wb0m_data_i[15]),
	.ck(clk));
   ms00f80 u3_u1_slv_dout_reg_16_ (.o(slv0_dout[16]),
	.d(wb0m_data_i[16]),
	.ck(clk));
   ms00f80 u3_u1_slv_dout_reg_17_ (.o(slv0_dout[17]),
	.d(wb0m_data_i[17]),
	.ck(clk));
   ms00f80 u3_u1_slv_dout_reg_18_ (.o(slv0_dout[18]),
	.d(wb0m_data_i[18]),
	.ck(clk));
   ms00f80 u3_u1_slv_dout_reg_19_ (.o(slv0_dout[19]),
	.d(wb0m_data_i[19]),
	.ck(clk));
   ms00f80 u3_u1_slv_dout_reg_20_ (.o(slv0_dout[20]),
	.d(wb0m_data_i[20]),
	.ck(clk));
   ms00f80 u3_u1_slv_dout_reg_21_ (.o(slv0_dout[21]),
	.d(wb0m_data_i[21]),
	.ck(clk));
   ms00f80 u3_u1_slv_dout_reg_22_ (.o(slv0_dout[22]),
	.d(wb0m_data_i[22]),
	.ck(clk));
   ms00f80 u3_u1_slv_dout_reg_23_ (.o(slv0_dout[23]),
	.d(wb0m_data_i[23]),
	.ck(clk));
   ms00f80 u3_u1_slv_dout_reg_24_ (.o(slv0_dout[24]),
	.d(wb0m_data_i[24]),
	.ck(clk));
   ms00f80 u3_u1_slv_dout_reg_25_ (.o(slv0_dout[25]),
	.d(wb0m_data_i[25]),
	.ck(clk));
   ms00f80 u3_u1_slv_dout_reg_26_ (.o(slv0_dout[26]),
	.d(wb0m_data_i[26]),
	.ck(clk));
   ms00f80 u3_u1_slv_dout_reg_27_ (.o(slv0_dout[27]),
	.d(wb0m_data_i[27]),
	.ck(clk));
   ms00f80 u3_u1_slv_dout_reg_28_ (.o(slv0_dout[28]),
	.d(wb0m_data_i[28]),
	.ck(clk));
   ms00f80 u3_u1_slv_dout_reg_29_ (.o(slv0_dout[29]),
	.d(wb0m_data_i[29]),
	.ck(clk));
   ms00f80 u3_u1_slv_dout_reg_30_ (.o(slv0_dout[30]),
	.d(wb0m_data_i[30]),
	.ck(clk));
   ms00f80 u3_u1_slv_dout_reg_31_ (.o(slv0_dout[31]),
	.d(wb0m_data_i[31]),
	.ck(clk));
   ms00f80 u3_u1_slv_re_reg (.o(slv0_re),
	.d(u3_u1_N3),
	.ck(clk));
   ms00f80 u3_u1_rf_ack_reg (.o(u3_u1_rf_ack),
	.d(u3_u1_N5),
	.ck(clk));
   ms00f80 u3_u1_slv_we_reg (.o(slv0_we),
	.d(u3_u1_N4),
	.ck(clk));
   ms00f80 u3_u1_slv_adr_reg_2_ (.o(slv0_adr[2]),
	.d(wb0_addr_i[2]),
	.ck(clk));
   ms00f80 u3_u1_slv_adr_reg_3_ (.o(slv0_adr[3]),
	.d(wb0_addr_i[3]),
	.ck(clk));
   ms00f80 u3_u1_slv_adr_reg_4_ (.o(slv0_adr[4]),
	.d(wb0_addr_i[4]),
	.ck(clk));
   ms00f80 u3_u1_slv_adr_reg_5_ (.o(slv0_adr[5]),
	.d(wb0_addr_i[5]),
	.ck(clk));
   ms00f80 u3_u1_slv_adr_reg_6_ (.o(slv0_adr[6]),
	.d(wb0_addr_i[6]),
	.ck(clk));
   ms00f80 u3_u1_slv_adr_reg_7_ (.o(slv0_adr[7]),
	.d(wb0_addr_i[7]),
	.ck(clk));
   ms00f80 u3_u1_slv_adr_reg_8_ (.o(slv0_adr[8]),
	.d(wb0_addr_i[8]),
	.ck(clk));
   ms00f80 u3_u1_slv_adr_reg_9_ (.o(slv0_adr[9]),
	.d(wb0_addr_i[9]),
	.ck(clk));
   ms00f80 u0_wb_rf_dout_reg_31_ (.o(slv0_din[31]),
	.d(u0_N3074),
	.ck(clk));
   ms00f80 u0_intb_o_reg (.o(intb_o),
	.d(n2466),
	.ck(clk));
   ms00f80 u0_inta_o_reg (.o(inta_o),
	.d(n2465),
	.ck(clk));
   ms00f80 u0_wb_rf_dout_reg_1_ (.o(slv0_din[1]),
	.d(n2464),
	.ck(clk));
   ms00f80 u0_wb_rf_dout_reg_2_ (.o(slv0_din[2]),
	.d(n2463),
	.ck(clk));
   ms00f80 u0_wb_rf_dout_reg_3_ (.o(slv0_din[3]),
	.d(n2462),
	.ck(clk));
   ms00f80 u0_wb_rf_dout_reg_4_ (.o(slv0_din[4]),
	.d(n2461),
	.ck(clk));
   ms00f80 u0_wb_rf_dout_reg_5_ (.o(slv0_din[5]),
	.d(n2460),
	.ck(clk));
   ms00f80 u0_wb_rf_dout_reg_6_ (.o(slv0_din[6]),
	.d(n2459),
	.ck(clk));
   ms00f80 u0_wb_rf_dout_reg_7_ (.o(slv0_din[7]),
	.d(n2458),
	.ck(clk));
   ms00f80 u0_wb_rf_dout_reg_8_ (.o(slv0_din[8]),
	.d(n2457),
	.ck(clk));
   ms00f80 u0_wb_rf_dout_reg_9_ (.o(slv0_din[9]),
	.d(n2456),
	.ck(clk));
   ms00f80 u0_wb_rf_dout_reg_10_ (.o(slv0_din[10]),
	.d(n2455),
	.ck(clk));
   ms00f80 u0_wb_rf_dout_reg_11_ (.o(slv0_din[11]),
	.d(n2454),
	.ck(clk));
   ms00f80 u0_wb_rf_dout_reg_12_ (.o(slv0_din[12]),
	.d(n2453),
	.ck(clk));
   ms00f80 u0_wb_rf_dout_reg_13_ (.o(slv0_din[13]),
	.d(n2452),
	.ck(clk));
   ms00f80 u0_wb_rf_dout_reg_14_ (.o(slv0_din[14]),
	.d(n2451),
	.ck(clk));
   ms00f80 u0_wb_rf_dout_reg_15_ (.o(slv0_din[15]),
	.d(n2450),
	.ck(clk));
   ms00f80 u0_wb_rf_dout_reg_16_ (.o(slv0_din[16]),
	.d(n2449),
	.ck(clk));
   ms00f80 u0_wb_rf_dout_reg_17_ (.o(slv0_din[17]),
	.d(n2448),
	.ck(clk));
   ms00f80 u0_wb_rf_dout_reg_18_ (.o(slv0_din[18]),
	.d(FE_OCPN674_n2186),
	.ck(clk));
   ms00f80 u0_wb_rf_dout_reg_19_ (.o(slv0_din[19]),
	.d(n2446),
	.ck(clk));
   ms00f80 u0_wb_rf_dout_reg_20_ (.o(slv0_din[20]),
	.d(n2445),
	.ck(clk));
   ms00f80 u0_wb_rf_dout_reg_21_ (.o(slv0_din[21]),
	.d(n2444),
	.ck(clk));
   ms00f80 u0_wb_rf_dout_reg_22_ (.o(slv0_din[22]),
	.d(n2443),
	.ck(clk));
   ms00f80 u0_wb_rf_dout_reg_23_ (.o(slv0_din[23]),
	.d(n2442),
	.ck(clk));
   ms00f80 u0_wb_rf_dout_reg_24_ (.o(slv0_din[24]),
	.d(n2441),
	.ck(clk));
   ms00f80 u0_wb_rf_dout_reg_25_ (.o(slv0_din[25]),
	.d(n2440),
	.ck(clk));
   ms00f80 u0_wb_rf_dout_reg_26_ (.o(slv0_din[26]),
	.d(n2439),
	.ck(clk));
   ms00f80 u0_wb_rf_dout_reg_27_ (.o(slv0_din[27]),
	.d(n2438),
	.ck(clk));
   ms00f80 u0_wb_rf_dout_reg_28_ (.o(slv0_din[28]),
	.d(n2437),
	.ck(clk));
   ms00f80 u0_wb_rf_dout_reg_29_ (.o(slv0_din[29]),
	.d(n2436),
	.ck(clk));
   ms00f80 u0_wb_rf_dout_reg_30_ (.o(slv0_din[30]),
	.d(n2435),
	.ck(clk));
   ms00f80 u0_wb_rf_dout_reg_0_ (.o(slv0_din[0]),
	.d(n2434),
	.ck(clk));
   ms00f80 u4_u1_slv_re_reg (.o(slv1_re),
	.d(u4_u1_N3),
	.ck(clk));
   ms00f80 u4_u1_rf_ack_reg (.o(u4_u1_rf_ack),
	.d(n893),
	.ck(clk));
   ms00f80 u4_u1_slv_we_reg (.o(slv1_we),
	.d(u4_u1_N4),
	.ck(clk));
   ms00f80 u3_u0_mast_dout_reg_0_ (.o(de_csr[0]),
	.d(n831),
	.ck(clk));
   ms00f80 u3_u0_mast_dout_reg_1_ (.o(de_csr[1]),
	.d(n830),
	.ck(clk));
   ms00f80 u3_u0_mast_dout_reg_2_ (.o(de_csr[2]),
	.d(n829),
	.ck(clk));
   ms00f80 u3_u0_mast_dout_reg_3_ (.o(de_csr[3]),
	.d(n828),
	.ck(clk));
   ms00f80 u3_u0_mast_dout_reg_4_ (.o(de_csr[4]),
	.d(n827),
	.ck(clk));
   ms00f80 u3_u0_mast_dout_reg_5_ (.o(de_csr[5]),
	.d(n826),
	.ck(clk));
   ms00f80 u3_u0_mast_dout_reg_6_ (.o(de_csr[6]),
	.d(n825),
	.ck(clk));
   ms00f80 u3_u0_mast_dout_reg_7_ (.o(de_csr[7]),
	.d(n824),
	.ck(clk));
   ms00f80 u3_u0_mast_dout_reg_8_ (.o(de_csr[8]),
	.d(n823),
	.ck(clk));
   ms00f80 u3_u0_mast_dout_reg_9_ (.o(de_csr[9]),
	.d(n822),
	.ck(clk));
   ms00f80 u3_u0_mast_dout_reg_10_ (.o(de_csr[10]),
	.d(n821),
	.ck(clk));
   ms00f80 u3_u0_mast_dout_reg_11_ (.o(de_csr[11]),
	.d(n820),
	.ck(clk));
   ms00f80 u3_u0_mast_dout_reg_12_ (.o(de_csr[12]),
	.d(n819),
	.ck(clk));
   ms00f80 u3_u0_mast_dout_reg_13_ (.o(de_csr[13]),
	.d(n818),
	.ck(clk));
   ms00f80 u3_u0_mast_dout_reg_14_ (.o(de_csr[14]),
	.d(n817),
	.ck(clk));
   ms00f80 u3_u0_mast_dout_reg_15_ (.o(de_csr[15]),
	.d(n816),
	.ck(clk));
   ms00f80 u3_u0_mast_dout_reg_16_ (.o(de_csr[16]),
	.d(n815),
	.ck(clk));
   ms00f80 u3_u0_mast_dout_reg_17_ (.o(de_csr[17]),
	.d(n814),
	.ck(clk));
   ms00f80 u3_u0_mast_dout_reg_18_ (.o(de_csr[18]),
	.d(n813),
	.ck(clk));
   ms00f80 u3_u0_mast_dout_reg_19_ (.o(de_csr[19]),
	.d(n812),
	.ck(clk));
   ms00f80 u3_u0_mast_dout_reg_20_ (.o(de_csr[20]),
	.d(n811),
	.ck(clk));
   ms00f80 u3_u0_mast_dout_reg_21_ (.o(de_csr[21]),
	.d(n810),
	.ck(clk));
   ms00f80 u3_u0_mast_dout_reg_22_ (.o(de_csr[22]),
	.d(n809),
	.ck(clk));
   ms00f80 u3_u0_mast_dout_reg_23_ (.o(de_csr[23]),
	.d(n808),
	.ck(clk));
   ms00f80 u3_u0_mast_dout_reg_24_ (.o(de_csr[24]),
	.d(n807),
	.ck(clk));
   ms00f80 u3_u0_mast_dout_reg_25_ (.o(de_csr[25]),
	.d(n806),
	.ck(clk));
   ms00f80 u3_u0_mast_dout_reg_26_ (.o(de_csr[26]),
	.d(n805),
	.ck(clk));
   ms00f80 u3_u0_mast_dout_reg_27_ (.o(de_csr[27]),
	.d(n804),
	.ck(clk));
   ms00f80 u3_u0_mast_dout_reg_28_ (.o(de_csr[28]),
	.d(n803),
	.ck(clk));
   ms00f80 u3_u0_mast_dout_reg_29_ (.o(de_csr[29]),
	.d(n802),
	.ck(clk));
   ms00f80 u3_u0_mast_dout_reg_30_ (.o(de_csr[30]),
	.d(n801),
	.ck(clk));
   ms00f80 u3_u0_mast_dout_reg_31_ (.o(de_csr[31]),
	.d(n800),
	.ck(clk));
   ms00f80 u0_u0_ch_csr_r3_reg_2_ (.o(ch0_csr[19]),
	.d(n767),
	.ck(clk));
   ms00f80 u0_u0_ch_csr_r3_reg_1_ (.o(ch0_csr[18]),
	.d(n766),
	.ck(clk));
   ms00f80 u0_u0_ch_csr_r3_reg_0_ (.o(ch0_csr[17]),
	.d(n765),
	.ck(clk));
   ms00f80 u0_u0_rest_en_reg (.o(ch0_csr[16]),
	.d(n764),
	.ck(clk));
   ms00f80 u0_u0_ch_csr_r2_reg_2_ (.o(ch0_csr[15]),
	.d(n763),
	.ck(clk));
   ms00f80 u0_u0_ch_csr_r2_reg_1_ (.o(ch0_csr[14]),
	.d(n762),
	.ck(clk));
   ms00f80 u0_u0_ch_csr_r2_reg_0_ (.o(ch0_csr[13]),
	.d(n761),
	.ck(clk));
   ms00f80 u0_u0_ch_csr_r_reg_8_ (.o(ch0_csr[8]),
	.d(n760),
	.ck(clk));
   ms00f80 u0_u0_ch_csr_r_reg_7_ (.o(ch0_csr[7]),
	.d(n759),
	.ck(clk));
   ms00f80 u0_u0_ch_csr_r_reg_6_ (.o(ch0_csr[6]),
	.d(n758),
	.ck(clk));
   ms00f80 u0_u0_ch_csr_r_reg_5_ (.o(ch0_csr[5]),
	.d(n757),
	.ck(clk));
   ms00f80 u0_u0_ch_chk_sz_r_reg_0_ (.o(ch0_txsz[16]),
	.d(n756),
	.ck(clk));
   ms00f80 u0_u0_ch_chk_sz_r_reg_1_ (.o(ch0_txsz[17]),
	.d(n755),
	.ck(clk));
   ms00f80 u0_u0_ch_chk_sz_r_reg_2_ (.o(ch0_txsz[18]),
	.d(n754),
	.ck(clk));
   ms00f80 u0_u0_ch_chk_sz_r_reg_3_ (.o(ch0_txsz[19]),
	.d(n753),
	.ck(clk));
   ms00f80 u0_u0_ch_chk_sz_r_reg_4_ (.o(ch0_txsz[20]),
	.d(n752),
	.ck(clk));
   ms00f80 u0_u0_ch_chk_sz_r_reg_5_ (.o(ch0_txsz[21]),
	.d(n751),
	.ck(clk));
   ms00f80 u0_u0_ch_chk_sz_r_reg_6_ (.o(ch0_txsz[22]),
	.d(n750),
	.ck(clk));
   ms00f80 u0_u0_ch_chk_sz_r_reg_7_ (.o(ch0_txsz[23]),
	.d(n749),
	.ck(clk));
   ms00f80 u0_u0_ch_chk_sz_r_reg_8_ (.o(ch0_txsz[24]),
	.d(n748),
	.ck(clk));
   ms00f80 u0_u0_ch_chk_sz_r_reg_9_ (.o(ch0_txsz[25]),
	.d(n747),
	.ck(clk));
   ms00f80 u0_u0_ch_chk_sz_r_reg_10_ (.o(ch0_txsz[26]),
	.d(n746),
	.ck(clk));
   ms00f80 u0_u0_ch_sz_inf_reg (.o(ch0_txsz[15]),
	.d(n745),
	.ck(clk));
   ms00f80 u0_u0_ch_tot_sz_r_reg_0_ (.o(ch0_txsz[0]),
	.d(n742),
	.ck(clk));
   ms00f80 u0_u0_ch_csr_r_reg_1_ (.o(ch0_csr[1]),
	.d(n734),
	.ck(clk));
   ms00f80 u0_u0_ch_csr_r_reg_2_ (.o(ch0_csr[2]),
	.d(n733),
	.ck(clk));
   ms00f80 u0_u0_ch_csr_r_reg_3_ (.o(ch0_csr[3]),
	.d(n732),
	.ck(clk));
   ms00f80 u0_u0_ch_csr_r_reg_4_ (.o(ch0_csr[4]),
	.d(n731),
	.ck(clk));
   ms00f80 u0_u0_ch_adr0_r_reg_29_ (.o(ch0_adr0[31]),
	.d(n721),
	.ck(clk));
   ms00f80 u0_u0_ch_adr0_r_reg_28_ (.o(ch0_adr0[30]),
	.d(n719),
	.ck(clk));
   ms00f80 u0_u0_ch_adr0_r_reg_27_ (.o(ch0_adr0[29]),
	.d(n717),
	.ck(clk));
   ms00f80 u0_u0_ch_adr0_r_reg_26_ (.o(ch0_adr0[28]),
	.d(n715),
	.ck(clk));
   ms00f80 u0_u0_ch_adr0_r_reg_25_ (.o(ch0_adr0[27]),
	.d(n713),
	.ck(clk));
   ms00f80 u0_u0_ch_adr0_r_reg_24_ (.o(ch0_adr0[26]),
	.d(n711),
	.ck(clk));
   ms00f80 u0_u0_ch_adr0_r_reg_23_ (.o(ch0_adr0[25]),
	.d(n709),
	.ck(clk));
   ms00f80 u0_u0_ch_adr0_r_reg_22_ (.o(ch0_adr0[24]),
	.d(n707),
	.ck(clk));
   ms00f80 u0_u0_ch_adr0_r_reg_21_ (.o(ch0_adr0[23]),
	.d(n705),
	.ck(clk));
   ms00f80 u0_u0_ch_adr0_r_reg_20_ (.o(ch0_adr0[22]),
	.d(n703),
	.ck(clk));
   ms00f80 u0_u0_ch_adr0_r_reg_19_ (.o(ch0_adr0[21]),
	.d(n701),
	.ck(clk));
   ms00f80 u0_u0_ch_adr0_r_reg_18_ (.o(ch0_adr0[20]),
	.d(n699),
	.ck(clk));
   ms00f80 u0_u0_ch_adr0_r_reg_17_ (.o(ch0_adr0[19]),
	.d(n697),
	.ck(clk));
   ms00f80 u0_u0_ch_adr0_r_reg_16_ (.o(ch0_adr0[18]),
	.d(n695),
	.ck(clk));
   ms00f80 u0_u0_ch_adr0_r_reg_15_ (.o(ch0_adr0[17]),
	.d(n693),
	.ck(clk));
   ms00f80 u0_u0_ch_adr0_r_reg_14_ (.o(ch0_adr0[16]),
	.d(n691),
	.ck(clk));
   ms00f80 u0_u0_ch_adr0_r_reg_13_ (.o(ch0_adr0[15]),
	.d(n689),
	.ck(clk));
   ms00f80 u0_u0_ch_adr0_r_reg_12_ (.o(ch0_adr0[14]),
	.d(n687),
	.ck(clk));
   ms00f80 u0_u0_ch_adr0_r_reg_11_ (.o(ch0_adr0[13]),
	.d(n685),
	.ck(clk));
   ms00f80 u0_u0_ch_adr0_r_reg_10_ (.o(ch0_adr0[12]),
	.d(n683),
	.ck(clk));
   ms00f80 u0_u0_ch_adr0_r_reg_9_ (.o(ch0_adr0[11]),
	.d(n681),
	.ck(clk));
   ms00f80 u0_u0_ch_adr0_r_reg_8_ (.o(ch0_adr0[10]),
	.d(n679),
	.ck(clk));
   ms00f80 u0_u0_ch_adr0_r_reg_7_ (.o(ch0_adr0[9]),
	.d(n677),
	.ck(clk));
   ms00f80 u0_u0_ch_adr0_r_reg_6_ (.o(ch0_adr0[8]),
	.d(n675),
	.ck(clk));
   ms00f80 u0_u0_ch_adr0_r_reg_5_ (.o(ch0_adr0[7]),
	.d(n673),
	.ck(clk));
   ms00f80 u0_u0_ch_adr0_r_reg_4_ (.o(ch0_adr0[6]),
	.d(n671),
	.ck(clk));
   ms00f80 u0_u0_ch_adr0_r_reg_3_ (.o(ch0_adr0[5]),
	.d(n669),
	.ck(clk));
   ms00f80 u0_u0_ch_adr0_r_reg_2_ (.o(ch0_adr0[4]),
	.d(n667),
	.ck(clk));
   ms00f80 u0_u0_ch_adr0_r_reg_1_ (.o(ch0_adr0[3]),
	.d(n665),
	.ck(clk));
   ms00f80 u0_u0_ch_adr0_r_reg_0_ (.o(ch0_adr0[2]),
	.d(n663),
	.ck(clk));
   ms00f80 u0_u0_ch_tot_sz_r_reg_11_ (.o(ch0_txsz[11]),
	.d(n661),
	.ck(clk));
   ms00f80 u0_u0_ch_tot_sz_r_reg_10_ (.o(ch0_txsz[10]),
	.d(n659),
	.ck(clk));
   ms00f80 u0_u0_ch_tot_sz_r_reg_9_ (.o(ch0_txsz[9]),
	.d(n657),
	.ck(clk));
   ms00f80 u0_u0_ch_tot_sz_r_reg_8_ (.o(ch0_txsz[8]),
	.d(n655),
	.ck(clk));
   ms00f80 u0_u0_ch_tot_sz_r_reg_7_ (.o(ch0_txsz[7]),
	.d(n653),
	.ck(clk));
   ms00f80 u0_u0_ch_tot_sz_r_reg_6_ (.o(ch0_txsz[6]),
	.d(n651),
	.ck(clk));
   ms00f80 u0_u0_ch_tot_sz_r_reg_5_ (.o(ch0_txsz[5]),
	.d(n649),
	.ck(clk));
   ms00f80 u0_u0_ch_tot_sz_r_reg_4_ (.o(ch0_txsz[4]),
	.d(n647),
	.ck(clk));
   ms00f80 u0_u0_ch_tot_sz_r_reg_3_ (.o(ch0_txsz[3]),
	.d(n645),
	.ck(clk));
   ms00f80 u0_u0_ch_tot_sz_r_reg_2_ (.o(ch0_txsz[2]),
	.d(n643),
	.ck(clk));
   ms00f80 u0_u0_ch_tot_sz_r_reg_1_ (.o(ch0_txsz[1]),
	.d(n641),
	.ck(clk));
   ms00f80 u0_u0_ch_adr1_r_reg_29_ (.o(ch0_adr1[31]),
	.d(n639),
	.ck(clk));
   ms00f80 u0_u0_ch_adr1_r_reg_28_ (.o(ch0_adr1[30]),
	.d(n637),
	.ck(clk));
   ms00f80 u0_u0_ch_adr1_r_reg_27_ (.o(ch0_adr1[29]),
	.d(n635),
	.ck(clk));
   ms00f80 u0_u0_ch_adr1_r_reg_26_ (.o(ch0_adr1[28]),
	.d(n633),
	.ck(clk));
   ms00f80 u0_u0_ch_adr1_r_reg_25_ (.o(ch0_adr1[27]),
	.d(n631),
	.ck(clk));
   ms00f80 u0_u0_ch_adr1_r_reg_24_ (.o(ch0_adr1[26]),
	.d(n629),
	.ck(clk));
   ms00f80 u0_u0_ch_adr1_r_reg_23_ (.o(ch0_adr1[25]),
	.d(n627),
	.ck(clk));
   ms00f80 u0_u0_ch_adr1_r_reg_22_ (.o(ch0_adr1[24]),
	.d(n625),
	.ck(clk));
   ms00f80 u0_u0_ch_adr1_r_reg_21_ (.o(ch0_adr1[23]),
	.d(n623),
	.ck(clk));
   ms00f80 u0_u0_ch_adr1_r_reg_20_ (.o(ch0_adr1[22]),
	.d(n621),
	.ck(clk));
   ms00f80 u0_u0_ch_adr1_r_reg_19_ (.o(ch0_adr1[21]),
	.d(n619),
	.ck(clk));
   ms00f80 u0_u0_ch_adr1_r_reg_18_ (.o(ch0_adr1[20]),
	.d(n617),
	.ck(clk));
   ms00f80 u0_u0_ch_adr1_r_reg_17_ (.o(ch0_adr1[19]),
	.d(n615),
	.ck(clk));
   ms00f80 u0_u0_ch_adr1_r_reg_16_ (.o(ch0_adr1[18]),
	.d(n613),
	.ck(clk));
   ms00f80 u0_u0_ch_adr1_r_reg_15_ (.o(ch0_adr1[17]),
	.d(n611),
	.ck(clk));
   ms00f80 u0_u0_ch_adr1_r_reg_14_ (.o(ch0_adr1[16]),
	.d(n609),
	.ck(clk));
   ms00f80 u0_u0_ch_adr1_r_reg_13_ (.o(ch0_adr1[15]),
	.d(n607),
	.ck(clk));
   ms00f80 u0_u0_ch_adr1_r_reg_12_ (.o(ch0_adr1[14]),
	.d(n605),
	.ck(clk));
   ms00f80 u0_u0_ch_adr1_r_reg_11_ (.o(ch0_adr1[13]),
	.d(n603),
	.ck(clk));
   ms00f80 u0_u0_ch_adr1_r_reg_10_ (.o(ch0_adr1[12]),
	.d(n601),
	.ck(clk));
   ms00f80 u0_u0_ch_adr1_r_reg_9_ (.o(ch0_adr1[11]),
	.d(n599),
	.ck(clk));
   ms00f80 u0_u0_ch_adr1_r_reg_8_ (.o(ch0_adr1[10]),
	.d(n597),
	.ck(clk));
   ms00f80 u0_u0_ch_adr1_r_reg_7_ (.o(ch0_adr1[9]),
	.d(n595),
	.ck(clk));
   ms00f80 u0_u0_ch_adr1_r_reg_6_ (.o(ch0_adr1[8]),
	.d(n593),
	.ck(clk));
   ms00f80 u0_u0_ch_adr1_r_reg_5_ (.o(ch0_adr1[7]),
	.d(n591),
	.ck(clk));
   ms00f80 u0_u0_ch_adr1_r_reg_4_ (.o(ch0_adr1[6]),
	.d(n589),
	.ck(clk));
   ms00f80 u0_u0_ch_adr1_r_reg_3_ (.o(ch0_adr1[5]),
	.d(n587),
	.ck(clk));
   ms00f80 u0_u0_ch_adr1_r_reg_2_ (.o(ch0_adr1[4]),
	.d(n585),
	.ck(clk));
   ms00f80 u0_u0_ch_adr1_r_reg_1_ (.o(ch0_adr1[3]),
	.d(n583),
	.ck(clk));
   ms00f80 u0_u0_ch_adr1_r_reg_0_ (.o(ch0_adr1[2]),
	.d(n581),
	.ck(clk));
   ms00f80 u0_u0_ch_done_reg (.o(ch0_csr[11]),
	.d(n571),
	.ck(clk));
   ms00f80 u0_u0_ch_csr_r_reg_0_ (.o(ch0_csr[0]),
	.d(n570),
	.ck(clk));
   ms00f80 u0_u0_int_src_r_reg_1_ (.o(ch0_csr[21]),
	.d(n560),
	.ck(clk));
   ms00f80 u0_int_maskb_r_reg_30_ (.o(u0_int_maskb_30_),
	.d(n559),
	.ck(clk));
   ms00f80 u0_int_maskb_r_reg_29_ (.o(u0_int_maskb_29_),
	.d(n558),
	.ck(clk));
   ms00f80 u0_int_maskb_r_reg_28_ (.o(u0_int_maskb_28_),
	.d(n557),
	.ck(clk));
   ms00f80 u0_int_maskb_r_reg_27_ (.o(u0_int_maskb_27_),
	.d(n556),
	.ck(clk));
   ms00f80 u0_int_maskb_r_reg_26_ (.o(u0_int_maskb_26_),
	.d(n555),
	.ck(clk));
   ms00f80 u0_int_maskb_r_reg_25_ (.o(u0_int_maskb_25_),
	.d(n554),
	.ck(clk));
   ms00f80 u0_int_maskb_r_reg_24_ (.o(u0_int_maskb_24_),
	.d(n553),
	.ck(clk));
   ms00f80 u0_int_maskb_r_reg_23_ (.o(u0_int_maskb_23_),
	.d(n552),
	.ck(clk));
   ms00f80 u0_int_maskb_r_reg_22_ (.o(u0_int_maskb_22_),
	.d(n551),
	.ck(clk));
   ms00f80 u0_int_maskb_r_reg_21_ (.o(u0_int_maskb_21_),
	.d(n550),
	.ck(clk));
   ms00f80 u0_int_maskb_r_reg_20_ (.o(u0_int_maskb_20_),
	.d(n549),
	.ck(clk));
   ms00f80 u0_int_maskb_r_reg_19_ (.o(u0_int_maskb_19_),
	.d(n548),
	.ck(clk));
   ms00f80 u0_int_maskb_r_reg_18_ (.o(u0_int_maskb_18_),
	.d(n547),
	.ck(clk));
   ms00f80 u0_int_maskb_r_reg_17_ (.o(u0_int_maskb_17_),
	.d(n546),
	.ck(clk));
   ms00f80 u0_int_maskb_r_reg_16_ (.o(u0_int_maskb_16_),
	.d(n545),
	.ck(clk));
   ms00f80 u0_int_maskb_r_reg_15_ (.o(u0_int_maskb_15_),
	.d(n544),
	.ck(clk));
   ms00f80 u0_int_maskb_r_reg_14_ (.o(u0_int_maskb_14_),
	.d(n543),
	.ck(clk));
   ms00f80 u0_int_maskb_r_reg_13_ (.o(u0_int_maskb_13_),
	.d(n542),
	.ck(clk));
   ms00f80 u0_int_maskb_r_reg_12_ (.o(u0_int_maskb_12_),
	.d(n541),
	.ck(clk));
   ms00f80 u0_int_maskb_r_reg_11_ (.o(u0_int_maskb_11_),
	.d(n540),
	.ck(clk));
   ms00f80 u0_int_maskb_r_reg_10_ (.o(u0_int_maskb_10_),
	.d(n539),
	.ck(clk));
   ms00f80 u0_int_maskb_r_reg_9_ (.o(u0_int_maskb_9_),
	.d(n538),
	.ck(clk));
   ms00f80 u0_int_maskb_r_reg_8_ (.o(u0_int_maskb_8_),
	.d(n537),
	.ck(clk));
   ms00f80 u0_int_maskb_r_reg_7_ (.o(u0_int_maskb_7_),
	.d(n536),
	.ck(clk));
   ms00f80 u0_int_maskb_r_reg_6_ (.o(u0_int_maskb_6_),
	.d(n535),
	.ck(clk));
   ms00f80 u0_int_maskb_r_reg_5_ (.o(u0_int_maskb_5_),
	.d(n534),
	.ck(clk));
   ms00f80 u0_int_maskb_r_reg_4_ (.o(u0_int_maskb_4_),
	.d(n533),
	.ck(clk));
   ms00f80 u0_int_maskb_r_reg_3_ (.o(u0_int_maskb_3_),
	.d(n532),
	.ck(clk));
   ms00f80 u0_int_maskb_r_reg_2_ (.o(u0_int_maskb_2_),
	.d(n531),
	.ck(clk));
   ms00f80 u0_int_maskb_r_reg_1_ (.o(u0_int_maskb_1_),
	.d(n530),
	.ck(clk));
   ms00f80 u0_int_maskb_r_reg_0_ (.o(u0_int_maskb_0_),
	.d(n529),
	.ck(clk));
   ms00f80 u0_int_maska_r_reg_0_ (.o(u0_int_maska_0_),
	.d(n528),
	.ck(clk));
   ms00f80 u0_int_maska_r_reg_1_ (.o(u0_int_maska_1_),
	.d(n527),
	.ck(clk));
   ms00f80 u0_int_maska_r_reg_2_ (.o(u0_int_maska_2_),
	.d(n526),
	.ck(clk));
   ms00f80 u0_int_maska_r_reg_3_ (.o(u0_int_maska_3_),
	.d(n525),
	.ck(clk));
   ms00f80 u0_int_maska_r_reg_4_ (.o(u0_int_maska_4_),
	.d(n524),
	.ck(clk));
   ms00f80 u0_int_maska_r_reg_5_ (.o(u0_int_maska_5_),
	.d(n523),
	.ck(clk));
   ms00f80 u0_int_maska_r_reg_6_ (.o(u0_int_maska_6_),
	.d(n522),
	.ck(clk));
   ms00f80 u0_int_maska_r_reg_7_ (.o(u0_int_maska_7_),
	.d(n521),
	.ck(clk));
   ms00f80 u0_int_maska_r_reg_8_ (.o(u0_int_maska_8_),
	.d(n520),
	.ck(clk));
   ms00f80 u0_int_maska_r_reg_9_ (.o(u0_int_maska_9_),
	.d(n519),
	.ck(clk));
   ms00f80 u0_int_maska_r_reg_10_ (.o(u0_int_maska_10_),
	.d(n518),
	.ck(clk));
   ms00f80 u0_int_maska_r_reg_11_ (.o(u0_int_maska_11_),
	.d(n517),
	.ck(clk));
   ms00f80 u0_int_maska_r_reg_12_ (.o(u0_int_maska_12_),
	.d(n516),
	.ck(clk));
   ms00f80 u0_int_maska_r_reg_13_ (.o(u0_int_maska_13_),
	.d(n515),
	.ck(clk));
   ms00f80 u0_int_maska_r_reg_14_ (.o(u0_int_maska_14_),
	.d(n514),
	.ck(clk));
   ms00f80 u0_int_maska_r_reg_15_ (.o(u0_int_maska_15_),
	.d(n513),
	.ck(clk));
   ms00f80 u0_int_maska_r_reg_16_ (.o(u0_int_maska_16_),
	.d(n512),
	.ck(clk));
   ms00f80 u0_int_maska_r_reg_17_ (.o(u0_int_maska_17_),
	.d(n511),
	.ck(clk));
   ms00f80 u0_int_maska_r_reg_18_ (.o(u0_int_maska_18_),
	.d(n510),
	.ck(clk));
   ms00f80 u0_int_maska_r_reg_19_ (.o(u0_int_maska_19_),
	.d(n509),
	.ck(clk));
   ms00f80 u0_int_maska_r_reg_20_ (.o(u0_int_maska_20_),
	.d(n508),
	.ck(clk));
   ms00f80 u0_int_maska_r_reg_21_ (.o(u0_int_maska_21_),
	.d(n507),
	.ck(clk));
   ms00f80 u0_int_maska_r_reg_22_ (.o(u0_int_maska_22_),
	.d(n506),
	.ck(clk));
   ms00f80 u0_int_maska_r_reg_23_ (.o(u0_int_maska_23_),
	.d(n505),
	.ck(clk));
   ms00f80 u0_int_maska_r_reg_24_ (.o(u0_int_maska_24_),
	.d(n504),
	.ck(clk));
   ms00f80 u0_int_maska_r_reg_25_ (.o(u0_int_maska_25_),
	.d(n503),
	.ck(clk));
   ms00f80 u0_int_maska_r_reg_26_ (.o(u0_int_maska_26_),
	.d(n502),
	.ck(clk));
   ms00f80 u0_int_maska_r_reg_27_ (.o(u0_int_maska_27_),
	.d(n501),
	.ck(clk));
   ms00f80 u0_int_maska_r_reg_28_ (.o(u0_int_maska_28_),
	.d(n500),
	.ck(clk));
   ms00f80 u0_int_maska_r_reg_29_ (.o(u0_int_maska_29_),
	.d(n499),
	.ck(clk));
   ms00f80 u0_int_maska_r_reg_30_ (.o(u0_int_maska_30_),
	.d(n498),
	.ck(clk));
   no02m08 U1746 (.o(n2254),
	.b(n1425),
	.a(n2253));
   in01s01 U1747 (.o(n2253),
	.a(u0_int_maskb_23_));
   no02s06 U1748 (.o(n2297),
	.b(n2296),
	.a(n1425));
   in01s01 U1749 (.o(n2296),
	.a(u0_int_maskb_26_));
   ao22s08 U1750 (.o(n1873),
	.d(slv0_adr[4]),
	.c(u0_int_maskb_0_),
	.b(u0_int_maska_0_),
	.a(FE_OCPN139_slv0_adr_2_));
   no02s02 U1751 (.o(n1528),
	.b(FE_OCPN78_n2056),
	.a(ch0_csr[11]));
   in01s03 U1752 (.o(n1975),
	.a(ch0_csr[6]));
   na02m20 U1754 (.o(n1940),
	.b(FE_OCPN511_slv0_adr_3_),
	.a(slv0_adr[4]));
   in01f20 U1755 (.o(n1557),
	.a(n1581));
   na02m06 U1756 (.o(n1552),
	.b(FE_OCPN544_n2159),
	.a(u0_int_maskb_1_));
   na02f03 U1757 (.o(n1551),
	.b(n2343),
	.a(u0_int_maska_1_));
   na02s02 U1758 (.o(n1636),
	.b(wb0_addr_i[0]),
	.a(wb1_cyc_o));
   na02s02 U1759 (.o(n1631),
	.b(wb0_we_i),
	.a(wb1_cyc_o));
   na02s01 U1760 (.o(n1667),
	.b(wb0_addr_i[18]),
	.a(FE_OCPN661_wb1_cyc_o));
   na02s02 U1761 (.o(n1665),
	.b(wb0_addr_i[17]),
	.a(FE_OCPN651_wb1_cyc_o));
   na02s02 U1762 (.o(n1637),
	.b(wb0_addr_i[1]),
	.a(wb1_cyc_o));
   na02s01 U1763 (.o(n1697),
	.b(wb0s_data_i[9]),
	.a(FE_OCPN277_wb0_cyc_o));
   na02s01 U1764 (.o(n1693),
	.b(wb0s_data_i[5]),
	.a(FE_OCPN277_wb0_cyc_o));
   na02s01 U1765 (.o(n1692),
	.b(wb0s_data_i[4]),
	.a(n1414));
   na02s01 U1766 (.o(n1691),
	.b(wb0s_data_i[3]),
	.a(FE_RN_17));
   na02s01 U1767 (.o(n1688),
	.b(wb0s_data_i[0]),
	.a(FE_RN_17));
   na02s01 U1768 (.o(n1713),
	.b(wb0s_data_i[25]),
	.a(FE_OCPN277_wb0_cyc_o));
   na02s01 U1769 (.o(n1706),
	.b(wb0s_data_i[18]),
	.a(FE_OCPN277_wb0_cyc_o));
   na02s01 U1770 (.o(n1705),
	.b(wb0s_data_i[17]),
	.a(n1414));
   na02s02 U1771 (.o(n1704),
	.b(wb0s_data_i[16]),
	.a(wb0_cyc_o));
   na02s01 U1772 (.o(n1701),
	.b(wb0s_data_i[13]),
	.a(FE_OCPN284_wb0_cyc_o));
   na02s01 U1773 (.o(n1836),
	.b(wb1_we_i),
	.a(FE_RN_17));
   na02s01 U1774 (.o(n1729),
	.b(u4_u1_rf_ack),
	.a(n1442));
   na02s01 U1775 (.o(n1720),
	.b(wb0_rty_i),
	.a(FE_OCPN277_wb0_cyc_o));
   na02s01 U1776 (.o(n1719),
	.b(wb0s_data_i[31]),
	.a(FE_OCPN277_wb0_cyc_o));
   na02s01 U1777 (.o(n1718),
	.b(wb0s_data_i[30]),
	.a(FE_OCPN277_wb0_cyc_o));
   na02s01 U1778 (.o(n1716),
	.b(wb0s_data_i[28]),
	.a(FE_RN_17));
   na02s02 U1779 (.o(n1843),
	.b(wb1_addr_i[2]),
	.a(wb0_cyc_o));
   na02s01 U1780 (.o(n1842),
	.b(wb1_addr_i[1]),
	.a(FE_OCPN277_wb0_cyc_o));
   na02s01 U1781 (.o(n1841),
	.b(wb1_addr_i[0]),
	.a(FE_OCPN284_wb0_cyc_o));
   no02s01 U1782 (.o(n1839),
	.b(wb1_sel_i[2]),
	.a(n1442));
   na02s01 U1783 (.o(n1857),
	.b(wb1_addr_i[16]),
	.a(n1414));
   na02s01 U1784 (.o(n2389),
	.b(wb1m_data_i[9]),
	.a(FE_OCPN277_wb0_cyc_o));
   na02s01 U1785 (.o(n2388),
	.b(FE_OCPN528_n1597),
	.a(de_csr[9]));
   in01s01 U1786 (.o(n1765),
	.a(de_csr[9]));
   no02s20 U1787 (.o(n1414),
	.b(n1725),
	.a(n2364));
   in01s10 U1788 (.o(n2364),
	.a(wb1_cyc_i));
   na02s01 U1789 (.o(n2418),
	.b(FE_OCPN528_n1597),
	.a(de_csr[24]));
   in01s01 U1790 (.o(n1810),
	.a(de_csr[24]));
   in01s01 U1791 (.o(n2252),
	.a(slv0_dout[23]));
   in01s01 U1792 (.o(n2249),
	.a(u0_int_maska_23_));
   in01s01 U1794 (.o(n2267),
	.a(slv0_dout[24]));
   in01s01 U1795 (.o(n2264),
	.a(u0_int_maska_24_));
   in01s02 U1796 (.o(n2278),
	.a(u0_int_maska_25_));
   in01s01 U1797 (.o(n2292),
	.a(u0_int_maska_26_));
   in01s01 U1798 (.o(n2310),
	.a(u0_int_maska_27_));
   in01s01 U1799 (.o(n2320),
	.a(u0_int_maska_28_));
   in01s01 U1800 (.o(n2330),
	.a(u0_int_maska_29_));
   in01s01 U1801 (.o(n2340),
	.a(u0_int_maska_30_));
   in01s02 U1802 (.o(n2005),
	.a(slv0_dout[8]));
   in01s01 U1803 (.o(n2002),
	.a(u0_int_maska_8_));
   in01m01 U1804 (.o(n2023),
	.a(slv0_dout[9]));
   in01s01 U1805 (.o(n2021),
	.a(u0_int_maska_9_));
   in01s02 U1806 (.o(n2037),
	.a(slv0_dout[10]));
   in01s01 U1807 (.o(n2034),
	.a(u0_int_maska_10_));
   in01s02 U1808 (.o(n2054),
	.a(slv0_dout[11]));
   in01s01 U1809 (.o(n2050),
	.a(u0_int_maska_11_));
   in01s01 U1810 (.o(n2074),
	.a(slv0_dout[12]));
   in01s01 U1811 (.o(n2073),
	.a(u0_int_maska_12_));
   in01s01 U1812 (.o(n2088),
	.a(slv0_dout[13]));
   in01s01 U1813 (.o(n2087),
	.a(u0_int_maska_13_));
   in01s02 U1814 (.o(n2104),
	.a(slv0_dout[14]));
   in01s01 U1815 (.o(n2103),
	.a(u0_int_maska_14_));
   in01s02 U1816 (.o(n2120),
	.a(slv0_dout[15]));
   in01s01 U1817 (.o(n2116),
	.a(u0_int_maska_15_));
   in01s01 U1818 (.o(n2134),
	.a(u0_int_maska_16_));
   in01s01 U1819 (.o(n2152),
	.a(u0_int_maska_17_));
   in01s01 U1820 (.o(n2174),
	.a(u0_int_maska_18_));
   in01s01 U1821 (.o(n2191),
	.a(u0_int_maska_19_));
   in01s03 U1822 (.o(n2211),
	.a(slv0_dout[20]));
   in01s01 U1823 (.o(n2210),
	.a(u0_int_maska_20_));
   in01s03 U1824 (.o(n2222),
	.a(slv0_dout[21]));
   in01s01 U1825 (.o(n2221),
	.a(u0_int_maska_21_));
   in01s01 U1826 (.o(n2234),
	.a(u0_int_maska_22_));
   in01s01 U1827 (.o(n1974),
	.a(slv0_dout[6]));
   na02f40 U1828 (.o(n1591),
	.b(n1522),
	.a(FE_OCPN552_n1424));
   in01s01 U1830 (.o(n1969),
	.a(u0_int_maskb_6_));
   in01s01 U1832 (.o(n1956),
	.a(slv0_dout[5]));
   in01s01 U1833 (.o(n1954),
	.a(u0_int_maskb_5_));
   oa22m02 U1834 (.o(n533),
	.d(n1935),
	.c(n1591),
	.b(n1472),
	.a(FE_OCPN385_n1579));
   in01s01 U1835 (.o(n1472),
	.a(u0_int_maskb_4_));
   oa12s02 U1836 (.o(n532),
	.c(n1914),
	.b(FE_RN_18),
	.a(n1910));
   in01s02 U1837 (.o(n1895),
	.a(u0_int_maskb_2_));
   na02m04 U1838 (.o(n1887),
	.b(FE_OCPN384_n1579),
	.a(slv0_dout[2]));
   oa12s02 U1839 (.o(n530),
	.c(n1883),
	.b(FE_RN_18),
	.a(n1535));
   na02s04 U1840 (.o(n1535),
	.b(u0_int_maskb_1_),
	.a(FE_RN_18));
   oa12f02 U1841 (.o(n529),
	.c(FE_OCPN385_n1579),
	.b(n1876),
	.a(n1614));
   in01s02 U1842 (.o(n1876),
	.a(u0_int_maskb_0_));
   na02f04 U1843 (.o(n1614),
	.b(FE_OCPN618_n1591),
	.a(slv0_dout[0]));
   in01s01 U1844 (.o(n1875),
	.a(u0_int_maska_0_));
   na02s04 U1845 (.o(n1628),
	.b(n1426),
	.a(slv0_dout[0]));
   oa12s02 U1847 (.o(n527),
	.c(n1883),
	.b(FE_OCPN540_n1595),
	.a(n1563));
   in01s02 U1848 (.o(n1563),
	.a(n1541));
   no02s04 U1849 (.o(n1541),
	.b(n1426),
	.a(n1542));
   in01s01 U1850 (.o(n1542),
	.a(u0_int_maska_1_));
   in01s02 U1852 (.o(n1894),
	.a(u0_int_maska_2_));
   na02s04 U1853 (.o(n1911),
	.b(u0_int_maska_3_),
	.a(FE_OCPN537_n1595));
   na02m06 U1854 (.o(n1934),
	.b(u0_int_maska_4_),
	.a(FE_OCPN539_n1595));
   in01s01 U1855 (.o(n1955),
	.a(u0_int_maska_5_));
   na02m20 U1857 (.o(n1580),
	.b(n1562),
	.a(FE_OCPN163_n2346));
   oa22m04 U1858 (.o(n522),
	.d(FE_OCPN676_n1580),
	.c(n1970),
	.b(FE_OCPN538_n1595),
	.a(n1974));
   in01s01 U1859 (.o(n1970),
	.a(u0_int_maska_6_));
   in01s01 U1860 (.o(n1989),
	.a(slv0_dout[7]));
   in01s01 U1861 (.o(n1985),
	.a(u0_int_maska_7_));
   in01s01 U1862 (.o(n1943),
	.a(ch0_adr1[4]));
   in01s01 U1863 (.o(n1935),
	.a(slv0_dout[4]));
   in01s01 U1864 (.o(n1920),
	.a(ch0_adr1[3]));
   in01s01 U1865 (.o(n1488),
	.a(slv0_dout[2]));
   in01s01 U1866 (.o(n1898),
	.a(ch0_adr1[2]));
   in01s01 U1867 (.o(n1527),
	.a(n1528));
   no02s08 U1868 (.o(n1524),
	.b(FE_OCPN365_n2194),
	.a(n1525));
   in01s01 U1869 (.o(n1525),
	.a(slv0_dout[0]));
   na02s01 U1870 (.o(n1638),
	.b(ch0_csr[0]),
	.a(FE_OCPN79_n2056));
   oa12s04 U1871 (.o(n560),
	.c(n2072),
	.b(n2223),
	.a(FE_OCPN79_n2056));
   in01s02 U1872 (.o(n2223),
	.a(ch0_csr[21]));
   no02s08 U1873 (.o(n2072),
	.b(n2156),
	.a(n1622));
   in01s02 U1874 (.o(n1622),
	.a(slv0_re));
   in01s01 U1878 (.o(n2339),
	.a(u0_int_maskb_30_));
   in01s02 U1879 (.o(n2332),
	.a(slv0_dout[29]));
   na02f08 U1882 (.o(n1579),
	.b(n1484),
	.a(FE_OCPN163_n2346));
   in01s01 U1883 (.o(n2329),
	.a(u0_int_maskb_29_));
   in01s02 U1884 (.o(n2322),
	.a(slv0_dout[28]));
   in01s01 U1885 (.o(n2319),
	.a(u0_int_maskb_28_));
   in01s01 U1886 (.o(n2309),
	.a(u0_int_maskb_27_));
   in01s01 U1887 (.o(n2295),
	.a(slv0_dout[26]));
   in01s01 U1888 (.o(n2281),
	.a(slv0_dout[25]));
   in01s01 U1889 (.o(n2282),
	.a(u0_int_maskb_25_));
   in01s01 U1890 (.o(n2268),
	.a(u0_int_maskb_24_));
   in01s02 U1891 (.o(n2237),
	.a(slv0_dout[22]));
   in01s01 U1892 (.o(n2238),
	.a(u0_int_maskb_22_));
   in01s02 U1893 (.o(n1914),
	.a(slv0_dout[3]));
   na02f06 U1894 (.o(n1912),
	.b(ch0_txsz[3]),
	.a(FE_RN_9));
   na02s02 U1895 (.o(n1889),
	.b(ch0_txsz[2]),
	.a(FE_RN_9));
   in01s02 U1896 (.o(n1883),
	.a(slv0_dout[1]));
   na02s03 U1897 (.o(n1881),
	.b(ch0_txsz[1]),
	.a(FE_RN_9));
   in01s01 U1898 (.o(n1687),
	.a(ch0_adr1[31]));
   in01s02 U1899 (.o(n2342),
	.a(slv0_dout[30]));
   oa12f02 U1900 (.o(n635),
	.c(FE_OCPN179_n1521),
	.b(n2334),
	.a(n1685));
   in01s01 U1901 (.o(n2334),
	.a(ch0_adr1[29]));
   in01s01 U1902 (.o(n2324),
	.a(ch0_adr1[28]));
   in01s02 U1903 (.o(n2312),
	.a(slv0_dout[27]));
   in01m01 U1904 (.o(n2314),
	.a(ch0_adr1[27]));
   in01s01 U1905 (.o(n2300),
	.a(ch0_adr1[26]));
   in01s01 U1906 (.o(n2284),
	.a(ch0_adr1[25]));
   in01s01 U1907 (.o(n2270),
	.a(ch0_adr1[24]));
   na02f03 U1908 (.o(n1677),
	.b(FE_OCPN178_n1521),
	.a(slv0_dout[24]));
   in01s01 U1909 (.o(n2256),
	.a(ch0_adr1[23]));
   in01s02 U1910 (.o(n2240),
	.a(ch0_adr1[22]));
   na02s02 U1912 (.o(n675),
	.b(n2003),
	.a(n1534));
   in01s01 U1913 (.o(n1987),
	.a(ch0_adr0[7]));
   na02s04 U1914 (.o(n1986),
	.b(slv0_dout[7]),
	.a(n1573));
   in01s01 U1915 (.o(n1972),
	.a(ch0_adr0[6]));
   in01s01 U1916 (.o(n1953),
	.a(ch0_adr0[5]));
   in01s01 U1917 (.o(n1933),
	.a(ch0_adr0[4]));
   in01s01 U1918 (.o(n1916),
	.a(ch0_adr0[3]));
   in01s01 U1919 (.o(n1904),
	.a(ch0_adr0[2]));
   oa12s02 U1920 (.o(n655),
	.c(n2005),
	.b(n1513),
	.a(n2004));
   oa12m02 U1921 (.o(n746),
	.c(n2295),
	.b(n1513),
	.a(n2294));
   na02m40 U1923 (.o(n1890),
	.b(n1544),
	.a(n1545));
   in01s01 U1925 (.o(n2369),
	.a(ch0_csr[2]));
   oa12s02 U1927 (.o(n732),
	.c(FE_OCPN363_n2194),
	.b(n1914),
	.a(n1913));
   na02s03 U1928 (.o(n1913),
	.b(ch0_csr[3]),
	.a(FE_OCPN363_n2194));
   oa12f02 U1929 (.o(n731),
	.c(FE_OCPN367_n2194),
	.b(n1937),
	.a(n1936));
   in01s01 U1930 (.o(n1937),
	.a(ch0_csr[4]));
   na02m06 U1931 (.o(n1936),
	.b(slv0_dout[4]),
	.a(FE_OCPN367_n2194));
   in01s01 U1932 (.o(n2358),
	.a(ch0_adr0[31]));
   in01s01 U1933 (.o(n2302),
	.a(ch0_adr0[26]));
   in01s01 U1934 (.o(n2286),
	.a(ch0_adr0[25]));
   in01s01 U1935 (.o(n2272),
	.a(ch0_adr0[24]));
   oa12s01 U1936 (.o(n808),
	.c(FE_OFN427_wb0_ack_i),
	.b(n1807),
	.a(n2478));
   in01s01 U1937 (.o(n1807),
	.a(de_csr[23]));
   oa12s01 U1938 (.o(n807),
	.c(wb0_ack_i),
	.b(n1810),
	.a(n2477));
   oa12s01 U1939 (.o(n806),
	.c(FE_OFN427_wb0_ack_i),
	.b(n1813),
	.a(n2476));
   in01s01 U1940 (.o(n1813),
	.a(de_csr[25]));
   oa12s01 U1941 (.o(n805),
	.c(wb0_ack_i),
	.b(n1816),
	.a(n2475));
   oa12s01 U1942 (.o(n804),
	.c(FE_OFN427_wb0_ack_i),
	.b(n1819),
	.a(n2474));
   in01s01 U1943 (.o(n1819),
	.a(de_csr[27]));
   oa12s01 U1944 (.o(n803),
	.c(wb0_ack_i),
	.b(n1822),
	.a(n2473));
   in01s01 U1945 (.o(n1822),
	.a(de_csr[28]));
   oa12s01 U1946 (.o(n802),
	.c(FE_OFN427_wb0_ack_i),
	.b(n1825),
	.a(n2472));
   in01s01 U1947 (.o(n1825),
	.a(de_csr[29]));
   oa12s01 U1948 (.o(n801),
	.c(FE_OFN427_wb0_ack_i),
	.b(n1828),
	.a(n2471));
   in01s01 U1949 (.o(n1828),
	.a(de_csr[30]));
   oa12s01 U1950 (.o(n800),
	.c(FE_OFN427_wb0_ack_i),
	.b(n1831),
	.a(n2470));
   in01s01 U1951 (.o(n1831),
	.a(de_csr[31]));
   oa12m02 U1952 (.o(n767),
	.c(FE_OCPN368_n2194),
	.b(n2199),
	.a(n2193));
   in01s01 U1953 (.o(n2199),
	.a(ch0_csr[19]));
   in01s01 U1954 (.o(n2182),
	.a(ch0_csr[18]));
   in01s01 U1955 (.o(n2157),
	.a(ch0_csr[17]));
   in01s01 U1956 (.o(n2140),
	.a(ch0_csr[16]));
   in01s01 U1957 (.o(n2122),
	.a(ch0_csr[15]));
   in01s01 U1959 (.o(n2110),
	.a(ch0_csr[14]));
   in01s01 U1960 (.o(n1762),
	.a(de_csr[8]));
   oa12s01 U1961 (.o(n822),
	.c(FE_OFN427_wb0_ack_i),
	.b(n1765),
	.a(n2492));
   oa12s01 U1962 (.o(n821),
	.c(wb0_ack_i),
	.b(n1768),
	.a(n2491));
   in01s01 U1963 (.o(n1768),
	.a(de_csr[10]));
   oa12s01 U1964 (.o(n820),
	.c(wb0_ack_i),
	.b(n1771),
	.a(n2490));
   in01s01 U1965 (.o(n1774),
	.a(de_csr[12]));
   in01s01 U1966 (.o(n1777),
	.a(de_csr[13]));
   in01s01 U1967 (.o(n1780),
	.a(de_csr[14]));
   in01s01 U1968 (.o(n1783),
	.a(de_csr[15]));
   in01s01 U1969 (.o(n1786),
	.a(de_csr[16]));
   in01s01 U1970 (.o(n1789),
	.a(de_csr[17]));
   oa12s01 U1971 (.o(n813),
	.c(FE_OFN427_wb0_ack_i),
	.b(n1792),
	.a(n2483));
   in01s01 U1972 (.o(n1792),
	.a(de_csr[18]));
   oa12s01 U1973 (.o(n812),
	.c(wb0_ack_i),
	.b(n1795),
	.a(n2482));
   oa12s01 U1974 (.o(n811),
	.c(FE_OFN427_wb0_ack_i),
	.b(n1798),
	.a(n2481));
   in01s01 U1975 (.o(n1798),
	.a(de_csr[20]));
   oa12s01 U1976 (.o(n810),
	.c(FE_OFN427_wb0_ack_i),
	.b(n1801),
	.a(n2480));
   in01s01 U1977 (.o(n1801),
	.a(de_csr[21]));
   no02s06 U1979 (.o(n1496),
	.b(n2355),
	.a(n1497));
   in01f10 U1980 (.o(n2355),
	.a(n2241));
   no02s06 U1981 (.o(n1497),
	.b(FE_OCPN562_n2357),
	.a(n2326));
   in01s01 U1982 (.o(n2326),
	.a(ch0_adr0[28]));
   no02m04 U1983 (.o(n1499),
	.b(n2355),
	.a(n1500));
   in01s01 U1984 (.o(n2347),
	.a(ch0_adr1[30]));
   no02f04 U1985 (.o(n1502),
	.b(n2355),
	.a(n1503));
   in01s04 U1986 (.o(n1554),
	.a(n1555));
   no04s02 U1987 (.o(u4_u1_N3),
	.d(wb1_we_i),
	.c(n1723),
	.b(slv1_re),
	.a(n1724));
   no02s02 U1988 (.o(n1727),
	.b(u4_u1_rf_ack),
	.a(n1722));
   in01s01 U1989 (.o(n893),
	.a(n1728));
   in01s01 U1991 (.o(u4_u1_N4),
	.a(n1726));
   oa12s01 U1992 (.o(n831),
	.c(wb0_ack_i),
	.b(n1730),
	.a(n2501));
   in01s01 U1993 (.o(n1730),
	.a(de_csr[0]));
   oa12s01 U1994 (.o(n830),
	.c(wb0_ack_i),
	.b(n1741),
	.a(n2500));
   in01s01 U1995 (.o(n1741),
	.a(de_csr[1]));
   oa12s01 U1996 (.o(n829),
	.c(wb0_ack_i),
	.b(n1744),
	.a(n2499));
   in01s01 U1997 (.o(n1744),
	.a(de_csr[2]));
   oa12s01 U1998 (.o(n828),
	.c(wb0_ack_i),
	.b(n1747),
	.a(n2498));
   in01s01 U1999 (.o(n1747),
	.a(de_csr[3]));
   in01s01 U2000 (.o(n1753),
	.a(de_csr[5]));
   in01s01 U2001 (.o(n1756),
	.a(de_csr[6]));
   in01s01 U2002 (.o(n1759),
	.a(de_csr[7]));
   na02m02 U2003 (.o(u0_N3074),
	.b(n1489),
	.a(n1491));
   na02s04 U2004 (.o(n1491),
	.b(ch0_adr1[31]),
	.a(n2356));
   no02f04 U2005 (.o(n1489),
	.b(n2355),
	.a(n1490));
   no02m02 U2006 (.o(n1490),
	.b(FE_OCPN565_n2357),
	.a(n2358));
   na02f20 U2007 (.o(n1474),
	.b(n1940),
	.a(n1939));
   no02s01 U2008 (.o(n2466),
	.b(n1872),
	.a(n1876));
   na02s02 U2009 (.o(n1872),
	.b(ch0_csr[21]),
	.a(ch0_csr[18]));
   no02s01 U2010 (.o(n2465),
	.b(n1417),
	.a(n1875));
   na02s01 U2011 (.o(n1417),
	.b(ch0_csr[21]),
	.a(ch0_csr[18]));
   in01s01 U2012 (.o(n1884),
	.a(ch0_csr[1]));
   ao22f04 U2013 (.o(n1549),
	.d(n2304),
	.c(ch0_txsz[1]),
	.b(FE_OCPN163_n2346),
	.a(n1550));
   na02s08 U2018 (.o(n1946),
	.b(ch0_adr0[4]),
	.a(n1416));
   na02s08 U2020 (.o(n1964),
	.b(ch0_adr0[5]),
	.a(n1416));
   no02f08 U2021 (.o(n1998),
	.b(FE_OCPN673_n1577),
	.a(n1996));
   na02s06 U2022 (.o(n1997),
	.b(ch0_adr0[7]),
	.a(n1416));
   na02m04 U2023 (.o(n2015),
	.b(ch0_adr0[8]),
	.a(n1416));
   no02f08 U2025 (.o(n2031),
	.b(FE_OCPN673_n1577),
	.a(n2028));
   na02s06 U2026 (.o(n2030),
	.b(ch0_adr0[9]),
	.a(n1416));
   na02s06 U2027 (.o(n2029),
	.b(ch0_txsz[9]),
	.a(n2304));
   in01s03 U2029 (.o(n2047),
	.a(n2039));
   in01s01 U2030 (.o(n2038),
	.a(ch0_txsz[10]));
   no02f06 U2031 (.o(n2046),
	.b(FE_OCPN673_n1577),
	.a(n2044));
   na02m04 U2032 (.o(n2045),
	.b(ch0_adr0[10]),
	.a(n1416));
   na02s06 U2034 (.o(n2080),
	.b(ch0_adr0[12]),
	.a(n2165));
   in01s01 U2035 (.o(wb1_sel_o[1]),
	.a(n1633));
   in01s01 U2036 (.o(wb1_sel_o[0]),
	.a(n1632));
   na02m01 U2037 (.o(wb1_addr_o[16]),
	.b(wb1_cyc_o),
	.a(n1663));
   na02s02 U2038 (.o(n1663),
	.b(wb0_addr_i[16]),
	.a(FE_OCPN651_wb1_cyc_o));
   na02s02 U2040 (.o(n1662),
	.b(wb0_addr_i[15]),
	.a(FE_OCPN651_wb1_cyc_o));
   na02s02 U2041 (.o(wb1_addr_o[13]),
	.b(wb1_cyc_o),
	.a(n1660));
   na02s02 U2042 (.o(n1660),
	.b(wb0_addr_i[13]),
	.a(FE_OCPN651_wb1_cyc_o));
   na02s01 U2043 (.o(wb1_addr_o[12]),
	.b(wb1_cyc_o),
	.a(n1658));
   na02s02 U2044 (.o(n1658),
	.b(wb0_addr_i[12]),
	.a(FE_OCPN651_wb1_cyc_o));
   na02m01 U2045 (.o(wb1_addr_o[11]),
	.b(wb1_cyc_o),
	.a(n1656));
   na02s02 U2046 (.o(n1656),
	.b(wb0_addr_i[11]),
	.a(FE_OCPN651_wb1_cyc_o));
   na02s02 U2047 (.o(wb1_addr_o[10]),
	.b(wb1_cyc_o),
	.a(n1654));
   na02s02 U2048 (.o(n1654),
	.b(wb0_addr_i[10]),
	.a(FE_OCPN651_wb1_cyc_o));
   oa12s01 U2049 (.o(wb1_addr_o[9]),
	.c(n1653),
	.b(FE_OCPN656_wb1_cyc_o),
	.a(wb1_cyc_o));
   in01s01 U2050 (.o(n1653),
	.a(wb0_addr_i[9]));
   in01s01 U2051 (.o(n1652),
	.a(wb0_addr_i[8]));
   in01s01 U2052 (.o(n1651),
	.a(wb0_addr_i[7]));
   oa12s01 U2053 (.o(wb1_addr_o[6]),
	.c(n1649),
	.b(FE_OCPN658_wb1_cyc_o),
	.a(wb1_cyc_o));
   in01s01 U2054 (.o(n1649),
	.a(wb0_addr_i[6]));
   oa12s01 U2055 (.o(wb1_addr_o[5]),
	.c(n1647),
	.b(FE_OCPN656_wb1_cyc_o),
	.a(wb1_cyc_o));
   in01s01 U2056 (.o(n1647),
	.a(wb0_addr_i[5]));
   in01s01 U2057 (.o(n1645),
	.a(wb0_addr_i[4]));
   in01s01 U2058 (.o(n1643),
	.a(wb0_addr_i[3]));
   in01s01 U2059 (.o(n1641),
	.a(wb0_addr_i[2]));
   na02s01 U2060 (.o(wb1_addr_o[31]),
	.b(n1735),
	.a(wb1_cyc_o));
   na02s01 U2061 (.o(wb1_addr_o[28]),
	.b(n1733),
	.a(wb1_cyc_o));
   na02s01 U2062 (.o(wb1_addr_o[27]),
	.b(wb1_cyc_o),
	.a(n1683));
   na02s02 U2063 (.o(wb1_addr_o[26]),
	.b(wb1_cyc_o),
	.a(n1682));
   na02s02 U2064 (.o(n1682),
	.b(wb0_addr_i[26]),
	.a(FE_OCPN666_wb1_cyc_o));
   na02s01 U2067 (.o(wb1_addr_o[24]),
	.b(wb1_cyc_o),
	.a(n1678));
   na02s01 U2068 (.o(n1678),
	.b(wb0_addr_i[24]),
	.a(FE_OCPN661_wb1_cyc_o));
   na02s02 U2069 (.o(wb1_addr_o[23]),
	.b(wb1_cyc_o),
	.a(n1676));
   na02s02 U2070 (.o(n1676),
	.b(wb0_addr_i[23]),
	.a(FE_OCPN666_wb1_cyc_o));
   na02s02 U2071 (.o(n1674),
	.b(wb0_addr_i[22]),
	.a(FE_OCPN642_wb1_cyc_o));
   na02s01 U2072 (.o(wb1_addr_o[21]),
	.b(wb1_cyc_o),
	.a(n1673));
   na02s02 U2073 (.o(n1673),
	.b(wb0_addr_i[21]),
	.a(FE_OCPN651_wb1_cyc_o));
   na02s01 U2074 (.o(wb1_addr_o[20]),
	.b(wb1_cyc_o),
	.a(n1671));
   na02s01 U2075 (.o(n1671),
	.b(wb0_addr_i[20]),
	.a(FE_OCPN661_wb1_cyc_o));
   na02s01 U2076 (.o(wb1_addr_o[19]),
	.b(wb1_cyc_o),
	.a(n1669));
   na02s01 U2077 (.o(n1669),
	.b(wb0_addr_i[19]),
	.a(FE_OCPN659_wb1_cyc_o));
   in01s01 U2078 (.o(wb1m_data_o[14]),
	.a(n1702));
   na02s01 U2079 (.o(n1702),
	.b(wb0s_data_i[14]),
	.a(FE_OCPN284_wb0_cyc_o));
   in01s01 U2080 (.o(wb1m_data_o[10]),
	.a(n1698));
   na02s01 U2081 (.o(n1698),
	.b(wb0s_data_i[10]),
	.a(n1414));
   in01s01 U2082 (.o(wb1m_data_o[8]),
	.a(n1696));
   in01s01 U2083 (.o(wb1m_data_o[7]),
	.a(n1695));
   na02s01 U2084 (.o(n1695),
	.b(wb0s_data_i[7]),
	.a(FE_OCPN277_wb0_cyc_o));
   in01s01 U2085 (.o(wb1m_data_o[6]),
	.a(n1694));
   na02s01 U2086 (.o(n1694),
	.b(wb0s_data_i[6]),
	.a(FE_OCPN277_wb0_cyc_o));
   in01s01 U2087 (.o(wb1m_data_o[2]),
	.a(n1690));
   na02s01 U2088 (.o(n1690),
	.b(wb0s_data_i[2]),
	.a(FE_RN_17));
   in01s01 U2089 (.o(wb1m_data_o[23]),
	.a(n1711));
   in01s01 U2090 (.o(wb1m_data_o[22]),
	.a(n1710));
   na02s01 U2091 (.o(n1710),
	.b(wb0s_data_i[22]),
	.a(FE_OCPN277_wb0_cyc_o));
   in01s01 U2092 (.o(wb1m_data_o[21]),
	.a(n1709));
   na02s01 U2093 (.o(n1709),
	.b(wb0s_data_i[21]),
	.a(n1414));
   in01s01 U2094 (.o(wb1m_data_o[20]),
	.a(n1708));
   na02s01 U2095 (.o(n1708),
	.b(wb0s_data_i[20]),
	.a(n1414));
   na02s01 U2096 (.o(wb0_addr_o[15]),
	.b(n1414),
	.a(n1856));
   na02s01 U2097 (.o(wb0_addr_o[14]),
	.b(n1414),
	.a(n1855));
   na02s01 U2098 (.o(n1855),
	.b(wb1_addr_i[14]),
	.a(n1414));
   na02s01 U2099 (.o(wb0_addr_o[13]),
	.b(n1414),
	.a(n1854));
   na02s01 U2100 (.o(wb0_addr_o[12]),
	.b(n1414),
	.a(n1853));
   na02s01 U2101 (.o(n1853),
	.b(wb1_addr_i[12]),
	.a(FE_OCPN277_wb0_cyc_o));
   na02s01 U2102 (.o(wb0_addr_o[11]),
	.b(FE_OCPN284_wb0_cyc_o),
	.a(n1852));
   na02s01 U2103 (.o(wb0_addr_o[10]),
	.b(FE_OCPN284_wb0_cyc_o),
	.a(n1851));
   na02s01 U2104 (.o(wb0_addr_o[9]),
	.b(FE_OCPN284_wb0_cyc_o),
	.a(n1850));
   na02s01 U2105 (.o(n1850),
	.b(wb1_addr_i[9]),
	.a(FE_RN_17));
   na02s01 U2106 (.o(wb0_addr_o[8]),
	.b(FE_OCPN284_wb0_cyc_o),
	.a(n1849));
   na02s01 U2107 (.o(wb0_addr_o[7]),
	.b(n1414),
	.a(n1848));
   na02m01 U2108 (.o(wb0_addr_o[6]),
	.b(n1414),
	.a(n1847));
   na02s02 U2109 (.o(n1847),
	.b(wb1_addr_i[6]),
	.a(FE_OCPN284_wb0_cyc_o));
   na02s01 U2110 (.o(wb0_addr_o[5]),
	.b(n1414),
	.a(n1846));
   na02s01 U2111 (.o(n1846),
	.b(wb1_addr_i[5]),
	.a(FE_RN_17));
   na02s01 U2112 (.o(wb0_addr_o[4]),
	.b(n1414),
	.a(n1845));
   na02s01 U2113 (.o(wb0_addr_o[3]),
	.b(n1414),
	.a(n1844));
   na02s01 U2114 (.o(wb0_addr_o[30]),
	.b(n2368),
	.a(FE_RN_17));
   na02s01 U2115 (.o(wb0_addr_o[29]),
	.b(n2366),
	.a(FE_RN_17));
   na02s01 U2116 (.o(wb0_addr_o[28]),
	.b(n2365),
	.a(n1414));
   na02s02 U2117 (.o(wb0_addr_o[27]),
	.b(wb0_cyc_o),
	.a(n1868));
   na02s02 U2118 (.o(wb0_addr_o[26]),
	.b(wb0_cyc_o),
	.a(n1867));
   na02s02 U2119 (.o(n1867),
	.b(wb1_addr_i[26]),
	.a(wb0_cyc_o));
   na02s01 U2120 (.o(wb0_addr_o[25]),
	.b(FE_OCPN284_wb0_cyc_o),
	.a(n1866));
   na02s01 U2121 (.o(wb0_addr_o[24]),
	.b(n1414),
	.a(n1865));
   na02s01 U2122 (.o(wb0_addr_o[23]),
	.b(n1414),
	.a(n1864));
   na02s01 U2123 (.o(n1864),
	.b(wb1_addr_i[23]),
	.a(FE_RN_17));
   na02s01 U2125 (.o(wb0_addr_o[22]),
	.b(n1414),
	.a(n1863));
   na02s01 U2126 (.o(n1863),
	.b(wb1_addr_i[22]),
	.a(FE_RN_17));
   na02s01 U2127 (.o(wb0_addr_o[21]),
	.b(FE_OCPN284_wb0_cyc_o),
	.a(n1862));
   na02s01 U2128 (.o(wb0_addr_o[20]),
	.b(FE_OCPN284_wb0_cyc_o),
	.a(n1861));
   na02s01 U2129 (.o(n1861),
	.b(wb1_addr_i[20]),
	.a(n1414));
   na02s02 U2130 (.o(wb0_addr_o[19]),
	.b(FE_OCPN277_wb0_cyc_o),
	.a(n1860));
   na02s01 U2131 (.o(wb0_addr_o[18]),
	.b(FE_OCPN284_wb0_cyc_o),
	.a(n1859));
   na02s01 U2132 (.o(wb0_addr_o[17]),
	.b(FE_OCPN284_wb0_cyc_o),
	.a(n1858));
   na02s01 U2133 (.o(n1858),
	.b(wb1_addr_i[17]),
	.a(n1414));
   na02s02 U2134 (.o(wb0s_data_o[8]),
	.b(n2386),
	.a(n2387));
   na02s02 U2135 (.o(n2387),
	.b(wb1m_data_i[8]),
	.a(wb0_cyc_o));
   na02s02 U2136 (.o(wb0s_data_o[7]),
	.b(n2384),
	.a(n2385));
   na02s01 U2137 (.o(n2385),
	.b(wb1m_data_i[7]),
	.a(FE_OCPN277_wb0_cyc_o));
   na02s01 U2138 (.o(wb0s_data_o[6]),
	.b(n2382),
	.a(n2383));
   na02s01 U2139 (.o(n2383),
	.b(wb1m_data_i[6]),
	.a(FE_OCPN277_wb0_cyc_o));
   na02s01 U2140 (.o(wb0s_data_o[5]),
	.b(n2380),
	.a(n2381));
   na02s01 U2141 (.o(n2381),
	.b(wb1m_data_i[5]),
	.a(n1414));
   na02s01 U2142 (.o(wb0s_data_o[4]),
	.b(n2378),
	.a(n2379));
   na02s01 U2143 (.o(n2379),
	.b(wb1m_data_i[4]),
	.a(n1414));
   na02s01 U2144 (.o(wb0s_data_o[3]),
	.b(n2376),
	.a(n2377));
   na02s01 U2145 (.o(n2377),
	.b(wb1m_data_i[3]),
	.a(FE_RN_17));
   na02s01 U2146 (.o(wb0s_data_o[2]),
	.b(n2374),
	.a(n2375));
   na02s01 U2147 (.o(wb0s_data_o[1]),
	.b(n2372),
	.a(n2373));
   na02s01 U2148 (.o(n2373),
	.b(wb1m_data_i[1]),
	.a(FE_RN_17));
   na02s01 U2149 (.o(wb0s_data_o[0]),
	.b(n2370),
	.a(n2371));
   na02s01 U2150 (.o(n2371),
	.b(wb1m_data_i[0]),
	.a(FE_RN_17));
   in01s20 U2151 (.o(n1732),
	.a(wb0_cyc_i));
   oa12s01 U2152 (.o(wb0m_data_o[31]),
	.c(n2360),
	.b(FE_OCPN658_wb1_cyc_o),
	.a(n2359));
   na02s01 U2153 (.o(n2359),
	.b(slv0_din[31]),
	.a(FE_OCPN630_wb1_cyc_o));
   na02s01 U2154 (.o(n2351),
	.b(slv0_din[30]),
	.a(FE_OCPN657_wb1_cyc_o));
   na02s01 U2155 (.o(wb0s_data_o[23]),
	.b(n2416),
	.a(n2417));
   na02s01 U2157 (.o(n2416),
	.b(FE_OCPN528_n1597),
	.a(de_csr[23]));
   na02s01 U2158 (.o(wb0s_data_o[22]),
	.b(n2414),
	.a(n2415));
   na02s01 U2159 (.o(n2415),
	.b(wb1m_data_i[22]),
	.a(FE_OCPN277_wb0_cyc_o));
   na02s01 U2160 (.o(n2414),
	.b(FE_OCPN528_n1597),
	.a(de_csr[22]));
   in01s01 U2161 (.o(n1804),
	.a(de_csr[22]));
   na02s01 U2162 (.o(wb0s_data_o[21]),
	.b(n2412),
	.a(n2413));
   na02s01 U2163 (.o(wb0s_data_o[20]),
	.b(n2410),
	.a(n2411));
   na02s01 U2164 (.o(n2410),
	.b(FE_OCPN528_n1597),
	.a(de_csr[20]));
   na02s01 U2165 (.o(wb0s_data_o[19]),
	.b(n2408),
	.a(n2409));
   na02s01 U2166 (.o(n2409),
	.b(wb1m_data_i[19]),
	.a(FE_RN_17));
   na02s01 U2167 (.o(n2408),
	.b(FE_OCPN528_n1597),
	.a(de_csr[19]));
   na02s01 U2168 (.o(wb0s_data_o[18]),
	.b(n2406),
	.a(n2407));
   na02s01 U2169 (.o(n2407),
	.b(wb1m_data_i[18]),
	.a(FE_OCPN277_wb0_cyc_o));
   na02s01 U2170 (.o(wb0s_data_o[17]),
	.b(n2404),
	.a(n2405));
   na02s02 U2171 (.o(n2405),
	.b(wb1m_data_i[17]),
	.a(FE_OCPN284_wb0_cyc_o));
   na02m01 U2172 (.o(wb0s_data_o[16]),
	.b(n2402),
	.a(n2403));
   na02s02 U2173 (.o(n2403),
	.b(wb1m_data_i[16]),
	.a(wb0_cyc_o));
   na02s02 U2174 (.o(wb0s_data_o[15]),
	.b(n2400),
	.a(n2401));
   na02s02 U2175 (.o(n2401),
	.b(wb1m_data_i[15]),
	.a(wb0_cyc_o));
   na02s01 U2176 (.o(wb0s_data_o[14]),
	.b(n2398),
	.a(n2399));
   na02s01 U2177 (.o(n2399),
	.b(wb1m_data_i[14]),
	.a(FE_OCPN284_wb0_cyc_o));
   na02s01 U2178 (.o(n2398),
	.b(FE_OCPN528_n1597),
	.a(de_csr[14]));
   na02s01 U2179 (.o(wb0s_data_o[13]),
	.b(n2396),
	.a(n2397));
   na02s01 U2180 (.o(n2396),
	.b(FE_OCPN528_n1597),
	.a(de_csr[13]));
   na02s01 U2181 (.o(wb0s_data_o[12]),
	.b(n2394),
	.a(n2395));
   na02s01 U2182 (.o(n2395),
	.b(wb1m_data_i[12]),
	.a(FE_RN_17));
   na02s01 U2183 (.o(wb0s_data_o[11]),
	.b(n2392),
	.a(n2393));
   na02s01 U2184 (.o(n2393),
	.b(wb1m_data_i[11]),
	.a(FE_RN_17));
   na02s01 U2185 (.o(wb0s_data_o[10]),
	.b(n2390),
	.a(n2391));
   na02s01 U2186 (.o(wb0s_data_o[31]),
	.b(n2432),
	.a(n2433));
   na02s02 U2187 (.o(n2432),
	.b(FE_OCPN528_n1597),
	.a(de_csr[31]));
   no02s20 U2188 (.o(FE_OCPN277_wb0_cyc_o),
	.b(n1725),
	.a(n2364));
   na02s01 U2190 (.o(wb0s_data_o[30]),
	.b(n2430),
	.a(n2431));
   na02s01 U2191 (.o(n2430),
	.b(FE_OCPN528_n1597),
	.a(de_csr[30]));
   na02s01 U2192 (.o(wb0s_data_o[29]),
	.b(n2428),
	.a(n2429));
   na02s01 U2193 (.o(wb0s_data_o[28]),
	.b(n2426),
	.a(n2427));
   na02s01 U2194 (.o(n2426),
	.b(FE_OCPN528_n1597),
	.a(de_csr[28]));
   na02s01 U2195 (.o(wb0s_data_o[27]),
	.b(n2424),
	.a(n2425));
   na02s02 U2196 (.o(n2424),
	.b(FE_OCPN528_n1597),
	.a(de_csr[27]));
   na02s01 U2197 (.o(wb0s_data_o[26]),
	.b(n2422),
	.a(n2423));
   na02s01 U2198 (.o(n2423),
	.b(wb1m_data_i[26]),
	.a(FE_RN_17));
   na02s01 U2199 (.o(n2422),
	.b(FE_OCPN528_n1597),
	.a(de_csr[26]));
   na02s01 U2200 (.o(wb0s_data_o[25]),
	.b(n2420),
	.a(n2421));
   na02s01 U2201 (.o(n2420),
	.b(FE_OCPN528_n1597),
	.a(de_csr[25]));
   no02f10 U2202 (.o(n2011),
	.b(n1425),
	.a(n2010));
   in01s04 U2203 (.o(n1623),
	.a(ndnr_0_));
   na03m10 U2204 (.o(n1558),
	.c(n1557),
	.b(ch0_csr[0]),
	.a(n1543));
   no02m06 U2205 (.o(n1905),
	.b(n1904),
	.a(FE_OCPN561_n2357));
   in01s02 U2206 (.o(n1442),
	.a(n1414));
   na02s03 U2209 (.o(n1910),
	.b(u0_int_maskb_3_),
	.a(FE_RN_18));
   in01s01 U2210 (.o(n2105),
	.a(u0_int_maskb_14_));
   in01s01 U2211 (.o(n2052),
	.a(ch0_adr0[11]));
   in01f04 U2212 (.o(n2153),
	.a(n1532));
   in01s02 U2213 (.o(n2201),
	.a(ch0_txsz[19]));
   in01s02 U2214 (.o(n1990),
	.a(ch0_csr[7]));
   in01s01 U2215 (.o(n1816),
	.a(de_csr[26]));
   in01s01 U2216 (.o(n1795),
	.a(de_csr[19]));
   in01s01 U2217 (.o(n1771),
	.a(de_csr[11]));
   in01s01 U2218 (.o(n1750),
	.a(de_csr[4]));
   na02s02 U2219 (.o(n1630),
	.b(wb0_stb_i),
	.a(wb1_cyc_o));
   na02s01 U2220 (.o(n1661),
	.b(wb0_addr_i[14]),
	.a(FE_OCPN661_wb1_cyc_o));
   na02s01 U2221 (.o(n1696),
	.b(wb0s_data_i[8]),
	.a(n1414));
   na02s01 U2222 (.o(n1711),
	.b(wb0s_data_i[23]),
	.a(n1414));
   na02s02 U2223 (.o(n1740),
	.b(wb0m_data_i[0]),
	.a(FE_OCPN666_wb1_cyc_o));
   na02s02 U2224 (.o(n1763),
	.b(de_csr[8]),
	.a(FE_RN_1));
   na02s02 U2225 (.o(n1785),
	.b(wb0m_data_i[15]),
	.a(FE_OCPN651_wb1_cyc_o));
   na02s01 U2226 (.o(n1845),
	.b(wb1_addr_i[4]),
	.a(n1414));
   na02s02 U2227 (.o(n1860),
	.b(wb1_addr_i[19]),
	.a(wb0_cyc_o));
   na02s01 U2228 (.o(n2114),
	.b(slv0_din[14]),
	.a(FE_OCPN626_wb1_cyc_o));
   na02s02 U2229 (.o(n2382),
	.b(FE_OCPN528_n1597),
	.a(de_csr[6]));
   na02s01 U2230 (.o(n2412),
	.b(FE_OCPN528_n1597),
	.a(de_csr[21]));
   na02s01 U2231 (.o(n2428),
	.b(FE_OCPN528_n1597),
	.a(de_csr[29]));
   oa22f02 U2233 (.o(n536),
	.d(FE_RN_13),
	.c(n1992),
	.b(n1591),
	.a(n1989));
   oa12f02 U2234 (.o(n587),
	.c(FE_OCPN179_n1521),
	.b(n1961),
	.a(n1646));
   oa12m01 U2235 (.o(n647),
	.c(n1935),
	.b(n1513),
	.a(n1931));
   oa12s01 U2236 (.o(n809),
	.c(FE_OFN427_wb0_ack_i),
	.b(n1804),
	.a(n2479));
   no03s02 U2237 (.o(u3_u1_N4),
	.c(n1610),
	.b(n1611),
	.a(n1612));
   na02s01 U2238 (.o(wb1_addr_o[18]),
	.b(wb1_cyc_o),
	.a(n1667));
   in01s01 U2239 (.o(wb1m_data_o[0]),
	.a(n1688));
   in01s01 U2240 (.o(wb1m_data_o[18]),
	.a(n1706));
   oa12s01 U2241 (.o(wb1_ack_o),
	.c(n1607),
	.b(n1438),
	.a(n1729));
   na02s02 U2242 (.o(wb0_addr_o[2]),
	.b(wb0_cyc_o),
	.a(n1843));
   na02s01 U2243 (.o(wb0_addr_o[16]),
	.b(FE_OCPN284_wb0_cyc_o),
	.a(n1857));
   na02s01 U2244 (.o(wb0s_data_o[9]),
	.b(n2388),
	.a(n2389));
   na02s01 U2245 (.o(wb0s_data_o[24]),
	.b(n2418),
	.a(n2419));
   no02f40 U2247 (.o(n1595),
	.b(n1626),
	.a(n2346));
   in01s03 U2248 (.o(n1874),
	.a(n1621));
   na02s20 U2249 (.o(n1737),
	.b(n1735),
	.a(n1736));
   no02s06 U2250 (.o(n1878),
	.b(n1872),
	.a(n1873));
   no02f10 U2251 (.o(n2041),
	.b(n1425),
	.a(n2040));
   in01m20 U2252 (.o(n2225),
	.a(n2200));
   na02s02 U2253 (.o(n1888),
	.b(n1426),
	.a(slv0_dout[2]));
   in01s01 U2254 (.o(n2190),
	.a(u0_int_maskb_19_));
   na02s04 U2255 (.o(n2056),
	.b(n1624),
	.a(n1975));
   in01m01 U2256 (.o(n1978),
	.a(ch0_adr1[6]));
   na02s03 U2258 (.o(n1686),
	.b(FE_OCPN176_n1521),
	.a(slv0_dout[31]));
   in01s01 U2259 (.o(n2071),
	.a(ch0_adr0[12]));
   in01s01 U2260 (.o(n2154),
	.a(ch0_adr0[17]));
   no02f04 U2261 (.o(n2289),
	.b(n2355),
	.a(n2285));
   na02m06 U2262 (.o(n1980),
	.b(ch0_adr0[6]),
	.a(n1416));
   na02f80 U2263 (.o(n2156),
	.b(n1557),
	.a(n1543));
   na02s02 U2264 (.o(n1700),
	.b(wb0s_data_i[12]),
	.a(FE_OCPN284_wb0_cyc_o));
   na02s01 U2265 (.o(n1715),
	.b(wb0s_data_i[27]),
	.a(FE_OCPN277_wb0_cyc_o));
   na02s01 U2266 (.o(n1745),
	.b(de_csr[2]),
	.a(FE_RN_1));
   na02s02 U2267 (.o(n1767),
	.b(wb0m_data_i[9]),
	.a(FE_OCPN642_wb1_cyc_o));
   na02s02 U2268 (.o(n1790),
	.b(de_csr[17]),
	.a(FE_RN_1));
   na02s01 U2269 (.o(n1835),
	.b(wb1_stb_i),
	.a(FE_RN_17));
   na02s01 U2270 (.o(n1848),
	.b(wb1_addr_i[7]),
	.a(FE_RN_17));
   na02s01 U2271 (.o(n1862),
	.b(wb1_addr_i[21]),
	.a(FE_RN_17));
   na02s01 U2272 (.o(n1885),
	.b(slv0_din[1]),
	.a(FE_OCPN626_wb1_cyc_o));
   na02s02 U2273 (.o(n2018),
	.b(slv0_din[8]),
	.a(FE_OCPN629_wb1_cyc_o));
   na02s02 U2274 (.o(n2132),
	.b(slv0_din[15]),
	.a(FE_OCPN629_wb1_cyc_o));
   na02s01 U2275 (.o(n2397),
	.b(wb1m_data_i[13]),
	.a(n1414));
   na02s01 U2276 (.o(n2427),
	.b(wb1m_data_i[28]),
	.a(n1414));
   oa12s02 U2277 (.o(n617),
	.c(n2211),
	.b(n1521),
	.a(n1670));
   na02f02 U2278 (.o(n2453),
	.b(n2080),
	.a(n2081));
   no02s01 U2279 (.o(u1_N1032),
	.b(dma_req_i[0]),
	.a(n2469));
   oa12s01 U2280 (.o(wb1_addr_o[2]),
	.c(n1641),
	.b(FE_OCPN658_wb1_cyc_o),
	.a(wb1_cyc_o));
   na02s01 U2281 (.o(wb1_addr_o[17]),
	.b(wb1_cyc_o),
	.a(n1665));
   in01s01 U2282 (.o(wb1m_data_o[17]),
	.a(n1705));
   na02s02 U2283 (.o(wb1s_data_o[25]),
	.b(n1814),
	.a(n1815));
   na02s01 U2284 (.o(wb0_addr_o[31]),
	.b(n2367),
	.a(n1414));
   na02s02 U2285 (.o(wb1s_data_o[6]),
	.b(n1757),
	.a(n1758));
   na02s02 U2286 (.o(wb1s_data_o[7]),
	.b(n1760),
	.a(n1761));
   no02m10 U2287 (.o(n1924),
	.b(n1923),
	.a(FE_OCPN481_n2343));
   oa12s02 U2288 (.o(wb0m_data_o[4]),
	.c(n1950),
	.b(FE_OCPN656_wb1_cyc_o),
	.a(n1949));
   na02s02 U2289 (.o(wb1s_data_o[24]),
	.b(n1811),
	.a(n1812));
   na02m01 U2290 (.o(wb1s_data_o[26]),
	.b(n1817),
	.a(n1818));
   na02s02 U2291 (.o(wb1s_data_o[27]),
	.b(n1820),
	.a(n1821));
   na02s10 U2292 (.o(n2215),
	.b(n2225),
	.a(ch0_txsz[20]));
   na02f08 U2294 (.o(n2197),
	.b(ch0_adr0[19]),
	.a(FE_OCPN559_n2357));
   ao12f04 U2296 (.o(n1479),
	.c(n2304),
	.b(ch0_txsz[0]),
	.a(n1480));
   no02m04 U2298 (.o(n2259),
	.b(FE_OCPN566_n2357),
	.a(n2258));
   oa22f08 U2299 (.o(n1428),
	.d(FE_OCPN126_FE_RN_),
	.c(n2278),
	.b(n2282),
	.a(n1425));
   na03s40 U2300 (.o(n1576),
	.c(FE_OCPN512_slv0_adr_3_),
	.b(FE_OCPN669_slv0_adr_4_),
	.a(FE_OCPN139_slv0_adr_2_));
   ao12f02 U2305 (.o(n2260),
	.c(ch0_txsz[23]),
	.b(n2304),
	.a(n2259));
   no02f20 U2306 (.o(n1416),
	.b(n1425),
	.a(n1923));
   na02m40 U2307 (.o(n1923),
	.b(n1901),
	.a(FE_RN_2));
   no02m10 U2308 (.o(n2165),
	.b(n1425),
	.a(n1923));
   na02s04 U2309 (.o(n2119),
	.b(ch0_txsz[15]),
	.a(FE_RN_9));
   na02s04 U2310 (.o(n2155),
	.b(ch0_txsz[17]),
	.a(FE_RN_9));
   na02s02 U2311 (.o(n2266),
	.b(ch0_txsz[24]),
	.a(n1510));
   na02s02 U2312 (.o(n2171),
	.b(ch0_txsz[18]),
	.a(n1510));
   na02s04 U2313 (.o(n2036),
	.b(ch0_txsz[10]),
	.a(FE_RN_9));
   ao22f04 U2315 (.o(n2198),
	.d(n2356),
	.c(ch0_adr1[19]),
	.b(n1494),
	.a(FE_OCPN163_n2346));
   no02f04 U2316 (.o(n2306),
	.b(n2355),
	.a(n2301));
   na02f20 U2317 (.o(n2241),
	.b(n1473),
	.a(n1474));
   na02f06 U2318 (.o(n1418),
	.b(n2241),
	.a(n2197));
   na03f06 U2320 (.o(n1469),
	.c(n1470),
	.b(n1492),
	.a(n2241));
   in01s20 U2321 (.o(n1544),
	.a(slv0_adr[7]));
   in01s40 U2322 (.o(n1545),
	.a(slv0_adr[6]));
   ao12f04 U2323 (.o(n2214),
	.c(n2212),
	.b(n2213),
	.a(FE_OCPN169_n2346));
   na02f04 U2324 (.o(n2203),
	.b(n1419),
	.a(n2198));
   in01f04 U2325 (.o(n1419),
	.a(n1418));
   na02f20 U2328 (.o(n1577),
	.b(n1495),
	.a(n2179));
   ao12f20 U2329 (.o(n2179),
	.c(n1939),
	.b(n1940),
	.a(FE_OCPN106_slv0_adr_2_));
   no02s04 U2330 (.o(n2039),
	.b(n2200),
	.a(n2038));
   oa22m06 U2331 (.o(n2184),
	.d(n2156),
	.c(n2182),
	.b(n2200),
	.a(n2183));
   no02f20 U2334 (.o(n2194),
	.b(n2178),
	.a(n1615));
   oa12s02 U2335 (.o(wb0m_data_o[10]),
	.c(n2049),
	.b(FE_OCPN656_wb1_cyc_o),
	.a(n2048));
   na02s02 U2337 (.o(n2169),
	.b(slv0_din[17]),
	.a(FE_OCPN626_wb1_cyc_o));
   na02s02 U2338 (.o(n1755),
	.b(wb0m_data_i[5]),
	.a(FE_OCPN666_wb1_cyc_o));
   na02s04 U2339 (.o(n1752),
	.b(wb0m_data_i[4]),
	.a(FE_OCPN642_wb1_cyc_o));
   na02s02 U2341 (.o(n1815),
	.b(wb0m_data_i[25]),
	.a(FE_OCPN642_wb1_cyc_o));
   na02s02 U2342 (.o(n1809),
	.b(wb0m_data_i[23]),
	.a(FE_OCPN642_wb1_cyc_o));
   na02s02 U2343 (.o(n1806),
	.b(wb0m_data_i[22]),
	.a(FE_OCPN666_wb1_cyc_o));
   na02s01 U2344 (.o(n1797),
	.b(wb0m_data_i[19]),
	.a(FE_OCPN643_wb1_cyc_o));
   na02s06 U2349 (.o(n2193),
	.b(slv0_dout[19]),
	.a(FE_OCPN368_n2194));
   no02f40 U2350 (.o(n1522),
	.b(n2346),
	.a(FE_OCPN554_n1529));
   na02f80 U2352 (.o(n1424),
	.b(FE_OCPN514_slv0_adr_3_),
	.a(n1613));
   na02f80 U2353 (.o(n1425),
	.b(FE_OCPN610_slv0_adr_3_),
	.a(n1613));
   na02f40 U2354 (.o(n2159),
	.b(slv0_adr[3]),
	.a(n1613));
   no02f80 U2355 (.o(n1613),
	.b(slv0_adr[2]),
	.a(slv0_adr[4]));
   na04f40 U2358 (.o(n2357),
	.d(n1613),
	.c(FE_RN_16),
	.b(n1477),
	.a(FE_RN_4));
   no02m10 U2359 (.o(n2125),
	.b(n2159),
	.a(n2124));
   no02m08 U2360 (.o(n2076),
	.b(n2159),
	.a(n2075));
   no02m10 U2361 (.o(n2143),
	.b(n2159),
	.a(n2142));
   no02m10 U2362 (.o(n1993),
	.b(n2159),
	.a(n1992));
   oa22f08 U2363 (.o(n1919),
	.d(FE_OCPN126_FE_RN_),
	.c(n1917),
	.b(n1918),
	.a(n1424));
   no02f10 U2364 (.o(n2090),
	.b(n1424),
	.a(n2089));
   no02m20 U2365 (.o(n1484),
	.b(n1425),
	.a(FE_OCPN547_n1529));
   oa22m06 U2366 (.o(n512),
	.d(FE_OCPN676_n1580),
	.c(n2134),
	.b(FE_OCPN539_n1595),
	.a(n2138));
   oa22f04 U2367 (.o(n511),
	.d(FE_OCPN676_n1580),
	.c(n2152),
	.b(FE_OCPN539_n1595),
	.a(n1533));
   oa22m04 U2368 (.o(n498),
	.d(FE_OCPN676_n1580),
	.c(n2340),
	.b(FE_OCPN538_n1595),
	.a(n2342));
   oa22m04 U2369 (.o(n523),
	.d(FE_OCPN676_n1580),
	.c(n1955),
	.b(FE_OCPN538_n1595),
	.a(n1956));
   oa22m04 U2370 (.o(n520),
	.d(FE_OCPN676_n1580),
	.c(n2002),
	.b(FE_OCPN539_n1595),
	.a(n2005));
   oa22s04 U2371 (.o(n519),
	.d(FE_OCPN675_n1580),
	.c(n2021),
	.b(FE_OCPN538_n1595),
	.a(n2023));
   oa22f04 U2373 (.o(n517),
	.d(FE_OCPN676_n1580),
	.c(n2050),
	.b(FE_OCPN540_n1595),
	.a(n2054));
   oa22f04 U2374 (.o(n516),
	.d(FE_OCPN676_n1580),
	.c(n2073),
	.b(FE_OCPN540_n1595),
	.a(n2074));
   oa22m04 U2375 (.o(n515),
	.d(FE_OCPN676_n1580),
	.c(n2087),
	.b(n2088),
	.a(FE_OCPN540_n1595));
   oa22m04 U2376 (.o(n514),
	.d(FE_OCPN676_n1580),
	.c(n2103),
	.b(FE_OCPN540_n1595),
	.a(n2104));
   oa22s02 U2377 (.o(n513),
	.d(FE_OCPN675_n1580),
	.c(n2116),
	.b(FE_OCPN539_n1595),
	.a(n2120));
   oa22m04 U2378 (.o(n510),
	.d(FE_OCPN676_n1580),
	.c(n2174),
	.b(FE_OCPN538_n1595),
	.a(n2175));
   oa22m04 U2380 (.o(n508),
	.d(FE_OCPN676_n1580),
	.c(n2210),
	.b(FE_OCPN538_n1595),
	.a(n2211));
   oa22f04 U2381 (.o(n507),
	.d(FE_OCPN676_n1580),
	.c(n2221),
	.b(FE_OCPN538_n1595),
	.a(n2222));
   oa22m04 U2382 (.o(n506),
	.d(FE_OCPN676_n1580),
	.c(n2234),
	.b(FE_OCPN538_n1595),
	.a(n2237));
   oa22m04 U2383 (.o(n505),
	.d(FE_OCPN676_n1580),
	.c(n2249),
	.b(FE_OCPN538_n1595),
	.a(n2252));
   oa22f04 U2384 (.o(n504),
	.d(FE_OCPN676_n1580),
	.c(n2264),
	.b(FE_OCPN538_n1595),
	.a(n2267));
   oa22s04 U2385 (.o(n502),
	.d(FE_OCPN676_n1580),
	.c(n2292),
	.b(FE_OCPN538_n1595),
	.a(n2295));
   oa22f04 U2386 (.o(n501),
	.d(FE_OCPN676_n1580),
	.c(n2310),
	.b(FE_OCPN538_n1595),
	.a(n2312));
   oa22s04 U2387 (.o(n500),
	.d(FE_OCPN676_n1580),
	.c(n2320),
	.b(FE_OCPN538_n1595),
	.a(n2322));
   oa22m04 U2388 (.o(n499),
	.d(FE_OCPN676_n1580),
	.c(n2330),
	.b(FE_OCPN538_n1595),
	.a(n2332));
   oa22f04 U2389 (.o(n503),
	.d(FE_OCPN676_n1580),
	.c(n2278),
	.b(FE_OCPN538_n1595),
	.a(n2281));
   no02m10 U2390 (.o(n1426),
	.b(n1626),
	.a(n2346));
   na02m40 U2391 (.o(n1900),
	.b(FE_RN_16),
	.a(slv0_adr[5]));
   in01s01 U2393 (.o(n2243),
	.a(ch0_adr0[22]));
   na02f20 U2396 (.o(n1476),
	.b(slv0_adr[5]),
	.a(FE_RN_4));
   in01s02 U2401 (.o(n1438),
	.a(FE_RN_17));
   in01s02 U2404 (.o(n2089),
	.a(u0_int_maskb_13_));
   no02s03 U2405 (.o(n1624),
	.b(ch0_csr[7]),
	.a(n1623));
   in01m01 U2406 (.o(n1961),
	.a(ch0_adr1[5]));
   in01s01 U2407 (.o(n1995),
	.a(ch0_adr1[7]));
   in01m01 U2408 (.o(n2013),
	.a(ch0_adr1[8]));
   in01s02 U2409 (.o(n2027),
	.a(ch0_adr1[9]));
   in01m01 U2410 (.o(n2043),
	.a(ch0_adr1[10]));
   in01s01 U2411 (.o(n2063),
	.a(ch0_adr1[11]));
   in01s01 U2412 (.o(n2092),
	.a(ch0_adr1[13]));
   in01s01 U2413 (.o(n2108),
	.a(ch0_adr1[14]));
   in01s02 U2414 (.o(n2127),
	.a(ch0_adr1[15]));
   in01s02 U2415 (.o(n2145),
	.a(ch0_adr1[16]));
   in01s02 U2416 (.o(n2163),
	.a(ch0_adr1[17]));
   in01s03 U2417 (.o(n2175),
	.a(slv0_dout[18]));
   in01s01 U2418 (.o(n1957),
	.a(ch0_csr[5]));
   in01s01 U2419 (.o(n2008),
	.a(ch0_csr[8]));
   in01s01 U2420 (.o(n1607),
	.a(wb0_ack_i));
   na02s02 U2421 (.o(n1722),
	.b(wb1_stb_i),
	.a(wb1_cyc_i));
   in01s01 U2422 (.o(n2350),
	.a(ch0_adr0[30]));
   in01s01 U2423 (.o(n2336),
	.a(ch0_adr0[29]));
   in01s01 U2424 (.o(n2316),
	.a(ch0_adr0[27]));
   na02s04 U2425 (.o(n2213),
	.b(u0_int_maskb_20_),
	.a(n1566));
   na02s08 U2426 (.o(n2212),
	.b(u0_int_maska_20_),
	.a(FE_OCPN124_FE_RN_));
   na02m04 U2427 (.o(n2180),
	.b(ch0_adr0[18]),
	.a(FE_OCPN560_n2357));
   in01s01 U2428 (.o(n2183),
	.a(ch0_txsz[18]));
   na02m20 U2429 (.o(n2200),
	.b(n2343),
	.a(n2007));
   in01s02 U2430 (.o(n2078),
	.a(ch0_adr1[12]));
   ao22f08 U2431 (.o(n1977),
	.d(n2343),
	.c(u0_int_maska_6_),
	.b(n1566),
	.a(u0_int_maskb_6_));
   no02m08 U2432 (.o(n1944),
	.b(FE_OCPN670_n2356),
	.a(n1943));
   na02s08 U2433 (.o(n1942),
	.b(u0_int_maskb_4_),
	.a(n1566));
   na02m08 U2434 (.o(n1941),
	.b(u0_int_maska_4_),
	.a(FE_OCPN124_FE_RN_));
   in01s04 U2435 (.o(n1926),
	.a(n1925));
   in01f10 U2436 (.o(n1477),
	.a(n1478));
   no02s02 U2437 (.o(n1609),
	.b(u3_u1_rf_ack),
	.a(n1608));
   oa12s02 U2438 (.o(n641),
	.c(n1883),
	.b(n1513),
	.a(n1881));
   in01s01 U2439 (.o(n2025),
	.a(ch0_adr0[9]));
   in01s01 U2440 (.o(n2101),
	.a(ch0_adr0[14]));
   oa12s02 U2441 (.o(n745),
	.c(n2120),
	.b(n1513),
	.a(n2119));
   oa12s02 U2442 (.o(n748),
	.c(n2267),
	.b(n1513),
	.a(n2266));
   oa12f02 U2443 (.o(n756),
	.c(n2138),
	.b(n1513),
	.a(n2137));
   in01s20 U2444 (.o(n1531),
	.a(n1890));
   na02f40 U2445 (.o(n1939),
	.b(FE_OCPN669_slv0_adr_4_),
	.a(FE_OCPN611_slv0_adr_3_));
   na02s20 U2446 (.o(n1733),
	.b(wb0_addr_i[28]),
	.a(wb0_cyc_i));
   na02s40 U2447 (.o(n1734),
	.b(wb0_addr_i[29]),
	.a(wb0_cyc_i));
   na02s10 U2448 (.o(n1736),
	.b(wb0_addr_i[30]),
	.a(wb0_cyc_i));
   na02s20 U2449 (.o(n1735),
	.b(wb0_cyc_i),
	.a(wb0_addr_i[31]));
   na02s10 U2450 (.o(n2365),
	.b(wb1_cyc_i),
	.a(wb1_addr_i[28]));
   na02s20 U2451 (.o(n2366),
	.b(wb1_addr_i[29]),
	.a(wb1_cyc_i));
   na02s20 U2452 (.o(n2368),
	.b(wb1_addr_i[30]),
	.a(wb1_cyc_i));
   na02s20 U2453 (.o(n2367),
	.b(wb1_addr_i[31]),
	.a(wb1_cyc_i));
   in01s02 U2457 (.o(n1992),
	.a(u0_int_maskb_7_));
   in01s02 U2458 (.o(n2010),
	.a(u0_int_maskb_8_));
   in01s02 U2459 (.o(n2040),
	.a(u0_int_maskb_10_));
   in01s01 U2460 (.o(n2060),
	.a(u0_int_maskb_11_));
   in01s02 U2461 (.o(n2075),
	.a(u0_int_maskb_12_));
   in01s02 U2462 (.o(n2124),
	.a(u0_int_maskb_15_));
   in01s02 U2463 (.o(n2142),
	.a(u0_int_maskb_16_));
   in01s02 U2464 (.o(n2160),
	.a(u0_int_maskb_17_));
   no02f20 U2467 (.o(n1523),
	.b(slv0_adr[4]),
	.a(n1529));
   no04f80 U2468 (.o(n1537),
	.d(FE_OCPN513_slv0_adr_3_),
	.c(FE_OCPN139_slv0_adr_2_),
	.b(n1529),
	.a(FE_OCPN617_slv0_adr_5_));
   in01s02 U2470 (.o(n2192),
	.a(slv0_dout[19]));
   in01s01 U2471 (.o(n2258),
	.a(ch0_adr0[23]));
   in01s02 U2473 (.o(n1533),
	.a(slv0_dout[17]));
   in01s02 U2474 (.o(n2138),
	.a(slv0_dout[16]));
   in01s04 U2478 (.o(n1480),
	.a(n1558));
   na02s06 U2479 (.o(n1555),
	.b(n1877),
	.a(n1878));
   na02s08 U2480 (.o(n1877),
	.b(slv0_adr[4]),
	.a(n1874));
   no02s06 U2481 (.o(n1556),
	.b(n1875),
	.a(FE_RN_7));
   ao12f06 U2482 (.o(n2255),
	.c(FE_OCPN124_FE_RN_),
	.b(u0_int_maska_23_),
	.a(n2254));
   na02m06 U2483 (.o(n2226),
	.b(u0_int_maska_21_),
	.a(FE_OCPN124_FE_RN_));
   na02s06 U2484 (.o(n2227),
	.b(u0_int_maskb_21_),
	.a(n1566));
   no02f10 U2485 (.o(n2224),
	.b(n2156),
	.a(n2223));
   in01s01 U2486 (.o(n2094),
	.a(ch0_csr[13]));
   in01s01 U2488 (.o(n1918),
	.a(u0_int_maskb_3_));
   in01s01 U2489 (.o(n1917),
	.a(u0_int_maska_3_));
   no02s04 U2491 (.o(n1633),
	.b(wb0_sel_i[1]),
	.a(FE_OCPN658_wb1_cyc_o));
   na02s01 U2492 (.o(wb1_addr_o[14]),
	.b(wb1_cyc_o),
	.a(n1661));
   na02s02 U2493 (.o(wb1_addr_o[15]),
	.b(wb1_cyc_o),
	.a(n1662));
   na02s02 U2494 (.o(n1683),
	.b(wb0_addr_i[27]),
	.a(FE_OCPN651_wb1_cyc_o));
   na02s01 U2495 (.o(n1699),
	.b(wb0s_data_i[11]),
	.a(FE_RN_17));
   na02s01 U2496 (.o(n1703),
	.b(wb0s_data_i[15]),
	.a(n1414));
   na02s01 U2497 (.o(n1714),
	.b(wb0s_data_i[26]),
	.a(FE_RN_17));
   na02s01 U2498 (.o(n1717),
	.b(wb0s_data_i[29]),
	.a(n1414));
   na02s06 U2500 (.o(n1751),
	.b(de_csr[4]),
	.a(FE_RN_12));
   na02s02 U2501 (.o(n1754),
	.b(de_csr[5]),
	.a(FE_RN_12));
   na02s02 U2502 (.o(n1758),
	.b(wb0m_data_i[6]),
	.a(FE_OCPN642_wb1_cyc_o));
   na02s02 U2503 (.o(n1761),
	.b(wb0m_data_i[7]),
	.a(FE_OCPN642_wb1_cyc_o));
   na02s02 U2504 (.o(n1764),
	.b(wb0m_data_i[8]),
	.a(FE_OCPN651_wb1_cyc_o));
   na02s02 U2505 (.o(n1766),
	.b(de_csr[9]),
	.a(FE_RN_12));
   na02s02 U2506 (.o(n1769),
	.b(de_csr[10]),
	.a(FE_RN_1));
   na02s02 U2507 (.o(n1770),
	.b(wb0m_data_i[10]),
	.a(FE_OCPN666_wb1_cyc_o));
   na02s02 U2508 (.o(n1772),
	.b(de_csr[11]),
	.a(FE_RN_1));
   na02s02 U2509 (.o(n1773),
	.b(wb0m_data_i[11]),
	.a(FE_OCPN643_wb1_cyc_o));
   na02s02 U2510 (.o(n1775),
	.b(de_csr[12]),
	.a(FE_RN_1));
   na02s02 U2511 (.o(n1776),
	.b(wb0m_data_i[12]),
	.a(FE_OCPN666_wb1_cyc_o));
   na02s02 U2512 (.o(n1778),
	.b(de_csr[13]),
	.a(FE_RN_1));
   na02s02 U2513 (.o(n1779),
	.b(wb0m_data_i[13]),
	.a(FE_OCPN666_wb1_cyc_o));
   na02s02 U2514 (.o(n1781),
	.b(de_csr[14]),
	.a(FE_RN_1));
   na02s01 U2515 (.o(n1782),
	.b(wb0m_data_i[14]),
	.a(FE_OCPN643_wb1_cyc_o));
   na02s02 U2516 (.o(n1784),
	.b(de_csr[15]),
	.a(FE_RN_11));
   na02s02 U2517 (.o(n1787),
	.b(de_csr[16]),
	.a(FE_RN_11));
   na02s02 U2518 (.o(n1788),
	.b(wb0m_data_i[16]),
	.a(FE_OCPN651_wb1_cyc_o));
   na02s02 U2519 (.o(n1791),
	.b(wb0m_data_i[17]),
	.a(FE_OCPN651_wb1_cyc_o));
   na02m01 U2520 (.o(wb1s_data_o[19]),
	.b(n1796),
	.a(n1797));
   na02s01 U2521 (.o(n1796),
	.b(de_csr[19]),
	.a(FE_RN_1));
   na02s02 U2522 (.o(n1799),
	.b(de_csr[20]),
	.a(n1832));
   na02s02 U2523 (.o(n1800),
	.b(wb0m_data_i[20]),
	.a(FE_OCPN666_wb1_cyc_o));
   na02s02 U2524 (.o(n1802),
	.b(de_csr[21]),
	.a(n1832));
   na02s02 U2525 (.o(n1803),
	.b(wb0m_data_i[21]),
	.a(FE_OCPN642_wb1_cyc_o));
   na02s02 U2526 (.o(wb1s_data_o[22]),
	.b(n1805),
	.a(n1806));
   na02s02 U2527 (.o(n1805),
	.b(de_csr[22]),
	.a(n1832));
   na02s02 U2528 (.o(wb1s_data_o[23]),
	.b(n1808),
	.a(n1809));
   na02s02 U2529 (.o(n1808),
	.b(de_csr[23]),
	.a(FE_RN_12));
   na02s02 U2530 (.o(n1814),
	.b(de_csr[25]),
	.a(n1832));
   no02s01 U2531 (.o(n1837),
	.b(wb1_sel_i[0]),
	.a(n1438));
   no02s01 U2532 (.o(n1838),
	.b(wb1_sel_i[1]),
	.a(n1438));
   no02s01 U2533 (.o(n1840),
	.b(wb1_sel_i[3]),
	.a(n1438));
   na02s01 U2534 (.o(n1844),
	.b(wb1_addr_i[3]),
	.a(FE_RN_17));
   na02s02 U2535 (.o(n1849),
	.b(wb1_addr_i[8]),
	.a(FE_OCPN284_wb0_cyc_o));
   na02s02 U2536 (.o(n1851),
	.b(wb1_addr_i[10]),
	.a(FE_OCPN284_wb0_cyc_o));
   na02s01 U2537 (.o(n1852),
	.b(wb1_addr_i[11]),
	.a(FE_RN_17));
   na02s02 U2538 (.o(n1854),
	.b(wb1_addr_i[13]),
	.a(FE_OCPN284_wb0_cyc_o));
   na02s02 U2539 (.o(n1859),
	.b(wb1_addr_i[18]),
	.a(FE_OCPN284_wb0_cyc_o));
   na02s01 U2540 (.o(n1865),
	.b(wb1_addr_i[24]),
	.a(FE_RN_17));
   na02s02 U2541 (.o(n1866),
	.b(wb1_addr_i[25]),
	.a(FE_OCPN284_wb0_cyc_o));
   na02s02 U2542 (.o(n1868),
	.b(wb1_addr_i[27]),
	.a(wb0_cyc_o));
   oa12s01 U2543 (.o(wb0m_data_o[1]),
	.c(n1886),
	.b(FE_OCPN656_wb1_cyc_o),
	.a(n1885));
   oa12s02 U2544 (.o(wb0m_data_o[2]),
	.c(n1909),
	.b(FE_OCPN656_wb1_cyc_o),
	.a(n1908));
   na02s03 U2545 (.o(n1908),
	.b(slv0_din[2]),
	.a(FE_OCPN626_wb1_cyc_o));
   na02s02 U2546 (.o(n1949),
	.b(slv0_din[4]),
	.a(FE_OCPN629_wb1_cyc_o));
   oa12s02 U2547 (.o(wb0m_data_o[5]),
	.c(n1968),
	.b(FE_OCPN633_wb1_cyc_o),
	.a(n1967));
   na02s03 U2548 (.o(n1967),
	.b(slv0_din[5]),
	.a(FE_OCPN627_wb1_cyc_o));
   na02s02 U2550 (.o(n2000),
	.b(slv0_din[7]),
	.a(FE_OCPN626_wb1_cyc_o));
   oa12s02 U2551 (.o(wb0m_data_o[8]),
	.c(n2019),
	.b(FE_OCPN658_wb1_cyc_o),
	.a(n2018));
   oa12s02 U2552 (.o(wb0m_data_o[9]),
	.c(n2033),
	.b(FE_OCPN633_wb1_cyc_o),
	.a(n2032));
   na02s02 U2553 (.o(n2032),
	.b(slv0_din[9]),
	.a(FE_OCPN627_wb1_cyc_o));
   oa12s02 U2554 (.o(wb0m_data_o[12]),
	.c(n2083),
	.b(FE_OCPN658_wb1_cyc_o),
	.a(n2082));
   na02s01 U2555 (.o(n2082),
	.b(slv0_din[12]),
	.a(FE_OCPN626_wb1_cyc_o));
   oa12s02 U2556 (.o(wb0m_data_o[13]),
	.c(n2099),
	.b(FE_OCPN656_wb1_cyc_o),
	.a(n2098));
   na02s01 U2557 (.o(n2098),
	.b(slv0_din[13]),
	.a(FE_OCPN626_wb1_cyc_o));
   oa12s01 U2558 (.o(wb0m_data_o[14]),
	.c(n2115),
	.b(FE_OCPN658_wb1_cyc_o),
	.a(n2114));
   oa12s02 U2559 (.o(wb0m_data_o[16]),
	.c(n2151),
	.b(FE_OCPN667_wb1_cyc_o),
	.a(n2150));
   na02s01 U2560 (.o(n2150),
	.b(slv0_din[16]),
	.a(FE_OCPN629_wb1_cyc_o));
   oa12s01 U2561 (.o(wb0m_data_o[20]),
	.c(n2217),
	.b(FE_OCPN658_wb1_cyc_o),
	.a(n2216));
   na02s01 U2562 (.o(n2216),
	.b(slv0_din[20]),
	.a(FE_OCPN626_wb1_cyc_o));
   oa12s02 U2563 (.o(wb0m_data_o[23]),
	.c(n2263),
	.b(FE_OCPN656_wb1_cyc_o),
	.a(n2262));
   na02s01 U2564 (.o(n2262),
	.b(slv0_din[23]),
	.a(FE_OCPN624_wb1_cyc_o));
   oa12s02 U2565 (.o(wb0m_data_o[27]),
	.c(n2318),
	.b(FE_OCPN667_wb1_cyc_o),
	.a(n2317));
   na02s01 U2566 (.o(n2317),
	.b(slv0_din[27]),
	.a(FE_OCPN630_wb1_cyc_o));
   na02s02 U2567 (.o(n2361),
	.b(wb1_rty_i),
	.a(wb1_cyc_o));
   na02s02 U2568 (.o(n2362),
	.b(wb1_err_i),
	.a(wb1_cyc_o));
   na02s01 U2569 (.o(n2375),
	.b(wb1m_data_i[2]),
	.a(FE_RN_17));
   na02s01 U2570 (.o(n2411),
	.b(wb1m_data_i[20]),
	.a(FE_OCPN277_wb0_cyc_o));
   na02s01 U2571 (.o(n2413),
	.b(wb1m_data_i[21]),
	.a(FE_OCPN277_wb0_cyc_o));
   na02s01 U2572 (.o(n2417),
	.b(wb1m_data_i[23]),
	.a(FE_OCPN277_wb0_cyc_o));
   na02s01 U2573 (.o(n2419),
	.b(wb1m_data_i[24]),
	.a(FE_RN_17));
   na02s01 U2574 (.o(n2421),
	.b(wb1m_data_i[25]),
	.a(FE_OCPN277_wb0_cyc_o));
   na02s01 U2575 (.o(n2429),
	.b(wb1m_data_i[29]),
	.a(FE_OCPN277_wb0_cyc_o));
   na02s01 U2576 (.o(n2431),
	.b(wb1m_data_i[30]),
	.a(FE_OCPN277_wb0_cyc_o));
   na02s01 U2577 (.o(n2433),
	.b(wb1m_data_i[31]),
	.a(FE_OCPN277_wb0_cyc_o));
   oa12s02 U2578 (.o(n525),
	.c(n1914),
	.b(FE_OCPN539_n1595),
	.a(n1911));
   oa22s02 U2580 (.o(n534),
	.d(FE_OCPN383_n1512),
	.c(n1954),
	.b(n1591),
	.a(n1956));
   oa22s02 U2581 (.o(n535),
	.d(FE_OCPN383_n1512),
	.c(n1969),
	.b(n1591),
	.a(n1974));
   oa22s04 U2582 (.o(n537),
	.d(FE_RN_13),
	.c(n2010),
	.b(n1591),
	.a(n2005));
   in01s01 U2584 (.o(n2020),
	.a(u0_int_maskb_9_));
   oa22m02 U2585 (.o(n539),
	.d(FE_RN_13),
	.c(n2040),
	.b(n1591),
	.a(n2037));
   oa22m02 U2586 (.o(n540),
	.d(FE_RN_13),
	.c(n2060),
	.b(n1591),
	.a(n2054));
   oa22m02 U2587 (.o(n541),
	.d(FE_RN_13),
	.c(n2075),
	.b(n1591),
	.a(n2074));
   oa22m02 U2588 (.o(n542),
	.d(FE_RN_13),
	.c(n2089),
	.b(n1591),
	.a(n2088));
   oa22m02 U2589 (.o(n543),
	.d(FE_RN_13),
	.c(n2105),
	.b(n1591),
	.a(n2104));
   oa22s02 U2590 (.o(n544),
	.d(FE_RN_13),
	.c(n2124),
	.b(n1591),
	.a(n2120));
   oa22m02 U2591 (.o(n545),
	.d(FE_RN_13),
	.c(n2142),
	.b(n1591),
	.a(n2138));
   oa22m02 U2592 (.o(n546),
	.d(FE_RN_13),
	.c(n2160),
	.b(n1591),
	.a(n1533));
   oa22m04 U2593 (.o(n547),
	.d(FE_OCPN383_n1512),
	.c(n2173),
	.b(n1579),
	.a(n2175));
   in01s01 U2594 (.o(n2173),
	.a(u0_int_maskb_18_));
   oa22m04 U2595 (.o(n548),
	.d(FE_OCPN383_n1512),
	.c(n2190),
	.b(n1579),
	.a(n2192));
   oa22m02 U2596 (.o(n549),
	.d(FE_OCPN383_n1512),
	.c(n2209),
	.b(n1579),
	.a(n2211));
   in01s01 U2597 (.o(n2209),
	.a(u0_int_maskb_20_));
   oa22m04 U2598 (.o(n550),
	.d(FE_OCPN383_n1512),
	.c(n2220),
	.b(n1579),
	.a(n2222));
   in01s01 U2599 (.o(n2220),
	.a(u0_int_maskb_21_));
   oa22m02 U2601 (.o(n552),
	.d(FE_OCPN383_n1512),
	.c(n2253),
	.b(n1591),
	.a(n2252));
   oa22m02 U2602 (.o(n553),
	.d(FE_OCPN383_n1512),
	.c(n2268),
	.b(n1579),
	.a(n2267));
   oa22s02 U2603 (.o(n554),
	.d(FE_OCPN383_n1512),
	.c(n2282),
	.b(n1591),
	.a(n2281));
   oa22s02 U2604 (.o(n555),
	.d(FE_OCPN383_n1512),
	.c(n2296),
	.b(n1591),
	.a(n2295));
   oa22m04 U2605 (.o(n556),
	.d(FE_OCPN383_n1512),
	.c(n2309),
	.b(n1579),
	.a(n2312));
   oa22s02 U2606 (.o(n557),
	.d(FE_OCPN383_n1512),
	.c(n2319),
	.b(FE_RN_18),
	.a(n2322));
   oa22m02 U2607 (.o(n558),
	.d(FE_OCPN383_n1512),
	.c(n2329),
	.b(FE_RN_18),
	.a(n2332));
   oa22m02 U2608 (.o(n559),
	.d(FE_OCPN383_n1512),
	.c(n2339),
	.b(n1591),
	.a(n2342));
   oa12f02 U2609 (.o(n570),
	.c(FE_OCPN367_n2194),
	.b(n1638),
	.a(n2055));
   in01s04 U2610 (.o(n2055),
	.a(n1524));
   no02s02 U2611 (.o(n571),
	.b(n1524),
	.a(n1526));
   no02s04 U2612 (.o(n1526),
	.b(FE_OCPN367_n2194),
	.a(n1527));
   oa12f04 U2613 (.o(n613),
	.c(n2175),
	.b(FE_OCPN462_n1521),
	.a(n1666));
   na02m08 U2614 (.o(n1672),
	.b(ch0_adr1[21]),
	.a(FE_OCPN462_n1521));
   na02f06 U2615 (.o(n1685),
	.b(FE_OCPN178_n1521),
	.a(slv0_dout[29]));
   oa12m02 U2616 (.o(n639),
	.c(FE_OCPN179_n1521),
	.b(n1687),
	.a(n1686));
   in01s01 U2617 (.o(n2085),
	.a(ch0_adr0[13]));
   na02s04 U2618 (.o(n2084),
	.b(slv0_dout[13]),
	.a(n1573));
   oa12s02 U2619 (.o(n733),
	.c(FE_OCPN367_n2194),
	.b(n2369),
	.a(n1731));
   na02s01 U2620 (.o(n1731),
	.b(slv0_dout[2]),
	.a(n2194));
   oa12f02 U2621 (.o(n753),
	.c(FE_OCPN619_n1513),
	.b(n2201),
	.a(n1564));
   na02m04 U2622 (.o(n1564),
	.b(FE_OCPN619_n1513),
	.a(slv0_dout[19]));
   oa12m02 U2623 (.o(n754),
	.c(n2175),
	.b(n1513),
	.a(n2171));
   oa12f02 U2624 (.o(n759),
	.c(FE_OCPN370_n2194),
	.b(n1990),
	.a(n1618));
   na02m06 U2625 (.o(n1618),
	.b(FE_OCPN370_n2194),
	.a(slv0_dout[7]));
   oa12m04 U2626 (.o(n761),
	.c(FE_OCPN370_n2194),
	.b(n2094),
	.a(n2086));
   na02s08 U2627 (.o(n2086),
	.b(FE_OCPN370_n2194),
	.a(slv0_dout[13]));
   oa12f02 U2628 (.o(n763),
	.c(FE_OCPN370_n2194),
	.b(n2122),
	.a(n2121));
   na02f06 U2629 (.o(n2121),
	.b(slv0_dout[15]),
	.a(FE_OCPN370_n2194));
   oa12f02 U2630 (.o(n764),
	.c(FE_OCPN370_n2194),
	.b(n2140),
	.a(n2139));
   na02f06 U2631 (.o(n2139),
	.b(slv0_dout[16]),
	.a(FE_OCPN370_n2194));
   oa12f02 U2632 (.o(n765),
	.c(FE_OCPN370_n2194),
	.b(n2157),
	.a(n1625));
   na02s08 U2633 (.o(n1625),
	.b(slv0_dout[17]),
	.a(FE_OCPN370_n2194));
   no02f02 U2634 (.o(n1503),
	.b(FE_OCPN565_n2357),
	.a(n2350));
   no02s04 U2635 (.o(n1500),
	.b(FE_OCPN566_n2357),
	.a(n2336));
   no02f08 U2636 (.o(n1505),
	.b(n2355),
	.a(n1506));
   no02s06 U2637 (.o(n1506),
	.b(FE_OCPN565_n2357),
	.a(n2316));
   ao12m04 U2638 (.o(n2305),
	.c(ch0_txsz[26]),
	.b(n2304),
	.a(n2303));
   ao12f04 U2639 (.o(n2288),
	.c(ch0_txsz[25]),
	.b(n2304),
	.a(n2287));
   oa22f06 U2640 (.o(n2285),
	.d(FE_OCPN663_n1428),
	.c(FE_OCPN169_n2346),
	.b(n2284),
	.a(FE_OCPN670_n2356));
   ao12f04 U2641 (.o(n2274),
	.c(ch0_txsz[24]),
	.b(n2304),
	.a(n2273));
   in01m02 U2644 (.o(n1560),
	.a(n2214));
   na02s04 U2646 (.o(n2166),
	.b(ch0_adr0[17]),
	.a(n2165));
   no02f08 U2647 (.o(n2148),
	.b(FE_OCPN673_n1577),
	.a(n2146));
   na02m06 U2648 (.o(n2147),
	.b(ch0_adr0[16]),
	.a(n2165));
   no02f06 U2649 (.o(n2130),
	.b(FE_OCPN673_n1577),
	.a(n2128));
   na02s08 U2650 (.o(n2129),
	.b(ch0_adr0[15]),
	.a(n2165));
   no02f08 U2651 (.o(n2111),
	.b(n2156),
	.a(n2110));
   no02f08 U2652 (.o(n1981),
	.b(FE_OCPN673_n1577),
	.a(n1979));
   ao12s01 U2654 (.o(u3_u1_N5),
	.c(FE_OCPN554_n1529),
	.b(n1622),
	.a(n1610));
   no04s02 U2655 (.o(u3_u1_N3),
	.d(slv0_re),
	.c(n1612),
	.b(wb0_we_i),
	.a(n1610));
   na02f80 U2659 (.o(n2346),
	.b(n1871),
	.a(FE_RN_4));
   oa12f02 U2661 (.o(n531),
	.c(FE_OCPN385_n1579),
	.b(n1895),
	.a(n1887));
   na02s01 U2665 (.o(wb1_addr_o[22]),
	.b(wb1_cyc_o),
	.a(n1674));
   in01s01 U2670 (.o(n1610),
	.a(n1609));
   oa12s01 U2671 (.o(wb0_ack_o),
	.c(n1605),
	.b(FE_OCPN658_wb1_cyc_o),
	.a(n2363));
   in01s01 U2672 (.o(wb1_stb_o),
	.a(n1630));
   in01s01 U2673 (.o(wb1_we_o),
	.a(n1631));
   in01s01 U2674 (.o(wb1_addr_o[0]),
	.a(n1636));
   in01s01 U2675 (.o(wb1_addr_o[1]),
	.a(n1637));
   oa22m08 U2676 (.o(n2202),
	.d(n2156),
	.c(n2199),
	.b(n2200),
	.a(n2201));
   oa12s02 U2680 (.o(wb0m_data_o[17]),
	.c(n2170),
	.b(FE_OCPN656_wb1_cyc_o),
	.a(n2169));
   oa12s02 U2681 (.o(wb1_addr_o[3]),
	.c(n1643),
	.b(FE_OCPN658_wb1_cyc_o),
	.a(wb1_cyc_o));
   in01s01 U2682 (.o(wb0_sel_o[0]),
	.a(n1837));
   in01s01 U2684 (.o(wb1_sel_o[2]),
	.a(n1634));
   in01s01 U2685 (.o(wb1_sel_o[3]),
	.a(n1635));
   oa12s02 U2686 (.o(wb0m_data_o[15]),
	.c(n2133),
	.b(FE_OCPN658_wb1_cyc_o),
	.a(n2132));
   na02s02 U2687 (.o(wb1s_data_o[15]),
	.b(n1784),
	.a(n1785));
   na02s02 U2688 (.o(wb1s_data_o[12]),
	.b(n1775),
	.a(n1776));
   na02s01 U2689 (.o(wb1s_data_o[14]),
	.b(n1781),
	.a(n1782));
   na02s02 U2690 (.o(wb1s_data_o[13]),
	.b(n1778),
	.a(n1779));
   in01s01 U2691 (.o(wb1m_data_o[9]),
	.a(n1697));
   in01s01 U2692 (.o(wb1m_data_o[27]),
	.a(n1715));
   in01s01 U2693 (.o(wb1m_data_o[30]),
	.a(n1718));
   in01s01 U2694 (.o(wb1m_data_o[5]),
	.a(n1693));
   in01s01 U2695 (.o(wb1m_data_o[31]),
	.a(n1719));
   na02s01 U2698 (.o(n2391),
	.b(wb1m_data_i[10]),
	.a(n1414));
   na02s01 U2699 (.o(n2482),
	.b(wb0s_data_i[19]),
	.a(wb0_ack_i));
   na02s01 U2700 (.o(n2483),
	.b(wb0s_data_i[18]),
	.a(FE_OFN427_wb0_ack_i));
   na02s01 U2701 (.o(n2484),
	.b(wb0s_data_i[17]),
	.a(wb0_ack_i));
   na02s01 U2702 (.o(n2485),
	.b(wb0s_data_i[16]),
	.a(wb0_ack_i));
   na02s01 U2703 (.o(n2486),
	.b(wb0s_data_i[15]),
	.a(wb0_ack_i));
   na02s01 U2704 (.o(n2487),
	.b(wb0s_data_i[14]),
	.a(wb0_ack_i));
   na02s01 U2705 (.o(n2488),
	.b(wb0s_data_i[13]),
	.a(wb0_ack_i));
   na02s01 U2706 (.o(n2489),
	.b(wb0s_data_i[12]),
	.a(wb0_ack_i));
   na02s01 U2707 (.o(n2490),
	.b(wb0s_data_i[11]),
	.a(wb0_ack_i));
   na02s01 U2708 (.o(n2491),
	.b(wb0s_data_i[10]),
	.a(wb0_ack_i));
   na02s01 U2709 (.o(n2492),
	.b(wb0s_data_i[9]),
	.a(FE_OFN427_wb0_ack_i));
   na02s01 U2710 (.o(n2493),
	.b(wb0s_data_i[8]),
	.a(wb0_ack_i));
   na02s01 U2711 (.o(n2494),
	.b(wb0s_data_i[7]),
	.a(wb0_ack_i));
   na02s01 U2712 (.o(n2495),
	.b(wb0s_data_i[6]),
	.a(wb0_ack_i));
   na02s01 U2713 (.o(n2496),
	.b(wb0s_data_i[5]),
	.a(FE_OFN427_wb0_ack_i));
   na02s01 U2714 (.o(n2497),
	.b(wb0s_data_i[4]),
	.a(wb0_ack_i));
   na02s01 U2715 (.o(n2498),
	.b(wb0s_data_i[3]),
	.a(wb0_ack_i));
   na02s01 U2716 (.o(n2499),
	.b(wb0s_data_i[2]),
	.a(wb0_ack_i));
   na02s01 U2717 (.o(n2500),
	.b(wb0s_data_i[1]),
	.a(wb0_ack_i));
   na02s01 U2718 (.o(n2501),
	.b(wb0s_data_i[0]),
	.a(wb0_ack_i));
   oa12m01 U2719 (.o(wb0m_data_o[30]),
	.c(n2352),
	.b(FE_OCPN667_wb1_cyc_o),
	.a(n2351));
   oa12s02 U2720 (.o(wb0m_data_o[3]),
	.c(n1930),
	.b(FE_OCPN656_wb1_cyc_o),
	.a(n1929));
   oa12s04 U2721 (.o(wb0m_data_o[11]),
	.c(n2069),
	.b(FE_OCPN668_wb1_cyc_o),
	.a(n2068));
   na02s02 U2722 (.o(wb1s_data_o[29]),
	.b(n1826),
	.a(n1827));
   na02s02 U2723 (.o(wb1s_data_o[30]),
	.b(n1829),
	.a(n1830));
   na02s02 U2724 (.o(wb1s_data_o[31]),
	.b(n1833),
	.a(n1834));
   na02s02 U2725 (.o(wb1s_data_o[28]),
	.b(n1823),
	.a(n1824));
   na02s01 U2726 (.o(wb1s_data_o[8]),
	.b(n1763),
	.a(n1764));
   na02s02 U2727 (.o(wb1s_data_o[9]),
	.b(n1766),
	.a(n1767));
   na02s02 U2728 (.o(wb1s_data_o[10]),
	.b(n1769),
	.a(n1770));
   na02s02 U2729 (.o(wb1s_data_o[11]),
	.b(n1772),
	.a(n1773));
   no02s04 U2730 (.o(n1632),
	.b(wb0_sel_i[0]),
	.a(FE_OCPN658_wb1_cyc_o));
   in01s01 U2731 (.o(wb0_rty_o),
	.a(n2361));
   in01s01 U2732 (.o(wb0_err_o),
	.a(n2362));
   no02s02 U2733 (.o(n1634),
	.b(wb0_sel_i[2]),
	.a(FE_OCPN633_wb1_cyc_o));
   no02s02 U2734 (.o(n1635),
	.b(wb0_sel_i[3]),
	.a(FE_OCPN633_wb1_cyc_o));
   in01s01 U2735 (.o(wb0_sel_o[1]),
	.a(n1838));
   in01s01 U2736 (.o(wb0_sel_o[2]),
	.a(n1839));
   in01s01 U2737 (.o(wb0_sel_o[3]),
	.a(n1840));
   in01s01 U2739 (.o(wb1m_data_o[25]),
	.a(n1713));
   in01s01 U2740 (.o(wb1m_data_o[26]),
	.a(n1714));
   in01s01 U2741 (.o(wb1m_data_o[28]),
	.a(n1716));
   in01s01 U2742 (.o(wb1m_data_o[29]),
	.a(n1717));
   in01s01 U2743 (.o(wb1_rty_o),
	.a(n1720));
   in01s01 U2744 (.o(wb1m_data_o[4]),
	.a(n1692));
   in01s01 U2745 (.o(wb0_addr_o[1]),
	.a(n1842));
   in01s01 U2746 (.o(wb1m_data_o[3]),
	.a(n1691));
   in01s01 U2747 (.o(wb0_addr_o[0]),
	.a(n1841));
   in01s01 U2748 (.o(wb0_stb_o),
	.a(n1835));
   in01s01 U2749 (.o(wb0_we_o),
	.a(n1836));
   in01s01 U2750 (.o(wb1m_data_o[11]),
	.a(n1699));
   in01s01 U2751 (.o(wb1m_data_o[16]),
	.a(n1704));
   in01s01 U2752 (.o(wb1m_data_o[15]),
	.a(n1703));
   in01s01 U2753 (.o(wb1m_data_o[13]),
	.a(n1701));
   in01s01 U2754 (.o(wb1m_data_o[12]),
	.a(n1700));
   in01s01 U2755 (.o(wb1m_data_o[1]),
	.a(n1689));
   in01s01 U2757 (.o(wb1_err_o),
	.a(n1721));
   in01s01 U2758 (.o(wb1m_data_o[19]),
	.a(n1707));
   in01s01 U2759 (.o(wb1m_data_o[24]),
	.a(n1712));
   na02s01 U2760 (.o(n1856),
	.b(wb1_addr_i[15]),
	.a(n1414));
   na02s01 U2761 (.o(n1721),
	.b(wb0_err_i),
	.a(n1414));
   na02s01 U2762 (.o(n1689),
	.b(wb0s_data_i[1]),
	.a(FE_RN_17));
   na02s01 U2763 (.o(n1707),
	.b(wb0s_data_i[19]),
	.a(n1414));
   na02s01 U2764 (.o(n1712),
	.b(wb0s_data_i[24]),
	.a(FE_RN_17));
   na02s01 U2765 (.o(n2425),
	.b(wb1m_data_i[27]),
	.a(FE_OCPN277_wb0_cyc_o));
   na02s01 U2766 (.o(n2481),
	.b(wb0s_data_i[20]),
	.a(FE_OFN427_wb0_ack_i));
   na02s01 U2767 (.o(n2480),
	.b(wb0s_data_i[21]),
	.a(FE_OFN427_wb0_ack_i));
   na02s01 U2768 (.o(n2479),
	.b(wb0s_data_i[22]),
	.a(FE_OFN427_wb0_ack_i));
   na02s01 U2769 (.o(n2478),
	.b(wb0s_data_i[23]),
	.a(FE_OFN427_wb0_ack_i));
   na02s01 U2770 (.o(n2476),
	.b(wb0s_data_i[25]),
	.a(FE_OFN427_wb0_ack_i));
   na02s01 U2771 (.o(n2474),
	.b(wb0s_data_i[27]),
	.a(FE_OFN427_wb0_ack_i));
   na02s01 U2772 (.o(n2472),
	.b(wb0s_data_i[29]),
	.a(FE_OFN427_wb0_ack_i));
   na02s01 U2773 (.o(n2471),
	.b(wb0s_data_i[30]),
	.a(FE_OFN427_wb0_ack_i));
   na02s01 U2774 (.o(n2470),
	.b(wb0s_data_i[31]),
	.a(FE_OFN427_wb0_ack_i));
   no02s01 U2776 (.o(n1574),
	.b(n1575),
	.a(n1607));
   no02s01 U2777 (.o(n1582),
	.b(n1583),
	.a(n1607));
   no02s01 U2778 (.o(n1584),
	.b(n1585),
	.a(n1607));
   in01s01 U2779 (.o(n1612),
	.a(n1629));
   in01m20 U2782 (.o(n1901),
	.a(n1900));
   no02f20 U2783 (.o(n1536),
	.b(FE_OCPN186_n1893),
	.a(n1468));
   in01s01 U2784 (.o(n1724),
	.a(n1727));
   na02s01 U2785 (.o(n1608),
	.b(wb0_stb_i),
	.a(wb0_cyc_i));
   oa12s02 U2786 (.o(wb0m_data_o[6]),
	.c(n1984),
	.b(FE_OCPN658_wb1_cyc_o),
	.a(n1983));
   oa12s01 U2787 (.o(wb0m_data_o[22]),
	.c(n2248),
	.b(FE_OCPN656_wb1_cyc_o),
	.a(n2247));
   oa12s01 U2788 (.o(wb0m_data_o[21]),
	.c(n2233),
	.b(FE_OCPN658_wb1_cyc_o),
	.a(n2232));
   oa12m01 U2789 (.o(wb0m_data_o[19]),
	.c(n2206),
	.b(FE_OCPN667_wb1_cyc_o),
	.a(n2205));
   no02f04 U2790 (.o(n2275),
	.b(n2355),
	.a(n2271));
   na02s06 U2791 (.o(n1517),
	.b(n1516),
	.a(ch0_adr0[22]));
   no02f04 U2792 (.o(n2081),
	.b(FE_OCPN672_n1577),
	.a(n2079));
   na02s02 U2793 (.o(wb1s_data_o[5]),
	.b(n1754),
	.a(n1755));
   na02s02 U2794 (.o(wb1s_data_o[16]),
	.b(n1787),
	.a(n1788));
   na02s02 U2795 (.o(wb1s_data_o[21]),
	.b(n1802),
	.a(n1803));
   na02s02 U2796 (.o(wb1s_data_o[0]),
	.b(n1739),
	.a(n1740));
   na02s02 U2797 (.o(wb1s_data_o[20]),
	.b(n1799),
	.a(n1800));
   na02s02 U2799 (.o(wb1s_data_o[4]),
	.b(n1751),
	.a(n1752));
   na02s02 U2800 (.o(wb1s_data_o[1]),
	.b(n1742),
	.a(n1743));
   na02s01 U2801 (.o(wb1s_data_o[17]),
	.b(n1790),
	.a(n1791));
   na02s02 U2802 (.o(wb1s_data_o[18]),
	.b(n1793),
	.a(n1794));
   na02s02 U2803 (.o(wb1s_data_o[2]),
	.b(n1745),
	.a(n1746));
   no02f08 U2804 (.o(n2095),
	.b(n2156),
	.a(n2094));
   ao12f04 U2808 (.o(n2228),
	.c(n2226),
	.b(n2227),
	.a(FE_OCPN169_n2346));
   ao12f08 U2809 (.o(n1963),
	.c(n1959),
	.b(n1960),
	.a(FE_RN_14));
   na02f10 U2810 (.o(n1493),
	.b(n2177),
	.a(n2176));
   in01f20 U2812 (.o(n1620),
	.a(n1619));
   no02f20 U2813 (.o(n2007),
	.b(FE_OCPN664_FE_RN_16),
	.a(n1476));
   na03m01 U2814 (.o(n1726),
	.c(n1727),
	.b(wb1_we_i),
	.a(n1725));
   in01s01 U2815 (.o(n2475),
	.a(n1582));
   in01s01 U2816 (.o(n2473),
	.a(n1584));
   in01s01 U2817 (.o(n2477),
	.a(n1574));
   in01s01 U2818 (.o(n1723),
	.a(n1725));
   in01s01 U2819 (.o(n2360),
	.a(wb1s_data_i[31]));
   in01s01 U2820 (.o(n2188),
	.a(wb1s_data_i[18]));
   in01s01 U2821 (.o(n2151),
	.a(wb1s_data_i[16]));
   in01s01 U2822 (.o(n2170),
	.a(wb1s_data_i[17]));
   in01s01 U2823 (.o(n2352),
	.a(wb1s_data_i[30]));
   in01s01 U2824 (.o(n2338),
	.a(wb1s_data_i[29]));
   in01s01 U2825 (.o(n2206),
	.a(wb1s_data_i[19]));
   in01s01 U2826 (.o(n1605),
	.a(wb1_ack_i));
   in01s01 U2827 (.o(n2217),
	.a(wb1s_data_i[20]));
   in01s01 U2828 (.o(n2328),
	.a(wb1s_data_i[28]));
   in01s01 U2829 (.o(n2233),
	.a(wb1s_data_i[21]));
   in01s01 U2830 (.o(n1585),
	.a(wb0s_data_i[28]));
   in01s01 U2831 (.o(n2318),
	.a(wb1s_data_i[27]));
   in01s01 U2832 (.o(n2248),
	.a(wb1s_data_i[22]));
   in01s01 U2833 (.o(n1583),
	.a(wb0s_data_i[26]));
   in01s01 U2834 (.o(n1575),
	.a(wb0s_data_i[24]));
   in01s01 U2835 (.o(n2263),
	.a(wb1s_data_i[23]));
   in01s01 U2836 (.o(n2308),
	.a(wb1s_data_i[26]));
   in01s01 U2837 (.o(n2277),
	.a(wb1s_data_i[24]));
   in01s01 U2839 (.o(n2001),
	.a(wb1s_data_i[7]));
   in01s01 U2840 (.o(n1984),
	.a(wb1s_data_i[6]));
   in01s01 U2841 (.o(n1968),
	.a(wb1s_data_i[5]));
   in01s01 U2842 (.o(n2469),
	.a(dma_nd_i[0]));
   in01s01 U2843 (.o(n1950),
	.a(wb1s_data_i[4]));
   in01s01 U2844 (.o(n1930),
	.a(wb1s_data_i[3]));
   in01s01 U2845 (.o(n1909),
	.a(wb1s_data_i[2]));
   in01s01 U2846 (.o(n1886),
	.a(wb1s_data_i[1]));
   in01s01 U2847 (.o(n1880),
	.a(wb1s_data_i[0]));
   in01s01 U2848 (.o(n1611),
	.a(wb0_we_i));
   in01s01 U2849 (.o(n2019),
	.a(wb1s_data_i[8]));
   in01s01 U2850 (.o(n2083),
	.a(wb1s_data_i[12]));
   in01s01 U2851 (.o(n2133),
	.a(wb1s_data_i[15]));
   in01s01 U2852 (.o(n2115),
	.a(wb1s_data_i[14]));
   in01s01 U2853 (.o(n2099),
	.a(wb1s_data_i[13]));
   in01s01 U2854 (.o(n2033),
	.a(wb1s_data_i[9]));
   in01s01 U2855 (.o(n2049),
	.a(wb1s_data_i[10]));
   in01s01 U2856 (.o(n2069),
	.a(wb1s_data_i[11]));
   na02f40 U2857 (.o(n1516),
	.b(FE_OCPN545_n2159),
	.a(n1467));
   in01f10 U2858 (.o(n1467),
	.a(n1891));
   no02m20 U2859 (.o(n1473),
	.b(FE_OCPN106_slv0_adr_2_),
	.a(n2178));
   no02f20 U2860 (.o(n1621),
	.b(slv0_adr[3]),
	.a(slv0_adr[2]));
   oa12s01 U2861 (.o(wb0m_data_o[0]),
	.c(n1880),
	.b(FE_OCPN658_wb1_cyc_o),
	.a(n1879));
   na02f08 U2862 (.o(n1959),
	.b(u0_int_maska_5_),
	.a(FE_OCPN124_FE_RN_));
   no02m40 U2864 (.o(FE_OCPN659_wb1_cyc_o),
	.b(n1629),
	.a(n1732));
   na02f10 U2865 (.o(n1468),
	.b(slv0_adr[4]),
	.a(FE_RN_16));
   na02s02 U2866 (.o(n2187),
	.b(slv0_din[18]),
	.a(FE_OCPN626_wb1_cyc_o));
   na02f40 U2867 (.o(n1581),
	.b(FE_OCPN669_slv0_adr_4_),
	.a(n1621));
   na02f20 U2868 (.o(n1615),
	.b(n1523),
	.a(n1621));
   oa12s02 U2869 (.o(n766),
	.c(FE_OCPN368_n2194),
	.b(n2182),
	.a(n1616));
   oa12m02 U2870 (.o(n762),
	.c(FE_OCPN370_n2194),
	.b(n2110),
	.a(n2102));
   na02s02 U2871 (.o(n2247),
	.b(slv0_din[22]),
	.a(FE_OCPN657_wb1_cyc_o));
   na02f40 U2872 (.o(n1891),
	.b(n1530),
	.a(n1531));
   na02f06 U2873 (.o(n1897),
	.b(FE_OCPN163_n2346),
	.a(n1896));
   ao12m06 U2874 (.o(n2077),
	.c(n2343),
	.b(u0_int_maska_12_),
	.a(n2076));
   no02f04 U2875 (.o(n2230),
	.b(n2228),
	.a(n1469));
   na02s06 U2876 (.o(n1470),
	.b(ch0_adr0[21]),
	.a(FE_OCPN560_n2357));
   oa12f06 U2877 (.o(n1899),
	.c(FE_OCPN671_n2356),
	.b(n1898),
	.a(n1897));
   na02f40 U2878 (.o(n1521),
	.b(n1536),
	.a(n1537));
   na02f20 U2879 (.o(n1553),
	.b(FE_RN_16),
	.a(FE_RN_4));
   no02f40 U2880 (.o(n2356),
	.b(n1553),
	.a(n1471));
   no03f80 U2881 (.o(n1619),
	.c(FE_OCPN617_slv0_adr_5_),
	.b(slv0_adr[7]),
	.a(slv0_adr[6]));
   no02f04 U2882 (.o(n2186),
	.b(n2184),
	.a(n2185));
   oa22f08 U2883 (.o(n2028),
	.d(n2026),
	.c(FE_RN_14),
	.b(n2027),
	.a(FE_OCPN670_n2356));
   na04f40 U2884 (.o(n1471),
	.d(slv0_adr[4]),
	.c(slv0_adr[5]),
	.b(FE_OCPN138_slv0_adr_2_),
	.a(FE_OCPN511_slv0_adr_3_));
   no02f40 U2885 (.o(n1543),
	.b(n1620),
	.a(FE_OCPN186_n1893));
   ao12f06 U2888 (.o(n2107),
	.c(n2343),
	.b(u0_int_maska_14_),
	.a(n2106));
   no02f04 U2889 (.o(n2204),
	.b(n2202),
	.a(n2203));
   na02f10 U2890 (.o(n2176),
	.b(u0_int_maska_18_),
	.a(FE_OCPN122_FE_RN_));
   na02f40 U2891 (.o(n2178),
	.b(FE_RN_4),
	.a(n1619));
   na02f20 U2892 (.o(n1478),
	.b(slv0_adr[3]),
	.a(slv0_adr[5]));
   oa12f02 U2893 (.o(n2434),
	.c(n1481),
	.b(FE_OCPN167_n2346),
	.a(n1479));
   no03f40 U2895 (.o(n1566),
	.c(FE_OCPN512_slv0_adr_3_),
	.b(slv0_adr[4]),
	.a(FE_OCPN139_slv0_adr_2_));
   na02f10 U2896 (.o(n2177),
	.b(n1566),
	.a(u0_int_maskb_18_));
   in01s80 U2899 (.o(n1529),
	.a(slv0_we));
   no02f40 U2901 (.o(n1573),
	.b(n1891),
	.a(n1424));
   na02s03 U2903 (.o(n1892),
	.b(slv0_dout[2]),
	.a(n1573));
   oa22s04 U2904 (.o(n631),
	.d(FE_OCPN179_n1521),
	.c(n2314),
	.b(FE_OCPN462_n1521),
	.a(n2312));
   oa22f02 U2905 (.o(n607),
	.d(FE_OCPN180_n1521),
	.c(n2127),
	.b(FE_OCPN463_n1521),
	.a(n2120));
   oa22f02 U2906 (.o(n597),
	.d(FE_OCPN180_n1521),
	.c(n2043),
	.b(FE_OCPN463_n1521),
	.a(n2037));
   oa22f02 U2907 (.o(n605),
	.d(FE_OCPN180_n1521),
	.c(n2108),
	.b(FE_OCPN463_n1521),
	.a(n2104));
   oa22m04 U2908 (.o(n637),
	.d(FE_OCPN179_n1521),
	.c(n2347),
	.b(FE_OCPN462_n1521),
	.a(n2342));
   oa22f04 U2909 (.o(n609),
	.d(FE_OCPN180_n1521),
	.c(n2145),
	.b(FE_OCPN463_n1521),
	.a(n2138));
   oa22m02 U2910 (.o(n581),
	.d(FE_OCPN180_n1521),
	.c(n1898),
	.b(FE_OCPN463_n1521),
	.a(n1488));
   oa22s04 U2911 (.o(n621),
	.d(FE_OCPN179_n1521),
	.c(n2240),
	.b(FE_OCPN462_n1521),
	.a(n2237));
   oa22m02 U2913 (.o(n595),
	.d(FE_OCPN179_n1521),
	.c(n2027),
	.b(FE_OCPN464_n1521),
	.a(n2023));
   ao12m08 U2914 (.o(n2144),
	.c(n2343),
	.b(u0_int_maska_16_),
	.a(n2143));
   oa12s02 U2915 (.o(n657),
	.c(n2023),
	.b(n1513),
	.a(n2022));
   oa12f01 U2916 (.o(n659),
	.c(n2037),
	.b(n1513),
	.a(n2036));
   oa12m02 U2917 (.o(n747),
	.c(n2281),
	.b(n1513),
	.a(n2280));
   oa12s02 U2918 (.o(n742),
	.c(n1525),
	.b(n1513),
	.a(n1870));
   oa12f01 U2919 (.o(n645),
	.c(n1914),
	.b(n1513),
	.a(n1912));
   oa12m02 U2920 (.o(n752),
	.c(n2211),
	.b(n1513),
	.a(n2207));
   oa12s02 U2921 (.o(n750),
	.c(n2237),
	.b(n1513),
	.a(n2236));
   oa12s02 U2923 (.o(n751),
	.c(n2222),
	.b(n1513),
	.a(n2218));
   oa12s02 U2924 (.o(n749),
	.c(n2252),
	.b(n1513),
	.a(n2251));
   oa12s02 U2925 (.o(n649),
	.c(n1956),
	.b(n1513),
	.a(n1951));
   oa12s02 U2926 (.o(n653),
	.c(n1989),
	.b(n1513),
	.a(n1988));
   oa12s02 U2927 (.o(n651),
	.c(n1974),
	.b(n1513),
	.a(n1973));
   na02f02 U2929 (.o(n2437),
	.b(n1496),
	.a(n1498));
   na02f02 U2930 (.o(n2436),
	.b(n1499),
	.a(n1501));
   na02f02 U2931 (.o(n2435),
	.b(n1502),
	.a(n1504));
   na02f04 U2932 (.o(n2438),
	.b(n1505),
	.a(n1507));
   ao22f08 U2933 (.o(n2026),
	.d(u0_int_maska_9_),
	.c(n2343),
	.b(u0_int_maskb_9_),
	.a(FE_OCPN544_n2159));
   na02m40 U2934 (.o(n1513),
	.b(n2343),
	.a(FE_RN_8));
   na02m06 U2935 (.o(n2006),
	.b(slv0_dout[8]),
	.a(FE_OCPN370_n2194));
   na02f06 U2936 (.o(n1494),
	.b(n2196),
	.a(n2195));
   na02s10 U2937 (.o(n1492),
	.b(ch0_adr1[21]),
	.a(n2356));
   ao22f08 U2939 (.o(n2181),
	.d(n2356),
	.c(ch0_adr1[18]),
	.b(n1493),
	.a(FE_OCPN163_n2346));
   ao12f06 U2941 (.o(n2096),
	.c(ch0_adr0[13]),
	.b(n1416),
	.a(n2095));
   in01m10 U2942 (.o(n1495),
	.a(n2178));
   in01m20 U2943 (.o(n1547),
	.a(slv0_adr[9]));
   in01m20 U2944 (.o(n1548),
	.a(slv0_adr[8]));
   na02f10 U2945 (.o(n1510),
	.b(FE_RN_8),
	.a(n2343));
   in01f02 U2946 (.o(n1498),
	.a(n2325));
   in01f02 U2947 (.o(n1501),
	.a(n2335));
   in01m02 U2948 (.o(n1504),
	.a(n2349));
   in01m02 U2949 (.o(n1507),
	.a(n2315));
   oa22f06 U2950 (.o(n1921),
	.d(FE_OCPN671_n2356),
	.c(n1920),
	.b(FE_OCPN167_n2346),
	.a(FE_OCPN80_n1919));
   no03f80 U2951 (.o(n1871),
	.c(slv0_adr[7]),
	.b(slv0_adr[5]),
	.a(slv0_adr[6]));
   na02s10 U2952 (.o(n1738),
	.b(n1733),
	.a(n1734));
   no02s10 U2953 (.o(n1832),
	.b(n1737),
	.a(n1738));
   na02s02 U2954 (.o(n1929),
	.b(slv0_din[3]),
	.a(FE_OCPN629_wb1_cyc_o));
   na02f08 U2956 (.o(n1668),
	.b(ch0_adr1[19]),
	.a(FE_OCPN462_n1521));
   no03f80 U2957 (.o(n2343),
	.c(FE_OCPN137_slv0_adr_2_),
	.b(slv0_adr[4]),
	.a(slv0_adr[3]));
   na02s01 U2958 (.o(n2232),
	.b(slv0_din[21]),
	.a(FE_OCPN627_wb1_cyc_o));
   na02s01 U2959 (.o(n2363),
	.b(u3_u1_rf_ack),
	.a(FE_OCPN628_wb1_cyc_o));
   na02s02 U2960 (.o(n1983),
	.b(slv0_din[6]),
	.a(FE_OCPN629_wb1_cyc_o));
   na02s02 U2962 (.o(n2048),
	.b(slv0_din[10]),
	.a(FE_OCPN629_wb1_cyc_o));
   ao12f06 U2963 (.o(n2112),
	.c(ch0_adr0[14]),
	.b(n1416),
	.a(n2111));
   na02m08 U2964 (.o(n1617),
	.b(slv0_dout[6]),
	.a(FE_OCPN370_n2194));
   na02f08 U2965 (.o(n2195),
	.b(u0_int_maska_19_),
	.a(FE_OCPN122_FE_RN_));
   na02s02 U2966 (.o(n2205),
	.b(slv0_din[19]),
	.a(FE_OCPN631_wb1_cyc_o));
   no02f08 U2967 (.o(n1962),
	.b(FE_OCPN670_n2356),
	.a(n1961));
   in01f02 U2968 (.o(n2446),
	.a(n2204));
   na02m06 U2969 (.o(n1639),
	.b(slv0_dout[5]),
	.a(FE_OCPN367_n2194));
   ao12f06 U2970 (.o(n1982),
	.c(ch0_txsz[6]),
	.b(n2304),
	.a(n1976));
   oa12s02 U2971 (.o(n689),
	.c(n1573),
	.b(n2118),
	.a(n2117));
   oa12s02 U2972 (.o(n683),
	.c(n1573),
	.b(n2071),
	.a(n2070));
   na02f08 U2973 (.o(n1666),
	.b(ch0_adr1[18]),
	.a(FE_OCPN462_n1521));
   oa12f04 U2974 (.o(n758),
	.c(FE_OCPN367_n2194),
	.b(n1975),
	.a(n1617));
   na02m10 U2975 (.o(n2250),
	.b(slv0_dout[23]),
	.a(FE_OCPN613_n1516));
   na02m06 U2976 (.o(n2293),
	.b(slv0_dout[26]),
	.a(FE_OCPN614_n1516));
   na02s10 U2977 (.o(n2279),
	.b(slv0_dout[25]),
	.a(FE_OCPN612_n1516));
   na02m04 U2978 (.o(n2265),
	.b(slv0_dout[24]),
	.a(FE_OCPN615_n1516));
   na02m08 U2979 (.o(n2353),
	.b(slv0_dout[31]),
	.a(FE_OCPN612_n1516));
   oa12f02 U2981 (.o(n760),
	.c(FE_OCPN370_n2194),
	.b(n2008),
	.a(n2006));
   oa12f02 U2982 (.o(n757),
	.c(FE_OCPN367_n2194),
	.b(n1957),
	.a(n1639));
   na02s02 U2983 (.o(n2068),
	.b(slv0_din[11]),
	.a(FE_OCPN626_wb1_cyc_o));
   oa12f02 U2984 (.o(n524),
	.c(n1935),
	.b(FE_OCPN538_n1595),
	.a(n1934));
   na02m08 U2985 (.o(n1960),
	.b(u0_int_maskb_5_),
	.a(n1566));
   na02f08 U2986 (.o(n2196),
	.b(u0_int_maskb_19_),
	.a(n1566));
   oa12m02 U2987 (.o(n661),
	.c(n2054),
	.b(n1513),
	.a(n2053));
   na02s04 U2988 (.o(n2053),
	.b(ch0_txsz[11]),
	.a(n1513));
   oa12s02 U2989 (.o(n687),
	.c(n1573),
	.b(n2101),
	.a(n2100));
   oa12m02 U2990 (.o(n667),
	.c(n1573),
	.b(n1933),
	.a(n1932));
   oa12m02 U2991 (.o(n691),
	.c(n1573),
	.b(n2136),
	.a(n2135));
   oa12s02 U2992 (.o(n685),
	.c(n1573),
	.b(n2085),
	.a(n2084));
   oa12s02 U2993 (.o(n681),
	.c(n1573),
	.b(n2052),
	.a(n2051));
   na02m02 U2994 (.o(n1515),
	.b(FE_OCPN480_n1573),
	.a(ch0_adr0[10]));
   na02s02 U2995 (.o(n679),
	.b(n2035),
	.a(n1515));
   oa12m02 U2997 (.o(n677),
	.c(n1573),
	.b(n2025),
	.a(n2024));
   oa12m02 U2998 (.o(n671),
	.c(n1573),
	.b(n1972),
	.a(n1971));
   oa12s02 U2999 (.o(n669),
	.c(n1573),
	.b(n1953),
	.a(n1952));
   oa12f01 U3000 (.o(n665),
	.c(n1573),
	.b(n1916),
	.a(n1915));
   ao12f06 U3002 (.o(n2168),
	.c(ch0_txsz[17]),
	.b(n2225),
	.a(n2158));
   ao12f06 U3003 (.o(n2149),
	.c(ch0_txsz[16]),
	.b(n2225),
	.a(n2141));
   ao12f06 U3004 (.o(n2131),
	.c(ch0_txsz[15]),
	.b(n2225),
	.a(n2123));
   ao12f06 U3005 (.o(n2231),
	.c(n2225),
	.b(ch0_txsz[21]),
	.a(n2224));
   ao12f06 U3006 (.o(n1948),
	.c(n2304),
	.b(ch0_txsz[4]),
	.a(n1938));
   ao12f06 U3007 (.o(n1966),
	.c(n2304),
	.b(ch0_txsz[5]),
	.a(n1958));
   ao12f06 U3008 (.o(n1999),
	.c(ch0_txsz[7]),
	.b(n2304),
	.a(n1991));
   ao12f06 U3009 (.o(n2017),
	.c(ch0_txsz[8]),
	.b(n2225),
	.a(n2009));
   na02m02 U3011 (.o(n703),
	.b(n2235),
	.a(n1517));
   oa22f08 U3013 (.o(n2257),
	.d(n2255),
	.c(FE_OCPN169_n2346),
	.b(n2256),
	.a(FE_OCPN670_n2356));
   ao12f06 U3014 (.o(n1945),
	.c(n1941),
	.b(n1942),
	.a(FE_RN_14));
   na02s06 U3016 (.o(n2137),
	.b(ch0_txsz[16]),
	.a(FE_RN_9));
   oa22f08 U3017 (.o(n1896),
	.d(FE_RN_7),
	.c(n1894),
	.b(n1895),
	.a(n1424));
   no02f40 U3018 (.o(n2304),
	.b(FE_OCPN129_n2007),
	.a(n1576));
   ao12f06 U3019 (.o(n1994),
	.c(n2343),
	.b(u0_int_maska_7_),
	.a(n1993));
   ao12f08 U3020 (.o(n2012),
	.c(n2343),
	.b(u0_int_maska_8_),
	.a(n2011));
   ao12f08 U3021 (.o(n2042),
	.c(n2343),
	.b(u0_int_maska_10_),
	.a(n2041));
   oa22f08 U3023 (.o(n2164),
	.d(n2162),
	.c(FE_OCPN170_n2346),
	.b(n2163),
	.a(FE_OCPN671_n2356));
   oa22m06 U3024 (.o(n2079),
	.d(n2077),
	.c(FE_OCPN170_n2346),
	.b(n2078),
	.a(FE_OCPN671_n2356));
   oa22f06 U3027 (.o(n2109),
	.d(n2107),
	.c(FE_OCPN170_n2346),
	.b(n2108),
	.a(FE_OCPN671_n2356));
   oa22f06 U3028 (.o(n2335),
	.d(n2333),
	.c(FE_OCPN169_n2346),
	.b(n2334),
	.a(FE_OCPN670_n2356));
   ao12f06 U3031 (.o(n2126),
	.c(n2343),
	.b(u0_int_maska_15_),
	.a(n2125));
   oa22f08 U3032 (.o(n2146),
	.d(n2144),
	.c(FE_RN_15),
	.b(n2145),
	.a(FE_OCPN671_n2356));
   ao12f08 U3033 (.o(n2162),
	.c(n2343),
	.b(u0_int_maska_17_),
	.a(n2161));
   na02f03 U3034 (.o(n1550),
	.b(n1551),
	.a(n1552));
   na02s06 U3035 (.o(n1925),
	.b(ch0_txsz[3]),
	.a(n1924));
   oa22f06 U3036 (.o(n2301),
	.d(n2299),
	.c(FE_OCPN169_n2346),
	.b(n2300),
	.a(FE_OCPN670_n2356));
   oa22f08 U3038 (.o(n2242),
	.d(n2239),
	.c(FE_OCPN169_n2346),
	.b(n2240),
	.a(FE_OCPN670_n2356));
   oa22f06 U3039 (.o(n2271),
	.d(n2269),
	.c(FE_OCPN169_n2346),
	.b(n2270),
	.a(FE_OCPN670_n2356));
   oa22f08 U3041 (.o(n2044),
	.d(n2042),
	.c(FE_OCPN171_n2346),
	.b(n2043),
	.a(FE_OCPN671_n2356));
   no02f06 U3042 (.o(n2097),
	.b(FE_OCPN673_n1577),
	.a(n2093));
   no02f04 U3043 (.o(n2113),
	.b(FE_OCPN672_n1577),
	.a(n2109));
   oa22f08 U3044 (.o(n2014),
	.d(n2012),
	.c(FE_RN_15),
	.b(n2013),
	.a(FE_OCPN671_n2356));
   oa22m04 U3045 (.o(n2315),
	.d(n2313),
	.c(FE_OCPN169_n2346),
	.b(n2314),
	.a(FE_OCPN670_n2356));
   oa22f08 U3046 (.o(n1996),
	.d(n1994),
	.c(FE_RN_15),
	.b(n1995),
	.a(FE_OCPN671_n2356));
   no02f04 U3047 (.o(n2261),
	.b(n2355),
	.a(n2257));
   no02f04 U3048 (.o(n2246),
	.b(n2355),
	.a(n2242));
   na02f04 U3049 (.o(n2452),
	.b(n2096),
	.a(n2097));
   na02f04 U3050 (.o(n2451),
	.b(n2112),
	.a(n2113));
   no02f06 U3051 (.o(n2167),
	.b(FE_OCPN672_n1577),
	.a(n2164));
   no02f06 U3052 (.o(n2016),
	.b(FE_OCPN673_n1577),
	.a(n2014));
   na02f02 U3054 (.o(n2442),
	.b(n2260),
	.a(n2261));
   na02f02 U3055 (.o(n2439),
	.b(n2305),
	.a(n2306));
   na02f02 U3056 (.o(n2440),
	.b(n2288),
	.a(n2289));
   na02f04 U3057 (.o(n2443),
	.b(n2245),
	.a(n2246));
   na02f02 U3058 (.o(n2441),
	.b(n2274),
	.a(n2275));
   na02f04 U3059 (.o(n2463),
	.b(n1906),
	.a(n1907));
   na02f02 U3060 (.o(n2462),
	.b(n1927),
	.a(n1928));
   na02f02 U3061 (.o(n2444),
	.b(n2230),
	.a(n2231));
   na03f06 U3063 (.o(n2457),
	.c(n2015),
	.b(n2016),
	.a(n2017));
   na03f06 U3065 (.o(n2458),
	.c(n1997),
	.b(n1998),
	.a(n1999));
   no02f20 U3072 (.o(n1562),
	.b(FE_RN_7),
	.a(FE_OCPN554_n1529));
   na02s01 U3075 (.o(wb1_addr_o[30]),
	.b(n1736),
	.a(wb1_cyc_o));
   na02s01 U3076 (.o(wb1_addr_o[29]),
	.b(n1734),
	.a(wb1_cyc_o));
   oa12s01 U3077 (.o(n819),
	.c(wb0_ack_i),
	.b(n1774),
	.a(n2489));
   oa12m02 U3078 (.o(n734),
	.c(n1883),
	.b(FE_OCPN363_n2194),
	.a(n1882));
   na02m02 U3079 (.o(n1882),
	.b(ch0_csr[1]),
	.a(FE_OCPN363_n2194));
   oa12s01 U3080 (.o(wb1_addr_o[4]),
	.c(n1645),
	.b(FE_OCPN656_wb1_cyc_o),
	.a(wb1_cyc_o));
   oa12s01 U3081 (.o(wb1_addr_o[7]),
	.c(n1651),
	.b(FE_OCPN658_wb1_cyc_o),
	.a(wb1_cyc_o));
   oa12f02 U3082 (.o(n615),
	.c(n2192),
	.b(FE_OCPN462_n1521),
	.a(n1668));
   na02s02 U3083 (.o(n1670),
	.b(ch0_adr1[20]),
	.a(n1521));
   oa12f02 U3084 (.o(n619),
	.c(n2222),
	.b(FE_OCPN462_n1521),
	.a(n1672));
   oa12m04 U3085 (.o(n697),
	.c(n2192),
	.b(FE_OCPN622_n1516),
	.a(n2189));
   na02s08 U3086 (.o(n2189),
	.b(ch0_adr0[19]),
	.a(n1516));
   oa12m02 U3087 (.o(n717),
	.c(n2332),
	.b(FE_OCPN620_n1516),
	.a(n2331));
   na02s04 U3088 (.o(n2331),
	.b(ch0_adr0[29]),
	.a(n1516));
   oa12m04 U3089 (.o(n715),
	.c(n2322),
	.b(FE_OCPN622_n1516),
	.a(n2321));
   na02s03 U3090 (.o(n2321),
	.b(ch0_adr0[28]),
	.a(n1516));
   oa12m04 U3091 (.o(n701),
	.c(n2222),
	.b(FE_OCPN622_n1516),
	.a(n2219));
   na02s06 U3092 (.o(n2219),
	.b(ch0_adr0[21]),
	.a(n1516));
   oa12f04 U3093 (.o(n713),
	.c(n2312),
	.b(FE_OCPN622_n1516),
	.a(n2311));
   na02s08 U3094 (.o(n2311),
	.b(ch0_adr0[27]),
	.a(n1516));
   oa12m04 U3095 (.o(n699),
	.c(n2211),
	.b(FE_OCPN622_n1516),
	.a(n2208));
   na02s06 U3096 (.o(n2208),
	.b(ch0_adr0[20]),
	.a(n1516));
   oa12f04 U3097 (.o(n719),
	.c(n2342),
	.b(FE_OCPN622_n1516),
	.a(n2341));
   na02s08 U3098 (.o(n2341),
	.b(ch0_adr0[30]),
	.a(n1516));
   oa12f04 U3099 (.o(n695),
	.c(n2175),
	.b(FE_OCPN622_n1516),
	.a(n2172));
   na02s06 U3100 (.o(n2172),
	.b(ch0_adr0[18]),
	.a(n1516));
   oa12s01 U3101 (.o(wb0m_data_o[28]),
	.c(n2328),
	.b(FE_OCPN658_wb1_cyc_o),
	.a(n2327));
   na02s01 U3102 (.o(n2327),
	.b(slv0_din[28]),
	.a(FE_OCPN631_wb1_cyc_o));
   oa12s01 U3103 (.o(wb0m_data_o[24]),
	.c(n2277),
	.b(FE_OCPN658_wb1_cyc_o),
	.a(n2276));
   na02s01 U3104 (.o(n2276),
	.b(slv0_din[24]),
	.a(FE_OCPN627_wb1_cyc_o));
   oa12s01 U3105 (.o(wb0m_data_o[18]),
	.c(n2188),
	.b(FE_OCPN658_wb1_cyc_o),
	.a(n2187));
   na02s02 U3106 (.o(n2378),
	.b(FE_OCPN528_n1597),
	.a(de_csr[4]));
   na02s01 U3107 (.o(n2390),
	.b(FE_OCPN528_n1597),
	.a(de_csr[10]));
   oa12s01 U3108 (.o(wb0m_data_o[26]),
	.c(n2308),
	.b(FE_OCPN658_wb1_cyc_o),
	.a(n2307));
   na02s01 U3109 (.o(n2307),
	.b(slv0_din[26]),
	.a(FE_OCPN626_wb1_cyc_o));
   na02s02 U3110 (.o(n1833),
	.b(de_csr[31]),
	.a(n1832));
   na02s02 U3111 (.o(n1834),
	.b(wb0m_data_i[31]),
	.a(FE_OCPN642_wb1_cyc_o));
   na02s02 U3112 (.o(n1826),
	.b(de_csr[29]),
	.a(FE_RN_12));
   na02s02 U3113 (.o(n1827),
	.b(wb0m_data_i[29]),
	.a(FE_OCPN666_wb1_cyc_o));
   na02s02 U3114 (.o(n1823),
	.b(de_csr[28]),
	.a(FE_RN_1));
   na02s02 U3115 (.o(n1824),
	.b(wb0m_data_i[28]),
	.a(FE_OCPN643_wb1_cyc_o));
   na02s02 U3116 (.o(n1820),
	.b(de_csr[27]),
	.a(n1832));
   na02s02 U3117 (.o(n1821),
	.b(wb0m_data_i[27]),
	.a(FE_OCPN666_wb1_cyc_o));
   na02s02 U3118 (.o(n1817),
	.b(de_csr[26]),
	.a(FE_RN_1));
   na02s01 U3119 (.o(n1818),
	.b(wb0m_data_i[26]),
	.a(FE_OCPN643_wb1_cyc_o));
   na02s08 U3120 (.o(n1811),
	.b(de_csr[24]),
	.a(FE_RN_1));
   na02s02 U3121 (.o(n1812),
	.b(wb0m_data_i[24]),
	.a(FE_OCPN642_wb1_cyc_o));
   na02s02 U3122 (.o(n1829),
	.b(de_csr[30]),
	.a(n1832));
   na02s03 U3123 (.o(n1830),
	.b(wb0m_data_i[30]),
	.a(FE_OCPN642_wb1_cyc_o));
   na02s01 U3124 (.o(n1739),
	.b(FE_RN_1),
	.a(de_csr[0]));
   na02s01 U3125 (.o(n1742),
	.b(de_csr[1]),
	.a(FE_RN_1));
   na02s02 U3126 (.o(n1743),
	.b(wb0m_data_i[1]),
	.a(FE_OCPN666_wb1_cyc_o));
   na02s02 U3127 (.o(n1793),
	.b(de_csr[18]),
	.a(n1832));
   na02s02 U3128 (.o(n1794),
	.b(wb0m_data_i[18]),
	.a(FE_OCPN642_wb1_cyc_o));
   na02s02 U3129 (.o(n1746),
	.b(wb0m_data_i[2]),
	.a(FE_OCPN643_wb1_cyc_o));
   na02s02 U3130 (.o(n1760),
	.b(de_csr[7]),
	.a(FE_RN_11));
   na02s04 U3131 (.o(n1757),
	.b(de_csr[6]),
	.a(FE_RN_12));
   na02s01 U3132 (.o(n2394),
	.b(FE_OCPN528_n1597),
	.a(de_csr[12]));
   oa12f02 U3133 (.o(n585),
	.c(FE_OCPN180_n1521),
	.b(n1943),
	.a(n1644));
   na02f06 U3134 (.o(n1644),
	.b(FE_OCPN178_n1521),
	.a(slv0_dout[4]));
   na02s01 U3136 (.o(n2370),
	.b(FE_OCPN528_n1597),
	.a(de_csr[0]));
   na02s01 U3137 (.o(n2374),
	.b(FE_OCPN528_n1597),
	.a(de_csr[2]));
   na02s02 U3138 (.o(n2384),
	.b(FE_OCPN528_n1597),
	.a(de_csr[7]));
   na02s01 U3139 (.o(n2372),
	.b(FE_OCPN528_n1597),
	.a(de_csr[1]));
   na02s01 U3140 (.o(n2376),
	.b(FE_OCPN528_n1597),
	.a(de_csr[3]));
   oa12s02 U3141 (.o(wb0m_data_o[29]),
	.c(n2338),
	.b(FE_OCPN667_wb1_cyc_o),
	.a(n2337));
   na02s02 U3142 (.o(n2337),
	.b(slv0_din[29]),
	.a(FE_OCPN627_wb1_cyc_o));
   na02s01 U3143 (.o(n2402),
	.b(FE_OCPN528_n1597),
	.a(de_csr[16]));
   oa12m02 U3144 (.o(n633),
	.c(FE_OCPN180_n1521),
	.b(n2324),
	.a(n1684));
   na02s10 U3145 (.o(n1684),
	.b(FE_OCPN176_n1521),
	.a(slv0_dout[28]));
   na02s03 U3146 (.o(n1879),
	.b(slv0_din[0]),
	.a(FE_OCPN629_wb1_cyc_o));
   na02s01 U3147 (.o(n2406),
	.b(FE_OCPN528_n1597),
	.a(de_csr[18]));
   na02s01 U3148 (.o(n2404),
	.b(FE_OCPN528_n1597),
	.a(de_csr[17]));
   na02s01 U3149 (.o(n2400),
	.b(FE_OCPN528_n1597),
	.a(de_csr[15]));
   na02s01 U3150 (.o(n2392),
	.b(FE_OCPN528_n1597),
	.a(de_csr[11]));
   na02s04 U3151 (.o(n2004),
	.b(ch0_txsz[8]),
	.a(FE_RN_9));
   na02s01 U3152 (.o(n2380),
	.b(FE_OCPN528_n1597),
	.a(de_csr[5]));
   na02s01 U3153 (.o(n2386),
	.b(FE_OCPN528_n1597),
	.a(de_csr[8]));
   na02s06 U3154 (.o(n2102),
	.b(slv0_dout[14]),
	.a(FE_OCPN370_n2194));
   oa12s01 U3155 (.o(n823),
	.c(wb0_ack_i),
	.b(n1762),
	.a(n2493));
   oa12s01 U3156 (.o(n824),
	.c(wb0_ack_i),
	.b(n1759),
	.a(n2494));
   oa12s01 U3157 (.o(n826),
	.c(FE_OFN427_wb0_ack_i),
	.b(n1753),
	.a(n2496));
   oa12s01 U3158 (.o(n825),
	.c(wb0_ack_i),
	.b(n1756),
	.a(n2495));
   oa12s01 U3159 (.o(n827),
	.c(wb0_ack_i),
	.b(n1750),
	.a(n2497));
   no02m04 U3160 (.o(n2303),
	.b(FE_OCPN562_n2357),
	.a(n2302));
   no02f06 U3161 (.o(n2287),
	.b(FE_OCPN566_n2357),
	.a(n2286));
   no02m06 U3162 (.o(n2244),
	.b(FE_OCPN566_n2357),
	.a(n2243));
   no02m06 U3163 (.o(n2273),
	.b(FE_OCPN562_n2357),
	.a(n2272));
   oa12f02 U3164 (.o(n625),
	.c(FE_OCPN179_n1521),
	.b(n2270),
	.a(n1677));
   na02m04 U3165 (.o(n2235),
	.b(slv0_dout[22]),
	.a(FE_OCPN613_n1516));
   oa12f02 U3166 (.o(n721),
	.c(FE_OCPN613_n1516),
	.b(n2358),
	.a(n2353));
   oa12m04 U3167 (.o(n705),
	.c(FE_OCPN613_n1516),
	.b(n2258),
	.a(n2250));
   oa12f02 U3168 (.o(n711),
	.c(FE_OCPN613_n1516),
	.b(n2302),
	.a(n2293));
   oa12f02 U3169 (.o(n709),
	.c(FE_OCPN613_n1516),
	.b(n2286),
	.a(n2279));
   oa12m02 U3170 (.o(n707),
	.c(FE_OCPN613_n1516),
	.b(n2272),
	.a(n2265));
   na02s04 U3171 (.o(n2035),
	.b(slv0_dout[10]),
	.a(n1573));
   na02s04 U3172 (.o(n2135),
	.b(slv0_dout[16]),
	.a(n1573));
   in01s01 U3173 (.o(n2136),
	.a(ch0_adr0[16]));
   na02s04 U3174 (.o(n2051),
	.b(slv0_dout[11]),
	.a(n1573));
   no02f08 U3176 (.o(n1976),
	.b(n2156),
	.a(n1975));
   no02f08 U3177 (.o(n1958),
	.b(n2156),
	.a(n1957));
   no02f08 U3178 (.o(n1938),
	.b(n2156),
	.a(n1937));
   oa12m02 U3179 (.o(n673),
	.c(n1573),
	.b(n1987),
	.a(n1986));
   na02s08 U3180 (.o(n2022),
	.b(ch0_txsz[9]),
	.a(FE_RN_9));
   na02m03 U3181 (.o(n1616),
	.b(slv0_dout[18]),
	.a(FE_OCPN368_n2194));
   ao22f04 U3182 (.o(n2323),
	.d(u0_int_maska_28_),
	.c(n2343),
	.b(u0_int_maskb_28_),
	.a(FE_OCPN544_n2159));
   no02f06 U3183 (.o(n1559),
	.b(n1876),
	.a(n1424));
   oa12m02 U3184 (.o(n755),
	.c(n1533),
	.b(n1513),
	.a(n2155));
   oa12f02 U3185 (.o(n589),
	.c(FE_OCPN179_n1521),
	.b(n1978),
	.a(n1648));
   na02f06 U3186 (.o(n1648),
	.b(FE_OCPN178_n1521),
	.a(slv0_dout[6]));
   na02f06 U3187 (.o(n1646),
	.b(FE_OCPN178_n1521),
	.a(slv0_dout[5]));
   oa12f04 U3188 (.o(n627),
	.c(FE_OCPN179_n1521),
	.b(n2284),
	.a(n1679));
   na02f08 U3189 (.o(n1679),
	.b(FE_OCPN178_n1521),
	.a(slv0_dout[25]));
   oa12m02 U3190 (.o(n623),
	.c(FE_OCPN179_n1521),
	.b(n2256),
	.a(n1675));
   na02s06 U3191 (.o(n1675),
	.b(FE_OCPN176_n1521),
	.a(slv0_dout[23]));
   na02s02 U3192 (.o(n2294),
	.b(ch0_txsz[26]),
	.a(n1510));
   na02s02 U3193 (.o(n2280),
	.b(ch0_txsz[25]),
	.a(n1510));
   na02s04 U3194 (.o(n1870),
	.b(ch0_txsz[0]),
	.a(FE_RN_9));
   no02f08 U3195 (.o(n2106),
	.b(n1425),
	.a(n2105));
   na02s06 U3196 (.o(n1971),
	.b(slv0_dout[6]),
	.a(n1573));
   na02m04 U3197 (.o(n1915),
	.b(slv0_dout[3]),
	.a(n1573));
   na02m03 U3198 (.o(n1952),
	.b(slv0_dout[5]),
	.a(n1573));
   oa12f02 U3199 (.o(n693),
	.c(n1573),
	.b(n2154),
	.a(n2153));
   no02f08 U3200 (.o(n1532),
	.b(FE_OCPN479_n1573),
	.a(n1533));
   na02m04 U3201 (.o(n2024),
	.b(slv0_dout[9]),
	.a(n1573));
   no02f10 U3203 (.o(n2161),
	.b(n1424),
	.a(n2160));
   no02f08 U3204 (.o(n2158),
	.b(n2156),
	.a(n2157));
   no02f08 U3205 (.o(n2009),
	.b(n2156),
	.a(n2008));
   no02f08 U3208 (.o(n2141),
	.b(n2156),
	.a(n2140));
   no02f08 U3209 (.o(n2123),
	.b(n2156),
	.a(n2122));
   na02s02 U3210 (.o(n2207),
	.b(ch0_txsz[20]),
	.a(n1510));
   na02s02 U3211 (.o(n2236),
	.b(ch0_txsz[22]),
	.a(n1510));
   na02s02 U3212 (.o(n2218),
	.b(ch0_txsz[21]),
	.a(n1510));
   na02s03 U3213 (.o(n2251),
	.b(ch0_txsz[23]),
	.a(n1510));
   na02s04 U3214 (.o(n1951),
	.b(ch0_txsz[5]),
	.a(FE_RN_9));
   na02s04 U3215 (.o(n1988),
	.b(ch0_txsz[7]),
	.a(FE_RN_9));
   na02s06 U3216 (.o(n1973),
	.b(ch0_txsz[6]),
	.a(FE_RN_9));
   na02s06 U3217 (.o(n1931),
	.b(ch0_txsz[4]),
	.a(FE_RN_9));
   ao22f04 U3218 (.o(n2333),
	.d(u0_int_maska_29_),
	.c(n2343),
	.b(u0_int_maskb_29_),
	.a(FE_OCPN544_n2159));
   ao22m08 U3219 (.o(n2345),
	.d(u0_int_maska_30_),
	.c(n2343),
	.b(u0_int_maskb_30_),
	.a(FE_OCPN544_n2159));
   ao22m04 U3220 (.o(n2313),
	.d(u0_int_maska_27_),
	.c(n2343),
	.b(u0_int_maskb_27_),
	.a(FE_OCPN544_n2159));
   na02s04 U3221 (.o(n2070),
	.b(slv0_dout[12]),
	.a(n1573));
   na02s04 U3222 (.o(n1932),
	.b(slv0_dout[4]),
	.a(n1573));
   na02s03 U3223 (.o(n2100),
	.b(slv0_dout[14]),
	.a(n1573));
   na02s06 U3224 (.o(n2117),
	.b(slv0_dout[15]),
	.a(n1573));
   in01s01 U3225 (.o(n2118),
	.a(ch0_adr0[15]));
   oa12f02 U3226 (.o(n603),
	.c(FE_OCPN180_n1521),
	.b(n2092),
	.a(n1659));
   na02s10 U3227 (.o(n1659),
	.b(FE_OCPN176_n1521),
	.a(slv0_dout[13]));
   oa12f02 U3228 (.o(n601),
	.c(FE_OCPN180_n1521),
	.b(n2078),
	.a(n1657));
   na02f06 U3229 (.o(n1657),
	.b(FE_OCPN178_n1521),
	.a(slv0_dout[12]));
   oa12f02 U3230 (.o(n599),
	.c(FE_OCPN180_n1521),
	.b(n2063),
	.a(n1655));
   na02m08 U3231 (.o(n1655),
	.b(FE_OCPN176_n1521),
	.a(slv0_dout[11]));
   oa12m02 U3232 (.o(n629),
	.c(FE_OCPN179_n1521),
	.b(n2300),
	.a(n1681));
   na02m06 U3233 (.o(n1681),
	.b(FE_OCPN176_n1521),
	.a(slv0_dout[26]));
   no02f10 U3234 (.o(n1991),
	.b(n2156),
	.a(n1990));
   oa12s02 U3235 (.o(n663),
	.c(n1573),
	.b(n1904),
	.a(n1892));
   oa12f02 U3236 (.o(n611),
	.c(FE_OCPN180_n1521),
	.b(n2163),
	.a(n1664));
   na02f06 U3237 (.o(n1664),
	.b(FE_OCPN178_n1521),
	.a(slv0_dout[17]));
   oa12f02 U3238 (.o(n591),
	.c(FE_OCPN180_n1521),
	.b(n1995),
	.a(n1650));
   na02m08 U3239 (.o(n1650),
	.b(FE_OCPN176_n1521),
	.a(slv0_dout[7]));
   oa12f02 U3240 (.o(n583),
	.c(FE_OCPN180_n1521),
	.b(n1920),
	.a(n1642));
   na02f08 U3241 (.o(n1642),
	.b(FE_OCPN178_n1521),
	.a(slv0_dout[3]));
   na02s04 U3242 (.o(n2003),
	.b(slv0_dout[8]),
	.a(n1573));
   na02s04 U3243 (.o(n1534),
	.b(FE_OCPN478_n1573),
	.a(ch0_adr0[8]));
   oa12s01 U3244 (.o(n818),
	.c(wb0_ack_i),
	.b(n1777),
	.a(n2488));
   oa12s01 U3245 (.o(n817),
	.c(wb0_ack_i),
	.b(n1780),
	.a(n2487));
   oa12s01 U3246 (.o(n816),
	.c(wb0_ack_i),
	.b(n1783),
	.a(n2486));
   oa12s01 U3247 (.o(n815),
	.c(wb0_ack_i),
	.b(n1786),
	.a(n2485));
   oa12s01 U3248 (.o(n814),
	.c(wb0_ack_i),
	.b(n1789),
	.a(n2484));
endmodule

