VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram45_1024x32
  FOREIGN fakeram45_1024x32 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 104.500 BY 317.800 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.365 0.070 1.435 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.165 0.070 4.235 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.965 0.070 7.035 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.765 0.070 9.835 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.565 0.070 12.635 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.365 0.070 15.435 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.165 0.070 18.235 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.765 0.070 23.835 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.565 0.070 26.635 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.365 0.070 29.435 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.165 0.070 32.235 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.965 0.070 35.035 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.765 0.070 37.835 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.565 0.070 40.635 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.365 0.070 43.435 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.165 0.070 46.235 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.965 0.070 49.035 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.765 0.070 51.835 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.565 0.070 54.635 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.365 0.070 57.435 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.165 0.070 60.235 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.965 0.070 63.035 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.765 0.070 65.835 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.565 0.070 68.635 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.365 0.070 71.435 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.165 0.070 74.235 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.965 0.070 77.035 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.765 0.070 79.835 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.565 0.070 82.635 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.365 0.070 85.435 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.165 0.070 88.235 ;
    END
  END w_mask_in[31]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.545 0.070 90.615 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.345 0.070 93.415 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.145 0.070 96.215 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.945 0.070 99.015 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.745 0.070 101.815 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.545 0.070 104.615 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.345 0.070 107.415 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.145 0.070 110.215 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.945 0.070 113.015 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.745 0.070 115.815 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.545 0.070 118.615 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.345 0.070 121.415 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.145 0.070 124.215 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.945 0.070 127.015 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.745 0.070 129.815 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 132.545 0.070 132.615 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 135.345 0.070 135.415 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 138.145 0.070 138.215 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 140.945 0.070 141.015 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 143.745 0.070 143.815 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 146.545 0.070 146.615 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 149.345 0.070 149.415 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 152.145 0.070 152.215 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 154.945 0.070 155.015 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 157.745 0.070 157.815 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 160.545 0.070 160.615 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 163.345 0.070 163.415 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 166.145 0.070 166.215 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 168.945 0.070 169.015 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 171.745 0.070 171.815 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 174.545 0.070 174.615 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 177.345 0.070 177.415 ;
    END
  END rd_out[31]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 179.725 0.070 179.795 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 182.525 0.070 182.595 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 185.325 0.070 185.395 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 188.125 0.070 188.195 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 190.925 0.070 190.995 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 193.725 0.070 193.795 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 196.525 0.070 196.595 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 199.325 0.070 199.395 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 202.125 0.070 202.195 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 204.925 0.070 204.995 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 207.725 0.070 207.795 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 210.525 0.070 210.595 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 213.325 0.070 213.395 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 216.125 0.070 216.195 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 218.925 0.070 218.995 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 221.725 0.070 221.795 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 224.525 0.070 224.595 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 227.325 0.070 227.395 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 230.125 0.070 230.195 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 232.925 0.070 232.995 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 235.725 0.070 235.795 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 238.525 0.070 238.595 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 241.325 0.070 241.395 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 244.125 0.070 244.195 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 246.925 0.070 246.995 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 249.725 0.070 249.795 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 252.525 0.070 252.595 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 255.325 0.070 255.395 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 258.125 0.070 258.195 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 260.925 0.070 260.995 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 263.725 0.070 263.795 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 266.525 0.070 266.595 ;
    END
  END wd_in[31]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 268.905 0.070 268.975 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 271.705 0.070 271.775 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 274.505 0.070 274.575 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 277.305 0.070 277.375 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 280.105 0.070 280.175 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 282.905 0.070 282.975 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 285.705 0.070 285.775 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 288.505 0.070 288.575 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 291.305 0.070 291.375 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 294.105 0.070 294.175 ;
    END
  END addr_in[9]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 296.485 0.070 296.555 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 299.285 0.070 299.355 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 302.085 0.070 302.155 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 316.400 ;
      RECT 3.500 1.400 3.780 316.400 ;
      RECT 5.740 1.400 6.020 316.400 ;
      RECT 7.980 1.400 8.260 316.400 ;
      RECT 10.220 1.400 10.500 316.400 ;
      RECT 12.460 1.400 12.740 316.400 ;
      RECT 14.700 1.400 14.980 316.400 ;
      RECT 16.940 1.400 17.220 316.400 ;
      RECT 19.180 1.400 19.460 316.400 ;
      RECT 21.420 1.400 21.700 316.400 ;
      RECT 23.660 1.400 23.940 316.400 ;
      RECT 25.900 1.400 26.180 316.400 ;
      RECT 28.140 1.400 28.420 316.400 ;
      RECT 30.380 1.400 30.660 316.400 ;
      RECT 32.620 1.400 32.900 316.400 ;
      RECT 34.860 1.400 35.140 316.400 ;
      RECT 37.100 1.400 37.380 316.400 ;
      RECT 39.340 1.400 39.620 316.400 ;
      RECT 41.580 1.400 41.860 316.400 ;
      RECT 43.820 1.400 44.100 316.400 ;
      RECT 46.060 1.400 46.340 316.400 ;
      RECT 48.300 1.400 48.580 316.400 ;
      RECT 50.540 1.400 50.820 316.400 ;
      RECT 52.780 1.400 53.060 316.400 ;
      RECT 55.020 1.400 55.300 316.400 ;
      RECT 57.260 1.400 57.540 316.400 ;
      RECT 59.500 1.400 59.780 316.400 ;
      RECT 61.740 1.400 62.020 316.400 ;
      RECT 63.980 1.400 64.260 316.400 ;
      RECT 66.220 1.400 66.500 316.400 ;
      RECT 68.460 1.400 68.740 316.400 ;
      RECT 70.700 1.400 70.980 316.400 ;
      RECT 72.940 1.400 73.220 316.400 ;
      RECT 75.180 1.400 75.460 316.400 ;
      RECT 77.420 1.400 77.700 316.400 ;
      RECT 79.660 1.400 79.940 316.400 ;
      RECT 81.900 1.400 82.180 316.400 ;
      RECT 84.140 1.400 84.420 316.400 ;
      RECT 86.380 1.400 86.660 316.400 ;
      RECT 88.620 1.400 88.900 316.400 ;
      RECT 90.860 1.400 91.140 316.400 ;
      RECT 93.100 1.400 93.380 316.400 ;
      RECT 95.340 1.400 95.620 316.400 ;
      RECT 97.580 1.400 97.860 316.400 ;
      RECT 99.820 1.400 100.100 316.400 ;
      RECT 102.060 1.400 102.340 316.400 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 316.400 ;
      RECT 4.620 1.400 4.900 316.400 ;
      RECT 6.860 1.400 7.140 316.400 ;
      RECT 9.100 1.400 9.380 316.400 ;
      RECT 11.340 1.400 11.620 316.400 ;
      RECT 13.580 1.400 13.860 316.400 ;
      RECT 15.820 1.400 16.100 316.400 ;
      RECT 18.060 1.400 18.340 316.400 ;
      RECT 20.300 1.400 20.580 316.400 ;
      RECT 22.540 1.400 22.820 316.400 ;
      RECT 24.780 1.400 25.060 316.400 ;
      RECT 27.020 1.400 27.300 316.400 ;
      RECT 29.260 1.400 29.540 316.400 ;
      RECT 31.500 1.400 31.780 316.400 ;
      RECT 33.740 1.400 34.020 316.400 ;
      RECT 35.980 1.400 36.260 316.400 ;
      RECT 38.220 1.400 38.500 316.400 ;
      RECT 40.460 1.400 40.740 316.400 ;
      RECT 42.700 1.400 42.980 316.400 ;
      RECT 44.940 1.400 45.220 316.400 ;
      RECT 47.180 1.400 47.460 316.400 ;
      RECT 49.420 1.400 49.700 316.400 ;
      RECT 51.660 1.400 51.940 316.400 ;
      RECT 53.900 1.400 54.180 316.400 ;
      RECT 56.140 1.400 56.420 316.400 ;
      RECT 58.380 1.400 58.660 316.400 ;
      RECT 60.620 1.400 60.900 316.400 ;
      RECT 62.860 1.400 63.140 316.400 ;
      RECT 65.100 1.400 65.380 316.400 ;
      RECT 67.340 1.400 67.620 316.400 ;
      RECT 69.580 1.400 69.860 316.400 ;
      RECT 71.820 1.400 72.100 316.400 ;
      RECT 74.060 1.400 74.340 316.400 ;
      RECT 76.300 1.400 76.580 316.400 ;
      RECT 78.540 1.400 78.820 316.400 ;
      RECT 80.780 1.400 81.060 316.400 ;
      RECT 83.020 1.400 83.300 316.400 ;
      RECT 85.260 1.400 85.540 316.400 ;
      RECT 87.500 1.400 87.780 316.400 ;
      RECT 89.740 1.400 90.020 316.400 ;
      RECT 91.980 1.400 92.260 316.400 ;
      RECT 94.220 1.400 94.500 316.400 ;
      RECT 96.460 1.400 96.740 316.400 ;
      RECT 98.700 1.400 98.980 316.400 ;
      RECT 100.940 1.400 101.220 316.400 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 104.500 317.800 ;
    LAYER metal2 ;
    RECT 0 0 104.500 317.800 ;
    LAYER metal3 ;
    RECT 0.070 0 104.500 317.800 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 4.165 ;
    RECT 0 4.235 0.070 6.965 ;
    RECT 0 7.035 0.070 9.765 ;
    RECT 0 9.835 0.070 12.565 ;
    RECT 0 12.635 0.070 15.365 ;
    RECT 0 15.435 0.070 18.165 ;
    RECT 0 18.235 0.070 20.965 ;
    RECT 0 21.035 0.070 23.765 ;
    RECT 0 23.835 0.070 26.565 ;
    RECT 0 26.635 0.070 29.365 ;
    RECT 0 29.435 0.070 32.165 ;
    RECT 0 32.235 0.070 34.965 ;
    RECT 0 35.035 0.070 37.765 ;
    RECT 0 37.835 0.070 40.565 ;
    RECT 0 40.635 0.070 43.365 ;
    RECT 0 43.435 0.070 46.165 ;
    RECT 0 46.235 0.070 48.965 ;
    RECT 0 49.035 0.070 51.765 ;
    RECT 0 51.835 0.070 54.565 ;
    RECT 0 54.635 0.070 57.365 ;
    RECT 0 57.435 0.070 60.165 ;
    RECT 0 60.235 0.070 62.965 ;
    RECT 0 63.035 0.070 65.765 ;
    RECT 0 65.835 0.070 68.565 ;
    RECT 0 68.635 0.070 71.365 ;
    RECT 0 71.435 0.070 74.165 ;
    RECT 0 74.235 0.070 76.965 ;
    RECT 0 77.035 0.070 79.765 ;
    RECT 0 79.835 0.070 82.565 ;
    RECT 0 82.635 0.070 85.365 ;
    RECT 0 85.435 0.070 88.165 ;
    RECT 0 88.235 0.070 90.545 ;
    RECT 0 90.615 0.070 93.345 ;
    RECT 0 93.415 0.070 96.145 ;
    RECT 0 96.215 0.070 98.945 ;
    RECT 0 99.015 0.070 101.745 ;
    RECT 0 101.815 0.070 104.545 ;
    RECT 0 104.615 0.070 107.345 ;
    RECT 0 107.415 0.070 110.145 ;
    RECT 0 110.215 0.070 112.945 ;
    RECT 0 113.015 0.070 115.745 ;
    RECT 0 115.815 0.070 118.545 ;
    RECT 0 118.615 0.070 121.345 ;
    RECT 0 121.415 0.070 124.145 ;
    RECT 0 124.215 0.070 126.945 ;
    RECT 0 127.015 0.070 129.745 ;
    RECT 0 129.815 0.070 132.545 ;
    RECT 0 132.615 0.070 135.345 ;
    RECT 0 135.415 0.070 138.145 ;
    RECT 0 138.215 0.070 140.945 ;
    RECT 0 141.015 0.070 143.745 ;
    RECT 0 143.815 0.070 146.545 ;
    RECT 0 146.615 0.070 149.345 ;
    RECT 0 149.415 0.070 152.145 ;
    RECT 0 152.215 0.070 154.945 ;
    RECT 0 155.015 0.070 157.745 ;
    RECT 0 157.815 0.070 160.545 ;
    RECT 0 160.615 0.070 163.345 ;
    RECT 0 163.415 0.070 166.145 ;
    RECT 0 166.215 0.070 168.945 ;
    RECT 0 169.015 0.070 171.745 ;
    RECT 0 171.815 0.070 174.545 ;
    RECT 0 174.615 0.070 177.345 ;
    RECT 0 177.415 0.070 179.725 ;
    RECT 0 179.795 0.070 182.525 ;
    RECT 0 182.595 0.070 185.325 ;
    RECT 0 185.395 0.070 188.125 ;
    RECT 0 188.195 0.070 190.925 ;
    RECT 0 190.995 0.070 193.725 ;
    RECT 0 193.795 0.070 196.525 ;
    RECT 0 196.595 0.070 199.325 ;
    RECT 0 199.395 0.070 202.125 ;
    RECT 0 202.195 0.070 204.925 ;
    RECT 0 204.995 0.070 207.725 ;
    RECT 0 207.795 0.070 210.525 ;
    RECT 0 210.595 0.070 213.325 ;
    RECT 0 213.395 0.070 216.125 ;
    RECT 0 216.195 0.070 218.925 ;
    RECT 0 218.995 0.070 221.725 ;
    RECT 0 221.795 0.070 224.525 ;
    RECT 0 224.595 0.070 227.325 ;
    RECT 0 227.395 0.070 230.125 ;
    RECT 0 230.195 0.070 232.925 ;
    RECT 0 232.995 0.070 235.725 ;
    RECT 0 235.795 0.070 238.525 ;
    RECT 0 238.595 0.070 241.325 ;
    RECT 0 241.395 0.070 244.125 ;
    RECT 0 244.195 0.070 246.925 ;
    RECT 0 246.995 0.070 249.725 ;
    RECT 0 249.795 0.070 252.525 ;
    RECT 0 252.595 0.070 255.325 ;
    RECT 0 255.395 0.070 258.125 ;
    RECT 0 258.195 0.070 260.925 ;
    RECT 0 260.995 0.070 263.725 ;
    RECT 0 263.795 0.070 266.525 ;
    RECT 0 266.595 0.070 268.905 ;
    RECT 0 268.975 0.070 271.705 ;
    RECT 0 271.775 0.070 274.505 ;
    RECT 0 274.575 0.070 277.305 ;
    RECT 0 277.375 0.070 280.105 ;
    RECT 0 280.175 0.070 282.905 ;
    RECT 0 282.975 0.070 285.705 ;
    RECT 0 285.775 0.070 288.505 ;
    RECT 0 288.575 0.070 291.305 ;
    RECT 0 291.375 0.070 294.105 ;
    RECT 0 294.175 0.070 296.485 ;
    RECT 0 296.555 0.070 299.285 ;
    RECT 0 299.355 0.070 302.085 ;
    RECT 0 302.155 0.070 317.800 ;
    LAYER metal4 ;
    RECT 0 0 104.500 1.400 ;
    RECT 0 316.400 104.500 317.800 ;
    RECT 0.000 1.400 1.260 316.400 ;
    RECT 1.540 1.400 2.380 316.400 ;
    RECT 2.660 1.400 3.500 316.400 ;
    RECT 3.780 1.400 4.620 316.400 ;
    RECT 4.900 1.400 5.740 316.400 ;
    RECT 6.020 1.400 6.860 316.400 ;
    RECT 7.140 1.400 7.980 316.400 ;
    RECT 8.260 1.400 9.100 316.400 ;
    RECT 9.380 1.400 10.220 316.400 ;
    RECT 10.500 1.400 11.340 316.400 ;
    RECT 11.620 1.400 12.460 316.400 ;
    RECT 12.740 1.400 13.580 316.400 ;
    RECT 13.860 1.400 14.700 316.400 ;
    RECT 14.980 1.400 15.820 316.400 ;
    RECT 16.100 1.400 16.940 316.400 ;
    RECT 17.220 1.400 18.060 316.400 ;
    RECT 18.340 1.400 19.180 316.400 ;
    RECT 19.460 1.400 20.300 316.400 ;
    RECT 20.580 1.400 21.420 316.400 ;
    RECT 21.700 1.400 22.540 316.400 ;
    RECT 22.820 1.400 23.660 316.400 ;
    RECT 23.940 1.400 24.780 316.400 ;
    RECT 25.060 1.400 25.900 316.400 ;
    RECT 26.180 1.400 27.020 316.400 ;
    RECT 27.300 1.400 28.140 316.400 ;
    RECT 28.420 1.400 29.260 316.400 ;
    RECT 29.540 1.400 30.380 316.400 ;
    RECT 30.660 1.400 31.500 316.400 ;
    RECT 31.780 1.400 32.620 316.400 ;
    RECT 32.900 1.400 33.740 316.400 ;
    RECT 34.020 1.400 34.860 316.400 ;
    RECT 35.140 1.400 35.980 316.400 ;
    RECT 36.260 1.400 37.100 316.400 ;
    RECT 37.380 1.400 38.220 316.400 ;
    RECT 38.500 1.400 39.340 316.400 ;
    RECT 39.620 1.400 40.460 316.400 ;
    RECT 40.740 1.400 41.580 316.400 ;
    RECT 41.860 1.400 42.700 316.400 ;
    RECT 42.980 1.400 43.820 316.400 ;
    RECT 44.100 1.400 44.940 316.400 ;
    RECT 45.220 1.400 46.060 316.400 ;
    RECT 46.340 1.400 47.180 316.400 ;
    RECT 47.460 1.400 48.300 316.400 ;
    RECT 48.580 1.400 49.420 316.400 ;
    RECT 49.700 1.400 50.540 316.400 ;
    RECT 50.820 1.400 51.660 316.400 ;
    RECT 51.940 1.400 52.780 316.400 ;
    RECT 53.060 1.400 53.900 316.400 ;
    RECT 54.180 1.400 55.020 316.400 ;
    RECT 55.300 1.400 56.140 316.400 ;
    RECT 56.420 1.400 57.260 316.400 ;
    RECT 57.540 1.400 58.380 316.400 ;
    RECT 58.660 1.400 59.500 316.400 ;
    RECT 59.780 1.400 60.620 316.400 ;
    RECT 60.900 1.400 61.740 316.400 ;
    RECT 62.020 1.400 62.860 316.400 ;
    RECT 63.140 1.400 63.980 316.400 ;
    RECT 64.260 1.400 65.100 316.400 ;
    RECT 65.380 1.400 66.220 316.400 ;
    RECT 66.500 1.400 67.340 316.400 ;
    RECT 67.620 1.400 68.460 316.400 ;
    RECT 68.740 1.400 69.580 316.400 ;
    RECT 69.860 1.400 70.700 316.400 ;
    RECT 70.980 1.400 71.820 316.400 ;
    RECT 72.100 1.400 72.940 316.400 ;
    RECT 73.220 1.400 74.060 316.400 ;
    RECT 74.340 1.400 75.180 316.400 ;
    RECT 75.460 1.400 76.300 316.400 ;
    RECT 76.580 1.400 77.420 316.400 ;
    RECT 77.700 1.400 78.540 316.400 ;
    RECT 78.820 1.400 79.660 316.400 ;
    RECT 79.940 1.400 80.780 316.400 ;
    RECT 81.060 1.400 81.900 316.400 ;
    RECT 82.180 1.400 83.020 316.400 ;
    RECT 83.300 1.400 84.140 316.400 ;
    RECT 84.420 1.400 85.260 316.400 ;
    RECT 85.540 1.400 86.380 316.400 ;
    RECT 86.660 1.400 87.500 316.400 ;
    RECT 87.780 1.400 88.620 316.400 ;
    RECT 88.900 1.400 89.740 316.400 ;
    RECT 90.020 1.400 90.860 316.400 ;
    RECT 91.140 1.400 91.980 316.400 ;
    RECT 92.260 1.400 93.100 316.400 ;
    RECT 93.380 1.400 94.220 316.400 ;
    RECT 94.500 1.400 95.340 316.400 ;
    RECT 95.620 1.400 96.460 316.400 ;
    RECT 96.740 1.400 97.580 316.400 ;
    RECT 97.860 1.400 98.700 316.400 ;
    RECT 98.980 1.400 99.820 316.400 ;
    RECT 100.100 1.400 100.940 316.400 ;
    RECT 101.220 1.400 102.060 316.400 ;
    RECT 102.340 1.400 104.500 316.400 ;
    LAYER OVERLAP ;
    RECT 0 0 104.500 317.800 ;
  END
END fakeram45_1024x32

END LIBRARY
