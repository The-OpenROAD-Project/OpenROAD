module top (clk,
    in1,
    in10,
    in2,
    in3,
    in4,
    in5,
    in6,
    in7,
    in8,
    in9,
    out2,
    out3,
    out4,
    out5,
    out1);
 input clk;
 input in1;
 input in10;
 input in2;
 input in3;
 input in4;
 input in5;
 input in6;
 input in7;
 input in8;
 input in9;
 output out2;
 output out3;
 output out4;
 output out5;
 output out1;

 wire sub1_out2;
 wire sub1_out1;
 wire n1;
 wire n2;
 wire n3;
 wire n4;
 wire n5;
 wire n6;
 wire reg1_q;
 wire reg2_q;

 AND2_X1 and1 (.A1(in6),
    .A2(in7),
    .ZN(n1));
 AOI21_X1 aoi1 (.A(n1),
    .B1(n2),
    .B2(sub1_out2),
    .ZN(out5));
 BUF_X1 b1 (.A(n5),
    .Z(n6));
 NAND2_X1 nand1 (.A1(sub1_out1),
    .A2(n3),
    .ZN(n4));
 NOR2_X1 nor1 (.A1(sub1_out2),
    .A2(in10),
    .ZN(n5));
 OR2_X1 or1 (.A1(in8),
    .A2(in9),
    .ZN(n2));
 DFF_X1 reg1 (.D(in1),
    .Q(reg1_q));
 DFF_X1 reg2 (.D(n3),
    .Q(reg2_q));
 XOR2_X1 xor1 (.A(reg1_q),
    .B(sub1_out1),
    .Z(n3));
 sub_module1 sub1_inst (.sub1_in1(in1),
    .sub1_in2(in2),
    .sub1_in3(in3),
    .sub1_in4(in4),
    .sub1_in5(in5),
    .sub1_out1(sub1_out1),
    .sub1_out2(sub1_out2));
 assign out2 = n4;
 assign out3 = n5;
 assign out4 = n6;
 assign out1 = reg2_q;
endmodule
module sub_module1 (sub1_in1,
    sub1_in2,
    sub1_in3,
    sub1_in4,
    sub1_in5,
    sub1_out1,
    sub1_out2);
 input sub1_in1;
 input sub1_in2;
 input sub1_in3;
 input sub1_in4;
 input sub1_in5;
 output sub1_out1;
 output sub1_out2;

 wire sub2_out2;
 wire sub2_out1;
 wire w1;
 wire w2;
 wire w3;

 BUF_X2 b1 (.A(sub1_in1),
    .Z(w1));
 BUF_X4 b2 (.A(sub1_in2),
    .Z(w2));
 BUF_X8 b3 (.A(w2),
    .Z(w3));
 OAI21_X1 oai_inst (.B1(w1),
    .ZN(sub1_out1));
 XNOR2_X1 xnor_inst (.A(sub2_out2),
    .B(sub1_in5),
    .ZN(sub1_out2));
 sub_module2 sub2_inst (.sub2_in1(sub1_in1),
    .sub2_in2(sub1_in2),
    .sub2_in3(sub1_in3),
    .sub2_in4(sub1_in4),
    .sub2_out1(sub2_out1),
    .sub2_out2(sub2_out2));
endmodule
module sub_module2 (sub2_in1,
    sub2_in2,
    sub2_in3,
    sub2_in4,
    sub2_out1,
    sub2_out2);
 input sub2_in1;
 input sub2_in2;
 input sub2_in3;
 input sub2_in4;
 output sub2_out1;
 output sub2_out2;

 wire w1;

 AND2_X1 and_inst (.A1(sub2_in1),
    .A2(sub2_in2),
    .ZN(w1));
 NOR2_X1 nor_inst (.A1(sub2_in3),
    .A2(sub2_in4),
    .ZN(sub2_out2));
 XOR2_X1 xor_inst (.A(w1),
    .B(sub2_in3),
    .Z(sub2_out1));
endmodule
