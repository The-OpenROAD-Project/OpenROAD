module io_constraints1 ( \io_1 , \io_2 , \io_3 );
  HM_100x100_1x1 MACRO_1 ( ) ;

  DFF_X1 _001_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _002_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _003_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _004_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _005_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _006_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _007_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _008_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _009_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _010_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _011_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _012_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _013_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _014_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _015_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _016_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _017_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _018_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _019_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _020_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _021_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _022_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _023_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _024_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _025_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _026_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _027_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _028_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _029_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _030_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _031_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _032_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _033_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _034_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _035_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _036_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _037_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _038_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _039_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _040_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _041_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _042_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _043_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _044_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _045_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _046_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _047_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _048_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _049_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _050_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _051_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _052_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _053_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _054_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _055_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _056_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _057_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _058_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _059_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _060_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _061_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _062_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _063_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _064_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _065_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _066_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _067_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _068_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _069_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _070_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _071_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _072_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _073_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _074_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _075_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _076_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _077_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _078_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _079_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _080_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _081_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _082_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _083_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _084_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _085_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _086_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _087_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _088_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _089_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _090_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _091_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _092_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _093_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _094_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _095_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _096_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _097_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _098_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _099_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _100_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _101_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _102_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _103_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _104_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _105_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _106_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _107_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _108_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _109_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _110_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _111_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _112_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _113_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _114_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _115_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _116_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _117_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _118_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _119_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _120_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _121_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _122_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _123_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _124_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _125_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _126_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _127_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _128_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _129_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _130_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _131_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _132_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _133_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _134_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _135_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _136_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _137_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _138_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _139_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _140_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _141_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _142_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _143_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _144_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _145_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _146_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _147_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _148_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _149_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _150_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _151_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _152_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _153_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _154_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _155_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _156_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _157_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _158_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _159_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _160_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _161_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _162_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _163_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _164_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _165_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _166_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _167_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _168_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _169_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _170_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _171_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _172_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _173_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _174_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _175_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _176_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _177_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _178_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _179_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _180_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _181_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _182_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _183_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _184_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _185_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _186_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _187_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _188_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _189_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _190_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _191_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _192_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _193_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _194_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _195_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _196_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _197_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _198_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _199_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _200_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _201_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _202_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _203_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _204_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _205_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _206_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _207_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _208_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _209_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _210_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _211_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _212_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _213_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _214_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _215_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _216_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _217_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _218_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _219_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _220_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _221_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _222_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _223_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _224_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _225_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _226_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _227_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _228_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _229_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _230_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _231_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _232_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _233_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _234_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _235_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _236_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _237_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _238_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _239_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _240_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _241_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _242_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _243_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _244_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _245_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _246_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _247_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _248_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _249_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _250_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _251_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _252_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _253_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _254_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _255_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _256_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _257_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _258_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _259_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _260_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _261_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _262_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _263_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _264_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _265_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _266_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _267_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _268_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _269_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _270_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _271_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _272_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _273_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _274_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _275_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _276_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _277_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _278_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _279_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _280_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _281_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _282_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _283_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _284_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _285_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _286_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _287_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _288_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _289_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _290_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _291_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _292_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _293_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _294_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _295_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _296_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _297_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _298_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _299_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _300_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _301_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _302_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _303_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _304_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _305_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _306_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _307_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _308_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _309_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _310_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _311_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _312_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _313_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _314_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _315_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _316_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _317_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _318_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _319_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _320_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _321_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _322_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _323_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _324_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _325_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _326_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _327_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _328_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _329_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _330_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _331_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _332_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _333_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _334_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _335_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _336_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _337_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _338_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _339_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _340_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _341_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _342_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _343_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _344_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _345_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _346_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _347_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _348_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _349_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _350_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _351_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _352_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _353_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _354_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _355_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _356_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _357_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _358_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _359_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _360_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _361_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _362_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _363_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _364_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _365_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _366_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _367_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _368_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _369_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _370_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _371_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _372_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _373_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _374_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _375_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _376_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _377_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _378_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _379_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _380_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _381_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _382_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _383_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _384_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _385_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _386_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _387_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _388_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _389_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _390_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _391_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _392_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _393_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _394_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _395_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _396_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _397_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _398_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _399_ ( .CK(), .D(), .Q(), .QN() );
  DFF_X1 _400_ ( .CK(), .D(), .Q(), .QN() );

  input io_1;
  input io_2;
  input io_3;
endmodule
