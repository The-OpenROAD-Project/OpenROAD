VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO h7
   CLASS BLOCK ;
   SIZE 344 BY 54 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   PIN FE_OFN1038_g64577_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 3.65 53.49 3.75 54 ;
      END
   END FE_OFN1038_g64577_p

   PIN FE_OFN1047_g64577_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 15.25 53.49 15.35 54 ;
      END
   END FE_OFN1047_g64577_p

   PIN FE_OFN1052_g64577_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 33.975 0.255 34.175 ;
      END
   END FE_OFN1052_g64577_p

   PIN FE_OFN1057_g64577_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 17.65 53.49 17.75 54 ;
      END
   END FE_OFN1057_g64577_p

   PIN FE_OFN1058_g64577_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 5.45 53.49 5.55 54 ;
      END
   END FE_OFN1058_g64577_p

   PIN g62724_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 32.625 0.51 32.725 ;
      END
   END g62724_db

   PIN g62724_sb
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 34.825 0.51 34.925 ;
      END
   END g62724_sb

   PIN g62776_sb
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 8.05 53.49 8.15 54 ;
      END
   END g62776_sb

   PIN g62799_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 2.05 53.49 2.15 54 ;
      END
   END g62799_db

   PIN g62805_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 5.65 53.49 5.75 54 ;
      END
   END g62805_da

   PIN g62806_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 30.45 53.49 30.55 54 ;
      END
   END g62806_da

   PIN g62813_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 3.05 53.49 3.15 54 ;
      END
   END g62813_db

   PIN g62817_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 1.85 53.49 1.95 54 ;
      END
   END g62817_da

   PIN g62826_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 24.225 0.51 24.325 ;
      END
   END g62826_db

   PIN g63015_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 24.45 53.49 24.55 54 ;
      END
   END g63015_da

   PIN g63072_sb
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 8.25 53.49 8.35 54 ;
      END
   END g63072_sb

   PIN g63105_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 3.85 53.49 3.95 54 ;
      END
   END g63105_db

   PIN g64152_sb
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 45.025 0.51 45.125 ;
      END
   END g64152_sb

   PIN g64158_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 30.625 0.51 30.725 ;
      END
   END g64158_da

   PIN g64184_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 42.025 0.51 42.125 ;
      END
   END g64184_da

   PIN g64211_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 3.25 53.49 3.35 54 ;
      END
   END g64211_db

   PIN g64235_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 44.025 0.51 44.125 ;
      END
   END g64235_da

   PIN g64235_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 45.225 0.51 45.325 ;
      END
   END g64235_db

   PIN g64273_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 14.85 53.49 14.95 54 ;
      END
   END g64273_da

   PIN g64273_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 15.45 53.49 15.55 54 ;
      END
   END g64273_db

   PIN g64313_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 7.05 53.49 7.15 54 ;
      END
   END g64313_da

   PIN g64313_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 45.425 0.51 45.525 ;
      END
   END g64313_db

   PIN n_14060
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 42.625 0.51 42.725 ;
      END
   END n_14060

   PIN n_14091
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 45.625 0.51 45.725 ;
      END
   END n_14091

   PIN n_14092
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 3.45 53.49 3.55 54 ;
      END
   END n_14092

   PIN n_14216
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 38.225 0.51 38.325 ;
      END
   END n_14216

   PIN n_14596
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 45.825 0.51 45.925 ;
      END
   END n_14596

   PIN n_14603
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 27.45 53.49 27.55 54 ;
      END
   END n_14603

   PIN n_14608
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 22.05 53.49 22.15 54 ;
      END
   END n_14608

   PIN n_14610
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 26.25 53.49 26.35 54 ;
      END
   END n_14610

   PIN n_14611
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 32.825 0.51 32.925 ;
      END
   END n_14611

   PIN n_16247
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 21.85 53.49 21.95 54 ;
      END
   END n_16247

   PIN n_16252
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 21.65 53.49 21.75 54 ;
      END
   END n_16252

   PIN n_3825
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 6.45 53.49 6.55 54 ;
      END
   END n_3825

   PIN n_3938
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 19.45 53.49 19.55 54 ;
      END
   END n_3938

   PIN n_3977
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 26.425 0.51 26.525 ;
      END
   END n_3977

   PIN n_3983
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 46.025 0.51 46.125 ;
      END
   END n_3983

   PIN n_4010
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 47.025 0.51 47.125 ;
      END
   END n_4010

   PIN n_4077
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 35.025 0.51 35.125 ;
      END
   END n_4077

   PIN n_5012
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 4.65 53.49 4.75 54 ;
      END
   END n_5012

   PIN n_5136
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 23.45 53.49 23.55 54 ;
      END
   END n_5136

   PIN n_5376
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 46.225 0.51 46.325 ;
      END
   END n_5376

   PIN pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__28__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 15.85 53.49 15.95 54 ;
      END
   END pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__28__Q

   PIN pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__28__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 8.45 53.49 8.55 54 ;
      END
   END pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__28__Q

   PIN pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__15__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 5.05 53.49 5.15 54 ;
      END
   END pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__15__Q

   PIN pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__18__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 43.825 0.51 43.925 ;
      END
   END pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__18__Q

   PIN pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__15__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 40.225 0.51 40.325 ;
      END
   END pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__15__Q

   PIN pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_51
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 99.05 53.49 99.15 54 ;
      END
   END pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_51

   PIN pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_63
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 73.85 53.49 73.95 54 ;
      END
   END pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_63

   PIN FE_OCP_RBN2037_FE_OCPN2000_n_13743
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 15.65 53.49 15.75 54 ;
      END
   END FE_OCP_RBN2037_FE_OCPN2000_n_13743

   PIN FE_OCP_RBN2086_FE_OFN1756_n_13997
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 32.6 53.745 32.8 54 ;
      END
   END FE_OCP_RBN2086_FE_OFN1756_n_13997

   PIN FE_OFN1015_g64577_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 11.45 53.49 11.55 54 ;
      END
   END FE_OFN1015_g64577_p

   PIN FE_OFN1027_g64577_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 37.775 0.255 37.975 ;
      END
   END FE_OFN1027_g64577_p

   PIN FE_OFN1034_g64577_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 11.2 53.745 11.4 54 ;
      END
   END FE_OFN1034_g64577_p

   PIN FE_OFN1043_g64577_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 33.65 53.49 33.75 54 ;
      END
   END FE_OFN1043_g64577_p

   PIN FE_OFN1046_g64577_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 34.2 53.745 34.4 54 ;
      END
   END FE_OFN1046_g64577_p

   PIN FE_OFN1054_g64577_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 32.2 53.745 32.4 54 ;
      END
   END FE_OFN1054_g64577_p

   PIN FE_OFN1464_n_13736
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 39.775 0.255 39.975 ;
      END
   END FE_OFN1464_n_13736

   PIN FE_OFN1465_n_13736
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 23.05 53.49 23.15 54 ;
      END
   END FE_OFN1465_n_13736

   PIN FE_OFN1466_n_13736
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 43.4 53.745 43.6 54 ;
      END
   END FE_OFN1466_n_13736

   PIN FE_OFN1469_n_13741
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 34.625 0.51 34.725 ;
      END
   END FE_OFN1469_n_13741

   PIN FE_OFN1470_n_13741
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 28.25 53.49 28.35 54 ;
      END
   END FE_OFN1470_n_13741

   PIN FE_OFN1471_n_13741
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 4.05 53.49 4.15 54 ;
      END
   END FE_OFN1471_n_13741

   PIN FE_OFN1478_n_13995
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 24.05 53.49 24.15 54 ;
      END
   END FE_OFN1478_n_13995

   PIN FE_OFN1479_n_13995
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 7.85 53.49 7.95 54 ;
      END
   END FE_OFN1479_n_13995

   PIN FE_OFN1522_n_4730
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 15.8 53.745 16 54 ;
      END
   END FE_OFN1522_n_4730

   PIN FE_OFN1523_n_4730
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 35.4 53.745 35.6 54 ;
      END
   END FE_OFN1523_n_4730

   PIN FE_OFN1524_n_4730
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 33.175 0.255 33.375 ;
      END
   END FE_OFN1524_n_4730

   PIN FE_OFN1557_n_4732
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 38.575 0.255 38.775 ;
      END
   END FE_OFN1557_n_4732

   PIN FE_OFN1558_n_4732
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 33.4 53.745 33.6 54 ;
      END
   END FE_OFN1558_n_4732

   PIN FE_OFN1559_n_4732
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 7.65 53.49 7.75 54 ;
      END
   END FE_OFN1559_n_4732

   PIN FE_OFN1581_n_16657
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 41.575 0.255 41.775 ;
      END
   END FE_OFN1581_n_16657

   PIN FE_OFN1583_n_16657
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 31.8 53.745 32 54 ;
      END
   END FE_OFN1583_n_16657

   PIN FE_OFN1584_n_16657
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 39.375 0.255 39.575 ;
      END
   END FE_OFN1584_n_16657

   PIN FE_OFN1612_n_4740
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 40.575 0.255 40.775 ;
      END
   END FE_OFN1612_n_4740

   PIN FE_OFN1613_n_4740
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 5.25 53.49 5.35 54 ;
      END
   END FE_OFN1613_n_4740

   PIN FE_OFN1614_n_4740
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 6.25 53.49 6.35 54 ;
      END
   END FE_OFN1614_n_4740

   PIN FE_OFN1757_n_13997
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 7.25 53.49 7.35 54 ;
      END
   END FE_OFN1757_n_13997

   PIN FE_OFN1761_n_14054
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 4.25 53.49 4.35 54 ;
      END
   END FE_OFN1761_n_14054

   PIN FE_OFN1762_n_14054
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 42.975 0.255 43.175 ;
      END
   END FE_OFN1762_n_14054

   PIN FE_OFN1764_n_14054
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 12.05 53.49 12.15 54 ;
      END
   END FE_OFN1764_n_14054

   PIN FE_OFN1770_n_13800
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 8.85 53.49 8.95 54 ;
      END
   END FE_OFN1770_n_13800

   PIN FE_OFN1771_n_13800
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 11.65 53.49 11.75 54 ;
      END
   END FE_OFN1771_n_13800

   PIN FE_OFN1772_n_13800
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 31.625 0.51 31.725 ;
      END
   END FE_OFN1772_n_13800

   PIN FE_OFN1776_n_13971
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 33.8 53.745 34 54 ;
      END
   END FE_OFN1776_n_13971

   PIN FE_OFN1777_n_13971
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 32.45 53.49 32.55 54 ;
      END
   END FE_OFN1777_n_13971

   PIN FE_OFN854_n_4736
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 15.05 53.49 15.15 54 ;
      END
   END FE_OFN854_n_4736

   PIN FE_OFN855_n_4736
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 33 53.745 33.2 54 ;
      END
   END FE_OFN855_n_4736

   PIN FE_OFN859_n_4734
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 6.85 53.49 6.95 54 ;
      END
   END FE_OFN859_n_4734

   PIN FE_OFN860_n_4734
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 38.975 0.255 39.175 ;
      END
   END FE_OFN860_n_4734

   PIN FE_OFN868_n_4725
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 28.175 0.255 28.375 ;
      END
   END FE_OFN868_n_4725

   PIN FE_OFN951_n_4725
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 31.05 53.49 31.15 54 ;
      END
   END FE_OFN951_n_4725

   PIN FE_OFN952_n_4725
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 37.375 0.255 37.575 ;
      END
   END FE_OFN952_n_4725

   PIN FE_OFN975_n_4727
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 24.2 53.745 24.4 54 ;
      END
   END FE_OFN975_n_4727

   PIN FE_OFN976_n_4727
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 43 53.745 43.2 54 ;
      END
   END FE_OFN976_n_4727

   PIN g62803_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 2.85 53.49 2.95 54 ;
      END
   END g62803_da

   PIN g62805_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 6.05 53.49 6.15 54 ;
      END
   END g62805_sb

   PIN g62862_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 4.45 53.49 4.55 54 ;
      END
   END g62862_sb

   PIN g63015_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 24.85 53.49 24.95 54 ;
      END
   END g63015_sb

   PIN g63057_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 22.85 53.49 22.95 54 ;
      END
   END g63057_sb

   PIN g63058_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 16.45 53.49 16.55 54 ;
      END
   END g63058_da

   PIN g63072_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 44.825 0.51 44.925 ;
      END
   END g63072_da

   PIN g63122_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 4.85 53.49 4.95 54 ;
      END
   END g63122_da

   PIN g64078_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 34.425 0.51 34.525 ;
      END
   END g64078_da

   PIN g64158_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 30.425 0.51 30.525 ;
      END
   END g64158_sb

   PIN g64217_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 30.05 53.49 30.15 54 ;
      END
   END g64217_db

   PIN g64217_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 29.25 53.49 29.35 54 ;
      END
   END g64217_sb

   PIN g64296_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 26.225 0.51 26.325 ;
      END
   END g64296_db

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 43.375 0.255 43.575 ;
      END
   END ispd_clk

   PIN n_13891
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 44.625 0.51 44.725 ;
      END
   END n_13891

   PIN n_13901
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 31.175 0.255 31.375 ;
      END
   END n_13901

   PIN n_13987
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 26.85 53.49 26.95 54 ;
      END
   END n_13987

   PIN n_13993
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 19.05 53.49 19.15 54 ;
      END
   END n_13993

   PIN n_14001
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 13.65 53.49 13.75 54 ;
      END
   END n_14001

   PIN n_14458
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 27.25 53.49 27.35 54 ;
      END
   END n_14458

   PIN n_14472
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 11.85 53.49 11.95 54 ;
      END
   END n_14472

   PIN n_14594
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 100.05 53.49 100.15 54 ;
      END
   END n_14594

   PIN n_14956
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 32.425 0.51 32.525 ;
      END
   END n_14956

   PIN n_16244
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 22.65 53.49 22.75 54 ;
      END
   END n_16244

   PIN n_16621
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 27.65 53.49 27.75 54 ;
      END
   END n_16621

   PIN n_3923
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 14.65 53.49 14.75 54 ;
      END
   END n_3923

   PIN n_3958
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 2.25 53.49 2.35 54 ;
      END
   END n_3958

   PIN n_4013
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 44.425 0.51 44.525 ;
      END
   END n_4013

   PIN n_5351
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 41.025 0.51 41.125 ;
      END
   END n_5351

   PIN n_5371
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 7.45 53.49 7.55 54 ;
      END
   END n_5371

   PIN n_5388
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 42.425 0.51 42.525 ;
      END
   END n_5388

   PIN pci_target_unit_fifos_pciw_addr_data_in_128
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 6.65 53.49 6.75 54 ;
      END
   END pci_target_unit_fifos_pciw_addr_data_in_128

   PIN pci_target_unit_fifos_pciw_addr_data_in_132
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 30.825 0.51 30.925 ;
      END
   END pci_target_unit_fifos_pciw_addr_data_in_132

   PIN pci_target_unit_fifos_pciw_addr_data_in_133
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 32.85 53.49 32.95 54 ;
      END
   END pci_target_unit_fifos_pciw_addr_data_in_133

   PIN pci_target_unit_fifos_pciw_addr_data_in_134
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 12.25 53.49 12.35 54 ;
      END
   END pci_target_unit_fifos_pciw_addr_data_in_134

   PIN pci_target_unit_fifos_pciw_addr_data_in_135
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 35.25 53.49 35.35 54 ;
      END
   END pci_target_unit_fifos_pciw_addr_data_in_135

   PIN pci_target_unit_fifos_pciw_addr_data_in_136
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 16.85 53.49 16.95 54 ;
      END
   END pci_target_unit_fifos_pciw_addr_data_in_136

   PIN pci_target_unit_fifos_pciw_addr_data_in_138
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 26.65 53.49 26.75 54 ;
      END
   END pci_target_unit_fifos_pciw_addr_data_in_138

   PIN pci_target_unit_fifos_pciw_addr_data_in_141
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 32.25 53.49 32.35 54 ;
      END
   END pci_target_unit_fifos_pciw_addr_data_in_141

   PIN pci_target_unit_fifos_pciw_addr_data_in_142
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 41.225 0.51 41.325 ;
      END
   END pci_target_unit_fifos_pciw_addr_data_in_142

   PIN pci_target_unit_fifos_pciw_addr_data_in_148
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 14.45 53.49 14.55 54 ;
      END
   END pci_target_unit_fifos_pciw_addr_data_in_148

   PIN pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__13__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 24.25 53.49 24.35 54 ;
      END
   END pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__13__Q

   PIN pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__16__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 21.45 53.49 21.55 54 ;
      END
   END pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__16__Q

   PIN pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__13__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 23.25 53.49 23.35 54 ;
      END
   END pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__13__Q

   PIN pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__22__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 5.85 53.49 5.95 54 ;
      END
   END pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__22__Q

   PIN pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__8__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 46.825 0.51 46.925 ;
      END
   END pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__8__Q

   PIN pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__8__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 46.625 0.51 46.725 ;
      END
   END pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__8__Q

   PIN pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__12__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 30.225 0.51 30.325 ;
      END
   END pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__12__Q

   PIN pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__17__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 2.45 53.49 2.55 54 ;
      END
   END pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__17__Q

   PIN pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__28__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 44.225 0.51 44.325 ;
      END
   END pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__28__Q

   PIN pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__14__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 5.05 53.49 5.15 54 ;
      END
   END pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__14__Q

   PIN pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__21__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 28.45 53.49 28.55 54 ;
      END
   END pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__21__Q

   PIN pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__28__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 46.425 0.51 46.525 ;
      END
   END pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__28__Q

   PIN pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__13__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 33.625 0.51 33.725 ;
      END
   END pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__13__Q

   PIN pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__22__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 2.65 53.49 2.75 54 ;
      END
   END pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__22__Q

   PIN pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__12__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 29.225 0.51 29.325 ;
      END
   END pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__12__Q

   PIN pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__13__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 32.225 0.51 32.325 ;
      END
   END pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__13__Q

   PIN pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__15__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 42.225 0.51 42.325 ;
      END
   END pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__15__Q

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 344 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 344 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 344 8.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 11.745 344 12.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 15.745 344 16.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 19.745 344 20.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 23.745 344 24.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 27.745 344 28.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 31.745 344 32.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 35.745 344 36.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 39.745 344 40.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 43.745 344 44.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 47.745 344 48.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 51.745 344 52.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 344 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 344 6.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 9.745 344 10.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 13.745 344 14.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 17.745 344 18.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 21.745 344 22.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 25.745 344 26.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 29.745 344 30.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 33.745 344 34.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 37.745 344 38.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 41.745 344 42.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 45.745 344 46.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 49.745 344 50.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 53.745 344 54.255 ;
      END
   END vdd

   OBS
      LAYER metal1 ;
         RECT 0 0 344 54 ;
   END
   OBS
      LAYER metal2 ;
         RECT 0 0 344 54 ;
   END
   OBS
      LAYER metal3 ;
         RECT 0 0 344 54 ;
   END
   OBS
      LAYER metal4 ;
         RECT 0 0 344 54 ;
   END
   OBS
      LAYER metal5 ;
         RECT 0 0 344 54 ;
   END
END h7

MACRO h8
   CLASS BLOCK ;
   SIZE 358.4 BY 50 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   PIN FE_OCP_RBN2089_FE_OFN1433_n_12042
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 26.9 0.51 27 ;
      END
   END FE_OCP_RBN2089_FE_OFN1433_n_12042

   PIN FE_OCP_RBN2094_FE_OCPN1856_n_12030
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 20.05 49.49 20.15 50 ;
      END
   END FE_OCP_RBN2094_FE_OCPN1856_n_12030

   PIN FE_OFN1124_n_6935
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 19.45 49.49 19.55 50 ;
      END
   END FE_OFN1124_n_6935

   PIN FE_OFN1204_n_4097
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 54 49.745 54.2 50 ;
      END
   END FE_OFN1204_n_4097

   PIN FE_OFN1205_n_4097
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 24.85 49.49 24.95 50 ;
      END
   END FE_OFN1205_n_4097

   PIN FE_OFN1206_n_4097
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 35.4 49.745 35.6 50 ;
      END
   END FE_OFN1206_n_4097

   PIN FE_OFN1207_n_4097
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 36.85 0.255 37.05 ;
      END
   END FE_OFN1207_n_4097

   PIN FE_OFN1238_n_6436
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 23.45 49.49 23.55 50 ;
      END
   END FE_OFN1238_n_6436

   PIN FE_OFN1450_n_10780
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 14.25 49.49 14.35 50 ;
      END
   END FE_OFN1450_n_10780

   PIN FE_OFN1723_n_16317
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 25.5 0.51 25.6 ;
      END
   END FE_OFN1723_n_16317

   PIN FE_OFN647_n_4460
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 32.05 49.49 32.15 50 ;
      END
   END FE_OFN647_n_4460

   PIN FE_OFN652_n_4417
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 29.2 0 29.4 0.255 ;
      END
   END FE_OFN652_n_4417

   PIN FE_OFN658_n_4438
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 22.25 49.49 22.35 50 ;
      END
   END FE_OFN658_n_4438

   PIN FE_RN_199_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 17.25 0 17.35 0.51 ;
      END
   END FE_RN_199_0

   PIN FE_RN_216_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 21.65 49.49 21.75 50 ;
      END
   END FE_RN_216_0

   PIN g54587_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 26.05 49.49 26.15 50 ;
      END
   END g54587_p

   PIN g62336_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 19.25 49.49 19.35 50 ;
      END
   END g62336_da

   PIN g62386_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 16.65 49.49 16.75 50 ;
      END
   END g62386_db

   PIN g62426_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 23.25 49.49 23.35 50 ;
      END
   END g62426_db

   PIN g62540_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 21.85 49.49 21.95 50 ;
      END
   END g62540_db

   PIN g62582_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 26.1 0.51 26.2 ;
      END
   END g62582_da

   PIN g62675_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 22.45 49.49 22.55 50 ;
      END
   END g62675_da

   PIN g62685_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 49.05 49.49 49.15 50 ;
      END
   END g62685_da

   PIN g62980_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 70.45 49.49 70.55 50 ;
      END
   END g62980_da

   PIN g62980_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 71.25 49.49 71.35 50 ;
      END
   END g62980_db

   PIN g64765_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 18.65 49.49 18.75 50 ;
      END
   END g64765_db

   PIN g64908_sb
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 27.85 49.49 27.95 50 ;
      END
   END g64908_sb

   PIN g64949_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 28.1 0.51 28.2 ;
      END
   END g64949_da

   PIN g64974_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 14.85 49.49 14.95 50 ;
      END
   END g64974_db

   PIN g64993_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 21.7 0.51 21.8 ;
      END
   END g64993_db

   PIN g65004_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 31.1 0.51 31.2 ;
      END
   END g65004_db

   PIN g65047_sb
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 18.85 49.49 18.95 50 ;
      END
   END g65047_sb

   PIN g65328_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 15.25 49.49 15.35 50 ;
      END
   END g65328_db

   PIN g65394_sb
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 72.85 49.49 72.95 50 ;
      END
   END g65394_sb

   PIN n_11898
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 16.85 49.49 16.95 50 ;
      END
   END n_11898

   PIN n_11899
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 15.65 49.49 15.75 50 ;
      END
   END n_11899

   PIN n_11988
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 26.3 0.51 26.4 ;
      END
   END n_11988

   PIN n_12002
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 28.3 0.51 28.4 ;
      END
   END n_12002

   PIN n_12011
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 30.9 0.51 31 ;
      END
   END n_12011

   PIN n_12041
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 60.05 49.49 60.15 50 ;
      END
   END n_12041

   PIN n_12049
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 70.85 49.49 70.95 50 ;
      END
   END n_12049

   PIN n_12052
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 27.45 49.49 27.55 50 ;
      END
   END n_12052

   PIN n_12089
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 31.5 0.51 31.6 ;
      END
   END n_12089

   PIN n_12102
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 48.05 49.49 48.15 50 ;
      END
   END n_12102

   PIN n_12118
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 56.25 49.49 56.35 50 ;
      END
   END n_12118

   PIN n_12196
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 24.25 49.49 24.35 50 ;
      END
   END n_12196

   PIN n_12351
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 15.85 49.49 15.95 50 ;
      END
   END n_12351

   PIN n_12406
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 29.7 0.51 29.8 ;
      END
   END n_12406

   PIN n_12427
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 43.85 49.49 43.95 50 ;
      END
   END n_12427

   PIN n_12449
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 30.7 0.51 30.8 ;
      END
   END n_12449

   PIN n_12459
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 26.5 0.51 26.6 ;
      END
   END n_12459

   PIN n_12473
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 14.65 49.49 14.75 50 ;
      END
   END n_12473

   PIN n_12483
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 40.05 49.49 40.15 50 ;
      END
   END n_12483

   PIN n_12492
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 28.5 0.51 28.6 ;
      END
   END n_12492

   PIN n_12746
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 38.05 49.49 38.15 50 ;
      END
   END n_12746

   PIN n_12749
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 65.25 49.49 65.35 50 ;
      END
   END n_12749

   PIN n_12817
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 47.85 49.49 47.95 50 ;
      END
   END n_12817

   PIN n_12886
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 30.5 0.51 30.6 ;
      END
   END n_12886

   PIN n_12934
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 48.25 49.49 48.35 50 ;
      END
   END n_12934

   PIN n_13128
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 26.7 0.51 26.8 ;
      END
   END n_13128

   PIN n_13139
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 17.05 49.49 17.15 50 ;
      END
   END n_13139

   PIN n_14311
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 28.05 49.49 28.15 50 ;
      END
   END n_14311

   PIN n_14314
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 28.65 49.49 28.75 50 ;
      END
   END n_14314

   PIN n_14381
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 25.45 49.49 25.55 50 ;
      END
   END n_14381

   PIN n_16409
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 62.25 49.49 62.35 50 ;
      END
   END n_16409

   PIN n_3744
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 38.6 49.745 38.8 50 ;
      END
   END n_3744

   PIN n_3749
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 20.85 49.49 20.95 50 ;
      END
   END n_3749

   PIN n_3761
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 23.65 49.49 23.75 50 ;
      END
   END n_3761

   PIN n_4473
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 17.25 49.49 17.35 50 ;
      END
   END n_4473

   PIN n_4478
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 32.45 49.49 32.55 50 ;
      END
   END n_4478

   PIN n_5975
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 16.05 49.49 16.15 50 ;
      END
   END n_5975

   PIN n_6231
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 27.85 0 27.95 0.51 ;
      END
   END n_6231

   PIN n_6348
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 20.45 49.49 20.55 50 ;
      END
   END n_6348

   PIN n_6935
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 23.85 49.49 23.95 50 ;
      END
   END n_6935

   PIN parchk_pci_ad_out_in_1179
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 36.25 49.49 36.35 50 ;
      END
   END parchk_pci_ad_out_in_1179

   PIN parchk_pci_ad_out_in_1181
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 25.25 49.49 25.35 50 ;
      END
   END parchk_pci_ad_out_in_1181

   PIN parchk_pci_ad_out_in_1182
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 39.05 49.49 39.15 50 ;
      END
   END parchk_pci_ad_out_in_1182

   PIN wbs_wbb3_2_wbb2_dat_o_i_105
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 14.85 0 14.95 0.51 ;
      END
   END wbs_wbb3_2_wbb2_dat_o_i_105

   PIN wbs_wbb3_2_wbb2_dat_o_i_116
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 18.85 0 18.95 0.51 ;
      END
   END wbs_wbb3_2_wbb2_dat_o_i_116

   PIN wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__18__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 22.65 49.49 22.75 50 ;
      END
   END wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__18__Q

   PIN wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__37__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 35.05 49.49 35.15 50 ;
      END
   END wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__37__Q

   PIN wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__11__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 62.85 49.49 62.95 50 ;
      END
   END wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__11__Q

   PIN wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__26__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 29.25 49.49 29.35 50 ;
      END
   END wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__26__Q

   PIN wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__12__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 19.05 49.49 19.15 50 ;
      END
   END wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__12__Q

   PIN wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__6__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 14.45 49.49 14.55 50 ;
      END
   END wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__6__Q

   PIN wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__25__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 20.45 49.49 20.55 50 ;
      END
   END wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__25__Q

   PIN wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__26__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 34.85 49.49 34.95 50 ;
      END
   END wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__26__Q

   PIN wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__28__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 31.7 0.51 31.8 ;
      END
   END wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__28__Q

   PIN wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__28__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 19.9 0.51 20 ;
      END
   END wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__28__Q

   PIN wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__24__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 30.65 49.49 30.75 50 ;
      END
   END wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__24__Q

   PIN wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__5__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 45.45 49.49 45.55 50 ;
      END
   END wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__5__Q

   PIN wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__8__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 23.5 0.51 23.6 ;
      END
   END wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__8__Q

   PIN wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__11__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 40.25 49.49 40.35 50 ;
      END
   END wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__11__Q

   PIN FE_OCPN1856_n_12030
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 20.65 49.49 20.75 50 ;
      END
   END FE_OCPN1856_n_12030

   PIN FE_OCPN1857_n_12030
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 29.3 0.51 29.4 ;
      END
   END FE_OCPN1857_n_12030

   PIN FE_OCPN1885_FE_OFN1454_n_12028
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 64.4 49.745 64.6 50 ;
      END
   END FE_OCPN1885_FE_OFN1454_n_12028

   PIN FE_OFN1120_n_6935
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 69.6 49.745 69.8 50 ;
      END
   END FE_OFN1120_n_6935

   PIN FE_OFN1127_n_4090
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 24.05 49.49 24.15 50 ;
      END
   END FE_OFN1127_n_4090

   PIN FE_OFN1128_n_4090
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 19.45 0.255 19.65 ;
      END
   END FE_OFN1128_n_4090

   PIN FE_OFN1132_n_6356
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 52.8 49.745 53 50 ;
      END
   END FE_OFN1132_n_6356

   PIN FE_OFN1135_n_4151
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 31.45 0.255 31.65 ;
      END
   END FE_OFN1135_n_4151

   PIN FE_OFN1140_n_6886
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 60.85 49.49 60.95 50 ;
      END
   END FE_OFN1140_n_6886

   PIN FE_OFN1147_n_6391
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 20.25 0.255 20.45 ;
      END
   END FE_OFN1147_n_6391

   PIN FE_OFN1148_n_6391
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 40.45 0.255 40.65 ;
      END
   END FE_OFN1148_n_6391

   PIN FE_OFN1156_n_6391
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 71.8 49.745 72 50 ;
      END
   END FE_OFN1156_n_6391

   PIN FE_OFN1159_n_6391
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 54.8 0 55 0.255 ;
      END
   END FE_OFN1159_n_6391

   PIN FE_OFN1162_n_6391
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 38.2 49.745 38.4 50 ;
      END
   END FE_OFN1162_n_6391

   PIN FE_OFN1167_n_4092
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 23.2 0 23.4 0.255 ;
      END
   END FE_OFN1167_n_4092

   PIN FE_OFN1174_n_4093
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 16.65 0.255 16.85 ;
      END
   END FE_OFN1174_n_4093

   PIN FE_OFN1177_n_4143
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 38.65 49.49 38.75 50 ;
      END
   END FE_OFN1177_n_4143

   PIN FE_OFN1184_n_4143
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 38.85 0.255 39.05 ;
      END
   END FE_OFN1184_n_4143

   PIN FE_OFN1185_n_4143
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 37.8 49.745 38 50 ;
      END
   END FE_OFN1185_n_4143

   PIN FE_OFN1189_n_4095
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 36 0 36.2 0.255 ;
      END
   END FE_OFN1189_n_4095

   PIN FE_OFN1190_n_4095
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 56.6 49.745 56.8 50 ;
      END
   END FE_OFN1190_n_4095

   PIN FE_OFN1193_n_4095
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 33.4 0 33.6 0.255 ;
      END
   END FE_OFN1193_n_4095

   PIN FE_OFN1198_n_4096
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 32.85 0.255 33.05 ;
      END
   END FE_OFN1198_n_4096

   PIN FE_OFN119_n_12502
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 31.3 0.51 31.4 ;
      END
   END FE_OFN119_n_12502

   PIN FE_OFN1213_n_4098
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 40.2 0 40.4 0.255 ;
      END
   END FE_OFN1213_n_4098

   PIN FE_OFN1225_n_6624
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 38.45 0.255 38.65 ;
      END
   END FE_OFN1225_n_6624

   PIN FE_OFN1226_n_6624
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 39.4 0 39.6 0.255 ;
      END
   END FE_OFN1226_n_6624

   PIN FE_OFN1231_n_6624
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 36.4 0 36.6 0.255 ;
      END
   END FE_OFN1231_n_6624

   PIN FE_OFN1233_n_6624
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 59 49.745 59.2 50 ;
      END
   END FE_OFN1233_n_6624

   PIN FE_OFN1235_n_6436
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 25.85 49.49 25.95 50 ;
      END
   END FE_OFN1235_n_6436

   PIN FE_OFN130_n_12104
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 47.45 49.49 47.55 50 ;
      END
   END FE_OFN130_n_12104

   PIN FE_OFN1431_n_12104
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 16.25 49.49 16.35 50 ;
      END
   END FE_OFN1431_n_12104

   PIN FE_OFN1435_n_12042
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 73 49.745 73.2 50 ;
      END
   END FE_OFN1435_n_12042

   PIN FE_OFN1441_n_12502
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 28.45 49.49 28.55 50 ;
      END
   END FE_OFN1441_n_12502

   PIN FE_OFN1445_n_12502
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 70.8 49.745 71 50 ;
      END
   END FE_OFN1445_n_12502

   PIN FE_OFN1449_n_10780
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 21.25 49.49 21.35 50 ;
      END
   END FE_OFN1449_n_10780

   PIN FE_OFN1455_n_12028
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 37.25 0.255 37.45 ;
      END
   END FE_OFN1455_n_12028

   PIN FE_OFN1458_n_12306
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 24.45 49.49 24.55 50 ;
      END
   END FE_OFN1458_n_12306

   PIN FE_OFN1461_n_12306
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 17.85 49.49 17.95 50 ;
      END
   END FE_OFN1461_n_12306

   PIN FE_OFN1474_n_14995
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 39.25 49.49 39.35 50 ;
      END
   END FE_OFN1474_n_14995

   PIN FE_OFN1475_n_14995
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 15.05 49.49 15.15 50 ;
      END
   END FE_OFN1475_n_14995

   PIN FE_OFN1507_n_4460
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 31.45 49.49 31.55 50 ;
      END
   END FE_OFN1507_n_4460

   PIN FE_OFN1511_n_4460
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 30.05 0.255 30.25 ;
      END
   END FE_OFN1511_n_4460

   PIN FE_OFN1515_n_4677
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 16.2 0 16.4 0.255 ;
      END
   END FE_OFN1515_n_4677

   PIN FE_OFN1547_n_4501
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 37.65 0.255 37.85 ;
      END
   END FE_OFN1547_n_4501

   PIN FE_OFN1548_n_4501
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 35.25 49.49 35.35 50 ;
      END
   END FE_OFN1548_n_4501

   PIN FE_OFN1549_n_4501
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 54.6 49.745 54.8 50 ;
      END
   END FE_OFN1549_n_4501

   PIN FE_OFN1653_n_4868
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 37.4 49.745 37.6 50 ;
      END
   END FE_OFN1653_n_4868

   PIN FE_OFN1654_n_4868
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 12.6 49.745 12.8 50 ;
      END
   END FE_OFN1654_n_4868

   PIN FE_OFN1718_n_16317
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 26.45 49.49 26.55 50 ;
      END
   END FE_OFN1718_n_16317

   PIN FE_OFN1726_n_14987
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 44.05 49.49 44.15 50 ;
      END
   END FE_OFN1726_n_14987

   PIN FE_OFN1733_n_11019
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 26.25 0 26.35 0.51 ;
      END
   END FE_OFN1733_n_11019

   PIN FE_OFN1745_n_12086
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 32.5 0.51 32.6 ;
      END
   END FE_OFN1745_n_12086

   PIN FE_OFN1751_n_11027
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 29.5 0.51 29.6 ;
      END
   END FE_OFN1751_n_11027

   PIN FE_OFN1755_n_12681
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 16.65 0 16.75 0.51 ;
      END
   END FE_OFN1755_n_12681

   PIN FE_OFN1794_n_4508
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 31.05 0.255 31.25 ;
      END
   END FE_OFN1794_n_4508

   PIN FE_OFN1797_n_4508
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 39.85 0.255 40.05 ;
      END
   END FE_OFN1797_n_4508

   PIN FE_OFN1804_n_3741
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 27.45 0.255 27.65 ;
      END
   END FE_OFN1804_n_3741

   PIN FE_OFN1826_n_4490
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 57 49.745 57.2 50 ;
      END
   END FE_OFN1826_n_4490

   PIN FE_OFN325_g66125_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 23.05 49.49 23.15 50 ;
      END
   END FE_OFN325_g66125_p

   PIN FE_OFN589_n_4490
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 53.6 49.745 53.8 50 ;
      END
   END FE_OFN589_n_4490

   PIN FE_OFN590_n_4490
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 41.05 0.255 41.25 ;
      END
   END FE_OFN590_n_4490

   PIN FE_OFN591_n_4490
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 39 49.745 39.2 50 ;
      END
   END FE_OFN591_n_4490

   PIN FE_OFN595_n_4409
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 29.2 49.745 29.4 50 ;
      END
   END FE_OFN595_n_4409

   PIN FE_OFN596_n_4409
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 28.05 0.255 28.25 ;
      END
   END FE_OFN596_n_4409

   PIN FE_OFN597_n_4409
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 57.4 49.745 57.6 50 ;
      END
   END FE_OFN597_n_4409

   PIN FE_OFN599_n_4454
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 36.2 49.745 36.4 50 ;
      END
   END FE_OFN599_n_4454

   PIN FE_OFN600_n_4454
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 34.45 0.255 34.65 ;
      END
   END FE_OFN600_n_4454

   PIN FE_OFN607_n_4669
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 35.8 49.745 36 50 ;
      END
   END FE_OFN607_n_4669

   PIN FE_OFN612_n_4497
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 35.45 0.255 35.65 ;
      END
   END FE_OFN612_n_4497

   PIN FE_OFN613_n_4497
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 69.2 49.745 69.4 50 ;
      END
   END FE_OFN613_n_4497

   PIN FE_OFN614_n_4497
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 22.05 0.255 22.25 ;
      END
   END FE_OFN614_n_4497

   PIN FE_OFN626_n_4392
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 20.2 0 20.4 0.255 ;
      END
   END FE_OFN626_n_4392

   PIN FE_OFN629_n_4495
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 38.05 0.255 38.25 ;
      END
   END FE_OFN629_n_4495

   PIN FE_OFN631_n_4495
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 23.05 0.255 23.25 ;
      END
   END FE_OFN631_n_4495

   PIN FE_OFN634_n_4505
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 39.45 0.255 39.65 ;
      END
   END FE_OFN634_n_4505

   PIN FE_OFN635_n_4505
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 72.2 49.745 72.4 50 ;
      END
   END FE_OFN635_n_4505

   PIN FE_OFN636_n_4505
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 34.2 49.745 34.4 50 ;
      END
   END FE_OFN636_n_4505

   PIN FE_OFN649_n_4417
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 27.65 49.49 27.75 50 ;
      END
   END FE_OFN649_n_4417

   PIN FE_OFN654_n_4438
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 26.25 49.49 26.35 50 ;
      END
   END FE_OFN654_n_4438

   PIN FE_OFN656_n_4438
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 35.6 0 35.8 0.255 ;
      END
   END FE_OFN656_n_4438

   PIN FE_OFN967_n_4655
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 55 49.745 55.2 50 ;
      END
   END FE_OFN967_n_4655

   PIN FE_OFN968_n_4655
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 35 0 35.2 0.255 ;
      END
   END FE_OFN968_n_4655

   PIN FE_RN_203_0
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 17.65 49.49 17.75 50 ;
      END
   END FE_RN_203_0

   PIN g62336_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 19.85 49.49 19.95 50 ;
      END
   END g62336_sb

   PIN g62345_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 42.5 0.51 42.6 ;
      END
   END g62345_da

   PIN g62362_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 42.3 0.51 42.4 ;
      END
   END g62362_db

   PIN g62362_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 21.45 49.49 21.55 50 ;
      END
   END g62362_sb

   PIN g62389_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 33.25 49.49 33.35 50 ;
      END
   END g62389_db

   PIN g62389_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 32.25 49.49 32.35 50 ;
      END
   END g62389_sb

   PIN g62410_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 29.5 0.51 29.6 ;
      END
   END g62410_db

   PIN g62485_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 24.65 49.49 24.75 50 ;
      END
   END g62485_sb

   PIN g62547_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 47.65 49.49 47.75 50 ;
      END
   END g62547_db

   PIN g62601_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 42.1 0.51 42.2 ;
      END
   END g62601_sb

   PIN g62911_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 11.05 49.49 11.15 50 ;
      END
   END g62911_db

   PIN g62923_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 16.45 49.49 16.55 50 ;
      END
   END g62923_db

   PIN g62923_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 11.05 49.49 11.15 50 ;
      END
   END g62923_sb

   PIN g62953_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 10.85 49.49 10.95 50 ;
      END
   END g62953_db

   PIN g62980_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 71.05 49.49 71.15 50 ;
      END
   END g62980_sb

   PIN g63183_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 35.9 0.51 36 ;
      END
   END g63183_da

   PIN g64800_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 42.65 49.49 42.75 50 ;
      END
   END g64800_sb

   PIN g64906_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 50.85 49.49 50.95 50 ;
      END
   END g64906_sb

   PIN g64907_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 56.45 49.49 56.55 50 ;
      END
   END g64907_sb

   PIN g64908_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 25.05 49.49 25.15 50 ;
      END
   END g64908_da

   PIN g64949_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 27.9 0.51 28 ;
      END
   END g64949_sb

   PIN g65335_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 10.85 49.49 10.95 50 ;
      END
   END g65335_da

   PIN g65351_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 73.65 49.49 73.75 50 ;
      END
   END g65351_sb

   PIN g65381_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 29.65 49.49 29.75 50 ;
      END
   END g65381_db

   PIN g65394_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 72.25 49.49 72.35 50 ;
      END
   END g65394_da

   PIN g65394_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 72.45 49.49 72.55 50 ;
      END
   END g65394_db

   PIN g66098_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 31.05 49.49 31.15 50 ;
      END
   END g66098_p

   PIN g66128_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 21.05 49.49 21.15 50 ;
      END
   END g66128_p

   PIN g66134_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 10.65 49.49 10.75 50 ;
      END
   END g66134_p

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 20.25 49.49 20.35 50 ;
      END
   END ispd_clk

   PIN n_12001
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 26.5 0.51 26.6 ;
      END
   END n_12001

   PIN n_12010
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 30.65 0.255 30.85 ;
      END
   END n_12010

   PIN n_12042
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 10.65 49.49 10.75 50 ;
      END
   END n_12042

   PIN n_12105
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 38.45 49.49 38.55 50 ;
      END
   END n_12105

   PIN n_12356
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 33.3 0.51 33.4 ;
      END
   END n_12356

   PIN n_12403
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 19.25 0 19.35 0.51 ;
      END
   END n_12403

   PIN n_12433
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 49.85 49.49 49.95 50 ;
      END
   END n_12433

   PIN n_12458
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 28.5 0.51 28.6 ;
      END
   END n_12458

   PIN n_12612
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 25.9 0.51 26 ;
      END
   END n_12612

   PIN n_12645
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 32.1 0.51 32.2 ;
      END
   END n_12645

   PIN n_12685
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 62.45 49.49 62.55 50 ;
      END
   END n_12685

   PIN n_12695
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 18.45 49.49 18.55 50 ;
      END
   END n_12695

   PIN n_12865
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 32.3 0.51 32.4 ;
      END
   END n_12865

   PIN n_12866
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 25.7 0.51 25.8 ;
      END
   END n_12866

   PIN n_13058
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 10.45 49.49 10.55 50 ;
      END
   END n_13058

   PIN n_13144
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 19.85 0 19.95 0.51 ;
      END
   END n_13144

   PIN n_13402
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 16.05 0 16.15 0.51 ;
      END
   END n_13402

   PIN n_13760
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 28.25 49.49 28.35 50 ;
      END
   END n_13760

   PIN n_14309
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 40.85 49.49 40.95 50 ;
      END
   END n_14309

   PIN n_14313
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 29.05 49.49 29.15 50 ;
      END
   END n_14313

   PIN n_14317
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 36.85 49.49 36.95 50 ;
      END
   END n_14317

   PIN n_14353
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 41.9 0.51 42 ;
      END
   END n_14353

   PIN n_156
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 11.25 49.49 11.35 50 ;
      END
   END n_156

   PIN n_3464
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 12.2 49.745 12.4 50 ;
      END
   END n_3464

   PIN n_3752
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 51 49.745 51.2 50 ;
      END
   END n_3752

   PIN n_3755
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 56.2 49.745 56.4 50 ;
      END
   END n_3755

   PIN n_3770
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 70 49.745 70.2 50 ;
      END
   END n_3770

   PIN n_3774
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 72.6 49.745 72.8 50 ;
      END
   END n_3774

   PIN n_3777
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 11.8 49.745 12 50 ;
      END
   END n_3777

   PIN n_3785
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 18.25 49.49 18.35 50 ;
      END
   END n_3785

   PIN n_3792
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 55.4 49.745 55.6 50 ;
      END
   END n_3792

   PIN n_4308
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 31.9 0.51 32 ;
      END
   END n_4308

   PIN n_4357
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 15.05 0 15.15 0.51 ;
      END
   END n_4357

   PIN n_4373
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 17.45 49.49 17.55 50 ;
      END
   END n_4373

   PIN n_4442
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 22.45 0.255 22.65 ;
      END
   END n_4442

   PIN n_4444
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 49.2 49.745 49.4 50 ;
      END
   END n_4444

   PIN n_4450
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 37 49.745 37.2 50 ;
      END
   END n_4450

   PIN n_4452
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 36.6 49.745 36.8 50 ;
      END
   END n_4452

   PIN n_4465
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 34.2 0 34.4 0.255 ;
      END
   END n_4465

   PIN n_4476
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 34.6 0 34.8 0.255 ;
      END
   END n_4476

   PIN n_4479
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 11.4 49.745 11.6 50 ;
      END
   END n_4479

   PIN n_4488
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 55.8 49.745 56 50 ;
      END
   END n_4488

   PIN n_4493
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 18 0 18.2 0.255 ;
      END
   END n_4493

   PIN n_4645
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 32.05 0.255 32.25 ;
      END
   END n_4645

   PIN n_6189
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 19.65 49.49 19.75 50 ;
      END
   END n_6189

   PIN n_6232
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 53.2 49.745 53.4 50 ;
      END
   END n_6232

   PIN n_6287
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 41.45 0.255 41.65 ;
      END
   END n_6287

   PIN n_6319
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 30.4 49.745 30.6 50 ;
      END
   END n_6319

   PIN n_6388
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 15.85 0 15.95 0.51 ;
      END
   END n_6388

   PIN n_6645
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 13 49.745 13.2 50 ;
      END
   END n_6645

   PIN n_7631
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 28.85 49.49 28.95 50 ;
      END
   END n_7631

   PIN n_7671
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 25.65 49.49 25.75 50 ;
      END
   END n_7671

   PIN wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__0__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 18.05 49.49 18.15 50 ;
      END
   END wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__0__Q

   PIN wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__29__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 22.05 49.49 22.15 50 ;
      END
   END wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__29__Q

   PIN wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__8__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 10.45 49.49 10.55 50 ;
      END
   END wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__8__Q

   PIN wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__12__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 15.65 49.49 15.75 50 ;
      END
   END wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__12__Q

   PIN wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__21__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 48.85 49.49 48.95 50 ;
      END
   END wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__21__Q

   PIN wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__29__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 22.85 49.49 22.95 50 ;
      END
   END wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__29__Q

   PIN wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__30__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 63.45 49.49 63.55 50 ;
      END
   END wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__30__Q

   PIN wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__16__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 70.65 49.49 70.75 50 ;
      END
   END wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__16__Q

   PIN wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__14__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 21.5 0.51 21.6 ;
      END
   END wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__14__Q

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 358.4 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 358.4 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 358.4 8.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 11.745 358.4 12.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 15.745 358.4 16.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 19.745 358.4 20.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 23.745 358.4 24.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 27.745 358.4 28.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 31.745 358.4 32.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 35.745 358.4 36.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 39.745 358.4 40.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 43.745 358.4 44.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 47.745 358.4 48.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 358.4 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 358.4 6.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 9.745 358.4 10.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 13.745 358.4 14.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 17.745 358.4 18.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 21.745 358.4 22.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 25.745 358.4 26.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 29.745 358.4 30.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 33.745 358.4 34.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 37.745 358.4 38.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 41.745 358.4 42.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 45.745 358.4 46.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 49.745 358.4 50.255 ;
      END
   END vdd

   OBS
      LAYER metal1 ;
         RECT 0 0 358.4 50 ;
   END
   OBS
      LAYER metal2 ;
         RECT 0 0 358.4 50 ;
   END
   OBS
      LAYER metal3 ;
         RECT 0 0 358.4 50 ;
   END
   OBS
      LAYER metal4 ;
         RECT 0 0 358.4 50 ;
   END
   OBS
      LAYER metal5 ;
         RECT 0 0 358.4 50 ;
   END
END h8

MACRO hh4
   CLASS BLOCK ;
   SIZE 352.6 BY 160 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   PIN FE_OCP_RBN2106_n_9155
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 352.09 63.75 352.6 63.85 ;
      END
   END FE_OCP_RBN2106_n_9155

   PIN FE_OFN1262_n_8567
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 352.09 63.95 352.6 64.05 ;
      END
   END FE_OFN1262_n_8567

   PIN FE_OFN1316_n_8567
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 182.2 159.745 182.4 160 ;
      END
   END FE_OFN1316_n_8567

   PIN FE_OFN1334_n_9372
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 352.09 66.15 352.6 66.25 ;
      END
   END FE_OFN1334_n_9372

   PIN FE_OFN1336_n_9372
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 352.345 38.9 352.6 39.1 ;
      END
   END FE_OFN1336_n_9372

   PIN FE_OFN1337_n_9372
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 352.345 39.3 352.6 39.5 ;
      END
   END FE_OFN1337_n_9372

   PIN FE_OFN1340_n_9372
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 352.345 64.3 352.6 64.5 ;
      END
   END FE_OFN1340_n_9372

   PIN FE_OFN1498_n_9864
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 286.45 0 286.55 0.51 ;
      END
   END FE_OFN1498_n_9864

   PIN FE_OFN1499_n_9864
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 352.345 64.7 352.6 64.9 ;
      END
   END FE_OFN1499_n_9864

   PIN FE_OFN1537_n_9428
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 171.6 159.745 171.8 160 ;
      END
   END FE_OFN1537_n_9428

   PIN FE_OFN222_n_9844
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 352.345 13.3 352.6 13.5 ;
      END
   END FE_OFN222_n_9844

   PIN FE_OFN248_n_9114
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 352.345 138.7 352.6 138.9 ;
      END
   END FE_OFN248_n_9114

   PIN FE_OFN257_n_8969
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 261.85 159.49 261.95 160 ;
      END
   END FE_OFN257_n_8969

   PIN FE_OFN448_n_10853
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 352.09 65.15 352.6 65.25 ;
      END
   END FE_OFN448_n_10853

   PIN FE_OFN523_n_9690
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 289.2 0 289.4 0.255 ;
      END
   END FE_OFN523_n_9690

   PIN FE_OFN534_n_9864
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 131.8 0 132 0.255 ;
      END
   END FE_OFN534_n_9864

   PIN FE_OFN566_n_9692
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 352.345 65.5 352.6 65.7 ;
      END
   END FE_OFN566_n_9692

   PIN g57223_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 202.05 0 202.15 0.51 ;
      END
   END g57223_da

   PIN g57530_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 95.85 159.49 95.95 160 ;
      END
   END g57530_db

   PIN g57535_sb
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 82.85 0 82.95 0.51 ;
      END
   END g57535_sb

   PIN g57913_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 59.05 0 59.15 0.51 ;
      END
   END g57913_db

   PIN g58063_sb
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 24.45 0 24.55 0.51 ;
      END
   END g58063_sb

   PIN g58199_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 128.65 0 128.75 0.51 ;
      END
   END g58199_da

   PIN g58376_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 126.85 159.49 126.95 160 ;
      END
   END g58376_db

   PIN g58389_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 105.85 159.49 105.95 160 ;
      END
   END g58389_da

   PIN g58428_sb
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 159.05 159.49 159.15 160 ;
      END
   END g58428_sb

   PIN g58439_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 161.05 159.49 161.15 160 ;
      END
   END g58439_db

   PIN g58439_sb
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 164.45 159.49 164.55 160 ;
      END
   END g58439_sb

   PIN g58481_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 278.85 159.49 278.95 160 ;
      END
   END g58481_db

   PIN g58832_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 266.25 159.49 266.35 160 ;
      END
   END g58832_da

   PIN n_10185
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 231.05 0 231.15 0.51 ;
      END
   END n_10185

   PIN n_10627
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 257.45 0 257.55 0.51 ;
      END
   END n_10627

   PIN n_10753
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 138.35 0.51 138.45 ;
      END
   END n_10753

   PIN n_11005
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 265.45 0 265.55 0.51 ;
      END
   END n_11005

   PIN n_11236
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 166.85 0 166.95 0.51 ;
      END
   END n_11236

   PIN n_11410
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 321.45 0 321.55 0.51 ;
      END
   END n_11410

   PIN n_12573
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 176.65 0 176.75 0.51 ;
      END
   END n_12573

   PIN n_12578
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 278.45 0 278.55 0.51 ;
      END
   END n_12578

   PIN n_2933
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 352.09 113.35 352.6 113.45 ;
      END
   END n_2933

   PIN n_8714
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 78.65 159.49 78.75 160 ;
      END
   END n_8714

   PIN n_8884
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 223.8 159.745 224 160 ;
      END
   END n_8884

   PIN n_9228
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 232.25 159.49 232.35 160 ;
      END
   END n_9228

   PIN n_9419
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 98.25 159.49 98.35 160 ;
      END
   END n_9419

   PIN n_9440
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 118.25 0 118.35 0.51 ;
      END
   END n_9440

   PIN wbu_sel_in_312
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 238.25 0 238.35 0.51 ;
      END
   END wbu_sel_in_312

   PIN wishbone_slave_unit_del_sync_addr_out_reg_5__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 112.85 159.49 112.95 160 ;
      END
   END wishbone_slave_unit_del_sync_addr_out_reg_5__Q

   PIN wishbone_slave_unit_fifos_wbr_be_in_264
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 352.09 112.95 352.6 113.05 ;
      END
   END wishbone_slave_unit_fifos_wbr_be_in_264

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__16__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 298.45 0 298.55 0.51 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__16__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__31__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 352.09 90.15 352.6 90.25 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__31__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__33__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 80.45 159.49 80.55 160 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__33__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__10__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 275.45 0 275.55 0.51 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__10__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__22__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 186.45 0 186.55 0.51 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__22__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__20__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 89.55 0.51 89.65 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__20__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__5__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 89.35 0.51 89.45 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__5__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__27__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 220.85 0 220.95 0.51 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__27__Q

   PIN wishbone_slave_unit_pcim_if_wbw_addr_data_in_388
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 352.09 90.35 352.6 90.45 ;
      END
   END wishbone_slave_unit_pcim_if_wbw_addr_data_in_388

   PIN FE_OCPN1879_n_9991
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 138.55 0.51 138.65 ;
      END
   END FE_OCPN1879_n_9991

   PIN FE_OCPN1936_n_15566
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 257.6 0 257.8 0.255 ;
      END
   END FE_OCPN1936_n_15566

   PIN FE_OCP_RBN2104_n_9155
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 352.09 63.55 352.6 63.65 ;
      END
   END FE_OCP_RBN2104_n_9155

   PIN FE_OFN1251_n_16439
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 267.85 159.49 267.95 160 ;
      END
   END FE_OFN1251_n_16439

   PIN FE_OFN1253_n_8567
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 352.09 63.35 352.6 63.45 ;
      END
   END FE_OFN1253_n_8567

   PIN FE_OFN1282_n_8567
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 179.05 159.49 179.15 160 ;
      END
   END FE_OFN1282_n_8567

   PIN FE_OFN1285_n_8567
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 112.9 0.255 113.1 ;
      END
   END FE_OFN1285_n_8567

   PIN FE_OFN1287_n_8567
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 211.8 0 212 0.255 ;
      END
   END FE_OFN1287_n_8567

   PIN FE_OFN1289_n_8567
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 331 0 331.2 0.255 ;
      END
   END FE_OFN1289_n_8567

   PIN FE_OFN1296_n_8567
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 88.6 0 88.8 0.255 ;
      END
   END FE_OFN1296_n_8567

   PIN FE_OFN1298_n_8567
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 65.6 159.745 65.8 160 ;
      END
   END FE_OFN1298_n_8567

   PIN FE_OFN1308_n_8567
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 95.4 159.745 95.6 160 ;
      END
   END FE_OFN1308_n_8567

   PIN FE_OFN1315_n_8567
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 133.2 0 133.4 0.255 ;
      END
   END FE_OFN1315_n_8567

   PIN FE_OFN1341_n_9372
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 269.4 159.745 269.6 160 ;
      END
   END FE_OFN1341_n_9372

   PIN FE_OFN1377_n_10853
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 352.09 62.95 352.6 63.05 ;
      END
   END FE_OFN1377_n_10853

   PIN FE_OFN13_n_11877
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 255.2 0 255.4 0.255 ;
      END
   END FE_OFN13_n_11877

   PIN FE_OFN1400_n_10566
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 196.45 0 196.55 0.51 ;
      END
   END FE_OFN1400_n_10566

   PIN FE_OFN1496_n_9864
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 132.05 0 132.15 0.51 ;
      END
   END FE_OFN1496_n_9864

   PIN FE_OFN1497_n_9864
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 352.09 62.95 352.6 63.05 ;
      END
   END FE_OFN1497_n_9864

   PIN FE_OFN1534_n_9428
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 174.05 159.49 174.15 160 ;
      END
   END FE_OFN1534_n_9428

   PIN FE_OFN1541_n_9502
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 137.85 159.49 137.95 160 ;
      END
   END FE_OFN1541_n_9502

   PIN FE_OFN1572_n_9477
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 116.2 159.745 116.4 160 ;
      END
   END FE_OFN1572_n_9477

   PIN FE_OFN1632_n_9862
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 128 159.745 128.2 160 ;
      END
   END FE_OFN1632_n_9862

   PIN FE_OFN1687_n_15534
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 285.85 0 285.95 0.51 ;
      END
   END FE_OFN1687_n_15534

   PIN FE_OFN1692_n_16992
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 286.25 0 286.35 0.51 ;
      END
   END FE_OFN1692_n_16992

   PIN FE_OFN1713_n_9320
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 195.85 0 195.95 0.51 ;
      END
   END FE_OFN1713_n_9320

   PIN FE_OFN1807_n_9899
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 113.9 0.255 114.1 ;
      END
   END FE_OFN1807_n_9899

   PIN FE_OFN199_n_9228
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 161.25 159.49 161.35 160 ;
      END
   END FE_OFN199_n_9228

   PIN FE_OFN214_n_9856
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 117.4 0 117.6 0.255 ;
      END
   END FE_OFN214_n_9856

   PIN FE_OFN220_n_9846
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 128.4 159.745 128.6 160 ;
      END
   END FE_OFN220_n_9846

   PIN FE_OFN224_n_9122
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 137.4 159.745 137.6 160 ;
      END
   END FE_OFN224_n_9122

   PIN FE_OFN233_n_9876
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 108.6 0 108.8 0.255 ;
      END
   END FE_OFN233_n_9876

   PIN FE_OFN236_n_9834
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 171.2 159.745 171.4 160 ;
      END
   END FE_OFN236_n_9834

   PIN FE_OFN498_n_9697
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 196.2 159.745 196.4 160 ;
      END
   END FE_OFN498_n_9697

   PIN FE_OFN519_n_9690
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 289.45 0 289.55 0.51 ;
      END
   END FE_OFN519_n_9690

   PIN FE_OFN548_n_9502
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 152.6 159.745 152.8 160 ;
      END
   END FE_OFN548_n_9502

   PIN FE_OFN555_n_9902
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 162.2 0 162.4 0.255 ;
      END
   END FE_OFN555_n_9902

   PIN FE_OFN559_n_9531
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 109 0 109.2 0.255 ;
      END
   END FE_OFN559_n_9531

   PIN FE_OFN561_n_9692
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 352.09 63.15 352.6 63.25 ;
      END
   END FE_OFN561_n_9692

   PIN FE_OFN571_n_9694
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 165.2 159.745 165.4 160 ;
      END
   END FE_OFN571_n_9694

   PIN FE_OFN581_n_9904
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 88.9 0.255 89.1 ;
      END
   END FE_OFN581_n_9904

   PIN g57041_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 306.25 0 306.35 0.51 ;
      END
   END g57041_da

   PIN g57341_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 321.05 0 321.15 0.51 ;
      END
   END g57341_db

   PIN g58063_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 38.95 0.51 39.05 ;
      END
   END g58063_da

   PIN g58082_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 171.25 0 171.35 0.51 ;
      END
   END g58082_db

   PIN g58361_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 142.65 0 142.75 0.51 ;
      END
   END g58361_da

   PIN g58389_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 106.25 159.49 106.35 160 ;
      END
   END g58389_sb

   PIN g58393_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 118.45 0 118.55 0.51 ;
      END
   END g58393_da

   PIN g58428_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 98.45 159.49 98.55 160 ;
      END
   END g58428_da

   PIN g58829_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 210.85 159.49 210.95 160 ;
      END
   END g58829_db

   PIN g59091_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 78.85 159.49 78.95 160 ;
      END
   END g59091_da

   PIN g59091_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 79.05 159.49 79.15 160 ;
      END
   END g59091_db

   PIN g63585_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 244.45 0 244.55 0.51 ;
      END
   END g63585_da

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 251 0 251.2 0.255 ;
      END
   END ispd_clk

   PIN n_10051
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 160.65 0 160.75 0.51 ;
      END
   END n_10051

   PIN n_10054
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 166.05 0 166.15 0.51 ;
      END
   END n_10054

   PIN n_10057
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 165.05 0 165.15 0.51 ;
      END
   END n_10057

   PIN n_10314
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 111.45 159.49 111.55 160 ;
      END
   END n_10314

   PIN n_10693
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 138.75 0.51 138.85 ;
      END
   END n_10693

   PIN n_11223
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 276.45 0 276.55 0.51 ;
      END
   END n_11223

   PIN n_11264
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 352.09 89.95 352.6 90.05 ;
      END
   END n_11264

   PIN n_12153
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 278.65 0 278.75 0.51 ;
      END
   END n_12153

   PIN n_1252
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 352.09 89.75 352.6 89.85 ;
      END
   END n_1252

   PIN n_12825
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 352.09 89.55 352.6 89.65 ;
      END
   END n_12825

   PIN n_1340
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 352.09 89.35 352.6 89.45 ;
      END
   END n_1340

   PIN n_1342
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 352.09 89.15 352.6 89.25 ;
      END
   END n_1342

   PIN n_1354
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 352.09 88.95 352.6 89.05 ;
      END
   END n_1354

   PIN n_15568
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 258.25 0 258.35 0.51 ;
      END
   END n_15568

   PIN n_2401
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 352.09 113.15 352.6 113.25 ;
      END
   END n_2401

   PIN n_8605
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 251.65 159.49 251.75 160 ;
      END
   END n_8605

   PIN n_8831
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 231 159.745 231.2 160 ;
      END
   END n_8831

   PIN n_8832
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 245.05 159.49 245.15 160 ;
      END
   END n_8832

   PIN n_8927
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 231.25 0 231.35 0.51 ;
      END
   END n_8927

   PIN n_9116
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 279.05 159.49 279.15 160 ;
      END
   END n_9116

   PIN n_9269
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 165.65 0 165.75 0.51 ;
      END
   END n_9269

   PIN n_9372
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 352.09 65.95 352.6 66.05 ;
      END
   END n_9372

   PIN n_9407
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 92.85 0 92.95 0.51 ;
      END
   END n_9407

   PIN n_9586
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 314.85 0 314.95 0.51 ;
      END
   END n_9586

   PIN n_9844
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 313.85 0 313.95 0.51 ;
      END
   END n_9844

   PIN wbu_addr_in_254
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 303.25 159.49 303.35 160 ;
      END
   END wbu_addr_in_254

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__29__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 133.05 0 133.15 0.51 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__29__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__29__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 196.25 0 196.35 0.51 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__29__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__27__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 59.25 0 59.35 0.51 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__27__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__29__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 258.65 0 258.75 0.51 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__29__Q

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 352.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 352.6 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 352.6 8.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 11.745 352.6 12.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 15.745 352.6 16.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 19.745 352.6 20.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 23.745 352.6 24.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 27.745 352.6 28.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 31.745 352.6 32.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 35.745 352.6 36.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 39.745 352.6 40.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 43.745 352.6 44.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 47.745 352.6 48.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 51.745 352.6 52.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 55.745 352.6 56.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 59.745 352.6 60.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 63.745 352.6 64.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 67.745 352.6 68.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 71.745 352.6 72.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 75.745 352.6 76.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 79.745 352.6 80.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 83.745 352.6 84.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 87.745 352.6 88.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 91.745 352.6 92.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 95.745 352.6 96.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 99.745 352.6 100.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 103.745 352.6 104.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 107.745 352.6 108.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 111.745 352.6 112.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 115.745 352.6 116.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 119.745 352.6 120.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 123.745 352.6 124.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 127.745 352.6 128.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 131.745 352.6 132.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 135.745 352.6 136.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 139.745 352.6 140.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 143.745 352.6 144.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 147.745 352.6 148.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 151.745 352.6 152.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 155.745 352.6 156.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 159.745 352.6 160.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 352.6 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 352.6 6.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 9.745 352.6 10.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 13.745 352.6 14.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 17.745 352.6 18.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 21.745 352.6 22.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 25.745 352.6 26.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 29.745 352.6 30.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 33.745 352.6 34.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 37.745 352.6 38.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 41.745 352.6 42.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 45.745 352.6 46.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 49.745 352.6 50.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 53.745 352.6 54.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 57.745 352.6 58.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 61.745 352.6 62.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 65.745 352.6 66.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 69.745 352.6 70.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 73.745 352.6 74.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 77.745 352.6 78.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 81.745 352.6 82.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 85.745 352.6 86.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 89.745 352.6 90.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 93.745 352.6 94.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 97.745 352.6 98.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 101.745 352.6 102.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 105.745 352.6 106.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 109.745 352.6 110.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 113.745 352.6 114.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 117.745 352.6 118.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 121.745 352.6 122.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 125.745 352.6 126.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 129.745 352.6 130.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 133.745 352.6 134.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 137.745 352.6 138.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 141.745 352.6 142.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 145.745 352.6 146.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 149.745 352.6 150.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 153.745 352.6 154.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 157.745 352.6 158.255 ;
      END
   END vdd

   OBS
      LAYER metal1 ;
         RECT 0 0 352.6 160 ;
   END
   OBS
      LAYER metal2 ;
         RECT 0 0 352.6 160 ;
   END
   OBS
      LAYER metal3 ;
         RECT 0 0 352.6 160 ;
   END
   OBS
      LAYER metal4 ;
         RECT 0 0 352.6 160 ;
   END
   OBS
      LAYER metal5 ;
         RECT 0 0 352.6 160 ;
   END
END hh4

MACRO h5
   CLASS BLOCK ;
   SIZE 359 BY 154 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   PIN FE_OCPN1988_FE_OFN1264_n_8567
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 309.2 0 309.4 0.255 ;
      END
   END FE_OCPN1988_FE_OFN1264_n_8567

   PIN FE_OFN1299_n_8567
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 117.4 0 117.6 0.255 ;
      END
   END FE_OFN1299_n_8567

   PIN FE_OFN1504_n_9531
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 31.85 0 31.95 0.51 ;
      END
   END FE_OFN1504_n_9531

   PIN FE_OFN1675_n_10588
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 78.05 0 78.15 0.51 ;
      END
   END FE_OFN1675_n_10588

   PIN FE_OFN538_n_9895
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 90.9 0.255 91.1 ;
      END
   END FE_OFN538_n_9895

   PIN g57182_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 61.65 0 61.75 0.51 ;
      END
   END g57182_da

   PIN g57202_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 60.85 153.49 60.95 154 ;
      END
   END g57202_db

   PIN g57368_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 237.25 0 237.35 0.51 ;
      END
   END g57368_db

   PIN g57569_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 149.45 0 149.55 0.51 ;
      END
   END g57569_db

   PIN g57942_sb
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 71.65 0 71.75 0.51 ;
      END
   END g57942_sb

   PIN g58061_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 74.05 153.49 74.15 154 ;
      END
   END g58061_db

   PIN g58210_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 55.05 0 55.15 0.51 ;
      END
   END g58210_db

   PIN g58235_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 21.75 0.51 21.85 ;
      END
   END g58235_db

   PIN g58319_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 47.85 153.49 47.95 154 ;
      END
   END g58319_db

   PIN g58425_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 163.05 0 163.15 0.51 ;
      END
   END g58425_da

   PIN g61860_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 333.25 153.49 333.35 154 ;
      END
   END g61860_da

   PIN n_10554
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 57.55 0.51 57.65 ;
      END
   END n_10554

   PIN n_11097
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 163.45 153.49 163.55 154 ;
      END
   END n_11097

   PIN n_11198
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 358.49 57.15 359 57.25 ;
      END
   END n_11198

   PIN n_11261
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 358.49 57.35 359 57.45 ;
      END
   END n_11261

   PIN n_12158
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 189.45 0 189.55 0.51 ;
      END
   END n_12158

   PIN n_12530
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 109.05 153.49 109.15 154 ;
      END
   END n_12530

   PIN n_2151
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 159.85 153.49 159.95 154 ;
      END
   END n_2151

   PIN n_7842
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 338.25 0 338.35 0.51 ;
      END
   END n_7842

   PIN n_9878
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 57.75 0.51 57.85 ;
      END
   END n_9878

   PIN n_9971
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 256.85 0 256.95 0.51 ;
      END
   END n_9971

   PIN pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__8__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 139.65 153.49 139.75 154 ;
      END
   END pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__8__Q

   PIN pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__22__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 173.65 0 173.75 0.51 ;
      END
   END pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__22__Q

   PIN pci_target_unit_pcit_if_pcir_fifo_data_in_766
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 136.25 153.49 136.35 154 ;
      END
   END pci_target_unit_pcit_if_pcir_fifo_data_in_766

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__6__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 216.45 0 216.55 0.51 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__6__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__6__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 83.25 153.49 83.35 154 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__6__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__21__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 101.65 0 101.75 0.51 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__21__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__6__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 292.05 0 292.15 0.51 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__6__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__17__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 129.05 0 129.15 0.51 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__17__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__2__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 234.45 0 234.55 0.51 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__2__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__6__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 27.45 153.49 27.55 154 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__6__Q

   PIN FE_OCPN1987_FE_OFN1264_n_8567
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 308.65 0 308.75 0.51 ;
      END
   END FE_OCPN1987_FE_OFN1264_n_8567

   PIN FE_OCP_RBN2065_n_16572
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 173.45 0 173.55 0.51 ;
      END
   END FE_OCP_RBN2065_n_16572

   PIN FE_OFN1068_n_8176
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 358.49 90.95 359 91.05 ;
      END
   END FE_OFN1068_n_8176

   PIN FE_OFN1077_n_7845
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 329.2 0 329.4 0.255 ;
      END
   END FE_OFN1077_n_7845

   PIN FE_OFN1265_n_8567
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 358.745 57.7 359 57.9 ;
      END
   END FE_OFN1265_n_8567

   PIN FE_OFN1271_n_8567
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 90.5 0.255 90.7 ;
      END
   END FE_OFN1271_n_8567

   PIN FE_OFN1281_n_8567
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 64.4 0 64.6 0.255 ;
      END
   END FE_OFN1281_n_8567

   PIN FE_OFN1283_n_8567
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 117.65 0 117.75 0.51 ;
      END
   END FE_OFN1283_n_8567

   PIN FE_OFN1322_n_8567
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 237.6 0 237.8 0.255 ;
      END
   END FE_OFN1322_n_8567

   PIN FE_OFN1323_n_8567
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 274.8 0 275 0.255 ;
      END
   END FE_OFN1323_n_8567

   PIN FE_OFN1349_n_9163
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 113.85 153.49 113.95 154 ;
      END
   END FE_OFN1349_n_9163

   PIN FE_OFN1353_n_15558
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 147.85 0 147.95 0.51 ;
      END
   END FE_OFN1353_n_15558

   PIN FE_OFN1365_n_15587
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 257.45 0 257.55 0.51 ;
      END
   END FE_OFN1365_n_15587

   PIN FE_OFN1376_n_10853
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 57.35 0.51 57.45 ;
      END
   END FE_OFN1376_n_10853

   PIN FE_OFN1502_n_9531
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 32.05 0 32.15 0.51 ;
      END
   END FE_OFN1502_n_9531

   PIN FE_OFN1503_n_9531
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 301.45 153.49 301.55 154 ;
      END
   END FE_OFN1503_n_9531

   PIN FE_OFN1543_n_9502
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 358.745 126.9 359 127.1 ;
      END
   END FE_OFN1543_n_9502

   PIN FE_OFN1544_n_9502
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 49.2 153.745 49.4 154 ;
      END
   END FE_OFN1544_n_9502

   PIN FE_OFN1678_n_10588
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 57.15 0.51 57.25 ;
      END
   END FE_OFN1678_n_10588

   PIN FE_OFN1682_n_16891
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 258.05 0 258.15 0.51 ;
      END
   END FE_OFN1682_n_16891

   PIN FE_OFN1717_n_16637
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 113.25 153.49 113.35 154 ;
      END
   END FE_OFN1717_n_16637

   PIN FE_OFN1842_n_9828
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 301.2 153.745 301.4 154 ;
      END
   END FE_OFN1842_n_9828

   PIN FE_OFN222_n_9844
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 48.05 153.49 48.15 154 ;
      END
   END FE_OFN222_n_9844

   PIN FE_OFN239_n_9118
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 211.2 153.745 211.4 154 ;
      END
   END FE_OFN239_n_9118

   PIN FE_OFN521_n_9690
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 21.3 0.255 21.5 ;
      END
   END FE_OFN521_n_9690

   PIN FE_OFN535_n_9895
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 91.75 0.51 91.85 ;
      END
   END FE_OFN535_n_9895

   PIN FE_OFN536_n_9895
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 88.05 0 88.15 0.51 ;
      END
   END FE_OFN536_n_9895

   PIN FE_OFN551_n_9902
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 209.2 0 209.4 0.255 ;
      END
   END FE_OFN551_n_9902

   PIN FE_OFN568_n_9694
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 55.4 0 55.6 0.255 ;
      END
   END FE_OFN568_n_9694

   PIN FE_OFN579_n_9904
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 74.45 153.49 74.55 154 ;
      END
   END FE_OFN579_n_9904

   PIN FE_OFN680_n_8060
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 238.4 153.745 238.6 154 ;
      END
   END FE_OFN680_n_8060

   PIN g57065_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 91.55 0.51 91.65 ;
      END
   END g57065_db

   PIN g57353_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 82.25 0 82.35 0.51 ;
      END
   END g57353_da

   PIN g57473_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 358.49 56.95 359 57.05 ;
      END
   END g57473_db

   PIN g57932_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 56.95 0.51 57.05 ;
      END
   END g57932_da

   PIN g57942_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 91.35 0.51 91.45 ;
      END
   END g57942_da

   PIN g58425_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 163.45 0 163.55 0.51 ;
      END
   END g58425_sb

   PIN g61866_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 107.65 0 107.75 0.51 ;
      END
   END g61866_da

   PIN g62004_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 292.05 153.49 292.15 154 ;
      END
   END g62004_sb

   PIN g62027_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 338.65 0 338.75 0.51 ;
      END
   END g62027_db

   PIN g65976_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 318.05 0 318.15 0.51 ;
      END
   END g65976_da

   PIN g65976_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 318.25 0 318.35 0.51 ;
      END
   END g65976_db

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 102 0 102.2 0.255 ;
      END
   END ispd_clk

   PIN n_10151
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 190.25 0 190.35 0.51 ;
      END
   END n_10151

   PIN n_10154
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 190.05 0 190.15 0.51 ;
      END
   END n_10154

   PIN n_10381
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 291.05 0 291.15 0.51 ;
      END
   END n_10381

   PIN n_10414
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 217.45 0 217.55 0.51 ;
      END
   END n_10414

   PIN n_10426
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 28.45 153.49 28.55 154 ;
      END
   END n_10426

   PIN n_10588
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 78.25 0 78.35 0.51 ;
      END
   END n_10588

   PIN n_11040
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 110.65 153.49 110.75 154 ;
      END
   END n_11040

   PIN n_11041
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 110.05 153.49 110.15 154 ;
      END
   END n_11041

   PIN n_11572
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 130.05 0 130.15 0.51 ;
      END
   END n_11572

   PIN n_11773
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 109.65 153.49 109.75 154 ;
      END
   END n_11773

   PIN n_12548
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 137.25 153.49 137.35 154 ;
      END
   END n_12548

   PIN n_1851
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 333.45 153.49 333.55 154 ;
      END
   END n_1851

   PIN n_2053
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 189.2 153.745 189.4 154 ;
      END
   END n_2053

   PIN n_2299
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 173.2 153.745 173.4 154 ;
      END
   END n_2299

   PIN n_7853
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 140.65 153.49 140.75 154 ;
      END
   END n_7853

   PIN n_8407
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 129.2 0 129.4 0.255 ;
      END
   END n_8407

   PIN n_9307
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 189.65 0 189.75 0.51 ;
      END
   END n_9307

   PIN n_9744
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 61.85 0 61.95 0.51 ;
      END
   END n_9744

   PIN pci_target_unit_fifos_pcir_data_in_165
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 173.05 153.49 173.15 154 ;
      END
   END pci_target_unit_fifos_pcir_data_in_165

   PIN pci_target_unit_fifos_pcir_data_in_179
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 269.25 153.49 269.35 154 ;
      END
   END pci_target_unit_fifos_pcir_data_in_179

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__26__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 41.85 0 41.95 0.51 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__26__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__3__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 314.25 153.49 314.35 154 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__3__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__3__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 266.25 0 266.35 0.51 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__3__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__3__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 74.25 153.49 74.35 154 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__3__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__17__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 163.25 0 163.35 0.51 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__17__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__16__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 20.95 0.51 21.05 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__16__Q

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 359 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 359 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 359 8.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 11.745 359 12.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 15.745 359 16.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 19.745 359 20.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 23.745 359 24.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 27.745 359 28.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 31.745 359 32.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 35.745 359 36.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 39.745 359 40.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 43.745 359 44.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 47.745 359 48.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 51.745 359 52.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 55.745 359 56.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 59.745 359 60.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 63.745 359 64.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 67.745 359 68.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 71.745 359 72.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 75.745 359 76.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 79.745 359 80.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 83.745 359 84.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 87.745 359 88.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 91.745 359 92.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 95.745 359 96.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 99.745 359 100.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 103.745 359 104.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 107.745 359 108.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 111.745 359 112.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 115.745 359 116.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 119.745 359 120.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 123.745 359 124.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 127.745 359 128.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 131.745 359 132.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 135.745 359 136.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 139.745 359 140.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 143.745 359 144.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 147.745 359 148.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 151.745 359 152.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 359 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 359 6.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 9.745 359 10.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 13.745 359 14.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 17.745 359 18.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 21.745 359 22.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 25.745 359 26.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 29.745 359 30.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 33.745 359 34.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 37.745 359 38.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 41.745 359 42.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 45.745 359 46.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 49.745 359 50.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 53.745 359 54.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 57.745 359 58.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 61.745 359 62.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 65.745 359 66.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 69.745 359 70.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 73.745 359 74.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 77.745 359 78.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 81.745 359 82.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 85.745 359 86.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 89.745 359 90.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 93.745 359 94.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 97.745 359 98.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 101.745 359 102.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 105.745 359 106.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 109.745 359 110.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 113.745 359 114.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 117.745 359 118.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 121.745 359 122.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 125.745 359 126.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 129.745 359 130.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 133.745 359 134.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 137.745 359 138.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 141.745 359 142.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 145.745 359 146.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 149.745 359 150.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 153.745 359 154.255 ;
      END
   END vdd

   OBS
      LAYER metal1 ;
         RECT 0 0 359 154 ;
   END
   OBS
      LAYER metal2 ;
         RECT 0 0 359 154 ;
   END
   OBS
      LAYER metal3 ;
         RECT 0 0 359 154 ;
   END
   OBS
      LAYER metal4 ;
         RECT 0 0 359 154 ;
   END
   OBS
      LAYER metal5 ;
         RECT 0 0 359 154 ;
   END
END h5

MACRO h3
   CLASS BLOCK ;
   SIZE 356.4 BY 178 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   PIN FE_OFN1630_n_9862
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 85.85 177.49 85.95 178 ;
      END
   END FE_OFN1630_n_9862

   PIN FE_OFN199_n_9228
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 46.5 0.255 46.7 ;
      END
   END FE_OFN199_n_9228

   PIN FE_RN_189_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 100.25 0 100.35 0.51 ;
      END
   END FE_RN_189_0

   PIN g57181_sb
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 34.85 0 34.95 0.51 ;
      END
   END g57181_sb

   PIN g57242_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 173.45 0 173.55 0.51 ;
      END
   END g57242_db

   PIN g57370_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 81.65 0 81.75 0.51 ;
      END
   END g57370_da

   PIN g57404_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 175.05 177.49 175.15 178 ;
      END
   END g57404_db

   PIN g57508_sb
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 95.05 0 95.15 0.51 ;
      END
   END g57508_sb

   PIN g57581_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 123.85 0 123.95 0.51 ;
      END
   END g57581_db

   PIN g57909_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 15.35 0.51 15.45 ;
      END
   END g57909_da

   PIN g57912_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 222.85 0 222.95 0.51 ;
      END
   END g57912_db

   PIN g58049_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 45.95 0.51 46.05 ;
      END
   END g58049_da

   PIN g58066_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 74.95 0.51 75.05 ;
      END
   END g58066_da

   PIN g58066_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 277.85 0 277.95 0.51 ;
      END
   END g58066_db

   PIN g58107_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 75.65 177.49 75.75 178 ;
      END
   END g58107_da

   PIN g58339_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 227.85 177.49 227.95 178 ;
      END
   END g58339_da

   PIN g58434_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 134.65 0 134.75 0.51 ;
      END
   END g58434_da

   PIN g58437_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 184.85 0 184.95 0.51 ;
      END
   END g58437_da

   PIN n_10060
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 161.05 0 161.15 0.51 ;
      END
   END n_10060

   PIN n_10608
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 121.25 0 121.35 0.51 ;
      END
   END n_10608

   PIN n_11362
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 255.45 0 255.55 0.51 ;
      END
   END n_11362

   PIN n_11544
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 250.25 0 250.35 0.51 ;
      END
   END n_11544

   PIN n_11582
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 276.25 0 276.35 0.51 ;
      END
   END n_11582

   PIN n_12129
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 75.05 0 75.15 0.51 ;
      END
   END n_12129

   PIN n_12140
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 21.05 0 21.15 0.51 ;
      END
   END n_12140

   PIN n_9427
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 116.85 177.49 116.95 178 ;
      END
   END n_9427

   PIN n_9435
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 64.25 177.49 64.35 178 ;
      END
   END n_9435

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__35__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 102.95 0.51 103.05 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__35__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__8__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 233.85 177.49 233.95 178 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__8__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__0__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 313.05 0 313.15 0.51 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__0__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__33__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 171.25 177.49 171.35 178 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__33__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__35__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 45.45 177.49 45.55 178 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__35__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__14__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 150.25 177.49 150.35 178 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__14__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__32__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 202.85 0 202.95 0.51 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__32__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__20__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 100.05 177.49 100.15 178 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__20__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__35__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 56.05 0 56.15 0.51 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__35__Q

   PIN wishbone_slave_unit_pcim_if_wbw_addr_data_in_393
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 107.05 0 107.15 0.51 ;
      END
   END wishbone_slave_unit_pcim_if_wbw_addr_data_in_393

   PIN wishbone_slave_unit_pcim_if_wbw_addr_data_in_397
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 133.15 0.51 133.25 ;
      END
   END wishbone_slave_unit_pcim_if_wbw_addr_data_in_397

   PIN wishbone_slave_unit_pcim_if_wbw_addr_data_in_398
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 163.15 0.51 163.25 ;
      END
   END wishbone_slave_unit_pcim_if_wbw_addr_data_in_398

   PIN wishbone_slave_unit_pcim_if_wbw_addr_data_in_403
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 46.15 0.51 46.25 ;
      END
   END wishbone_slave_unit_pcim_if_wbw_addr_data_in_403

   PIN FE_OCPN1936_n_15566
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 57.2 0 57.4 0.255 ;
      END
   END FE_OCPN1936_n_15566

   PIN FE_OCP_RBN2062_n_16572
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 98.45 0 98.55 0.51 ;
      END
   END FE_OCP_RBN2062_n_16572

   PIN FE_OFN1257_n_8567
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 271 0 271.2 0.255 ;
      END
   END FE_OFN1257_n_8567

   PIN FE_OFN1273_n_8567
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 73.9 0.255 74.1 ;
      END
   END FE_OFN1273_n_8567

   PIN FE_OFN1274_n_8567
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 356.145 102.9 356.4 103.1 ;
      END
   END FE_OFN1274_n_8567

   PIN FE_OFN1285_n_8567
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 74.3 0.255 74.5 ;
      END
   END FE_OFN1285_n_8567

   PIN FE_OFN1286_n_8567
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 144.2 177.745 144.4 178 ;
      END
   END FE_OFN1286_n_8567

   PIN FE_OFN1288_n_8567
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 163.8 177.745 164 178 ;
      END
   END FE_OFN1288_n_8567

   PIN FE_OFN1289_n_8567
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 35 0 35.2 0.255 ;
      END
   END FE_OFN1289_n_8567

   PIN FE_OFN1292_n_8567
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 95.2 0 95.4 0.255 ;
      END
   END FE_OFN1292_n_8567

   PIN FE_OFN1308_n_8567
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 7.5 0.255 7.7 ;
      END
   END FE_OFN1308_n_8567

   PIN FE_OFN1311_n_8567
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 231 0 231.2 0.255 ;
      END
   END FE_OFN1311_n_8567

   PIN FE_OFN1312_n_8567
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 356.145 132.9 356.4 133.1 ;
      END
   END FE_OFN1312_n_8567

   PIN FE_OFN1319_n_8567
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 124.2 0 124.4 0.255 ;
      END
   END FE_OFN1319_n_8567

   PIN FE_OFN1320_n_8567
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 238.4 177.745 238.6 178 ;
      END
   END FE_OFN1320_n_8567

   PIN FE_OFN1354_n_15558
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 122.05 0 122.15 0.51 ;
      END
   END FE_OFN1354_n_15558

   PIN FE_OFN1355_n_15558
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 99.05 0 99.15 0.51 ;
      END
   END FE_OFN1355_n_15558

   PIN FE_OFN1367_n_15587
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 85.05 0 85.15 0.51 ;
      END
   END FE_OFN1367_n_15587

   PIN FE_OFN1368_n_15587
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 63.45 0 63.55 0.51 ;
      END
   END FE_OFN1368_n_15587

   PIN FE_OFN1378_n_10853
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 207.65 0 207.75 0.51 ;
      END
   END FE_OFN1378_n_10853

   PIN FE_OFN1505_n_9531
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 25.25 177.49 25.35 178 ;
      END
   END FE_OFN1505_n_9531

   PIN FE_OFN1537_n_9428
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 105.65 0 105.75 0.51 ;
      END
   END FE_OFN1537_n_9428

   PIN FE_OFN1538_n_9428
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 183 0 183.2 0.255 ;
      END
   END FE_OFN1538_n_9428

   PIN FE_OFN1565_n_9477
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 356.145 44.9 356.4 45.1 ;
      END
   END FE_OFN1565_n_9477

   PIN FE_OFN1629_n_9862
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 86.05 177.49 86.15 178 ;
      END
   END FE_OFN1629_n_9862

   PIN FE_OFN1677_n_10588
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 207.05 0 207.15 0.51 ;
      END
   END FE_OFN1677_n_10588

   PIN FE_OFN1685_n_16891
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 85.65 0 85.75 0.51 ;
      END
   END FE_OFN1685_n_16891

   PIN FE_OFN1688_n_15534
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 210.05 177.49 210.15 178 ;
      END
   END FE_OFN1688_n_15534

   PIN FE_OFN1693_n_16992
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 210.65 177.49 210.75 178 ;
      END
   END FE_OFN1693_n_16992

   PIN FE_OFN198_n_9228
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 45.75 0.51 45.85 ;
      END
   END FE_OFN198_n_9228

   PIN FE_OFN201_n_9140
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 263 177.745 263.2 178 ;
      END
   END FE_OFN201_n_9140

   PIN FE_OFN203_n_9865
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 356.145 45.3 356.4 45.5 ;
      END
   END FE_OFN203_n_9865

   PIN FE_OFN210_n_9858
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 239.25 0 239.35 0.51 ;
      END
   END FE_OFN210_n_9858

   PIN FE_OFN212_n_9124
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 145.4 0 145.6 0.255 ;
      END
   END FE_OFN212_n_9124

   PIN FE_OFN216_n_9889
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 14.9 0.255 15.1 ;
      END
   END FE_OFN216_n_9889

   PIN FE_OFN254_n_9868
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 82 177.745 82.2 178 ;
      END
   END FE_OFN254_n_9868

   PIN FE_OFN268_n_9884
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 45.3 0.255 45.5 ;
      END
   END FE_OFN268_n_9884

   PIN FE_OFN539_n_9895
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 356.145 74.7 356.4 74.9 ;
      END
   END FE_OFN539_n_9895

   PIN FE_OFN548_n_9502
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 219.2 0 219.4 0.255 ;
      END
   END FE_OFN548_n_9502

   PIN FE_OFN554_n_9902
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 231.4 0 231.6 0.255 ;
      END
   END FE_OFN554_n_9902

   PIN FE_OFN560_n_9531
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 82.4 177.745 82.6 178 ;
      END
   END FE_OFN560_n_9531

   PIN FE_OFN571_n_9694
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 15.7 0.255 15.9 ;
      END
   END FE_OFN571_n_9694

   PIN FE_OFN572_n_9694
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 274.8 177.745 275 178 ;
      END
   END FE_OFN572_n_9694

   PIN FE_OFN576_n_9687
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 103.3 0.255 103.5 ;
      END
   END FE_OFN576_n_9687

   PIN FE_OFN580_n_9904
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 278.2 0 278.4 0.255 ;
      END
   END FE_OFN580_n_9904

   PIN FE_OFN581_n_9904
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 75.2 0 75.4 0.255 ;
      END
   END FE_OFN581_n_9904

   PIN g57213_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 250.65 0 250.75 0.51 ;
      END
   END g57213_db

   PIN g57221_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 119.05 177.49 119.15 178 ;
      END
   END g57221_da

   PIN g57544_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 55.45 177.49 55.55 178 ;
      END
   END g57544_da

   PIN g57944_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 355.89 103.35 356.4 103.45 ;
      END
   END g57944_da

   PIN g58060_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 124.45 0 124.55 0.51 ;
      END
   END g58060_da

   PIN g58073_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 237.25 0 237.35 0.51 ;
      END
   END g58073_db

   PIN g58333_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 77.65 177.49 77.75 178 ;
      END
   END g58333_da

   PIN g58333_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 77.85 177.49 77.95 178 ;
      END
   END g58333_db

   PIN g58341_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 330.45 0 330.55 0.51 ;
      END
   END g58341_sb

   PIN g58402_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 64.65 177.49 64.75 178 ;
      END
   END g58402_db

   PIN g58438_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 201.05 0 201.15 0.51 ;
      END
   END g58438_db

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 46.9 0.255 47.1 ;
      END
   END ispd_clk

   PIN n_10002
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 21.65 0 21.75 0.51 ;
      END
   END n_10002

   PIN n_11259
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 234.85 177.49 234.95 178 ;
      END
   END n_11259

   PIN n_11337
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 162.85 177.49 162.95 178 ;
      END
   END n_11337

   PIN n_11516
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 186.25 177.49 186.35 178 ;
      END
   END n_11516

   PIN n_12841
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 44.95 0.51 45.05 ;
      END
   END n_12841

   PIN n_12847
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 162.95 0.51 163.05 ;
      END
   END n_12847

   PIN n_12848
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 132.95 0.51 133.05 ;
      END
   END n_12848

   PIN n_12852
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 108.05 0 108.15 0.51 ;
      END
   END n_12852

   PIN n_16840
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 21.25 0 21.35 0.51 ;
      END
   END n_16840

   PIN n_16841
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 22.25 0 22.35 0.51 ;
      END
   END n_16841

   PIN n_9551
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 245.25 0 245.35 0.51 ;
      END
   END n_9551

   PIN n_9726
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 259.85 0 259.95 0.51 ;
      END
   END n_9726

   PIN n_9868
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 182.85 0 182.95 0.51 ;
      END
   END n_9868

   PIN n_9908
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 74.75 0.51 74.85 ;
      END
   END n_9908

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__34__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 63.65 0 63.75 0.51 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__34__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__8__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 86.05 0 86.15 0.51 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__8__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__8__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 42.65 0 42.75 0.51 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__8__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__0__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 297.45 0 297.55 0.51 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__0__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__28__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 162.25 0 162.35 0.51 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__28__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__10__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 113.45 0 113.55 0.51 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__10__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__28__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 134.85 0 134.95 0.51 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__28__Q

   PIN wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__1__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 265.85 0 265.95 0.51 ;
      END
   END wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__1__Q

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 356.4 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 356.4 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 356.4 8.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 11.745 356.4 12.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 15.745 356.4 16.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 19.745 356.4 20.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 23.745 356.4 24.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 27.745 356.4 28.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 31.745 356.4 32.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 35.745 356.4 36.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 39.745 356.4 40.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 43.745 356.4 44.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 47.745 356.4 48.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 51.745 356.4 52.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 55.745 356.4 56.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 59.745 356.4 60.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 63.745 356.4 64.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 67.745 356.4 68.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 71.745 356.4 72.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 75.745 356.4 76.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 79.745 356.4 80.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 83.745 356.4 84.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 87.745 356.4 88.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 91.745 356.4 92.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 95.745 356.4 96.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 99.745 356.4 100.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 103.745 356.4 104.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 107.745 356.4 108.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 111.745 356.4 112.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 115.745 356.4 116.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 119.745 356.4 120.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 123.745 356.4 124.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 127.745 356.4 128.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 131.745 356.4 132.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 135.745 356.4 136.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 139.745 356.4 140.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 143.745 356.4 144.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 147.745 356.4 148.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 151.745 356.4 152.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 155.745 356.4 156.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 159.745 356.4 160.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 163.745 356.4 164.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 167.745 356.4 168.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 171.745 356.4 172.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 175.745 356.4 176.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 356.4 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 356.4 6.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 9.745 356.4 10.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 13.745 356.4 14.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 17.745 356.4 18.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 21.745 356.4 22.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 25.745 356.4 26.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 29.745 356.4 30.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 33.745 356.4 34.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 37.745 356.4 38.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 41.745 356.4 42.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 45.745 356.4 46.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 49.745 356.4 50.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 53.745 356.4 54.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 57.745 356.4 58.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 61.745 356.4 62.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 65.745 356.4 66.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 69.745 356.4 70.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 73.745 356.4 74.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 77.745 356.4 78.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 81.745 356.4 82.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 85.745 356.4 86.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 89.745 356.4 90.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 93.745 356.4 94.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 97.745 356.4 98.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 101.745 356.4 102.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 105.745 356.4 106.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 109.745 356.4 110.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 113.745 356.4 114.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 117.745 356.4 118.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 121.745 356.4 122.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 125.745 356.4 126.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 129.745 356.4 130.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 133.745 356.4 134.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 137.745 356.4 138.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 141.745 356.4 142.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 145.745 356.4 146.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 149.745 356.4 150.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 153.745 356.4 154.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 157.745 356.4 158.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 161.745 356.4 162.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 165.745 356.4 166.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 169.745 356.4 170.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 173.745 356.4 174.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 177.745 356.4 178.255 ;
      END
   END vdd

   OBS
      LAYER metal1 ;
         RECT 0 0 356.4 178 ;
   END
   OBS
      LAYER metal2 ;
         RECT 0 0 356.4 178 ;
   END
   OBS
      LAYER metal3 ;
         RECT 0 0 356.4 178 ;
   END
   OBS
      LAYER metal4 ;
         RECT 0 0 356.4 178 ;
   END
   OBS
      LAYER metal5 ;
         RECT 0 0 356.4 178 ;
   END
END h3

MACRO h2
   CLASS BLOCK ;
   SIZE 360.6 BY 178 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   PIN FE_OCP_RBN2122_n_16966
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 15.55 0.51 15.65 ;
      END
   END FE_OCP_RBN2122_n_16966

   PIN FE_OFN741_n_2678
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 225.85 0 225.95 0.51 ;
      END
   END FE_OFN741_n_2678

   PIN FE_OFN752_n_2547
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 55.65 0 55.75 0.51 ;
      END
   END FE_OFN752_n_2547

   PIN FE_RN_232_0
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 360.09 162.75 360.6 162.85 ;
      END
   END FE_RN_232_0

   PIN configuration_pci_err_addr_471
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 139.65 0 139.75 0.51 ;
      END
   END configuration_pci_err_addr_471

   PIN configuration_sync_cache_lsize_to_wb_bits_reg_3__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 360.09 45.15 360.6 45.25 ;
      END
   END configuration_sync_cache_lsize_to_wb_bits_reg_3__Q

   PIN g53255_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 46.65 0 46.75 0.51 ;
      END
   END g53255_p

   PIN g53301_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 110.85 177.49 110.95 178 ;
      END
   END g53301_p

   PIN g61965_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 162.55 0.51 162.65 ;
      END
   END g61965_da

   PIN g62827_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 56.65 177.49 56.75 178 ;
      END
   END g62827_da

   PIN g62837_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 132.95 0.51 133.05 ;
      END
   END g62837_da

   PIN g62837_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 133.15 0.51 133.25 ;
      END
   END g62837_db

   PIN g63077_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 87.85 0 87.95 0.51 ;
      END
   END g63077_da

   PIN g63080_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 72.55 0.51 72.65 ;
      END
   END g63080_db

   PIN g63568_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 37.65 177.49 37.75 178 ;
      END
   END g63568_db

   PIN g64259_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 45.15 0.51 45.25 ;
      END
   END g64259_db

   PIN g64259_sb
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 103.35 0.51 103.45 ;
      END
   END g64259_sb

   PIN g64301_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 61.05 177.49 61.15 178 ;
      END
   END g64301_db

   PIN g64332_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 42.95 0.51 43.05 ;
      END
   END g64332_db

   PIN g64332_sb
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 45.35 0.51 45.45 ;
      END
   END g64332_sb

   PIN g65212_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 293.65 0 293.75 0.51 ;
      END
   END g65212_da

   PIN g65234_sb
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 216.85 0 216.95 0.51 ;
      END
   END g65234_sb

   PIN g65240_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 181.65 0 181.75 0.51 ;
      END
   END g65240_db

   PIN g66184_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 360.09 103.95 360.6 104.05 ;
      END
   END g66184_p

   PIN g66726_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 360.09 14.95 360.6 15.05 ;
      END
   END g66726_p

   PIN n_10825
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 220.25 0 220.35 0.51 ;
      END
   END n_10825

   PIN n_1159
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 260.25 0 260.35 0.51 ;
      END
   END n_1159

   PIN n_1196
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 360.09 102.95 360.6 103.05 ;
      END
   END n_1196

   PIN n_13304
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 114.05 0 114.15 0.51 ;
      END
   END n_13304

   PIN n_13701
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 31.65 0 31.75 0.51 ;
      END
   END n_13701

   PIN n_13859
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 70.05 0 70.15 0.51 ;
      END
   END n_13859

   PIN n_13980
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 98.45 177.49 98.55 178 ;
      END
   END n_13980

   PIN n_14413
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 85.85 177.49 85.95 178 ;
      END
   END n_14413

   PIN n_14690
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 162.25 177.49 162.35 178 ;
      END
   END n_14690

   PIN n_14804
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 143.25 177.49 143.35 178 ;
      END
   END n_14804

   PIN n_1507
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 176.45 177.49 176.55 178 ;
      END
   END n_1507

   PIN n_1552
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 360.09 104.15 360.6 104.25 ;
      END
   END n_1552

   PIN n_15611
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 252.05 0 252.15 0.51 ;
      END
   END n_15611

   PIN n_16275
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 290.45 177.49 290.55 178 ;
      END
   END n_16275

   PIN n_16280
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 234.45 0 234.55 0.51 ;
      END
   END n_16280

   PIN n_16507
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 205.45 0 205.55 0.51 ;
      END
   END n_16507

   PIN n_16748
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 108.2 0 108.4 0.255 ;
      END
   END n_16748

   PIN n_16975
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 15.75 0.51 15.85 ;
      END
   END n_16975

   PIN n_177
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 284.65 0 284.75 0.51 ;
      END
   END n_177

   PIN n_2597
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 206.65 0 206.75 0.51 ;
      END
   END n_2597

   PIN n_2598
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 209.45 0 209.55 0.51 ;
      END
   END n_2598

   PIN n_2729
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 258.05 0 258.15 0.51 ;
      END
   END n_2729

   PIN n_2776
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 125.45 0 125.55 0.51 ;
      END
   END n_2776

   PIN n_3123
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 360.09 103.35 360.6 103.45 ;
      END
   END n_3123

   PIN n_3319
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 214.45 0 214.55 0.51 ;
      END
   END n_3319

   PIN n_3320
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 193.65 0 193.75 0.51 ;
      END
   END n_3320

   PIN n_8498
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 300.65 0 300.75 0.51 ;
      END
   END n_8498

   PIN n_8757
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 147.2 0 147.4 0.255 ;
      END
   END n_8757

   PIN n_8759
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 102.65 0 102.75 0.51 ;
      END
   END n_8759

   PIN n_8800
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 288.45 177.49 288.55 178 ;
      END
   END n_8800

   PIN n_8879
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 146.85 0 146.95 0.51 ;
      END
   END n_8879

   PIN n_9175
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 360.09 75.35 360.6 75.45 ;
      END
   END n_9175

   PIN pci_target_unit_fifos_pciw_addr_data_in_121
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 103.55 0.51 103.65 ;
      END
   END pci_target_unit_fifos_pciw_addr_data_in_121

   PIN pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__35__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 102.95 0.51 103.05 ;
      END
   END pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__35__Q

   PIN pci_target_unit_pcit_if_strd_bc_in
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 270.45 177.49 270.55 178 ;
      END
   END pci_target_unit_pcit_if_strd_bc_in

   PIN pci_target_unit_pcit_if_strd_bc_in_718
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 203.05 177.49 203.15 178 ;
      END
   END pci_target_unit_pcit_if_strd_bc_in_718

   PIN pci_target_unit_pcit_if_strd_bc_in_719
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 166.45 0 166.55 0.51 ;
      END
   END pci_target_unit_pcit_if_strd_bc_in_719

   PIN wbm_sel_o_0_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 68.55 0.51 68.65 ;
      END
   END wbm_sel_o_0_

   PIN wbm_sel_o_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 103.75 0.51 103.85 ;
      END
   END wbm_sel_o_3_

   PIN FE_OCP_RBN2123_n_16966
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 15.95 0.51 16.05 ;
      END
   END FE_OCP_RBN2123_n_16966

   PIN FE_OFN1017_g64577_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 72.1 0.255 72.3 ;
      END
   END FE_OFN1017_g64577_p

   PIN FE_OFN1019_g64577_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 101.6 177.745 101.8 178 ;
      END
   END FE_OFN1019_g64577_p

   PIN FE_OFN1112_n_3476
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 119.8 0 120 0.255 ;
      END
   END FE_OFN1112_n_3476

   PIN FE_OFN1463_n_13736
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 96.85 0 96.95 0.51 ;
      END
   END FE_OFN1463_n_13736

   PIN FE_OFN1520_n_4730
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 66.4 177.745 66.6 178 ;
      END
   END FE_OFN1520_n_4730

   PIN FE_OFN1776_n_13971
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 98.6 177.745 98.8 178 ;
      END
   END FE_OFN1776_n_13971

   PIN FE_OFN189_n_1193
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 301.25 177.49 301.35 178 ;
      END
   END FE_OFN189_n_1193

   PIN FE_OFN747_n_2678
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 186.4 0 186.6 0.255 ;
      END
   END FE_OFN747_n_2678

   PIN FE_OFN751_n_2547
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 55.85 0 55.95 0.51 ;
      END
   END FE_OFN751_n_2547

   PIN FE_OFN860_n_4734
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 133.7 0.255 133.9 ;
      END
   END FE_OFN860_n_4734

   PIN FE_OFN959_n_16760
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 110.45 0 110.55 0.51 ;
      END
   END FE_OFN959_n_16760

   PIN FE_OFN973_n_4727
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 44.5 0.255 44.7 ;
      END
   END FE_OFN973_n_4727

   PIN FE_RN_285_0
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 234.65 0 234.75 0.51 ;
      END
   END FE_RN_285_0

   PIN FE_RN_286_0
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 234.85 0 234.95 0.51 ;
      END
   END FE_RN_286_0

   PIN FE_RN_345_0
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 311.65 0 311.75 0.51 ;
      END
   END FE_RN_345_0

   PIN FE_RN_427_0
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 119.85 177.49 119.95 178 ;
      END
   END FE_RN_427_0

   PIN configuration_meta_cache_lsize_to_wb_bits_926
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 360.09 44.95 360.6 45.05 ;
      END
   END configuration_meta_cache_lsize_to_wb_bits_926

   PIN configuration_sync_cache_lsize_to_wb_bits_reg_2__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 244.65 0 244.75 0.51 ;
      END
   END configuration_sync_cache_lsize_to_wb_bits_reg_2__Q

   PIN g60615_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 158.45 0 158.55 0.51 ;
      END
   END g60615_db

   PIN g63564_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 161.45 177.49 161.55 178 ;
      END
   END g63564_sb

   PIN g65215_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 227.65 177.49 227.75 178 ;
      END
   END g65215_da

   PIN g65225_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 220.65 177.49 220.75 178 ;
      END
   END g65225_da

   PIN g65234_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 227.25 0 227.35 0.51 ;
      END
   END g65234_da

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 140 0 140.2 0.255 ;
      END
   END ispd_clk

   PIN n_1219
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 176.65 177.49 176.75 178 ;
      END
   END n_1219

   PIN n_1304
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 360.09 133.15 360.6 133.25 ;
      END
   END n_1304

   PIN n_13122
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 114.25 0 114.35 0.51 ;
      END
   END n_13122

   PIN n_13484
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 134.25 0 134.35 0.51 ;
      END
   END n_13484

   PIN n_1366
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 360.09 103.15 360.6 103.25 ;
      END
   END n_1366

   PIN n_13919
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 322.05 177.49 322.15 178 ;
      END
   END n_13919

   PIN n_13955
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 46.85 0 46.95 0.51 ;
      END
   END n_13955

   PIN n_13971
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 123.25 177.49 123.35 178 ;
      END
   END n_13971

   PIN n_1435
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 360.09 75.15 360.6 75.25 ;
      END
   END n_1435

   PIN n_14529
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 301.05 177.49 301.15 178 ;
      END
   END n_14529

   PIN n_14829
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 134.05 0 134.15 0.51 ;
      END
   END n_14829

   PIN n_14837
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 102.85 0 102.95 0.51 ;
      END
   END n_14837

   PIN n_14895
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 133.65 0 133.75 0.51 ;
      END
   END n_14895

   PIN n_14897
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 72.75 0.51 72.85 ;
      END
   END n_14897

   PIN n_15114
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 32.25 0 32.35 0.51 ;
      END
   END n_15114

   PIN n_1513
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 279.45 0 279.55 0.51 ;
      END
   END n_1513

   PIN n_15292
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 323.45 0 323.55 0.51 ;
      END
   END n_15292

   PIN n_15302
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 258.45 0 258.55 0.51 ;
      END
   END n_15302

   PIN n_1551
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 360.09 103.75 360.6 103.85 ;
      END
   END n_1551

   PIN n_15607
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 278.85 0 278.95 0.51 ;
      END
   END n_15607

   PIN n_16205
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 32.45 0 32.55 0.51 ;
      END
   END n_16205

   PIN n_16331
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 360.09 103.55 360.6 103.65 ;
      END
   END n_16331

   PIN n_16738
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 108.45 0 108.55 0.51 ;
      END
   END n_16738

   PIN n_16966
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 15.35 0.51 15.45 ;
      END
   END n_16966

   PIN n_16970
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 15.15 0.51 15.25 ;
      END
   END n_16970

   PIN n_16974
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 14.95 0.51 15.05 ;
      END
   END n_16974

   PIN n_2031
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 258.25 0 258.35 0.51 ;
      END
   END n_2031

   PIN n_2301
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 360.345 74.1 360.6 74.3 ;
      END
   END n_2301

   PIN n_2337
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 302.85 0 302.95 0.51 ;
      END
   END n_2337

   PIN n_2353
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 297.85 0 297.95 0.51 ;
      END
   END n_2353

   PIN n_2599
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 176.65 0 176.75 0.51 ;
      END
   END n_2599

   PIN n_2675
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 293.85 0 293.95 0.51 ;
      END
   END n_2675

   PIN n_2677
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 167.45 0 167.55 0.51 ;
      END
   END n_2677

   PIN n_2678
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 268.65 0 268.75 0.51 ;
      END
   END n_2678

   PIN n_2730
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 125.65 0 125.75 0.51 ;
      END
   END n_2730

   PIN n_2779
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 360.09 74.95 360.6 75.05 ;
      END
   END n_2779

   PIN n_4592
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 162.75 0.51 162.85 ;
      END
   END n_4592

   PIN n_5092
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 103.15 0.51 103.25 ;
      END
   END n_5092

   PIN n_657
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 341.85 0 341.95 0.51 ;
      END
   END n_657

   PIN n_7698
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 360.09 132.95 360.6 133.05 ;
      END
   END n_7698

   PIN n_8487
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 332.85 0 332.95 0.51 ;
      END
   END n_8487

   PIN n_8538
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 298.25 0 298.35 0.51 ;
      END
   END n_8538

   PIN n_8819
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 279.25 0 279.35 0.51 ;
      END
   END n_8819

   PIN n_9178
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 318.85 177.49 318.95 178 ;
      END
   END n_9178

   PIN output_backup_trdy_out_reg_Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 192.65 0 192.75 0.51 ;
      END
   END output_backup_trdy_out_reg_Q

   PIN parchk_pci_ad_reg_in
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 263.65 177.49 263.75 178 ;
      END
   END parchk_pci_ad_reg_in

   PIN parchk_pci_ad_reg_in_1205
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 243.45 0 243.55 0.51 ;
      END
   END parchk_pci_ad_reg_in_1205

   PIN pci_target_unit_del_sync_bc_in
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 233.25 177.49 233.35 178 ;
      END
   END pci_target_unit_del_sync_bc_in

   PIN pci_target_unit_del_sync_be_out_reg_3__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 181.85 0 181.95 0.51 ;
      END
   END pci_target_unit_del_sync_be_out_reg_3__Q

   PIN pci_target_unit_fifos_pciw_addr_data_in_123
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 61.25 177.49 61.35 178 ;
      END
   END pci_target_unit_fifos_pciw_addr_data_in_123

   PIN pci_target_unit_fifos_pciw_addr_data_in_126
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 44.95 0.51 45.05 ;
      END
   END pci_target_unit_fifos_pciw_addr_data_in_126

   PIN pci_target_unit_fifos_pciw_cbe_in
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 43.15 0.51 43.25 ;
      END
   END pci_target_unit_fifos_pciw_cbe_in

   PIN pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__1__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 70.45 0 70.55 0.51 ;
      END
   END pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__1__Q

   PIN pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__32__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 56.85 0 56.95 0.51 ;
      END
   END pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__32__Q

   PIN pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__3__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 83.45 0 83.55 0.51 ;
      END
   END pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__3__Q

   PIN pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__6__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 96.65 0 96.75 0.51 ;
      END
   END pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__6__Q

   PIN pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__32__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 133.35 0.51 133.45 ;
      END
   END pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__32__Q

   PIN pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__3__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 75.65 177.49 75.75 178 ;
      END
   END pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__3__Q

   PIN pci_target_unit_pcit_if_req_req_pending_in
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 341.65 0 341.75 0.51 ;
      END
   END pci_target_unit_pcit_if_req_req_pending_in

   PIN pci_target_unit_pcit_if_strd_bc_in_717
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 290.25 177.49 290.35 178 ;
      END
   END pci_target_unit_pcit_if_strd_bc_in_717

   PIN pci_target_unit_wbm_sm_pciw_fifo_addr_data_in
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 124.65 177.49 124.75 178 ;
      END
   END pci_target_unit_wbm_sm_pciw_fifo_addr_data_in

   PIN pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_50
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 163.45 177.49 163.55 178 ;
      END
   END pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_50

   PIN pciu_cache_lsize_not_zero_in
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 205.85 0 205.95 0.51 ;
      END
   END pciu_cache_lsize_not_zero_in

   PIN wbm_adr_o_0_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 92.45 0 92.55 0.51 ;
      END
   END wbm_adr_o_0_

   PIN wbm_adr_o_1_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 122.55 0.51 122.65 ;
      END
   END wbm_adr_o_1_

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 360.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 360.6 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 360.6 8.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 11.745 360.6 12.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 15.745 360.6 16.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 19.745 360.6 20.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 23.745 360.6 24.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 27.745 360.6 28.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 31.745 360.6 32.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 35.745 360.6 36.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 39.745 360.6 40.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 43.745 360.6 44.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 47.745 360.6 48.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 51.745 360.6 52.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 55.745 360.6 56.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 59.745 360.6 60.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 63.745 360.6 64.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 67.745 360.6 68.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 71.745 360.6 72.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 75.745 360.6 76.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 79.745 360.6 80.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 83.745 360.6 84.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 87.745 360.6 88.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 91.745 360.6 92.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 95.745 360.6 96.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 99.745 360.6 100.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 103.745 360.6 104.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 107.745 360.6 108.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 111.745 360.6 112.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 115.745 360.6 116.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 119.745 360.6 120.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 123.745 360.6 124.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 127.745 360.6 128.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 131.745 360.6 132.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 135.745 360.6 136.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 139.745 360.6 140.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 143.745 360.6 144.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 147.745 360.6 148.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 151.745 360.6 152.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 155.745 360.6 156.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 159.745 360.6 160.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 163.745 360.6 164.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 167.745 360.6 168.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 171.745 360.6 172.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 175.745 360.6 176.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 360.6 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 360.6 6.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 9.745 360.6 10.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 13.745 360.6 14.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 17.745 360.6 18.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 21.745 360.6 22.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 25.745 360.6 26.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 29.745 360.6 30.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 33.745 360.6 34.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 37.745 360.6 38.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 41.745 360.6 42.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 45.745 360.6 46.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 49.745 360.6 50.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 53.745 360.6 54.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 57.745 360.6 58.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 61.745 360.6 62.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 65.745 360.6 66.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 69.745 360.6 70.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 73.745 360.6 74.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 77.745 360.6 78.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 81.745 360.6 82.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 85.745 360.6 86.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 89.745 360.6 90.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 93.745 360.6 94.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 97.745 360.6 98.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 101.745 360.6 102.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 105.745 360.6 106.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 109.745 360.6 110.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 113.745 360.6 114.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 117.745 360.6 118.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 121.745 360.6 122.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 125.745 360.6 126.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 129.745 360.6 130.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 133.745 360.6 134.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 137.745 360.6 138.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 141.745 360.6 142.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 145.745 360.6 146.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 149.745 360.6 150.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 153.745 360.6 154.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 157.745 360.6 158.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 161.745 360.6 162.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 165.745 360.6 166.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 169.745 360.6 170.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 173.745 360.6 174.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 177.745 360.6 178.255 ;
      END
   END vdd

   OBS
      LAYER metal1 ;
         RECT 0 0 360.6 178 ;
   END
   OBS
      LAYER metal2 ;
         RECT 0 0 360.6 178 ;
   END
   OBS
      LAYER metal3 ;
         RECT 0 0 360.6 178 ;
   END
   OBS
      LAYER metal4 ;
         RECT 0 0 360.6 178 ;
   END
   OBS
      LAYER metal5 ;
         RECT 0 0 360.6 178 ;
   END
END h2

MACRO ms00f80
   CLASS CORE ;
   SIZE 1.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN ck
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END ck

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.05 0.5 1.15 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.6 2.255 ;
      END
   END vdd

END ms00f80

MACRO in01f01
   CLASS CORE ;
   SIZE 0.4 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 0.4 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 0.4 2.255 ;
      END
   END vdd

END in01f01

MACRO no02f01
   CLASS CORE ;
   SIZE 0.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 0.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 0.8 2.255 ;
      END
   END vdd

END no02f01

MACRO na02f01
   CLASS CORE ;
   SIZE 0.8 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END b

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 0.8 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 0.8 2.255 ;
      END
   END vdd

END na02f01

MACRO ao12f01
   CLASS CORE ;
   SIZE 1.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
   END vdd

END ao12f01

MACRO na03f01
   CLASS CORE ;
   SIZE 1.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
   END vdd

END na03f01

MACRO oa12f01
   CLASS CORE ;
   SIZE 1.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
   END vdd

END oa12f01

MACRO na04m01
   CLASS CORE ;
   SIZE 1.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.6 2.255 ;
      END
   END vdd

END na04m01

MACRO no04s01
   CLASS CORE ;
   SIZE 1.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.6 2.255 ;
      END
   END vdd

END no04s01

MACRO no03m01
   CLASS CORE ;
   SIZE 1.2 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.2 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.2 2.255 ;
      END
   END vdd

END no03m01

MACRO ao22s01
   CLASS CORE ;
   SIZE 1.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.6 2.255 ;
      END
   END vdd

END ao22s01

MACRO oa22f01
   CLASS CORE ;
   SIZE 1.6 BY 2 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 1.35 0.95 1.55 1.05 ;
         LAYER metal2 ;
             RECT 1.25 0.5 1.35 1.05 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END d

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 1.6 0.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 1.6 2.255 ;
      END
   END vdd

END oa22f01

MACRO in01f01X2HE
   CLASS CORE ;
   SIZE 3.6 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 3.6 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.6 2.255 ;
      END
   END vdd

END in01f01X2HE

MACRO in01f01X2HO
   CLASS CORE ;
   SIZE 3.6 BY 4 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 3.6 4.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.6 2.255 ;
      END
   END vss

END in01f01X2HO

MACRO in01f01X3H
   CLASS CORE ;
   SIZE 3.6 BY 6 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 4.5 1.75 5.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 0.5 1.95 1.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 3.6 4.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.6 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 3.6 6.255 ;
      END
   END vdd

END in01f01X3H

MACRO in01f01X4HE
   CLASS CORE ;
   SIZE 3.6 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 4.5 1.95 5.5 ;
      END
   END a

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 3.6 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 3.6 8.255 ;
      END
   END vss

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.6 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 3.6 6.255 ;
      END
   END vdd

END in01f01X4HE

MACRO in01f01X4HO
   CLASS CORE ;
   SIZE 3.6 BY 8 ;
   ORIGIN 0 0 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.65 0.5 1.75 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.85 4.5 1.95 5.5 ;
      END
   END a

   PIN vdd
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT 
         LAYER metal1 ;
             RECT 0 -0.255 3.6 0.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 3.745 3.6 4.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 7.745 3.6 8.255 ;
      END
   END vdd

   PIN vss
      DIRECTION INOUT ;
      USE GROUND ;
      PORT 
         LAYER metal1 ;
             RECT 0 1.745 3.6 2.255 ;
      END
      PORT 
         LAYER metal1 ;
             RECT 0 5.745 3.6 6.255 ;
      END
   END vss

END in01f01X4HO

END LIBRARY
