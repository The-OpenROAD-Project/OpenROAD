VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MANUFACTURINGGRID 0.0025 ;

MACRO NOP
  ORIGIN 0 0 ;
  OBS
    LAYER metal1 DESIGNRULEWIDTH 0.065 ;
    WIDTH 0.03 ;
      PATH 0.05 0.59 0.07 0.59 ;
  END 
END NOP
END LIBRARY