# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_io__overlay_vssio_lvc
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 198 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 51.125000 1.270000 54.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.125000 75.000000 54.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 46.365000 1.270000 49.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 46.365000 75.000000 49.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 6.885000 1.270000 11.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 6.885000 75.000000 11.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 6.985000 1.270000 11.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 6.985000 75.000000 11.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 0.035000 1.270000 5.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 0.035000 75.000000 5.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 0.135000 1.270000 5.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 0.135000 75.000000 5.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 12.935000 0.965000 16.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035000 12.935000 75.000000 16.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 13.035000 0.965000 16.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 13.035000 75.000000 16.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 17.785000 1.270000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 68.035000 1.270000 93.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 17.785000 75.000000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 68.035000 75.000000 93.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 17.885000 1.270000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 68.035000 1.270000 92.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 17.885000 75.000000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 68.035000 75.000000 92.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 62.085000 1.270000 66.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 62.085000 75.000000 66.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 62.185000 1.270000 66.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 62.185000 75.000000 66.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 34.735000 1.270000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 45.735000 1.270000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 49.645000 1.270000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 54.405000 1.270000 54.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 34.735000 75.000000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 45.735000 75.000000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 49.645000 75.000000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 54.405000 75.000000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 34.840000 1.270000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 45.735000 1.270000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 34.840000 75.000000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 45.735000 75.000000 54.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 39.585000 1.270000 44.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 39.585000 75.000000 44.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 39.685000 1.270000 44.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 39.685000 75.000000 44.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.500000 171.195000 12.900000 198.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.500000 23.840000 24.400000 28.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755000 23.840000 74.290000 28.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.045000 171.195000 74.700000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 173.785000  1.270000 173.835000 ;
        RECT 0.000000 173.835000 12.900000 197.970000 ;
        RECT 0.000000 197.970000  1.270000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 23.835000 24.375000 28.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.780000 23.835000 75.000000 28.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 62.075000 173.835000 75.000000 197.970000 ;
        RECT 73.730000 173.785000 75.000000 173.835000 ;
        RECT 73.730000 197.970000 75.000000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 23.935000 1.270000 28.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 23.935000 75.000000 28.385000 ;
    END
    PORT
      LAYER via3 ;
        RECT  0.590000  23.910000  0.790000  24.110000 ;
        RECT  0.590000  24.340000  0.790000  24.540000 ;
        RECT  0.590000  24.770000  0.790000  24.970000 ;
        RECT  0.590000  25.200000  0.790000  25.400000 ;
        RECT  0.590000  25.630000  0.790000  25.830000 ;
        RECT  0.590000  26.060000  0.790000  26.260000 ;
        RECT  0.590000  26.490000  0.790000  26.690000 ;
        RECT  0.590000  26.920000  0.790000  27.120000 ;
        RECT  0.590000  27.350000  0.790000  27.550000 ;
        RECT  0.590000  27.780000  0.790000  27.980000 ;
        RECT  0.590000  28.210000  0.790000  28.410000 ;
        RECT  0.615000 173.900000  0.815000 174.100000 ;
        RECT  0.615000 174.300000  0.815000 174.500000 ;
        RECT  0.615000 174.700000  0.815000 174.900000 ;
        RECT  0.615000 175.100000  0.815000 175.300000 ;
        RECT  0.615000 175.500000  0.815000 175.700000 ;
        RECT  0.615000 175.900000  0.815000 176.100000 ;
        RECT  0.615000 176.300000  0.815000 176.500000 ;
        RECT  0.615000 176.700000  0.815000 176.900000 ;
        RECT  0.615000 177.100000  0.815000 177.300000 ;
        RECT  0.615000 177.500000  0.815000 177.700000 ;
        RECT  0.615000 177.900000  0.815000 178.100000 ;
        RECT  0.615000 178.300000  0.815000 178.500000 ;
        RECT  0.615000 178.700000  0.815000 178.900000 ;
        RECT  0.615000 179.100000  0.815000 179.300000 ;
        RECT  0.615000 179.500000  0.815000 179.700000 ;
        RECT  0.615000 179.900000  0.815000 180.100000 ;
        RECT  0.615000 180.300000  0.815000 180.500000 ;
        RECT  0.615000 180.700000  0.815000 180.900000 ;
        RECT  0.615000 181.100000  0.815000 181.300000 ;
        RECT  0.615000 181.505000  0.815000 181.705000 ;
        RECT  0.615000 181.910000  0.815000 182.110000 ;
        RECT  0.615000 182.315000  0.815000 182.515000 ;
        RECT  0.615000 182.720000  0.815000 182.920000 ;
        RECT  0.615000 183.125000  0.815000 183.325000 ;
        RECT  0.615000 183.530000  0.815000 183.730000 ;
        RECT  0.615000 183.935000  0.815000 184.135000 ;
        RECT  0.615000 184.340000  0.815000 184.540000 ;
        RECT  0.615000 184.745000  0.815000 184.945000 ;
        RECT  0.615000 185.150000  0.815000 185.350000 ;
        RECT  0.615000 185.555000  0.815000 185.755000 ;
        RECT  0.615000 185.960000  0.815000 186.160000 ;
        RECT  0.615000 186.365000  0.815000 186.565000 ;
        RECT  0.615000 186.770000  0.815000 186.970000 ;
        RECT  0.615000 187.175000  0.815000 187.375000 ;
        RECT  0.615000 187.580000  0.815000 187.780000 ;
        RECT  0.615000 187.985000  0.815000 188.185000 ;
        RECT  0.615000 188.390000  0.815000 188.590000 ;
        RECT  0.615000 188.795000  0.815000 188.995000 ;
        RECT  0.615000 189.200000  0.815000 189.400000 ;
        RECT  0.615000 189.605000  0.815000 189.805000 ;
        RECT  0.615000 190.010000  0.815000 190.210000 ;
        RECT  0.615000 190.415000  0.815000 190.615000 ;
        RECT  0.615000 190.820000  0.815000 191.020000 ;
        RECT  0.615000 191.225000  0.815000 191.425000 ;
        RECT  0.615000 191.630000  0.815000 191.830000 ;
        RECT  0.615000 192.035000  0.815000 192.235000 ;
        RECT  0.615000 192.440000  0.815000 192.640000 ;
        RECT  0.615000 192.845000  0.815000 193.045000 ;
        RECT  0.615000 193.250000  0.815000 193.450000 ;
        RECT  0.615000 193.655000  0.815000 193.855000 ;
        RECT  0.615000 194.060000  0.815000 194.260000 ;
        RECT  0.615000 194.465000  0.815000 194.665000 ;
        RECT  0.615000 194.870000  0.815000 195.070000 ;
        RECT  0.615000 195.275000  0.815000 195.475000 ;
        RECT  0.615000 195.680000  0.815000 195.880000 ;
        RECT  0.615000 196.085000  0.815000 196.285000 ;
        RECT  0.615000 196.490000  0.815000 196.690000 ;
        RECT  0.615000 196.895000  0.815000 197.095000 ;
        RECT  0.615000 197.300000  0.815000 197.500000 ;
        RECT  0.615000 197.705000  0.815000 197.905000 ;
        RECT  1.000000  23.910000  1.200000  24.110000 ;
        RECT  1.000000  24.340000  1.200000  24.540000 ;
        RECT  1.000000  24.770000  1.200000  24.970000 ;
        RECT  1.000000  25.200000  1.200000  25.400000 ;
        RECT  1.000000  25.630000  1.200000  25.830000 ;
        RECT  1.000000  26.060000  1.200000  26.260000 ;
        RECT  1.000000  26.490000  1.200000  26.690000 ;
        RECT  1.000000  26.920000  1.200000  27.120000 ;
        RECT  1.000000  27.350000  1.200000  27.550000 ;
        RECT  1.000000  27.780000  1.200000  27.980000 ;
        RECT  1.000000  28.210000  1.200000  28.410000 ;
        RECT  1.015000 173.900000  1.215000 174.100000 ;
        RECT  1.015000 174.300000  1.215000 174.500000 ;
        RECT  1.015000 174.700000  1.215000 174.900000 ;
        RECT  1.015000 175.100000  1.215000 175.300000 ;
        RECT  1.015000 175.500000  1.215000 175.700000 ;
        RECT  1.015000 175.900000  1.215000 176.100000 ;
        RECT  1.015000 176.300000  1.215000 176.500000 ;
        RECT  1.015000 176.700000  1.215000 176.900000 ;
        RECT  1.015000 177.100000  1.215000 177.300000 ;
        RECT  1.015000 177.500000  1.215000 177.700000 ;
        RECT  1.015000 177.900000  1.215000 178.100000 ;
        RECT  1.015000 178.300000  1.215000 178.500000 ;
        RECT  1.015000 178.700000  1.215000 178.900000 ;
        RECT  1.015000 179.100000  1.215000 179.300000 ;
        RECT  1.015000 179.500000  1.215000 179.700000 ;
        RECT  1.015000 179.900000  1.215000 180.100000 ;
        RECT  1.015000 180.300000  1.215000 180.500000 ;
        RECT  1.015000 180.700000  1.215000 180.900000 ;
        RECT  1.015000 181.100000  1.215000 181.300000 ;
        RECT  1.015000 181.505000  1.215000 181.705000 ;
        RECT  1.015000 181.910000  1.215000 182.110000 ;
        RECT  1.015000 182.315000  1.215000 182.515000 ;
        RECT  1.015000 182.720000  1.215000 182.920000 ;
        RECT  1.015000 183.125000  1.215000 183.325000 ;
        RECT  1.015000 183.530000  1.215000 183.730000 ;
        RECT  1.015000 183.935000  1.215000 184.135000 ;
        RECT  1.015000 184.340000  1.215000 184.540000 ;
        RECT  1.015000 184.745000  1.215000 184.945000 ;
        RECT  1.015000 185.150000  1.215000 185.350000 ;
        RECT  1.015000 185.555000  1.215000 185.755000 ;
        RECT  1.015000 185.960000  1.215000 186.160000 ;
        RECT  1.015000 186.365000  1.215000 186.565000 ;
        RECT  1.015000 186.770000  1.215000 186.970000 ;
        RECT  1.015000 187.175000  1.215000 187.375000 ;
        RECT  1.015000 187.580000  1.215000 187.780000 ;
        RECT  1.015000 187.985000  1.215000 188.185000 ;
        RECT  1.015000 188.390000  1.215000 188.590000 ;
        RECT  1.015000 188.795000  1.215000 188.995000 ;
        RECT  1.015000 189.200000  1.215000 189.400000 ;
        RECT  1.015000 189.605000  1.215000 189.805000 ;
        RECT  1.015000 190.010000  1.215000 190.210000 ;
        RECT  1.015000 190.415000  1.215000 190.615000 ;
        RECT  1.015000 190.820000  1.215000 191.020000 ;
        RECT  1.015000 191.225000  1.215000 191.425000 ;
        RECT  1.015000 191.630000  1.215000 191.830000 ;
        RECT  1.015000 192.035000  1.215000 192.235000 ;
        RECT  1.015000 192.440000  1.215000 192.640000 ;
        RECT  1.015000 192.845000  1.215000 193.045000 ;
        RECT  1.015000 193.250000  1.215000 193.450000 ;
        RECT  1.015000 193.655000  1.215000 193.855000 ;
        RECT  1.015000 194.060000  1.215000 194.260000 ;
        RECT  1.015000 194.465000  1.215000 194.665000 ;
        RECT  1.015000 194.870000  1.215000 195.070000 ;
        RECT  1.015000 195.275000  1.215000 195.475000 ;
        RECT  1.015000 195.680000  1.215000 195.880000 ;
        RECT  1.015000 196.085000  1.215000 196.285000 ;
        RECT  1.015000 196.490000  1.215000 196.690000 ;
        RECT  1.015000 196.895000  1.215000 197.095000 ;
        RECT  1.015000 197.300000  1.215000 197.500000 ;
        RECT  1.015000 197.705000  1.215000 197.905000 ;
        RECT  1.410000  23.910000  1.610000  24.110000 ;
        RECT  1.410000  24.340000  1.610000  24.540000 ;
        RECT  1.410000  24.770000  1.610000  24.970000 ;
        RECT  1.410000  25.200000  1.610000  25.400000 ;
        RECT  1.410000  25.630000  1.610000  25.830000 ;
        RECT  1.410000  26.060000  1.610000  26.260000 ;
        RECT  1.410000  26.490000  1.610000  26.690000 ;
        RECT  1.410000  26.920000  1.610000  27.120000 ;
        RECT  1.410000  27.350000  1.610000  27.550000 ;
        RECT  1.410000  27.780000  1.610000  27.980000 ;
        RECT  1.410000  28.210000  1.610000  28.410000 ;
        RECT  1.415000 173.900000  1.615000 174.100000 ;
        RECT  1.415000 174.300000  1.615000 174.500000 ;
        RECT  1.415000 174.700000  1.615000 174.900000 ;
        RECT  1.415000 175.100000  1.615000 175.300000 ;
        RECT  1.415000 175.500000  1.615000 175.700000 ;
        RECT  1.415000 175.900000  1.615000 176.100000 ;
        RECT  1.415000 176.300000  1.615000 176.500000 ;
        RECT  1.415000 176.700000  1.615000 176.900000 ;
        RECT  1.415000 177.100000  1.615000 177.300000 ;
        RECT  1.415000 177.500000  1.615000 177.700000 ;
        RECT  1.415000 177.900000  1.615000 178.100000 ;
        RECT  1.415000 178.300000  1.615000 178.500000 ;
        RECT  1.415000 178.700000  1.615000 178.900000 ;
        RECT  1.415000 179.100000  1.615000 179.300000 ;
        RECT  1.415000 179.500000  1.615000 179.700000 ;
        RECT  1.415000 179.900000  1.615000 180.100000 ;
        RECT  1.415000 180.300000  1.615000 180.500000 ;
        RECT  1.415000 180.700000  1.615000 180.900000 ;
        RECT  1.415000 181.100000  1.615000 181.300000 ;
        RECT  1.415000 181.505000  1.615000 181.705000 ;
        RECT  1.415000 181.910000  1.615000 182.110000 ;
        RECT  1.415000 182.315000  1.615000 182.515000 ;
        RECT  1.415000 182.720000  1.615000 182.920000 ;
        RECT  1.415000 183.125000  1.615000 183.325000 ;
        RECT  1.415000 183.530000  1.615000 183.730000 ;
        RECT  1.415000 183.935000  1.615000 184.135000 ;
        RECT  1.415000 184.340000  1.615000 184.540000 ;
        RECT  1.415000 184.745000  1.615000 184.945000 ;
        RECT  1.415000 185.150000  1.615000 185.350000 ;
        RECT  1.415000 185.555000  1.615000 185.755000 ;
        RECT  1.415000 185.960000  1.615000 186.160000 ;
        RECT  1.415000 186.365000  1.615000 186.565000 ;
        RECT  1.415000 186.770000  1.615000 186.970000 ;
        RECT  1.415000 187.175000  1.615000 187.375000 ;
        RECT  1.415000 187.580000  1.615000 187.780000 ;
        RECT  1.415000 187.985000  1.615000 188.185000 ;
        RECT  1.415000 188.390000  1.615000 188.590000 ;
        RECT  1.415000 188.795000  1.615000 188.995000 ;
        RECT  1.415000 189.200000  1.615000 189.400000 ;
        RECT  1.415000 189.605000  1.615000 189.805000 ;
        RECT  1.415000 190.010000  1.615000 190.210000 ;
        RECT  1.415000 190.415000  1.615000 190.615000 ;
        RECT  1.415000 190.820000  1.615000 191.020000 ;
        RECT  1.415000 191.225000  1.615000 191.425000 ;
        RECT  1.415000 191.630000  1.615000 191.830000 ;
        RECT  1.415000 192.035000  1.615000 192.235000 ;
        RECT  1.415000 192.440000  1.615000 192.640000 ;
        RECT  1.415000 192.845000  1.615000 193.045000 ;
        RECT  1.415000 193.250000  1.615000 193.450000 ;
        RECT  1.415000 193.655000  1.615000 193.855000 ;
        RECT  1.415000 194.060000  1.615000 194.260000 ;
        RECT  1.415000 194.465000  1.615000 194.665000 ;
        RECT  1.415000 194.870000  1.615000 195.070000 ;
        RECT  1.415000 195.275000  1.615000 195.475000 ;
        RECT  1.415000 195.680000  1.615000 195.880000 ;
        RECT  1.415000 196.085000  1.615000 196.285000 ;
        RECT  1.415000 196.490000  1.615000 196.690000 ;
        RECT  1.415000 196.895000  1.615000 197.095000 ;
        RECT  1.415000 197.300000  1.615000 197.500000 ;
        RECT  1.415000 197.705000  1.615000 197.905000 ;
        RECT  1.815000 173.900000  2.015000 174.100000 ;
        RECT  1.815000 174.300000  2.015000 174.500000 ;
        RECT  1.815000 174.700000  2.015000 174.900000 ;
        RECT  1.815000 175.100000  2.015000 175.300000 ;
        RECT  1.815000 175.500000  2.015000 175.700000 ;
        RECT  1.815000 175.900000  2.015000 176.100000 ;
        RECT  1.815000 176.300000  2.015000 176.500000 ;
        RECT  1.815000 176.700000  2.015000 176.900000 ;
        RECT  1.815000 177.100000  2.015000 177.300000 ;
        RECT  1.815000 177.500000  2.015000 177.700000 ;
        RECT  1.815000 177.900000  2.015000 178.100000 ;
        RECT  1.815000 178.300000  2.015000 178.500000 ;
        RECT  1.815000 178.700000  2.015000 178.900000 ;
        RECT  1.815000 179.100000  2.015000 179.300000 ;
        RECT  1.815000 179.500000  2.015000 179.700000 ;
        RECT  1.815000 179.900000  2.015000 180.100000 ;
        RECT  1.815000 180.300000  2.015000 180.500000 ;
        RECT  1.815000 180.700000  2.015000 180.900000 ;
        RECT  1.815000 181.100000  2.015000 181.300000 ;
        RECT  1.815000 181.505000  2.015000 181.705000 ;
        RECT  1.815000 181.910000  2.015000 182.110000 ;
        RECT  1.815000 182.315000  2.015000 182.515000 ;
        RECT  1.815000 182.720000  2.015000 182.920000 ;
        RECT  1.815000 183.125000  2.015000 183.325000 ;
        RECT  1.815000 183.530000  2.015000 183.730000 ;
        RECT  1.815000 183.935000  2.015000 184.135000 ;
        RECT  1.815000 184.340000  2.015000 184.540000 ;
        RECT  1.815000 184.745000  2.015000 184.945000 ;
        RECT  1.815000 185.150000  2.015000 185.350000 ;
        RECT  1.815000 185.555000  2.015000 185.755000 ;
        RECT  1.815000 185.960000  2.015000 186.160000 ;
        RECT  1.815000 186.365000  2.015000 186.565000 ;
        RECT  1.815000 186.770000  2.015000 186.970000 ;
        RECT  1.815000 187.175000  2.015000 187.375000 ;
        RECT  1.815000 187.580000  2.015000 187.780000 ;
        RECT  1.815000 187.985000  2.015000 188.185000 ;
        RECT  1.815000 188.390000  2.015000 188.590000 ;
        RECT  1.815000 188.795000  2.015000 188.995000 ;
        RECT  1.815000 189.200000  2.015000 189.400000 ;
        RECT  1.815000 189.605000  2.015000 189.805000 ;
        RECT  1.815000 190.010000  2.015000 190.210000 ;
        RECT  1.815000 190.415000  2.015000 190.615000 ;
        RECT  1.815000 190.820000  2.015000 191.020000 ;
        RECT  1.815000 191.225000  2.015000 191.425000 ;
        RECT  1.815000 191.630000  2.015000 191.830000 ;
        RECT  1.815000 192.035000  2.015000 192.235000 ;
        RECT  1.815000 192.440000  2.015000 192.640000 ;
        RECT  1.815000 192.845000  2.015000 193.045000 ;
        RECT  1.815000 193.250000  2.015000 193.450000 ;
        RECT  1.815000 193.655000  2.015000 193.855000 ;
        RECT  1.815000 194.060000  2.015000 194.260000 ;
        RECT  1.815000 194.465000  2.015000 194.665000 ;
        RECT  1.815000 194.870000  2.015000 195.070000 ;
        RECT  1.815000 195.275000  2.015000 195.475000 ;
        RECT  1.815000 195.680000  2.015000 195.880000 ;
        RECT  1.815000 196.085000  2.015000 196.285000 ;
        RECT  1.815000 196.490000  2.015000 196.690000 ;
        RECT  1.815000 196.895000  2.015000 197.095000 ;
        RECT  1.815000 197.300000  2.015000 197.500000 ;
        RECT  1.815000 197.705000  2.015000 197.905000 ;
        RECT  1.820000  23.910000  2.020000  24.110000 ;
        RECT  1.820000  24.340000  2.020000  24.540000 ;
        RECT  1.820000  24.770000  2.020000  24.970000 ;
        RECT  1.820000  25.200000  2.020000  25.400000 ;
        RECT  1.820000  25.630000  2.020000  25.830000 ;
        RECT  1.820000  26.060000  2.020000  26.260000 ;
        RECT  1.820000  26.490000  2.020000  26.690000 ;
        RECT  1.820000  26.920000  2.020000  27.120000 ;
        RECT  1.820000  27.350000  2.020000  27.550000 ;
        RECT  1.820000  27.780000  2.020000  27.980000 ;
        RECT  1.820000  28.210000  2.020000  28.410000 ;
        RECT  2.215000 173.900000  2.415000 174.100000 ;
        RECT  2.215000 174.300000  2.415000 174.500000 ;
        RECT  2.215000 174.700000  2.415000 174.900000 ;
        RECT  2.215000 175.100000  2.415000 175.300000 ;
        RECT  2.215000 175.500000  2.415000 175.700000 ;
        RECT  2.215000 175.900000  2.415000 176.100000 ;
        RECT  2.215000 176.300000  2.415000 176.500000 ;
        RECT  2.215000 176.700000  2.415000 176.900000 ;
        RECT  2.215000 177.100000  2.415000 177.300000 ;
        RECT  2.215000 177.500000  2.415000 177.700000 ;
        RECT  2.215000 177.900000  2.415000 178.100000 ;
        RECT  2.215000 178.300000  2.415000 178.500000 ;
        RECT  2.215000 178.700000  2.415000 178.900000 ;
        RECT  2.215000 179.100000  2.415000 179.300000 ;
        RECT  2.215000 179.500000  2.415000 179.700000 ;
        RECT  2.215000 179.900000  2.415000 180.100000 ;
        RECT  2.215000 180.300000  2.415000 180.500000 ;
        RECT  2.215000 180.700000  2.415000 180.900000 ;
        RECT  2.215000 181.100000  2.415000 181.300000 ;
        RECT  2.215000 181.505000  2.415000 181.705000 ;
        RECT  2.215000 181.910000  2.415000 182.110000 ;
        RECT  2.215000 182.315000  2.415000 182.515000 ;
        RECT  2.215000 182.720000  2.415000 182.920000 ;
        RECT  2.215000 183.125000  2.415000 183.325000 ;
        RECT  2.215000 183.530000  2.415000 183.730000 ;
        RECT  2.215000 183.935000  2.415000 184.135000 ;
        RECT  2.215000 184.340000  2.415000 184.540000 ;
        RECT  2.215000 184.745000  2.415000 184.945000 ;
        RECT  2.215000 185.150000  2.415000 185.350000 ;
        RECT  2.215000 185.555000  2.415000 185.755000 ;
        RECT  2.215000 185.960000  2.415000 186.160000 ;
        RECT  2.215000 186.365000  2.415000 186.565000 ;
        RECT  2.215000 186.770000  2.415000 186.970000 ;
        RECT  2.215000 187.175000  2.415000 187.375000 ;
        RECT  2.215000 187.580000  2.415000 187.780000 ;
        RECT  2.215000 187.985000  2.415000 188.185000 ;
        RECT  2.215000 188.390000  2.415000 188.590000 ;
        RECT  2.215000 188.795000  2.415000 188.995000 ;
        RECT  2.215000 189.200000  2.415000 189.400000 ;
        RECT  2.215000 189.605000  2.415000 189.805000 ;
        RECT  2.215000 190.010000  2.415000 190.210000 ;
        RECT  2.215000 190.415000  2.415000 190.615000 ;
        RECT  2.215000 190.820000  2.415000 191.020000 ;
        RECT  2.215000 191.225000  2.415000 191.425000 ;
        RECT  2.215000 191.630000  2.415000 191.830000 ;
        RECT  2.215000 192.035000  2.415000 192.235000 ;
        RECT  2.215000 192.440000  2.415000 192.640000 ;
        RECT  2.215000 192.845000  2.415000 193.045000 ;
        RECT  2.215000 193.250000  2.415000 193.450000 ;
        RECT  2.215000 193.655000  2.415000 193.855000 ;
        RECT  2.215000 194.060000  2.415000 194.260000 ;
        RECT  2.215000 194.465000  2.415000 194.665000 ;
        RECT  2.215000 194.870000  2.415000 195.070000 ;
        RECT  2.215000 195.275000  2.415000 195.475000 ;
        RECT  2.215000 195.680000  2.415000 195.880000 ;
        RECT  2.215000 196.085000  2.415000 196.285000 ;
        RECT  2.215000 196.490000  2.415000 196.690000 ;
        RECT  2.215000 196.895000  2.415000 197.095000 ;
        RECT  2.215000 197.300000  2.415000 197.500000 ;
        RECT  2.215000 197.705000  2.415000 197.905000 ;
        RECT  2.230000  23.910000  2.430000  24.110000 ;
        RECT  2.230000  24.340000  2.430000  24.540000 ;
        RECT  2.230000  24.770000  2.430000  24.970000 ;
        RECT  2.230000  25.200000  2.430000  25.400000 ;
        RECT  2.230000  25.630000  2.430000  25.830000 ;
        RECT  2.230000  26.060000  2.430000  26.260000 ;
        RECT  2.230000  26.490000  2.430000  26.690000 ;
        RECT  2.230000  26.920000  2.430000  27.120000 ;
        RECT  2.230000  27.350000  2.430000  27.550000 ;
        RECT  2.230000  27.780000  2.430000  27.980000 ;
        RECT  2.230000  28.210000  2.430000  28.410000 ;
        RECT  2.615000 173.900000  2.815000 174.100000 ;
        RECT  2.615000 174.300000  2.815000 174.500000 ;
        RECT  2.615000 174.700000  2.815000 174.900000 ;
        RECT  2.615000 175.100000  2.815000 175.300000 ;
        RECT  2.615000 175.500000  2.815000 175.700000 ;
        RECT  2.615000 175.900000  2.815000 176.100000 ;
        RECT  2.615000 176.300000  2.815000 176.500000 ;
        RECT  2.615000 176.700000  2.815000 176.900000 ;
        RECT  2.615000 177.100000  2.815000 177.300000 ;
        RECT  2.615000 177.500000  2.815000 177.700000 ;
        RECT  2.615000 177.900000  2.815000 178.100000 ;
        RECT  2.615000 178.300000  2.815000 178.500000 ;
        RECT  2.615000 178.700000  2.815000 178.900000 ;
        RECT  2.615000 179.100000  2.815000 179.300000 ;
        RECT  2.615000 179.500000  2.815000 179.700000 ;
        RECT  2.615000 179.900000  2.815000 180.100000 ;
        RECT  2.615000 180.300000  2.815000 180.500000 ;
        RECT  2.615000 180.700000  2.815000 180.900000 ;
        RECT  2.615000 181.100000  2.815000 181.300000 ;
        RECT  2.615000 181.505000  2.815000 181.705000 ;
        RECT  2.615000 181.910000  2.815000 182.110000 ;
        RECT  2.615000 182.315000  2.815000 182.515000 ;
        RECT  2.615000 182.720000  2.815000 182.920000 ;
        RECT  2.615000 183.125000  2.815000 183.325000 ;
        RECT  2.615000 183.530000  2.815000 183.730000 ;
        RECT  2.615000 183.935000  2.815000 184.135000 ;
        RECT  2.615000 184.340000  2.815000 184.540000 ;
        RECT  2.615000 184.745000  2.815000 184.945000 ;
        RECT  2.615000 185.150000  2.815000 185.350000 ;
        RECT  2.615000 185.555000  2.815000 185.755000 ;
        RECT  2.615000 185.960000  2.815000 186.160000 ;
        RECT  2.615000 186.365000  2.815000 186.565000 ;
        RECT  2.615000 186.770000  2.815000 186.970000 ;
        RECT  2.615000 187.175000  2.815000 187.375000 ;
        RECT  2.615000 187.580000  2.815000 187.780000 ;
        RECT  2.615000 187.985000  2.815000 188.185000 ;
        RECT  2.615000 188.390000  2.815000 188.590000 ;
        RECT  2.615000 188.795000  2.815000 188.995000 ;
        RECT  2.615000 189.200000  2.815000 189.400000 ;
        RECT  2.615000 189.605000  2.815000 189.805000 ;
        RECT  2.615000 190.010000  2.815000 190.210000 ;
        RECT  2.615000 190.415000  2.815000 190.615000 ;
        RECT  2.615000 190.820000  2.815000 191.020000 ;
        RECT  2.615000 191.225000  2.815000 191.425000 ;
        RECT  2.615000 191.630000  2.815000 191.830000 ;
        RECT  2.615000 192.035000  2.815000 192.235000 ;
        RECT  2.615000 192.440000  2.815000 192.640000 ;
        RECT  2.615000 192.845000  2.815000 193.045000 ;
        RECT  2.615000 193.250000  2.815000 193.450000 ;
        RECT  2.615000 193.655000  2.815000 193.855000 ;
        RECT  2.615000 194.060000  2.815000 194.260000 ;
        RECT  2.615000 194.465000  2.815000 194.665000 ;
        RECT  2.615000 194.870000  2.815000 195.070000 ;
        RECT  2.615000 195.275000  2.815000 195.475000 ;
        RECT  2.615000 195.680000  2.815000 195.880000 ;
        RECT  2.615000 196.085000  2.815000 196.285000 ;
        RECT  2.615000 196.490000  2.815000 196.690000 ;
        RECT  2.615000 196.895000  2.815000 197.095000 ;
        RECT  2.615000 197.300000  2.815000 197.500000 ;
        RECT  2.615000 197.705000  2.815000 197.905000 ;
        RECT  2.640000  23.910000  2.840000  24.110000 ;
        RECT  2.640000  24.340000  2.840000  24.540000 ;
        RECT  2.640000  24.770000  2.840000  24.970000 ;
        RECT  2.640000  25.200000  2.840000  25.400000 ;
        RECT  2.640000  25.630000  2.840000  25.830000 ;
        RECT  2.640000  26.060000  2.840000  26.260000 ;
        RECT  2.640000  26.490000  2.840000  26.690000 ;
        RECT  2.640000  26.920000  2.840000  27.120000 ;
        RECT  2.640000  27.350000  2.840000  27.550000 ;
        RECT  2.640000  27.780000  2.840000  27.980000 ;
        RECT  2.640000  28.210000  2.840000  28.410000 ;
        RECT  3.015000 173.900000  3.215000 174.100000 ;
        RECT  3.015000 174.300000  3.215000 174.500000 ;
        RECT  3.015000 174.700000  3.215000 174.900000 ;
        RECT  3.015000 175.100000  3.215000 175.300000 ;
        RECT  3.015000 175.500000  3.215000 175.700000 ;
        RECT  3.015000 175.900000  3.215000 176.100000 ;
        RECT  3.015000 176.300000  3.215000 176.500000 ;
        RECT  3.015000 176.700000  3.215000 176.900000 ;
        RECT  3.015000 177.100000  3.215000 177.300000 ;
        RECT  3.015000 177.500000  3.215000 177.700000 ;
        RECT  3.015000 177.900000  3.215000 178.100000 ;
        RECT  3.015000 178.300000  3.215000 178.500000 ;
        RECT  3.015000 178.700000  3.215000 178.900000 ;
        RECT  3.015000 179.100000  3.215000 179.300000 ;
        RECT  3.015000 179.500000  3.215000 179.700000 ;
        RECT  3.015000 179.900000  3.215000 180.100000 ;
        RECT  3.015000 180.300000  3.215000 180.500000 ;
        RECT  3.015000 180.700000  3.215000 180.900000 ;
        RECT  3.015000 181.100000  3.215000 181.300000 ;
        RECT  3.015000 181.505000  3.215000 181.705000 ;
        RECT  3.015000 181.910000  3.215000 182.110000 ;
        RECT  3.015000 182.315000  3.215000 182.515000 ;
        RECT  3.015000 182.720000  3.215000 182.920000 ;
        RECT  3.015000 183.125000  3.215000 183.325000 ;
        RECT  3.015000 183.530000  3.215000 183.730000 ;
        RECT  3.015000 183.935000  3.215000 184.135000 ;
        RECT  3.015000 184.340000  3.215000 184.540000 ;
        RECT  3.015000 184.745000  3.215000 184.945000 ;
        RECT  3.015000 185.150000  3.215000 185.350000 ;
        RECT  3.015000 185.555000  3.215000 185.755000 ;
        RECT  3.015000 185.960000  3.215000 186.160000 ;
        RECT  3.015000 186.365000  3.215000 186.565000 ;
        RECT  3.015000 186.770000  3.215000 186.970000 ;
        RECT  3.015000 187.175000  3.215000 187.375000 ;
        RECT  3.015000 187.580000  3.215000 187.780000 ;
        RECT  3.015000 187.985000  3.215000 188.185000 ;
        RECT  3.015000 188.390000  3.215000 188.590000 ;
        RECT  3.015000 188.795000  3.215000 188.995000 ;
        RECT  3.015000 189.200000  3.215000 189.400000 ;
        RECT  3.015000 189.605000  3.215000 189.805000 ;
        RECT  3.015000 190.010000  3.215000 190.210000 ;
        RECT  3.015000 190.415000  3.215000 190.615000 ;
        RECT  3.015000 190.820000  3.215000 191.020000 ;
        RECT  3.015000 191.225000  3.215000 191.425000 ;
        RECT  3.015000 191.630000  3.215000 191.830000 ;
        RECT  3.015000 192.035000  3.215000 192.235000 ;
        RECT  3.015000 192.440000  3.215000 192.640000 ;
        RECT  3.015000 192.845000  3.215000 193.045000 ;
        RECT  3.015000 193.250000  3.215000 193.450000 ;
        RECT  3.015000 193.655000  3.215000 193.855000 ;
        RECT  3.015000 194.060000  3.215000 194.260000 ;
        RECT  3.015000 194.465000  3.215000 194.665000 ;
        RECT  3.015000 194.870000  3.215000 195.070000 ;
        RECT  3.015000 195.275000  3.215000 195.475000 ;
        RECT  3.015000 195.680000  3.215000 195.880000 ;
        RECT  3.015000 196.085000  3.215000 196.285000 ;
        RECT  3.015000 196.490000  3.215000 196.690000 ;
        RECT  3.015000 196.895000  3.215000 197.095000 ;
        RECT  3.015000 197.300000  3.215000 197.500000 ;
        RECT  3.015000 197.705000  3.215000 197.905000 ;
        RECT  3.050000  23.910000  3.250000  24.110000 ;
        RECT  3.050000  24.340000  3.250000  24.540000 ;
        RECT  3.050000  24.770000  3.250000  24.970000 ;
        RECT  3.050000  25.200000  3.250000  25.400000 ;
        RECT  3.050000  25.630000  3.250000  25.830000 ;
        RECT  3.050000  26.060000  3.250000  26.260000 ;
        RECT  3.050000  26.490000  3.250000  26.690000 ;
        RECT  3.050000  26.920000  3.250000  27.120000 ;
        RECT  3.050000  27.350000  3.250000  27.550000 ;
        RECT  3.050000  27.780000  3.250000  27.980000 ;
        RECT  3.050000  28.210000  3.250000  28.410000 ;
        RECT  3.415000 173.900000  3.615000 174.100000 ;
        RECT  3.415000 174.300000  3.615000 174.500000 ;
        RECT  3.415000 174.700000  3.615000 174.900000 ;
        RECT  3.415000 175.100000  3.615000 175.300000 ;
        RECT  3.415000 175.500000  3.615000 175.700000 ;
        RECT  3.415000 175.900000  3.615000 176.100000 ;
        RECT  3.415000 176.300000  3.615000 176.500000 ;
        RECT  3.415000 176.700000  3.615000 176.900000 ;
        RECT  3.415000 177.100000  3.615000 177.300000 ;
        RECT  3.415000 177.500000  3.615000 177.700000 ;
        RECT  3.415000 177.900000  3.615000 178.100000 ;
        RECT  3.415000 178.300000  3.615000 178.500000 ;
        RECT  3.415000 178.700000  3.615000 178.900000 ;
        RECT  3.415000 179.100000  3.615000 179.300000 ;
        RECT  3.415000 179.500000  3.615000 179.700000 ;
        RECT  3.415000 179.900000  3.615000 180.100000 ;
        RECT  3.415000 180.300000  3.615000 180.500000 ;
        RECT  3.415000 180.700000  3.615000 180.900000 ;
        RECT  3.415000 181.100000  3.615000 181.300000 ;
        RECT  3.415000 181.505000  3.615000 181.705000 ;
        RECT  3.415000 181.910000  3.615000 182.110000 ;
        RECT  3.415000 182.315000  3.615000 182.515000 ;
        RECT  3.415000 182.720000  3.615000 182.920000 ;
        RECT  3.415000 183.125000  3.615000 183.325000 ;
        RECT  3.415000 183.530000  3.615000 183.730000 ;
        RECT  3.415000 183.935000  3.615000 184.135000 ;
        RECT  3.415000 184.340000  3.615000 184.540000 ;
        RECT  3.415000 184.745000  3.615000 184.945000 ;
        RECT  3.415000 185.150000  3.615000 185.350000 ;
        RECT  3.415000 185.555000  3.615000 185.755000 ;
        RECT  3.415000 185.960000  3.615000 186.160000 ;
        RECT  3.415000 186.365000  3.615000 186.565000 ;
        RECT  3.415000 186.770000  3.615000 186.970000 ;
        RECT  3.415000 187.175000  3.615000 187.375000 ;
        RECT  3.415000 187.580000  3.615000 187.780000 ;
        RECT  3.415000 187.985000  3.615000 188.185000 ;
        RECT  3.415000 188.390000  3.615000 188.590000 ;
        RECT  3.415000 188.795000  3.615000 188.995000 ;
        RECT  3.415000 189.200000  3.615000 189.400000 ;
        RECT  3.415000 189.605000  3.615000 189.805000 ;
        RECT  3.415000 190.010000  3.615000 190.210000 ;
        RECT  3.415000 190.415000  3.615000 190.615000 ;
        RECT  3.415000 190.820000  3.615000 191.020000 ;
        RECT  3.415000 191.225000  3.615000 191.425000 ;
        RECT  3.415000 191.630000  3.615000 191.830000 ;
        RECT  3.415000 192.035000  3.615000 192.235000 ;
        RECT  3.415000 192.440000  3.615000 192.640000 ;
        RECT  3.415000 192.845000  3.615000 193.045000 ;
        RECT  3.415000 193.250000  3.615000 193.450000 ;
        RECT  3.415000 193.655000  3.615000 193.855000 ;
        RECT  3.415000 194.060000  3.615000 194.260000 ;
        RECT  3.415000 194.465000  3.615000 194.665000 ;
        RECT  3.415000 194.870000  3.615000 195.070000 ;
        RECT  3.415000 195.275000  3.615000 195.475000 ;
        RECT  3.415000 195.680000  3.615000 195.880000 ;
        RECT  3.415000 196.085000  3.615000 196.285000 ;
        RECT  3.415000 196.490000  3.615000 196.690000 ;
        RECT  3.415000 196.895000  3.615000 197.095000 ;
        RECT  3.415000 197.300000  3.615000 197.500000 ;
        RECT  3.415000 197.705000  3.615000 197.905000 ;
        RECT  3.455000  23.910000  3.655000  24.110000 ;
        RECT  3.455000  24.340000  3.655000  24.540000 ;
        RECT  3.455000  24.770000  3.655000  24.970000 ;
        RECT  3.455000  25.200000  3.655000  25.400000 ;
        RECT  3.455000  25.630000  3.655000  25.830000 ;
        RECT  3.455000  26.060000  3.655000  26.260000 ;
        RECT  3.455000  26.490000  3.655000  26.690000 ;
        RECT  3.455000  26.920000  3.655000  27.120000 ;
        RECT  3.455000  27.350000  3.655000  27.550000 ;
        RECT  3.455000  27.780000  3.655000  27.980000 ;
        RECT  3.455000  28.210000  3.655000  28.410000 ;
        RECT  3.815000 173.900000  4.015000 174.100000 ;
        RECT  3.815000 174.300000  4.015000 174.500000 ;
        RECT  3.815000 174.700000  4.015000 174.900000 ;
        RECT  3.815000 175.100000  4.015000 175.300000 ;
        RECT  3.815000 175.500000  4.015000 175.700000 ;
        RECT  3.815000 175.900000  4.015000 176.100000 ;
        RECT  3.815000 176.300000  4.015000 176.500000 ;
        RECT  3.815000 176.700000  4.015000 176.900000 ;
        RECT  3.815000 177.100000  4.015000 177.300000 ;
        RECT  3.815000 177.500000  4.015000 177.700000 ;
        RECT  3.815000 177.900000  4.015000 178.100000 ;
        RECT  3.815000 178.300000  4.015000 178.500000 ;
        RECT  3.815000 178.700000  4.015000 178.900000 ;
        RECT  3.815000 179.100000  4.015000 179.300000 ;
        RECT  3.815000 179.500000  4.015000 179.700000 ;
        RECT  3.815000 179.900000  4.015000 180.100000 ;
        RECT  3.815000 180.300000  4.015000 180.500000 ;
        RECT  3.815000 180.700000  4.015000 180.900000 ;
        RECT  3.815000 181.100000  4.015000 181.300000 ;
        RECT  3.815000 181.505000  4.015000 181.705000 ;
        RECT  3.815000 181.910000  4.015000 182.110000 ;
        RECT  3.815000 182.315000  4.015000 182.515000 ;
        RECT  3.815000 182.720000  4.015000 182.920000 ;
        RECT  3.815000 183.125000  4.015000 183.325000 ;
        RECT  3.815000 183.530000  4.015000 183.730000 ;
        RECT  3.815000 183.935000  4.015000 184.135000 ;
        RECT  3.815000 184.340000  4.015000 184.540000 ;
        RECT  3.815000 184.745000  4.015000 184.945000 ;
        RECT  3.815000 185.150000  4.015000 185.350000 ;
        RECT  3.815000 185.555000  4.015000 185.755000 ;
        RECT  3.815000 185.960000  4.015000 186.160000 ;
        RECT  3.815000 186.365000  4.015000 186.565000 ;
        RECT  3.815000 186.770000  4.015000 186.970000 ;
        RECT  3.815000 187.175000  4.015000 187.375000 ;
        RECT  3.815000 187.580000  4.015000 187.780000 ;
        RECT  3.815000 187.985000  4.015000 188.185000 ;
        RECT  3.815000 188.390000  4.015000 188.590000 ;
        RECT  3.815000 188.795000  4.015000 188.995000 ;
        RECT  3.815000 189.200000  4.015000 189.400000 ;
        RECT  3.815000 189.605000  4.015000 189.805000 ;
        RECT  3.815000 190.010000  4.015000 190.210000 ;
        RECT  3.815000 190.415000  4.015000 190.615000 ;
        RECT  3.815000 190.820000  4.015000 191.020000 ;
        RECT  3.815000 191.225000  4.015000 191.425000 ;
        RECT  3.815000 191.630000  4.015000 191.830000 ;
        RECT  3.815000 192.035000  4.015000 192.235000 ;
        RECT  3.815000 192.440000  4.015000 192.640000 ;
        RECT  3.815000 192.845000  4.015000 193.045000 ;
        RECT  3.815000 193.250000  4.015000 193.450000 ;
        RECT  3.815000 193.655000  4.015000 193.855000 ;
        RECT  3.815000 194.060000  4.015000 194.260000 ;
        RECT  3.815000 194.465000  4.015000 194.665000 ;
        RECT  3.815000 194.870000  4.015000 195.070000 ;
        RECT  3.815000 195.275000  4.015000 195.475000 ;
        RECT  3.815000 195.680000  4.015000 195.880000 ;
        RECT  3.815000 196.085000  4.015000 196.285000 ;
        RECT  3.815000 196.490000  4.015000 196.690000 ;
        RECT  3.815000 196.895000  4.015000 197.095000 ;
        RECT  3.815000 197.300000  4.015000 197.500000 ;
        RECT  3.815000 197.705000  4.015000 197.905000 ;
        RECT  3.860000  23.910000  4.060000  24.110000 ;
        RECT  3.860000  24.340000  4.060000  24.540000 ;
        RECT  3.860000  24.770000  4.060000  24.970000 ;
        RECT  3.860000  25.200000  4.060000  25.400000 ;
        RECT  3.860000  25.630000  4.060000  25.830000 ;
        RECT  3.860000  26.060000  4.060000  26.260000 ;
        RECT  3.860000  26.490000  4.060000  26.690000 ;
        RECT  3.860000  26.920000  4.060000  27.120000 ;
        RECT  3.860000  27.350000  4.060000  27.550000 ;
        RECT  3.860000  27.780000  4.060000  27.980000 ;
        RECT  3.860000  28.210000  4.060000  28.410000 ;
        RECT  4.215000 173.900000  4.415000 174.100000 ;
        RECT  4.215000 174.300000  4.415000 174.500000 ;
        RECT  4.215000 174.700000  4.415000 174.900000 ;
        RECT  4.215000 175.100000  4.415000 175.300000 ;
        RECT  4.215000 175.500000  4.415000 175.700000 ;
        RECT  4.215000 175.900000  4.415000 176.100000 ;
        RECT  4.215000 176.300000  4.415000 176.500000 ;
        RECT  4.215000 176.700000  4.415000 176.900000 ;
        RECT  4.215000 177.100000  4.415000 177.300000 ;
        RECT  4.215000 177.500000  4.415000 177.700000 ;
        RECT  4.215000 177.900000  4.415000 178.100000 ;
        RECT  4.215000 178.300000  4.415000 178.500000 ;
        RECT  4.215000 178.700000  4.415000 178.900000 ;
        RECT  4.215000 179.100000  4.415000 179.300000 ;
        RECT  4.215000 179.500000  4.415000 179.700000 ;
        RECT  4.215000 179.900000  4.415000 180.100000 ;
        RECT  4.215000 180.300000  4.415000 180.500000 ;
        RECT  4.215000 180.700000  4.415000 180.900000 ;
        RECT  4.215000 181.100000  4.415000 181.300000 ;
        RECT  4.215000 181.505000  4.415000 181.705000 ;
        RECT  4.215000 181.910000  4.415000 182.110000 ;
        RECT  4.215000 182.315000  4.415000 182.515000 ;
        RECT  4.215000 182.720000  4.415000 182.920000 ;
        RECT  4.215000 183.125000  4.415000 183.325000 ;
        RECT  4.215000 183.530000  4.415000 183.730000 ;
        RECT  4.215000 183.935000  4.415000 184.135000 ;
        RECT  4.215000 184.340000  4.415000 184.540000 ;
        RECT  4.215000 184.745000  4.415000 184.945000 ;
        RECT  4.215000 185.150000  4.415000 185.350000 ;
        RECT  4.215000 185.555000  4.415000 185.755000 ;
        RECT  4.215000 185.960000  4.415000 186.160000 ;
        RECT  4.215000 186.365000  4.415000 186.565000 ;
        RECT  4.215000 186.770000  4.415000 186.970000 ;
        RECT  4.215000 187.175000  4.415000 187.375000 ;
        RECT  4.215000 187.580000  4.415000 187.780000 ;
        RECT  4.215000 187.985000  4.415000 188.185000 ;
        RECT  4.215000 188.390000  4.415000 188.590000 ;
        RECT  4.215000 188.795000  4.415000 188.995000 ;
        RECT  4.215000 189.200000  4.415000 189.400000 ;
        RECT  4.215000 189.605000  4.415000 189.805000 ;
        RECT  4.215000 190.010000  4.415000 190.210000 ;
        RECT  4.215000 190.415000  4.415000 190.615000 ;
        RECT  4.215000 190.820000  4.415000 191.020000 ;
        RECT  4.215000 191.225000  4.415000 191.425000 ;
        RECT  4.215000 191.630000  4.415000 191.830000 ;
        RECT  4.215000 192.035000  4.415000 192.235000 ;
        RECT  4.215000 192.440000  4.415000 192.640000 ;
        RECT  4.215000 192.845000  4.415000 193.045000 ;
        RECT  4.215000 193.250000  4.415000 193.450000 ;
        RECT  4.215000 193.655000  4.415000 193.855000 ;
        RECT  4.215000 194.060000  4.415000 194.260000 ;
        RECT  4.215000 194.465000  4.415000 194.665000 ;
        RECT  4.215000 194.870000  4.415000 195.070000 ;
        RECT  4.215000 195.275000  4.415000 195.475000 ;
        RECT  4.215000 195.680000  4.415000 195.880000 ;
        RECT  4.215000 196.085000  4.415000 196.285000 ;
        RECT  4.215000 196.490000  4.415000 196.690000 ;
        RECT  4.215000 196.895000  4.415000 197.095000 ;
        RECT  4.215000 197.300000  4.415000 197.500000 ;
        RECT  4.215000 197.705000  4.415000 197.905000 ;
        RECT  4.265000  23.910000  4.465000  24.110000 ;
        RECT  4.265000  24.340000  4.465000  24.540000 ;
        RECT  4.265000  24.770000  4.465000  24.970000 ;
        RECT  4.265000  25.200000  4.465000  25.400000 ;
        RECT  4.265000  25.630000  4.465000  25.830000 ;
        RECT  4.265000  26.060000  4.465000  26.260000 ;
        RECT  4.265000  26.490000  4.465000  26.690000 ;
        RECT  4.265000  26.920000  4.465000  27.120000 ;
        RECT  4.265000  27.350000  4.465000  27.550000 ;
        RECT  4.265000  27.780000  4.465000  27.980000 ;
        RECT  4.265000  28.210000  4.465000  28.410000 ;
        RECT  4.615000 173.900000  4.815000 174.100000 ;
        RECT  4.615000 174.300000  4.815000 174.500000 ;
        RECT  4.615000 174.700000  4.815000 174.900000 ;
        RECT  4.615000 175.100000  4.815000 175.300000 ;
        RECT  4.615000 175.500000  4.815000 175.700000 ;
        RECT  4.615000 175.900000  4.815000 176.100000 ;
        RECT  4.615000 176.300000  4.815000 176.500000 ;
        RECT  4.615000 176.700000  4.815000 176.900000 ;
        RECT  4.615000 177.100000  4.815000 177.300000 ;
        RECT  4.615000 177.500000  4.815000 177.700000 ;
        RECT  4.615000 177.900000  4.815000 178.100000 ;
        RECT  4.615000 178.300000  4.815000 178.500000 ;
        RECT  4.615000 178.700000  4.815000 178.900000 ;
        RECT  4.615000 179.100000  4.815000 179.300000 ;
        RECT  4.615000 179.500000  4.815000 179.700000 ;
        RECT  4.615000 179.900000  4.815000 180.100000 ;
        RECT  4.615000 180.300000  4.815000 180.500000 ;
        RECT  4.615000 180.700000  4.815000 180.900000 ;
        RECT  4.615000 181.100000  4.815000 181.300000 ;
        RECT  4.615000 181.505000  4.815000 181.705000 ;
        RECT  4.615000 181.910000  4.815000 182.110000 ;
        RECT  4.615000 182.315000  4.815000 182.515000 ;
        RECT  4.615000 182.720000  4.815000 182.920000 ;
        RECT  4.615000 183.125000  4.815000 183.325000 ;
        RECT  4.615000 183.530000  4.815000 183.730000 ;
        RECT  4.615000 183.935000  4.815000 184.135000 ;
        RECT  4.615000 184.340000  4.815000 184.540000 ;
        RECT  4.615000 184.745000  4.815000 184.945000 ;
        RECT  4.615000 185.150000  4.815000 185.350000 ;
        RECT  4.615000 185.555000  4.815000 185.755000 ;
        RECT  4.615000 185.960000  4.815000 186.160000 ;
        RECT  4.615000 186.365000  4.815000 186.565000 ;
        RECT  4.615000 186.770000  4.815000 186.970000 ;
        RECT  4.615000 187.175000  4.815000 187.375000 ;
        RECT  4.615000 187.580000  4.815000 187.780000 ;
        RECT  4.615000 187.985000  4.815000 188.185000 ;
        RECT  4.615000 188.390000  4.815000 188.590000 ;
        RECT  4.615000 188.795000  4.815000 188.995000 ;
        RECT  4.615000 189.200000  4.815000 189.400000 ;
        RECT  4.615000 189.605000  4.815000 189.805000 ;
        RECT  4.615000 190.010000  4.815000 190.210000 ;
        RECT  4.615000 190.415000  4.815000 190.615000 ;
        RECT  4.615000 190.820000  4.815000 191.020000 ;
        RECT  4.615000 191.225000  4.815000 191.425000 ;
        RECT  4.615000 191.630000  4.815000 191.830000 ;
        RECT  4.615000 192.035000  4.815000 192.235000 ;
        RECT  4.615000 192.440000  4.815000 192.640000 ;
        RECT  4.615000 192.845000  4.815000 193.045000 ;
        RECT  4.615000 193.250000  4.815000 193.450000 ;
        RECT  4.615000 193.655000  4.815000 193.855000 ;
        RECT  4.615000 194.060000  4.815000 194.260000 ;
        RECT  4.615000 194.465000  4.815000 194.665000 ;
        RECT  4.615000 194.870000  4.815000 195.070000 ;
        RECT  4.615000 195.275000  4.815000 195.475000 ;
        RECT  4.615000 195.680000  4.815000 195.880000 ;
        RECT  4.615000 196.085000  4.815000 196.285000 ;
        RECT  4.615000 196.490000  4.815000 196.690000 ;
        RECT  4.615000 196.895000  4.815000 197.095000 ;
        RECT  4.615000 197.300000  4.815000 197.500000 ;
        RECT  4.615000 197.705000  4.815000 197.905000 ;
        RECT  4.670000  23.910000  4.870000  24.110000 ;
        RECT  4.670000  24.340000  4.870000  24.540000 ;
        RECT  4.670000  24.770000  4.870000  24.970000 ;
        RECT  4.670000  25.200000  4.870000  25.400000 ;
        RECT  4.670000  25.630000  4.870000  25.830000 ;
        RECT  4.670000  26.060000  4.870000  26.260000 ;
        RECT  4.670000  26.490000  4.870000  26.690000 ;
        RECT  4.670000  26.920000  4.870000  27.120000 ;
        RECT  4.670000  27.350000  4.870000  27.550000 ;
        RECT  4.670000  27.780000  4.870000  27.980000 ;
        RECT  4.670000  28.210000  4.870000  28.410000 ;
        RECT  5.015000 173.900000  5.215000 174.100000 ;
        RECT  5.015000 174.300000  5.215000 174.500000 ;
        RECT  5.015000 174.700000  5.215000 174.900000 ;
        RECT  5.015000 175.100000  5.215000 175.300000 ;
        RECT  5.015000 175.500000  5.215000 175.700000 ;
        RECT  5.015000 175.900000  5.215000 176.100000 ;
        RECT  5.015000 176.300000  5.215000 176.500000 ;
        RECT  5.015000 176.700000  5.215000 176.900000 ;
        RECT  5.015000 177.100000  5.215000 177.300000 ;
        RECT  5.015000 177.500000  5.215000 177.700000 ;
        RECT  5.015000 177.900000  5.215000 178.100000 ;
        RECT  5.015000 178.300000  5.215000 178.500000 ;
        RECT  5.015000 178.700000  5.215000 178.900000 ;
        RECT  5.015000 179.100000  5.215000 179.300000 ;
        RECT  5.015000 179.500000  5.215000 179.700000 ;
        RECT  5.015000 179.900000  5.215000 180.100000 ;
        RECT  5.015000 180.300000  5.215000 180.500000 ;
        RECT  5.015000 180.700000  5.215000 180.900000 ;
        RECT  5.015000 181.100000  5.215000 181.300000 ;
        RECT  5.015000 181.505000  5.215000 181.705000 ;
        RECT  5.015000 181.910000  5.215000 182.110000 ;
        RECT  5.015000 182.315000  5.215000 182.515000 ;
        RECT  5.015000 182.720000  5.215000 182.920000 ;
        RECT  5.015000 183.125000  5.215000 183.325000 ;
        RECT  5.015000 183.530000  5.215000 183.730000 ;
        RECT  5.015000 183.935000  5.215000 184.135000 ;
        RECT  5.015000 184.340000  5.215000 184.540000 ;
        RECT  5.015000 184.745000  5.215000 184.945000 ;
        RECT  5.015000 185.150000  5.215000 185.350000 ;
        RECT  5.015000 185.555000  5.215000 185.755000 ;
        RECT  5.015000 185.960000  5.215000 186.160000 ;
        RECT  5.015000 186.365000  5.215000 186.565000 ;
        RECT  5.015000 186.770000  5.215000 186.970000 ;
        RECT  5.015000 187.175000  5.215000 187.375000 ;
        RECT  5.015000 187.580000  5.215000 187.780000 ;
        RECT  5.015000 187.985000  5.215000 188.185000 ;
        RECT  5.015000 188.390000  5.215000 188.590000 ;
        RECT  5.015000 188.795000  5.215000 188.995000 ;
        RECT  5.015000 189.200000  5.215000 189.400000 ;
        RECT  5.015000 189.605000  5.215000 189.805000 ;
        RECT  5.015000 190.010000  5.215000 190.210000 ;
        RECT  5.015000 190.415000  5.215000 190.615000 ;
        RECT  5.015000 190.820000  5.215000 191.020000 ;
        RECT  5.015000 191.225000  5.215000 191.425000 ;
        RECT  5.015000 191.630000  5.215000 191.830000 ;
        RECT  5.015000 192.035000  5.215000 192.235000 ;
        RECT  5.015000 192.440000  5.215000 192.640000 ;
        RECT  5.015000 192.845000  5.215000 193.045000 ;
        RECT  5.015000 193.250000  5.215000 193.450000 ;
        RECT  5.015000 193.655000  5.215000 193.855000 ;
        RECT  5.015000 194.060000  5.215000 194.260000 ;
        RECT  5.015000 194.465000  5.215000 194.665000 ;
        RECT  5.015000 194.870000  5.215000 195.070000 ;
        RECT  5.015000 195.275000  5.215000 195.475000 ;
        RECT  5.015000 195.680000  5.215000 195.880000 ;
        RECT  5.015000 196.085000  5.215000 196.285000 ;
        RECT  5.015000 196.490000  5.215000 196.690000 ;
        RECT  5.015000 196.895000  5.215000 197.095000 ;
        RECT  5.015000 197.300000  5.215000 197.500000 ;
        RECT  5.015000 197.705000  5.215000 197.905000 ;
        RECT  5.075000  23.910000  5.275000  24.110000 ;
        RECT  5.075000  24.340000  5.275000  24.540000 ;
        RECT  5.075000  24.770000  5.275000  24.970000 ;
        RECT  5.075000  25.200000  5.275000  25.400000 ;
        RECT  5.075000  25.630000  5.275000  25.830000 ;
        RECT  5.075000  26.060000  5.275000  26.260000 ;
        RECT  5.075000  26.490000  5.275000  26.690000 ;
        RECT  5.075000  26.920000  5.275000  27.120000 ;
        RECT  5.075000  27.350000  5.275000  27.550000 ;
        RECT  5.075000  27.780000  5.275000  27.980000 ;
        RECT  5.075000  28.210000  5.275000  28.410000 ;
        RECT  5.415000 173.900000  5.615000 174.100000 ;
        RECT  5.415000 174.300000  5.615000 174.500000 ;
        RECT  5.415000 174.700000  5.615000 174.900000 ;
        RECT  5.415000 175.100000  5.615000 175.300000 ;
        RECT  5.415000 175.500000  5.615000 175.700000 ;
        RECT  5.415000 175.900000  5.615000 176.100000 ;
        RECT  5.415000 176.300000  5.615000 176.500000 ;
        RECT  5.415000 176.700000  5.615000 176.900000 ;
        RECT  5.415000 177.100000  5.615000 177.300000 ;
        RECT  5.415000 177.500000  5.615000 177.700000 ;
        RECT  5.415000 177.900000  5.615000 178.100000 ;
        RECT  5.415000 178.300000  5.615000 178.500000 ;
        RECT  5.415000 178.700000  5.615000 178.900000 ;
        RECT  5.415000 179.100000  5.615000 179.300000 ;
        RECT  5.415000 179.500000  5.615000 179.700000 ;
        RECT  5.415000 179.900000  5.615000 180.100000 ;
        RECT  5.415000 180.300000  5.615000 180.500000 ;
        RECT  5.415000 180.700000  5.615000 180.900000 ;
        RECT  5.415000 181.100000  5.615000 181.300000 ;
        RECT  5.415000 181.505000  5.615000 181.705000 ;
        RECT  5.415000 181.910000  5.615000 182.110000 ;
        RECT  5.415000 182.315000  5.615000 182.515000 ;
        RECT  5.415000 182.720000  5.615000 182.920000 ;
        RECT  5.415000 183.125000  5.615000 183.325000 ;
        RECT  5.415000 183.530000  5.615000 183.730000 ;
        RECT  5.415000 183.935000  5.615000 184.135000 ;
        RECT  5.415000 184.340000  5.615000 184.540000 ;
        RECT  5.415000 184.745000  5.615000 184.945000 ;
        RECT  5.415000 185.150000  5.615000 185.350000 ;
        RECT  5.415000 185.555000  5.615000 185.755000 ;
        RECT  5.415000 185.960000  5.615000 186.160000 ;
        RECT  5.415000 186.365000  5.615000 186.565000 ;
        RECT  5.415000 186.770000  5.615000 186.970000 ;
        RECT  5.415000 187.175000  5.615000 187.375000 ;
        RECT  5.415000 187.580000  5.615000 187.780000 ;
        RECT  5.415000 187.985000  5.615000 188.185000 ;
        RECT  5.415000 188.390000  5.615000 188.590000 ;
        RECT  5.415000 188.795000  5.615000 188.995000 ;
        RECT  5.415000 189.200000  5.615000 189.400000 ;
        RECT  5.415000 189.605000  5.615000 189.805000 ;
        RECT  5.415000 190.010000  5.615000 190.210000 ;
        RECT  5.415000 190.415000  5.615000 190.615000 ;
        RECT  5.415000 190.820000  5.615000 191.020000 ;
        RECT  5.415000 191.225000  5.615000 191.425000 ;
        RECT  5.415000 191.630000  5.615000 191.830000 ;
        RECT  5.415000 192.035000  5.615000 192.235000 ;
        RECT  5.415000 192.440000  5.615000 192.640000 ;
        RECT  5.415000 192.845000  5.615000 193.045000 ;
        RECT  5.415000 193.250000  5.615000 193.450000 ;
        RECT  5.415000 193.655000  5.615000 193.855000 ;
        RECT  5.415000 194.060000  5.615000 194.260000 ;
        RECT  5.415000 194.465000  5.615000 194.665000 ;
        RECT  5.415000 194.870000  5.615000 195.070000 ;
        RECT  5.415000 195.275000  5.615000 195.475000 ;
        RECT  5.415000 195.680000  5.615000 195.880000 ;
        RECT  5.415000 196.085000  5.615000 196.285000 ;
        RECT  5.415000 196.490000  5.615000 196.690000 ;
        RECT  5.415000 196.895000  5.615000 197.095000 ;
        RECT  5.415000 197.300000  5.615000 197.500000 ;
        RECT  5.415000 197.705000  5.615000 197.905000 ;
        RECT  5.480000  23.910000  5.680000  24.110000 ;
        RECT  5.480000  24.340000  5.680000  24.540000 ;
        RECT  5.480000  24.770000  5.680000  24.970000 ;
        RECT  5.480000  25.200000  5.680000  25.400000 ;
        RECT  5.480000  25.630000  5.680000  25.830000 ;
        RECT  5.480000  26.060000  5.680000  26.260000 ;
        RECT  5.480000  26.490000  5.680000  26.690000 ;
        RECT  5.480000  26.920000  5.680000  27.120000 ;
        RECT  5.480000  27.350000  5.680000  27.550000 ;
        RECT  5.480000  27.780000  5.680000  27.980000 ;
        RECT  5.480000  28.210000  5.680000  28.410000 ;
        RECT  5.815000 173.900000  6.015000 174.100000 ;
        RECT  5.815000 174.300000  6.015000 174.500000 ;
        RECT  5.815000 174.700000  6.015000 174.900000 ;
        RECT  5.815000 175.100000  6.015000 175.300000 ;
        RECT  5.815000 175.500000  6.015000 175.700000 ;
        RECT  5.815000 175.900000  6.015000 176.100000 ;
        RECT  5.815000 176.300000  6.015000 176.500000 ;
        RECT  5.815000 176.700000  6.015000 176.900000 ;
        RECT  5.815000 177.100000  6.015000 177.300000 ;
        RECT  5.815000 177.500000  6.015000 177.700000 ;
        RECT  5.815000 177.900000  6.015000 178.100000 ;
        RECT  5.815000 178.300000  6.015000 178.500000 ;
        RECT  5.815000 178.700000  6.015000 178.900000 ;
        RECT  5.815000 179.100000  6.015000 179.300000 ;
        RECT  5.815000 179.500000  6.015000 179.700000 ;
        RECT  5.815000 179.900000  6.015000 180.100000 ;
        RECT  5.815000 180.300000  6.015000 180.500000 ;
        RECT  5.815000 180.700000  6.015000 180.900000 ;
        RECT  5.815000 181.100000  6.015000 181.300000 ;
        RECT  5.815000 181.505000  6.015000 181.705000 ;
        RECT  5.815000 181.910000  6.015000 182.110000 ;
        RECT  5.815000 182.315000  6.015000 182.515000 ;
        RECT  5.815000 182.720000  6.015000 182.920000 ;
        RECT  5.815000 183.125000  6.015000 183.325000 ;
        RECT  5.815000 183.530000  6.015000 183.730000 ;
        RECT  5.815000 183.935000  6.015000 184.135000 ;
        RECT  5.815000 184.340000  6.015000 184.540000 ;
        RECT  5.815000 184.745000  6.015000 184.945000 ;
        RECT  5.815000 185.150000  6.015000 185.350000 ;
        RECT  5.815000 185.555000  6.015000 185.755000 ;
        RECT  5.815000 185.960000  6.015000 186.160000 ;
        RECT  5.815000 186.365000  6.015000 186.565000 ;
        RECT  5.815000 186.770000  6.015000 186.970000 ;
        RECT  5.815000 187.175000  6.015000 187.375000 ;
        RECT  5.815000 187.580000  6.015000 187.780000 ;
        RECT  5.815000 187.985000  6.015000 188.185000 ;
        RECT  5.815000 188.390000  6.015000 188.590000 ;
        RECT  5.815000 188.795000  6.015000 188.995000 ;
        RECT  5.815000 189.200000  6.015000 189.400000 ;
        RECT  5.815000 189.605000  6.015000 189.805000 ;
        RECT  5.815000 190.010000  6.015000 190.210000 ;
        RECT  5.815000 190.415000  6.015000 190.615000 ;
        RECT  5.815000 190.820000  6.015000 191.020000 ;
        RECT  5.815000 191.225000  6.015000 191.425000 ;
        RECT  5.815000 191.630000  6.015000 191.830000 ;
        RECT  5.815000 192.035000  6.015000 192.235000 ;
        RECT  5.815000 192.440000  6.015000 192.640000 ;
        RECT  5.815000 192.845000  6.015000 193.045000 ;
        RECT  5.815000 193.250000  6.015000 193.450000 ;
        RECT  5.815000 193.655000  6.015000 193.855000 ;
        RECT  5.815000 194.060000  6.015000 194.260000 ;
        RECT  5.815000 194.465000  6.015000 194.665000 ;
        RECT  5.815000 194.870000  6.015000 195.070000 ;
        RECT  5.815000 195.275000  6.015000 195.475000 ;
        RECT  5.815000 195.680000  6.015000 195.880000 ;
        RECT  5.815000 196.085000  6.015000 196.285000 ;
        RECT  5.815000 196.490000  6.015000 196.690000 ;
        RECT  5.815000 196.895000  6.015000 197.095000 ;
        RECT  5.815000 197.300000  6.015000 197.500000 ;
        RECT  5.815000 197.705000  6.015000 197.905000 ;
        RECT  5.885000  23.910000  6.085000  24.110000 ;
        RECT  5.885000  24.340000  6.085000  24.540000 ;
        RECT  5.885000  24.770000  6.085000  24.970000 ;
        RECT  5.885000  25.200000  6.085000  25.400000 ;
        RECT  5.885000  25.630000  6.085000  25.830000 ;
        RECT  5.885000  26.060000  6.085000  26.260000 ;
        RECT  5.885000  26.490000  6.085000  26.690000 ;
        RECT  5.885000  26.920000  6.085000  27.120000 ;
        RECT  5.885000  27.350000  6.085000  27.550000 ;
        RECT  5.885000  27.780000  6.085000  27.980000 ;
        RECT  5.885000  28.210000  6.085000  28.410000 ;
        RECT  6.215000 173.900000  6.415000 174.100000 ;
        RECT  6.215000 174.300000  6.415000 174.500000 ;
        RECT  6.215000 174.700000  6.415000 174.900000 ;
        RECT  6.215000 175.100000  6.415000 175.300000 ;
        RECT  6.215000 175.500000  6.415000 175.700000 ;
        RECT  6.215000 175.900000  6.415000 176.100000 ;
        RECT  6.215000 176.300000  6.415000 176.500000 ;
        RECT  6.215000 176.700000  6.415000 176.900000 ;
        RECT  6.215000 177.100000  6.415000 177.300000 ;
        RECT  6.215000 177.500000  6.415000 177.700000 ;
        RECT  6.215000 177.900000  6.415000 178.100000 ;
        RECT  6.215000 178.300000  6.415000 178.500000 ;
        RECT  6.215000 178.700000  6.415000 178.900000 ;
        RECT  6.215000 179.100000  6.415000 179.300000 ;
        RECT  6.215000 179.500000  6.415000 179.700000 ;
        RECT  6.215000 179.900000  6.415000 180.100000 ;
        RECT  6.215000 180.300000  6.415000 180.500000 ;
        RECT  6.215000 180.700000  6.415000 180.900000 ;
        RECT  6.215000 181.100000  6.415000 181.300000 ;
        RECT  6.215000 181.505000  6.415000 181.705000 ;
        RECT  6.215000 181.910000  6.415000 182.110000 ;
        RECT  6.215000 182.315000  6.415000 182.515000 ;
        RECT  6.215000 182.720000  6.415000 182.920000 ;
        RECT  6.215000 183.125000  6.415000 183.325000 ;
        RECT  6.215000 183.530000  6.415000 183.730000 ;
        RECT  6.215000 183.935000  6.415000 184.135000 ;
        RECT  6.215000 184.340000  6.415000 184.540000 ;
        RECT  6.215000 184.745000  6.415000 184.945000 ;
        RECT  6.215000 185.150000  6.415000 185.350000 ;
        RECT  6.215000 185.555000  6.415000 185.755000 ;
        RECT  6.215000 185.960000  6.415000 186.160000 ;
        RECT  6.215000 186.365000  6.415000 186.565000 ;
        RECT  6.215000 186.770000  6.415000 186.970000 ;
        RECT  6.215000 187.175000  6.415000 187.375000 ;
        RECT  6.215000 187.580000  6.415000 187.780000 ;
        RECT  6.215000 187.985000  6.415000 188.185000 ;
        RECT  6.215000 188.390000  6.415000 188.590000 ;
        RECT  6.215000 188.795000  6.415000 188.995000 ;
        RECT  6.215000 189.200000  6.415000 189.400000 ;
        RECT  6.215000 189.605000  6.415000 189.805000 ;
        RECT  6.215000 190.010000  6.415000 190.210000 ;
        RECT  6.215000 190.415000  6.415000 190.615000 ;
        RECT  6.215000 190.820000  6.415000 191.020000 ;
        RECT  6.215000 191.225000  6.415000 191.425000 ;
        RECT  6.215000 191.630000  6.415000 191.830000 ;
        RECT  6.215000 192.035000  6.415000 192.235000 ;
        RECT  6.215000 192.440000  6.415000 192.640000 ;
        RECT  6.215000 192.845000  6.415000 193.045000 ;
        RECT  6.215000 193.250000  6.415000 193.450000 ;
        RECT  6.215000 193.655000  6.415000 193.855000 ;
        RECT  6.215000 194.060000  6.415000 194.260000 ;
        RECT  6.215000 194.465000  6.415000 194.665000 ;
        RECT  6.215000 194.870000  6.415000 195.070000 ;
        RECT  6.215000 195.275000  6.415000 195.475000 ;
        RECT  6.215000 195.680000  6.415000 195.880000 ;
        RECT  6.215000 196.085000  6.415000 196.285000 ;
        RECT  6.215000 196.490000  6.415000 196.690000 ;
        RECT  6.215000 196.895000  6.415000 197.095000 ;
        RECT  6.215000 197.300000  6.415000 197.500000 ;
        RECT  6.215000 197.705000  6.415000 197.905000 ;
        RECT  6.290000  23.910000  6.490000  24.110000 ;
        RECT  6.290000  24.340000  6.490000  24.540000 ;
        RECT  6.290000  24.770000  6.490000  24.970000 ;
        RECT  6.290000  25.200000  6.490000  25.400000 ;
        RECT  6.290000  25.630000  6.490000  25.830000 ;
        RECT  6.290000  26.060000  6.490000  26.260000 ;
        RECT  6.290000  26.490000  6.490000  26.690000 ;
        RECT  6.290000  26.920000  6.490000  27.120000 ;
        RECT  6.290000  27.350000  6.490000  27.550000 ;
        RECT  6.290000  27.780000  6.490000  27.980000 ;
        RECT  6.290000  28.210000  6.490000  28.410000 ;
        RECT  6.615000 173.900000  6.815000 174.100000 ;
        RECT  6.615000 174.300000  6.815000 174.500000 ;
        RECT  6.615000 174.700000  6.815000 174.900000 ;
        RECT  6.615000 175.100000  6.815000 175.300000 ;
        RECT  6.615000 175.500000  6.815000 175.700000 ;
        RECT  6.615000 175.900000  6.815000 176.100000 ;
        RECT  6.615000 176.300000  6.815000 176.500000 ;
        RECT  6.615000 176.700000  6.815000 176.900000 ;
        RECT  6.615000 177.100000  6.815000 177.300000 ;
        RECT  6.615000 177.500000  6.815000 177.700000 ;
        RECT  6.615000 177.900000  6.815000 178.100000 ;
        RECT  6.615000 178.300000  6.815000 178.500000 ;
        RECT  6.615000 178.700000  6.815000 178.900000 ;
        RECT  6.615000 179.100000  6.815000 179.300000 ;
        RECT  6.615000 179.500000  6.815000 179.700000 ;
        RECT  6.615000 179.900000  6.815000 180.100000 ;
        RECT  6.615000 180.300000  6.815000 180.500000 ;
        RECT  6.615000 180.700000  6.815000 180.900000 ;
        RECT  6.615000 181.100000  6.815000 181.300000 ;
        RECT  6.615000 181.505000  6.815000 181.705000 ;
        RECT  6.615000 181.910000  6.815000 182.110000 ;
        RECT  6.615000 182.315000  6.815000 182.515000 ;
        RECT  6.615000 182.720000  6.815000 182.920000 ;
        RECT  6.615000 183.125000  6.815000 183.325000 ;
        RECT  6.615000 183.530000  6.815000 183.730000 ;
        RECT  6.615000 183.935000  6.815000 184.135000 ;
        RECT  6.615000 184.340000  6.815000 184.540000 ;
        RECT  6.615000 184.745000  6.815000 184.945000 ;
        RECT  6.615000 185.150000  6.815000 185.350000 ;
        RECT  6.615000 185.555000  6.815000 185.755000 ;
        RECT  6.615000 185.960000  6.815000 186.160000 ;
        RECT  6.615000 186.365000  6.815000 186.565000 ;
        RECT  6.615000 186.770000  6.815000 186.970000 ;
        RECT  6.615000 187.175000  6.815000 187.375000 ;
        RECT  6.615000 187.580000  6.815000 187.780000 ;
        RECT  6.615000 187.985000  6.815000 188.185000 ;
        RECT  6.615000 188.390000  6.815000 188.590000 ;
        RECT  6.615000 188.795000  6.815000 188.995000 ;
        RECT  6.615000 189.200000  6.815000 189.400000 ;
        RECT  6.615000 189.605000  6.815000 189.805000 ;
        RECT  6.615000 190.010000  6.815000 190.210000 ;
        RECT  6.615000 190.415000  6.815000 190.615000 ;
        RECT  6.615000 190.820000  6.815000 191.020000 ;
        RECT  6.615000 191.225000  6.815000 191.425000 ;
        RECT  6.615000 191.630000  6.815000 191.830000 ;
        RECT  6.615000 192.035000  6.815000 192.235000 ;
        RECT  6.615000 192.440000  6.815000 192.640000 ;
        RECT  6.615000 192.845000  6.815000 193.045000 ;
        RECT  6.615000 193.250000  6.815000 193.450000 ;
        RECT  6.615000 193.655000  6.815000 193.855000 ;
        RECT  6.615000 194.060000  6.815000 194.260000 ;
        RECT  6.615000 194.465000  6.815000 194.665000 ;
        RECT  6.615000 194.870000  6.815000 195.070000 ;
        RECT  6.615000 195.275000  6.815000 195.475000 ;
        RECT  6.615000 195.680000  6.815000 195.880000 ;
        RECT  6.615000 196.085000  6.815000 196.285000 ;
        RECT  6.615000 196.490000  6.815000 196.690000 ;
        RECT  6.615000 196.895000  6.815000 197.095000 ;
        RECT  6.615000 197.300000  6.815000 197.500000 ;
        RECT  6.615000 197.705000  6.815000 197.905000 ;
        RECT  6.695000  23.910000  6.895000  24.110000 ;
        RECT  6.695000  24.340000  6.895000  24.540000 ;
        RECT  6.695000  24.770000  6.895000  24.970000 ;
        RECT  6.695000  25.200000  6.895000  25.400000 ;
        RECT  6.695000  25.630000  6.895000  25.830000 ;
        RECT  6.695000  26.060000  6.895000  26.260000 ;
        RECT  6.695000  26.490000  6.895000  26.690000 ;
        RECT  6.695000  26.920000  6.895000  27.120000 ;
        RECT  6.695000  27.350000  6.895000  27.550000 ;
        RECT  6.695000  27.780000  6.895000  27.980000 ;
        RECT  6.695000  28.210000  6.895000  28.410000 ;
        RECT  7.015000 173.900000  7.215000 174.100000 ;
        RECT  7.015000 174.300000  7.215000 174.500000 ;
        RECT  7.015000 174.700000  7.215000 174.900000 ;
        RECT  7.015000 175.100000  7.215000 175.300000 ;
        RECT  7.015000 175.500000  7.215000 175.700000 ;
        RECT  7.015000 175.900000  7.215000 176.100000 ;
        RECT  7.015000 176.300000  7.215000 176.500000 ;
        RECT  7.015000 176.700000  7.215000 176.900000 ;
        RECT  7.015000 177.100000  7.215000 177.300000 ;
        RECT  7.015000 177.500000  7.215000 177.700000 ;
        RECT  7.015000 177.900000  7.215000 178.100000 ;
        RECT  7.015000 178.300000  7.215000 178.500000 ;
        RECT  7.015000 178.700000  7.215000 178.900000 ;
        RECT  7.015000 179.100000  7.215000 179.300000 ;
        RECT  7.015000 179.500000  7.215000 179.700000 ;
        RECT  7.015000 179.900000  7.215000 180.100000 ;
        RECT  7.015000 180.300000  7.215000 180.500000 ;
        RECT  7.015000 180.700000  7.215000 180.900000 ;
        RECT  7.015000 181.100000  7.215000 181.300000 ;
        RECT  7.015000 181.505000  7.215000 181.705000 ;
        RECT  7.015000 181.910000  7.215000 182.110000 ;
        RECT  7.015000 182.315000  7.215000 182.515000 ;
        RECT  7.015000 182.720000  7.215000 182.920000 ;
        RECT  7.015000 183.125000  7.215000 183.325000 ;
        RECT  7.015000 183.530000  7.215000 183.730000 ;
        RECT  7.015000 183.935000  7.215000 184.135000 ;
        RECT  7.015000 184.340000  7.215000 184.540000 ;
        RECT  7.015000 184.745000  7.215000 184.945000 ;
        RECT  7.015000 185.150000  7.215000 185.350000 ;
        RECT  7.015000 185.555000  7.215000 185.755000 ;
        RECT  7.015000 185.960000  7.215000 186.160000 ;
        RECT  7.015000 186.365000  7.215000 186.565000 ;
        RECT  7.015000 186.770000  7.215000 186.970000 ;
        RECT  7.015000 187.175000  7.215000 187.375000 ;
        RECT  7.015000 187.580000  7.215000 187.780000 ;
        RECT  7.015000 187.985000  7.215000 188.185000 ;
        RECT  7.015000 188.390000  7.215000 188.590000 ;
        RECT  7.015000 188.795000  7.215000 188.995000 ;
        RECT  7.015000 189.200000  7.215000 189.400000 ;
        RECT  7.015000 189.605000  7.215000 189.805000 ;
        RECT  7.015000 190.010000  7.215000 190.210000 ;
        RECT  7.015000 190.415000  7.215000 190.615000 ;
        RECT  7.015000 190.820000  7.215000 191.020000 ;
        RECT  7.015000 191.225000  7.215000 191.425000 ;
        RECT  7.015000 191.630000  7.215000 191.830000 ;
        RECT  7.015000 192.035000  7.215000 192.235000 ;
        RECT  7.015000 192.440000  7.215000 192.640000 ;
        RECT  7.015000 192.845000  7.215000 193.045000 ;
        RECT  7.015000 193.250000  7.215000 193.450000 ;
        RECT  7.015000 193.655000  7.215000 193.855000 ;
        RECT  7.015000 194.060000  7.215000 194.260000 ;
        RECT  7.015000 194.465000  7.215000 194.665000 ;
        RECT  7.015000 194.870000  7.215000 195.070000 ;
        RECT  7.015000 195.275000  7.215000 195.475000 ;
        RECT  7.015000 195.680000  7.215000 195.880000 ;
        RECT  7.015000 196.085000  7.215000 196.285000 ;
        RECT  7.015000 196.490000  7.215000 196.690000 ;
        RECT  7.015000 196.895000  7.215000 197.095000 ;
        RECT  7.015000 197.300000  7.215000 197.500000 ;
        RECT  7.015000 197.705000  7.215000 197.905000 ;
        RECT  7.100000  23.910000  7.300000  24.110000 ;
        RECT  7.100000  24.340000  7.300000  24.540000 ;
        RECT  7.100000  24.770000  7.300000  24.970000 ;
        RECT  7.100000  25.200000  7.300000  25.400000 ;
        RECT  7.100000  25.630000  7.300000  25.830000 ;
        RECT  7.100000  26.060000  7.300000  26.260000 ;
        RECT  7.100000  26.490000  7.300000  26.690000 ;
        RECT  7.100000  26.920000  7.300000  27.120000 ;
        RECT  7.100000  27.350000  7.300000  27.550000 ;
        RECT  7.100000  27.780000  7.300000  27.980000 ;
        RECT  7.100000  28.210000  7.300000  28.410000 ;
        RECT  7.415000 173.900000  7.615000 174.100000 ;
        RECT  7.415000 174.300000  7.615000 174.500000 ;
        RECT  7.415000 174.700000  7.615000 174.900000 ;
        RECT  7.415000 175.100000  7.615000 175.300000 ;
        RECT  7.415000 175.500000  7.615000 175.700000 ;
        RECT  7.415000 175.900000  7.615000 176.100000 ;
        RECT  7.415000 176.300000  7.615000 176.500000 ;
        RECT  7.415000 176.700000  7.615000 176.900000 ;
        RECT  7.415000 177.100000  7.615000 177.300000 ;
        RECT  7.415000 177.500000  7.615000 177.700000 ;
        RECT  7.415000 177.900000  7.615000 178.100000 ;
        RECT  7.415000 178.300000  7.615000 178.500000 ;
        RECT  7.415000 178.700000  7.615000 178.900000 ;
        RECT  7.415000 179.100000  7.615000 179.300000 ;
        RECT  7.415000 179.500000  7.615000 179.700000 ;
        RECT  7.415000 179.900000  7.615000 180.100000 ;
        RECT  7.415000 180.300000  7.615000 180.500000 ;
        RECT  7.415000 180.700000  7.615000 180.900000 ;
        RECT  7.415000 181.100000  7.615000 181.300000 ;
        RECT  7.415000 181.505000  7.615000 181.705000 ;
        RECT  7.415000 181.910000  7.615000 182.110000 ;
        RECT  7.415000 182.315000  7.615000 182.515000 ;
        RECT  7.415000 182.720000  7.615000 182.920000 ;
        RECT  7.415000 183.125000  7.615000 183.325000 ;
        RECT  7.415000 183.530000  7.615000 183.730000 ;
        RECT  7.415000 183.935000  7.615000 184.135000 ;
        RECT  7.415000 184.340000  7.615000 184.540000 ;
        RECT  7.415000 184.745000  7.615000 184.945000 ;
        RECT  7.415000 185.150000  7.615000 185.350000 ;
        RECT  7.415000 185.555000  7.615000 185.755000 ;
        RECT  7.415000 185.960000  7.615000 186.160000 ;
        RECT  7.415000 186.365000  7.615000 186.565000 ;
        RECT  7.415000 186.770000  7.615000 186.970000 ;
        RECT  7.415000 187.175000  7.615000 187.375000 ;
        RECT  7.415000 187.580000  7.615000 187.780000 ;
        RECT  7.415000 187.985000  7.615000 188.185000 ;
        RECT  7.415000 188.390000  7.615000 188.590000 ;
        RECT  7.415000 188.795000  7.615000 188.995000 ;
        RECT  7.415000 189.200000  7.615000 189.400000 ;
        RECT  7.415000 189.605000  7.615000 189.805000 ;
        RECT  7.415000 190.010000  7.615000 190.210000 ;
        RECT  7.415000 190.415000  7.615000 190.615000 ;
        RECT  7.415000 190.820000  7.615000 191.020000 ;
        RECT  7.415000 191.225000  7.615000 191.425000 ;
        RECT  7.415000 191.630000  7.615000 191.830000 ;
        RECT  7.415000 192.035000  7.615000 192.235000 ;
        RECT  7.415000 192.440000  7.615000 192.640000 ;
        RECT  7.415000 192.845000  7.615000 193.045000 ;
        RECT  7.415000 193.250000  7.615000 193.450000 ;
        RECT  7.415000 193.655000  7.615000 193.855000 ;
        RECT  7.415000 194.060000  7.615000 194.260000 ;
        RECT  7.415000 194.465000  7.615000 194.665000 ;
        RECT  7.415000 194.870000  7.615000 195.070000 ;
        RECT  7.415000 195.275000  7.615000 195.475000 ;
        RECT  7.415000 195.680000  7.615000 195.880000 ;
        RECT  7.415000 196.085000  7.615000 196.285000 ;
        RECT  7.415000 196.490000  7.615000 196.690000 ;
        RECT  7.415000 196.895000  7.615000 197.095000 ;
        RECT  7.415000 197.300000  7.615000 197.500000 ;
        RECT  7.415000 197.705000  7.615000 197.905000 ;
        RECT  7.505000  23.910000  7.705000  24.110000 ;
        RECT  7.505000  24.340000  7.705000  24.540000 ;
        RECT  7.505000  24.770000  7.705000  24.970000 ;
        RECT  7.505000  25.200000  7.705000  25.400000 ;
        RECT  7.505000  25.630000  7.705000  25.830000 ;
        RECT  7.505000  26.060000  7.705000  26.260000 ;
        RECT  7.505000  26.490000  7.705000  26.690000 ;
        RECT  7.505000  26.920000  7.705000  27.120000 ;
        RECT  7.505000  27.350000  7.705000  27.550000 ;
        RECT  7.505000  27.780000  7.705000  27.980000 ;
        RECT  7.505000  28.210000  7.705000  28.410000 ;
        RECT  7.815000 173.900000  8.015000 174.100000 ;
        RECT  7.815000 174.300000  8.015000 174.500000 ;
        RECT  7.815000 174.700000  8.015000 174.900000 ;
        RECT  7.815000 175.100000  8.015000 175.300000 ;
        RECT  7.815000 175.500000  8.015000 175.700000 ;
        RECT  7.815000 175.900000  8.015000 176.100000 ;
        RECT  7.815000 176.300000  8.015000 176.500000 ;
        RECT  7.815000 176.700000  8.015000 176.900000 ;
        RECT  7.815000 177.100000  8.015000 177.300000 ;
        RECT  7.815000 177.500000  8.015000 177.700000 ;
        RECT  7.815000 177.900000  8.015000 178.100000 ;
        RECT  7.815000 178.300000  8.015000 178.500000 ;
        RECT  7.815000 178.700000  8.015000 178.900000 ;
        RECT  7.815000 179.100000  8.015000 179.300000 ;
        RECT  7.815000 179.500000  8.015000 179.700000 ;
        RECT  7.815000 179.900000  8.015000 180.100000 ;
        RECT  7.815000 180.300000  8.015000 180.500000 ;
        RECT  7.815000 180.700000  8.015000 180.900000 ;
        RECT  7.815000 181.100000  8.015000 181.300000 ;
        RECT  7.815000 181.505000  8.015000 181.705000 ;
        RECT  7.815000 181.910000  8.015000 182.110000 ;
        RECT  7.815000 182.315000  8.015000 182.515000 ;
        RECT  7.815000 182.720000  8.015000 182.920000 ;
        RECT  7.815000 183.125000  8.015000 183.325000 ;
        RECT  7.815000 183.530000  8.015000 183.730000 ;
        RECT  7.815000 183.935000  8.015000 184.135000 ;
        RECT  7.815000 184.340000  8.015000 184.540000 ;
        RECT  7.815000 184.745000  8.015000 184.945000 ;
        RECT  7.815000 185.150000  8.015000 185.350000 ;
        RECT  7.815000 185.555000  8.015000 185.755000 ;
        RECT  7.815000 185.960000  8.015000 186.160000 ;
        RECT  7.815000 186.365000  8.015000 186.565000 ;
        RECT  7.815000 186.770000  8.015000 186.970000 ;
        RECT  7.815000 187.175000  8.015000 187.375000 ;
        RECT  7.815000 187.580000  8.015000 187.780000 ;
        RECT  7.815000 187.985000  8.015000 188.185000 ;
        RECT  7.815000 188.390000  8.015000 188.590000 ;
        RECT  7.815000 188.795000  8.015000 188.995000 ;
        RECT  7.815000 189.200000  8.015000 189.400000 ;
        RECT  7.815000 189.605000  8.015000 189.805000 ;
        RECT  7.815000 190.010000  8.015000 190.210000 ;
        RECT  7.815000 190.415000  8.015000 190.615000 ;
        RECT  7.815000 190.820000  8.015000 191.020000 ;
        RECT  7.815000 191.225000  8.015000 191.425000 ;
        RECT  7.815000 191.630000  8.015000 191.830000 ;
        RECT  7.815000 192.035000  8.015000 192.235000 ;
        RECT  7.815000 192.440000  8.015000 192.640000 ;
        RECT  7.815000 192.845000  8.015000 193.045000 ;
        RECT  7.815000 193.250000  8.015000 193.450000 ;
        RECT  7.815000 193.655000  8.015000 193.855000 ;
        RECT  7.815000 194.060000  8.015000 194.260000 ;
        RECT  7.815000 194.465000  8.015000 194.665000 ;
        RECT  7.815000 194.870000  8.015000 195.070000 ;
        RECT  7.815000 195.275000  8.015000 195.475000 ;
        RECT  7.815000 195.680000  8.015000 195.880000 ;
        RECT  7.815000 196.085000  8.015000 196.285000 ;
        RECT  7.815000 196.490000  8.015000 196.690000 ;
        RECT  7.815000 196.895000  8.015000 197.095000 ;
        RECT  7.815000 197.300000  8.015000 197.500000 ;
        RECT  7.815000 197.705000  8.015000 197.905000 ;
        RECT  7.910000  23.910000  8.110000  24.110000 ;
        RECT  7.910000  24.340000  8.110000  24.540000 ;
        RECT  7.910000  24.770000  8.110000  24.970000 ;
        RECT  7.910000  25.200000  8.110000  25.400000 ;
        RECT  7.910000  25.630000  8.110000  25.830000 ;
        RECT  7.910000  26.060000  8.110000  26.260000 ;
        RECT  7.910000  26.490000  8.110000  26.690000 ;
        RECT  7.910000  26.920000  8.110000  27.120000 ;
        RECT  7.910000  27.350000  8.110000  27.550000 ;
        RECT  7.910000  27.780000  8.110000  27.980000 ;
        RECT  7.910000  28.210000  8.110000  28.410000 ;
        RECT  8.215000 173.900000  8.415000 174.100000 ;
        RECT  8.215000 174.300000  8.415000 174.500000 ;
        RECT  8.215000 174.700000  8.415000 174.900000 ;
        RECT  8.215000 175.100000  8.415000 175.300000 ;
        RECT  8.215000 175.500000  8.415000 175.700000 ;
        RECT  8.215000 175.900000  8.415000 176.100000 ;
        RECT  8.215000 176.300000  8.415000 176.500000 ;
        RECT  8.215000 176.700000  8.415000 176.900000 ;
        RECT  8.215000 177.100000  8.415000 177.300000 ;
        RECT  8.215000 177.500000  8.415000 177.700000 ;
        RECT  8.215000 177.900000  8.415000 178.100000 ;
        RECT  8.215000 178.300000  8.415000 178.500000 ;
        RECT  8.215000 178.700000  8.415000 178.900000 ;
        RECT  8.215000 179.100000  8.415000 179.300000 ;
        RECT  8.215000 179.500000  8.415000 179.700000 ;
        RECT  8.215000 179.900000  8.415000 180.100000 ;
        RECT  8.215000 180.300000  8.415000 180.500000 ;
        RECT  8.215000 180.700000  8.415000 180.900000 ;
        RECT  8.215000 181.100000  8.415000 181.300000 ;
        RECT  8.215000 181.505000  8.415000 181.705000 ;
        RECT  8.215000 181.910000  8.415000 182.110000 ;
        RECT  8.215000 182.315000  8.415000 182.515000 ;
        RECT  8.215000 182.720000  8.415000 182.920000 ;
        RECT  8.215000 183.125000  8.415000 183.325000 ;
        RECT  8.215000 183.530000  8.415000 183.730000 ;
        RECT  8.215000 183.935000  8.415000 184.135000 ;
        RECT  8.215000 184.340000  8.415000 184.540000 ;
        RECT  8.215000 184.745000  8.415000 184.945000 ;
        RECT  8.215000 185.150000  8.415000 185.350000 ;
        RECT  8.215000 185.555000  8.415000 185.755000 ;
        RECT  8.215000 185.960000  8.415000 186.160000 ;
        RECT  8.215000 186.365000  8.415000 186.565000 ;
        RECT  8.215000 186.770000  8.415000 186.970000 ;
        RECT  8.215000 187.175000  8.415000 187.375000 ;
        RECT  8.215000 187.580000  8.415000 187.780000 ;
        RECT  8.215000 187.985000  8.415000 188.185000 ;
        RECT  8.215000 188.390000  8.415000 188.590000 ;
        RECT  8.215000 188.795000  8.415000 188.995000 ;
        RECT  8.215000 189.200000  8.415000 189.400000 ;
        RECT  8.215000 189.605000  8.415000 189.805000 ;
        RECT  8.215000 190.010000  8.415000 190.210000 ;
        RECT  8.215000 190.415000  8.415000 190.615000 ;
        RECT  8.215000 190.820000  8.415000 191.020000 ;
        RECT  8.215000 191.225000  8.415000 191.425000 ;
        RECT  8.215000 191.630000  8.415000 191.830000 ;
        RECT  8.215000 192.035000  8.415000 192.235000 ;
        RECT  8.215000 192.440000  8.415000 192.640000 ;
        RECT  8.215000 192.845000  8.415000 193.045000 ;
        RECT  8.215000 193.250000  8.415000 193.450000 ;
        RECT  8.215000 193.655000  8.415000 193.855000 ;
        RECT  8.215000 194.060000  8.415000 194.260000 ;
        RECT  8.215000 194.465000  8.415000 194.665000 ;
        RECT  8.215000 194.870000  8.415000 195.070000 ;
        RECT  8.215000 195.275000  8.415000 195.475000 ;
        RECT  8.215000 195.680000  8.415000 195.880000 ;
        RECT  8.215000 196.085000  8.415000 196.285000 ;
        RECT  8.215000 196.490000  8.415000 196.690000 ;
        RECT  8.215000 196.895000  8.415000 197.095000 ;
        RECT  8.215000 197.300000  8.415000 197.500000 ;
        RECT  8.215000 197.705000  8.415000 197.905000 ;
        RECT  8.315000  23.910000  8.515000  24.110000 ;
        RECT  8.315000  24.340000  8.515000  24.540000 ;
        RECT  8.315000  24.770000  8.515000  24.970000 ;
        RECT  8.315000  25.200000  8.515000  25.400000 ;
        RECT  8.315000  25.630000  8.515000  25.830000 ;
        RECT  8.315000  26.060000  8.515000  26.260000 ;
        RECT  8.315000  26.490000  8.515000  26.690000 ;
        RECT  8.315000  26.920000  8.515000  27.120000 ;
        RECT  8.315000  27.350000  8.515000  27.550000 ;
        RECT  8.315000  27.780000  8.515000  27.980000 ;
        RECT  8.315000  28.210000  8.515000  28.410000 ;
        RECT  8.615000 173.900000  8.815000 174.100000 ;
        RECT  8.615000 174.300000  8.815000 174.500000 ;
        RECT  8.615000 174.700000  8.815000 174.900000 ;
        RECT  8.615000 175.100000  8.815000 175.300000 ;
        RECT  8.615000 175.500000  8.815000 175.700000 ;
        RECT  8.615000 175.900000  8.815000 176.100000 ;
        RECT  8.615000 176.300000  8.815000 176.500000 ;
        RECT  8.615000 176.700000  8.815000 176.900000 ;
        RECT  8.615000 177.100000  8.815000 177.300000 ;
        RECT  8.615000 177.500000  8.815000 177.700000 ;
        RECT  8.615000 177.900000  8.815000 178.100000 ;
        RECT  8.615000 178.300000  8.815000 178.500000 ;
        RECT  8.615000 178.700000  8.815000 178.900000 ;
        RECT  8.615000 179.100000  8.815000 179.300000 ;
        RECT  8.615000 179.500000  8.815000 179.700000 ;
        RECT  8.615000 179.900000  8.815000 180.100000 ;
        RECT  8.615000 180.300000  8.815000 180.500000 ;
        RECT  8.615000 180.700000  8.815000 180.900000 ;
        RECT  8.615000 181.100000  8.815000 181.300000 ;
        RECT  8.615000 181.505000  8.815000 181.705000 ;
        RECT  8.615000 181.910000  8.815000 182.110000 ;
        RECT  8.615000 182.315000  8.815000 182.515000 ;
        RECT  8.615000 182.720000  8.815000 182.920000 ;
        RECT  8.615000 183.125000  8.815000 183.325000 ;
        RECT  8.615000 183.530000  8.815000 183.730000 ;
        RECT  8.615000 183.935000  8.815000 184.135000 ;
        RECT  8.615000 184.340000  8.815000 184.540000 ;
        RECT  8.615000 184.745000  8.815000 184.945000 ;
        RECT  8.615000 185.150000  8.815000 185.350000 ;
        RECT  8.615000 185.555000  8.815000 185.755000 ;
        RECT  8.615000 185.960000  8.815000 186.160000 ;
        RECT  8.615000 186.365000  8.815000 186.565000 ;
        RECT  8.615000 186.770000  8.815000 186.970000 ;
        RECT  8.615000 187.175000  8.815000 187.375000 ;
        RECT  8.615000 187.580000  8.815000 187.780000 ;
        RECT  8.615000 187.985000  8.815000 188.185000 ;
        RECT  8.615000 188.390000  8.815000 188.590000 ;
        RECT  8.615000 188.795000  8.815000 188.995000 ;
        RECT  8.615000 189.200000  8.815000 189.400000 ;
        RECT  8.615000 189.605000  8.815000 189.805000 ;
        RECT  8.615000 190.010000  8.815000 190.210000 ;
        RECT  8.615000 190.415000  8.815000 190.615000 ;
        RECT  8.615000 190.820000  8.815000 191.020000 ;
        RECT  8.615000 191.225000  8.815000 191.425000 ;
        RECT  8.615000 191.630000  8.815000 191.830000 ;
        RECT  8.615000 192.035000  8.815000 192.235000 ;
        RECT  8.615000 192.440000  8.815000 192.640000 ;
        RECT  8.615000 192.845000  8.815000 193.045000 ;
        RECT  8.615000 193.250000  8.815000 193.450000 ;
        RECT  8.615000 193.655000  8.815000 193.855000 ;
        RECT  8.615000 194.060000  8.815000 194.260000 ;
        RECT  8.615000 194.465000  8.815000 194.665000 ;
        RECT  8.615000 194.870000  8.815000 195.070000 ;
        RECT  8.615000 195.275000  8.815000 195.475000 ;
        RECT  8.615000 195.680000  8.815000 195.880000 ;
        RECT  8.615000 196.085000  8.815000 196.285000 ;
        RECT  8.615000 196.490000  8.815000 196.690000 ;
        RECT  8.615000 196.895000  8.815000 197.095000 ;
        RECT  8.615000 197.300000  8.815000 197.500000 ;
        RECT  8.615000 197.705000  8.815000 197.905000 ;
        RECT  8.720000  23.910000  8.920000  24.110000 ;
        RECT  8.720000  24.340000  8.920000  24.540000 ;
        RECT  8.720000  24.770000  8.920000  24.970000 ;
        RECT  8.720000  25.200000  8.920000  25.400000 ;
        RECT  8.720000  25.630000  8.920000  25.830000 ;
        RECT  8.720000  26.060000  8.920000  26.260000 ;
        RECT  8.720000  26.490000  8.920000  26.690000 ;
        RECT  8.720000  26.920000  8.920000  27.120000 ;
        RECT  8.720000  27.350000  8.920000  27.550000 ;
        RECT  8.720000  27.780000  8.920000  27.980000 ;
        RECT  8.720000  28.210000  8.920000  28.410000 ;
        RECT  9.015000 173.900000  9.215000 174.100000 ;
        RECT  9.015000 174.300000  9.215000 174.500000 ;
        RECT  9.015000 174.700000  9.215000 174.900000 ;
        RECT  9.015000 175.100000  9.215000 175.300000 ;
        RECT  9.015000 175.500000  9.215000 175.700000 ;
        RECT  9.015000 175.900000  9.215000 176.100000 ;
        RECT  9.015000 176.300000  9.215000 176.500000 ;
        RECT  9.015000 176.700000  9.215000 176.900000 ;
        RECT  9.015000 177.100000  9.215000 177.300000 ;
        RECT  9.015000 177.500000  9.215000 177.700000 ;
        RECT  9.015000 177.900000  9.215000 178.100000 ;
        RECT  9.015000 178.300000  9.215000 178.500000 ;
        RECT  9.015000 178.700000  9.215000 178.900000 ;
        RECT  9.015000 179.100000  9.215000 179.300000 ;
        RECT  9.015000 179.500000  9.215000 179.700000 ;
        RECT  9.015000 179.900000  9.215000 180.100000 ;
        RECT  9.015000 180.300000  9.215000 180.500000 ;
        RECT  9.015000 180.700000  9.215000 180.900000 ;
        RECT  9.015000 181.100000  9.215000 181.300000 ;
        RECT  9.015000 181.505000  9.215000 181.705000 ;
        RECT  9.015000 181.910000  9.215000 182.110000 ;
        RECT  9.015000 182.315000  9.215000 182.515000 ;
        RECT  9.015000 182.720000  9.215000 182.920000 ;
        RECT  9.015000 183.125000  9.215000 183.325000 ;
        RECT  9.015000 183.530000  9.215000 183.730000 ;
        RECT  9.015000 183.935000  9.215000 184.135000 ;
        RECT  9.015000 184.340000  9.215000 184.540000 ;
        RECT  9.015000 184.745000  9.215000 184.945000 ;
        RECT  9.015000 185.150000  9.215000 185.350000 ;
        RECT  9.015000 185.555000  9.215000 185.755000 ;
        RECT  9.015000 185.960000  9.215000 186.160000 ;
        RECT  9.015000 186.365000  9.215000 186.565000 ;
        RECT  9.015000 186.770000  9.215000 186.970000 ;
        RECT  9.015000 187.175000  9.215000 187.375000 ;
        RECT  9.015000 187.580000  9.215000 187.780000 ;
        RECT  9.015000 187.985000  9.215000 188.185000 ;
        RECT  9.015000 188.390000  9.215000 188.590000 ;
        RECT  9.015000 188.795000  9.215000 188.995000 ;
        RECT  9.015000 189.200000  9.215000 189.400000 ;
        RECT  9.015000 189.605000  9.215000 189.805000 ;
        RECT  9.015000 190.010000  9.215000 190.210000 ;
        RECT  9.015000 190.415000  9.215000 190.615000 ;
        RECT  9.015000 190.820000  9.215000 191.020000 ;
        RECT  9.015000 191.225000  9.215000 191.425000 ;
        RECT  9.015000 191.630000  9.215000 191.830000 ;
        RECT  9.015000 192.035000  9.215000 192.235000 ;
        RECT  9.015000 192.440000  9.215000 192.640000 ;
        RECT  9.015000 192.845000  9.215000 193.045000 ;
        RECT  9.015000 193.250000  9.215000 193.450000 ;
        RECT  9.015000 193.655000  9.215000 193.855000 ;
        RECT  9.015000 194.060000  9.215000 194.260000 ;
        RECT  9.015000 194.465000  9.215000 194.665000 ;
        RECT  9.015000 194.870000  9.215000 195.070000 ;
        RECT  9.015000 195.275000  9.215000 195.475000 ;
        RECT  9.015000 195.680000  9.215000 195.880000 ;
        RECT  9.015000 196.085000  9.215000 196.285000 ;
        RECT  9.015000 196.490000  9.215000 196.690000 ;
        RECT  9.015000 196.895000  9.215000 197.095000 ;
        RECT  9.015000 197.300000  9.215000 197.500000 ;
        RECT  9.015000 197.705000  9.215000 197.905000 ;
        RECT  9.125000  23.910000  9.325000  24.110000 ;
        RECT  9.125000  24.340000  9.325000  24.540000 ;
        RECT  9.125000  24.770000  9.325000  24.970000 ;
        RECT  9.125000  25.200000  9.325000  25.400000 ;
        RECT  9.125000  25.630000  9.325000  25.830000 ;
        RECT  9.125000  26.060000  9.325000  26.260000 ;
        RECT  9.125000  26.490000  9.325000  26.690000 ;
        RECT  9.125000  26.920000  9.325000  27.120000 ;
        RECT  9.125000  27.350000  9.325000  27.550000 ;
        RECT  9.125000  27.780000  9.325000  27.980000 ;
        RECT  9.125000  28.210000  9.325000  28.410000 ;
        RECT  9.415000 173.900000  9.615000 174.100000 ;
        RECT  9.415000 174.300000  9.615000 174.500000 ;
        RECT  9.415000 174.700000  9.615000 174.900000 ;
        RECT  9.415000 175.100000  9.615000 175.300000 ;
        RECT  9.415000 175.500000  9.615000 175.700000 ;
        RECT  9.415000 175.900000  9.615000 176.100000 ;
        RECT  9.415000 176.300000  9.615000 176.500000 ;
        RECT  9.415000 176.700000  9.615000 176.900000 ;
        RECT  9.415000 177.100000  9.615000 177.300000 ;
        RECT  9.415000 177.500000  9.615000 177.700000 ;
        RECT  9.415000 177.900000  9.615000 178.100000 ;
        RECT  9.415000 178.300000  9.615000 178.500000 ;
        RECT  9.415000 178.700000  9.615000 178.900000 ;
        RECT  9.415000 179.100000  9.615000 179.300000 ;
        RECT  9.415000 179.500000  9.615000 179.700000 ;
        RECT  9.415000 179.900000  9.615000 180.100000 ;
        RECT  9.415000 180.300000  9.615000 180.500000 ;
        RECT  9.415000 180.700000  9.615000 180.900000 ;
        RECT  9.415000 181.100000  9.615000 181.300000 ;
        RECT  9.415000 181.505000  9.615000 181.705000 ;
        RECT  9.415000 181.910000  9.615000 182.110000 ;
        RECT  9.415000 182.315000  9.615000 182.515000 ;
        RECT  9.415000 182.720000  9.615000 182.920000 ;
        RECT  9.415000 183.125000  9.615000 183.325000 ;
        RECT  9.415000 183.530000  9.615000 183.730000 ;
        RECT  9.415000 183.935000  9.615000 184.135000 ;
        RECT  9.415000 184.340000  9.615000 184.540000 ;
        RECT  9.415000 184.745000  9.615000 184.945000 ;
        RECT  9.415000 185.150000  9.615000 185.350000 ;
        RECT  9.415000 185.555000  9.615000 185.755000 ;
        RECT  9.415000 185.960000  9.615000 186.160000 ;
        RECT  9.415000 186.365000  9.615000 186.565000 ;
        RECT  9.415000 186.770000  9.615000 186.970000 ;
        RECT  9.415000 187.175000  9.615000 187.375000 ;
        RECT  9.415000 187.580000  9.615000 187.780000 ;
        RECT  9.415000 187.985000  9.615000 188.185000 ;
        RECT  9.415000 188.390000  9.615000 188.590000 ;
        RECT  9.415000 188.795000  9.615000 188.995000 ;
        RECT  9.415000 189.200000  9.615000 189.400000 ;
        RECT  9.415000 189.605000  9.615000 189.805000 ;
        RECT  9.415000 190.010000  9.615000 190.210000 ;
        RECT  9.415000 190.415000  9.615000 190.615000 ;
        RECT  9.415000 190.820000  9.615000 191.020000 ;
        RECT  9.415000 191.225000  9.615000 191.425000 ;
        RECT  9.415000 191.630000  9.615000 191.830000 ;
        RECT  9.415000 192.035000  9.615000 192.235000 ;
        RECT  9.415000 192.440000  9.615000 192.640000 ;
        RECT  9.415000 192.845000  9.615000 193.045000 ;
        RECT  9.415000 193.250000  9.615000 193.450000 ;
        RECT  9.415000 193.655000  9.615000 193.855000 ;
        RECT  9.415000 194.060000  9.615000 194.260000 ;
        RECT  9.415000 194.465000  9.615000 194.665000 ;
        RECT  9.415000 194.870000  9.615000 195.070000 ;
        RECT  9.415000 195.275000  9.615000 195.475000 ;
        RECT  9.415000 195.680000  9.615000 195.880000 ;
        RECT  9.415000 196.085000  9.615000 196.285000 ;
        RECT  9.415000 196.490000  9.615000 196.690000 ;
        RECT  9.415000 196.895000  9.615000 197.095000 ;
        RECT  9.415000 197.300000  9.615000 197.500000 ;
        RECT  9.415000 197.705000  9.615000 197.905000 ;
        RECT  9.530000  23.910000  9.730000  24.110000 ;
        RECT  9.530000  24.340000  9.730000  24.540000 ;
        RECT  9.530000  24.770000  9.730000  24.970000 ;
        RECT  9.530000  25.200000  9.730000  25.400000 ;
        RECT  9.530000  25.630000  9.730000  25.830000 ;
        RECT  9.530000  26.060000  9.730000  26.260000 ;
        RECT  9.530000  26.490000  9.730000  26.690000 ;
        RECT  9.530000  26.920000  9.730000  27.120000 ;
        RECT  9.530000  27.350000  9.730000  27.550000 ;
        RECT  9.530000  27.780000  9.730000  27.980000 ;
        RECT  9.530000  28.210000  9.730000  28.410000 ;
        RECT  9.815000 173.900000 10.015000 174.100000 ;
        RECT  9.815000 174.300000 10.015000 174.500000 ;
        RECT  9.815000 174.700000 10.015000 174.900000 ;
        RECT  9.815000 175.100000 10.015000 175.300000 ;
        RECT  9.815000 175.500000 10.015000 175.700000 ;
        RECT  9.815000 175.900000 10.015000 176.100000 ;
        RECT  9.815000 176.300000 10.015000 176.500000 ;
        RECT  9.815000 176.700000 10.015000 176.900000 ;
        RECT  9.815000 177.100000 10.015000 177.300000 ;
        RECT  9.815000 177.500000 10.015000 177.700000 ;
        RECT  9.815000 177.900000 10.015000 178.100000 ;
        RECT  9.815000 178.300000 10.015000 178.500000 ;
        RECT  9.815000 178.700000 10.015000 178.900000 ;
        RECT  9.815000 179.100000 10.015000 179.300000 ;
        RECT  9.815000 179.500000 10.015000 179.700000 ;
        RECT  9.815000 179.900000 10.015000 180.100000 ;
        RECT  9.815000 180.300000 10.015000 180.500000 ;
        RECT  9.815000 180.700000 10.015000 180.900000 ;
        RECT  9.815000 181.100000 10.015000 181.300000 ;
        RECT  9.815000 181.505000 10.015000 181.705000 ;
        RECT  9.815000 181.910000 10.015000 182.110000 ;
        RECT  9.815000 182.315000 10.015000 182.515000 ;
        RECT  9.815000 182.720000 10.015000 182.920000 ;
        RECT  9.815000 183.125000 10.015000 183.325000 ;
        RECT  9.815000 183.530000 10.015000 183.730000 ;
        RECT  9.815000 183.935000 10.015000 184.135000 ;
        RECT  9.815000 184.340000 10.015000 184.540000 ;
        RECT  9.815000 184.745000 10.015000 184.945000 ;
        RECT  9.815000 185.150000 10.015000 185.350000 ;
        RECT  9.815000 185.555000 10.015000 185.755000 ;
        RECT  9.815000 185.960000 10.015000 186.160000 ;
        RECT  9.815000 186.365000 10.015000 186.565000 ;
        RECT  9.815000 186.770000 10.015000 186.970000 ;
        RECT  9.815000 187.175000 10.015000 187.375000 ;
        RECT  9.815000 187.580000 10.015000 187.780000 ;
        RECT  9.815000 187.985000 10.015000 188.185000 ;
        RECT  9.815000 188.390000 10.015000 188.590000 ;
        RECT  9.815000 188.795000 10.015000 188.995000 ;
        RECT  9.815000 189.200000 10.015000 189.400000 ;
        RECT  9.815000 189.605000 10.015000 189.805000 ;
        RECT  9.815000 190.010000 10.015000 190.210000 ;
        RECT  9.815000 190.415000 10.015000 190.615000 ;
        RECT  9.815000 190.820000 10.015000 191.020000 ;
        RECT  9.815000 191.225000 10.015000 191.425000 ;
        RECT  9.815000 191.630000 10.015000 191.830000 ;
        RECT  9.815000 192.035000 10.015000 192.235000 ;
        RECT  9.815000 192.440000 10.015000 192.640000 ;
        RECT  9.815000 192.845000 10.015000 193.045000 ;
        RECT  9.815000 193.250000 10.015000 193.450000 ;
        RECT  9.815000 193.655000 10.015000 193.855000 ;
        RECT  9.815000 194.060000 10.015000 194.260000 ;
        RECT  9.815000 194.465000 10.015000 194.665000 ;
        RECT  9.815000 194.870000 10.015000 195.070000 ;
        RECT  9.815000 195.275000 10.015000 195.475000 ;
        RECT  9.815000 195.680000 10.015000 195.880000 ;
        RECT  9.815000 196.085000 10.015000 196.285000 ;
        RECT  9.815000 196.490000 10.015000 196.690000 ;
        RECT  9.815000 196.895000 10.015000 197.095000 ;
        RECT  9.815000 197.300000 10.015000 197.500000 ;
        RECT  9.815000 197.705000 10.015000 197.905000 ;
        RECT  9.935000  23.910000 10.135000  24.110000 ;
        RECT  9.935000  24.340000 10.135000  24.540000 ;
        RECT  9.935000  24.770000 10.135000  24.970000 ;
        RECT  9.935000  25.200000 10.135000  25.400000 ;
        RECT  9.935000  25.630000 10.135000  25.830000 ;
        RECT  9.935000  26.060000 10.135000  26.260000 ;
        RECT  9.935000  26.490000 10.135000  26.690000 ;
        RECT  9.935000  26.920000 10.135000  27.120000 ;
        RECT  9.935000  27.350000 10.135000  27.550000 ;
        RECT  9.935000  27.780000 10.135000  27.980000 ;
        RECT  9.935000  28.210000 10.135000  28.410000 ;
        RECT 10.215000 173.900000 10.415000 174.100000 ;
        RECT 10.215000 174.300000 10.415000 174.500000 ;
        RECT 10.215000 174.700000 10.415000 174.900000 ;
        RECT 10.215000 175.100000 10.415000 175.300000 ;
        RECT 10.215000 175.500000 10.415000 175.700000 ;
        RECT 10.215000 175.900000 10.415000 176.100000 ;
        RECT 10.215000 176.300000 10.415000 176.500000 ;
        RECT 10.215000 176.700000 10.415000 176.900000 ;
        RECT 10.215000 177.100000 10.415000 177.300000 ;
        RECT 10.215000 177.500000 10.415000 177.700000 ;
        RECT 10.215000 177.900000 10.415000 178.100000 ;
        RECT 10.215000 178.300000 10.415000 178.500000 ;
        RECT 10.215000 178.700000 10.415000 178.900000 ;
        RECT 10.215000 179.100000 10.415000 179.300000 ;
        RECT 10.215000 179.500000 10.415000 179.700000 ;
        RECT 10.215000 179.900000 10.415000 180.100000 ;
        RECT 10.215000 180.300000 10.415000 180.500000 ;
        RECT 10.215000 180.700000 10.415000 180.900000 ;
        RECT 10.215000 181.100000 10.415000 181.300000 ;
        RECT 10.215000 181.505000 10.415000 181.705000 ;
        RECT 10.215000 181.910000 10.415000 182.110000 ;
        RECT 10.215000 182.315000 10.415000 182.515000 ;
        RECT 10.215000 182.720000 10.415000 182.920000 ;
        RECT 10.215000 183.125000 10.415000 183.325000 ;
        RECT 10.215000 183.530000 10.415000 183.730000 ;
        RECT 10.215000 183.935000 10.415000 184.135000 ;
        RECT 10.215000 184.340000 10.415000 184.540000 ;
        RECT 10.215000 184.745000 10.415000 184.945000 ;
        RECT 10.215000 185.150000 10.415000 185.350000 ;
        RECT 10.215000 185.555000 10.415000 185.755000 ;
        RECT 10.215000 185.960000 10.415000 186.160000 ;
        RECT 10.215000 186.365000 10.415000 186.565000 ;
        RECT 10.215000 186.770000 10.415000 186.970000 ;
        RECT 10.215000 187.175000 10.415000 187.375000 ;
        RECT 10.215000 187.580000 10.415000 187.780000 ;
        RECT 10.215000 187.985000 10.415000 188.185000 ;
        RECT 10.215000 188.390000 10.415000 188.590000 ;
        RECT 10.215000 188.795000 10.415000 188.995000 ;
        RECT 10.215000 189.200000 10.415000 189.400000 ;
        RECT 10.215000 189.605000 10.415000 189.805000 ;
        RECT 10.215000 190.010000 10.415000 190.210000 ;
        RECT 10.215000 190.415000 10.415000 190.615000 ;
        RECT 10.215000 190.820000 10.415000 191.020000 ;
        RECT 10.215000 191.225000 10.415000 191.425000 ;
        RECT 10.215000 191.630000 10.415000 191.830000 ;
        RECT 10.215000 192.035000 10.415000 192.235000 ;
        RECT 10.215000 192.440000 10.415000 192.640000 ;
        RECT 10.215000 192.845000 10.415000 193.045000 ;
        RECT 10.215000 193.250000 10.415000 193.450000 ;
        RECT 10.215000 193.655000 10.415000 193.855000 ;
        RECT 10.215000 194.060000 10.415000 194.260000 ;
        RECT 10.215000 194.465000 10.415000 194.665000 ;
        RECT 10.215000 194.870000 10.415000 195.070000 ;
        RECT 10.215000 195.275000 10.415000 195.475000 ;
        RECT 10.215000 195.680000 10.415000 195.880000 ;
        RECT 10.215000 196.085000 10.415000 196.285000 ;
        RECT 10.215000 196.490000 10.415000 196.690000 ;
        RECT 10.215000 196.895000 10.415000 197.095000 ;
        RECT 10.215000 197.300000 10.415000 197.500000 ;
        RECT 10.215000 197.705000 10.415000 197.905000 ;
        RECT 10.340000  23.910000 10.540000  24.110000 ;
        RECT 10.340000  24.340000 10.540000  24.540000 ;
        RECT 10.340000  24.770000 10.540000  24.970000 ;
        RECT 10.340000  25.200000 10.540000  25.400000 ;
        RECT 10.340000  25.630000 10.540000  25.830000 ;
        RECT 10.340000  26.060000 10.540000  26.260000 ;
        RECT 10.340000  26.490000 10.540000  26.690000 ;
        RECT 10.340000  26.920000 10.540000  27.120000 ;
        RECT 10.340000  27.350000 10.540000  27.550000 ;
        RECT 10.340000  27.780000 10.540000  27.980000 ;
        RECT 10.340000  28.210000 10.540000  28.410000 ;
        RECT 10.615000 173.900000 10.815000 174.100000 ;
        RECT 10.615000 174.300000 10.815000 174.500000 ;
        RECT 10.615000 174.700000 10.815000 174.900000 ;
        RECT 10.615000 175.100000 10.815000 175.300000 ;
        RECT 10.615000 175.500000 10.815000 175.700000 ;
        RECT 10.615000 175.900000 10.815000 176.100000 ;
        RECT 10.615000 176.300000 10.815000 176.500000 ;
        RECT 10.615000 176.700000 10.815000 176.900000 ;
        RECT 10.615000 177.100000 10.815000 177.300000 ;
        RECT 10.615000 177.500000 10.815000 177.700000 ;
        RECT 10.615000 177.900000 10.815000 178.100000 ;
        RECT 10.615000 178.300000 10.815000 178.500000 ;
        RECT 10.615000 178.700000 10.815000 178.900000 ;
        RECT 10.615000 179.100000 10.815000 179.300000 ;
        RECT 10.615000 179.500000 10.815000 179.700000 ;
        RECT 10.615000 179.900000 10.815000 180.100000 ;
        RECT 10.615000 180.300000 10.815000 180.500000 ;
        RECT 10.615000 180.700000 10.815000 180.900000 ;
        RECT 10.615000 181.100000 10.815000 181.300000 ;
        RECT 10.615000 181.505000 10.815000 181.705000 ;
        RECT 10.615000 181.910000 10.815000 182.110000 ;
        RECT 10.615000 182.315000 10.815000 182.515000 ;
        RECT 10.615000 182.720000 10.815000 182.920000 ;
        RECT 10.615000 183.125000 10.815000 183.325000 ;
        RECT 10.615000 183.530000 10.815000 183.730000 ;
        RECT 10.615000 183.935000 10.815000 184.135000 ;
        RECT 10.615000 184.340000 10.815000 184.540000 ;
        RECT 10.615000 184.745000 10.815000 184.945000 ;
        RECT 10.615000 185.150000 10.815000 185.350000 ;
        RECT 10.615000 185.555000 10.815000 185.755000 ;
        RECT 10.615000 185.960000 10.815000 186.160000 ;
        RECT 10.615000 186.365000 10.815000 186.565000 ;
        RECT 10.615000 186.770000 10.815000 186.970000 ;
        RECT 10.615000 187.175000 10.815000 187.375000 ;
        RECT 10.615000 187.580000 10.815000 187.780000 ;
        RECT 10.615000 187.985000 10.815000 188.185000 ;
        RECT 10.615000 188.390000 10.815000 188.590000 ;
        RECT 10.615000 188.795000 10.815000 188.995000 ;
        RECT 10.615000 189.200000 10.815000 189.400000 ;
        RECT 10.615000 189.605000 10.815000 189.805000 ;
        RECT 10.615000 190.010000 10.815000 190.210000 ;
        RECT 10.615000 190.415000 10.815000 190.615000 ;
        RECT 10.615000 190.820000 10.815000 191.020000 ;
        RECT 10.615000 191.225000 10.815000 191.425000 ;
        RECT 10.615000 191.630000 10.815000 191.830000 ;
        RECT 10.615000 192.035000 10.815000 192.235000 ;
        RECT 10.615000 192.440000 10.815000 192.640000 ;
        RECT 10.615000 192.845000 10.815000 193.045000 ;
        RECT 10.615000 193.250000 10.815000 193.450000 ;
        RECT 10.615000 193.655000 10.815000 193.855000 ;
        RECT 10.615000 194.060000 10.815000 194.260000 ;
        RECT 10.615000 194.465000 10.815000 194.665000 ;
        RECT 10.615000 194.870000 10.815000 195.070000 ;
        RECT 10.615000 195.275000 10.815000 195.475000 ;
        RECT 10.615000 195.680000 10.815000 195.880000 ;
        RECT 10.615000 196.085000 10.815000 196.285000 ;
        RECT 10.615000 196.490000 10.815000 196.690000 ;
        RECT 10.615000 196.895000 10.815000 197.095000 ;
        RECT 10.615000 197.300000 10.815000 197.500000 ;
        RECT 10.615000 197.705000 10.815000 197.905000 ;
        RECT 10.745000  23.910000 10.945000  24.110000 ;
        RECT 10.745000  24.340000 10.945000  24.540000 ;
        RECT 10.745000  24.770000 10.945000  24.970000 ;
        RECT 10.745000  25.200000 10.945000  25.400000 ;
        RECT 10.745000  25.630000 10.945000  25.830000 ;
        RECT 10.745000  26.060000 10.945000  26.260000 ;
        RECT 10.745000  26.490000 10.945000  26.690000 ;
        RECT 10.745000  26.920000 10.945000  27.120000 ;
        RECT 10.745000  27.350000 10.945000  27.550000 ;
        RECT 10.745000  27.780000 10.945000  27.980000 ;
        RECT 10.745000  28.210000 10.945000  28.410000 ;
        RECT 11.015000 173.900000 11.215000 174.100000 ;
        RECT 11.015000 174.300000 11.215000 174.500000 ;
        RECT 11.015000 174.700000 11.215000 174.900000 ;
        RECT 11.015000 175.100000 11.215000 175.300000 ;
        RECT 11.015000 175.500000 11.215000 175.700000 ;
        RECT 11.015000 175.900000 11.215000 176.100000 ;
        RECT 11.015000 176.300000 11.215000 176.500000 ;
        RECT 11.015000 176.700000 11.215000 176.900000 ;
        RECT 11.015000 177.100000 11.215000 177.300000 ;
        RECT 11.015000 177.500000 11.215000 177.700000 ;
        RECT 11.015000 177.900000 11.215000 178.100000 ;
        RECT 11.015000 178.300000 11.215000 178.500000 ;
        RECT 11.015000 178.700000 11.215000 178.900000 ;
        RECT 11.015000 179.100000 11.215000 179.300000 ;
        RECT 11.015000 179.500000 11.215000 179.700000 ;
        RECT 11.015000 179.900000 11.215000 180.100000 ;
        RECT 11.015000 180.300000 11.215000 180.500000 ;
        RECT 11.015000 180.700000 11.215000 180.900000 ;
        RECT 11.015000 181.100000 11.215000 181.300000 ;
        RECT 11.015000 181.505000 11.215000 181.705000 ;
        RECT 11.015000 181.910000 11.215000 182.110000 ;
        RECT 11.015000 182.315000 11.215000 182.515000 ;
        RECT 11.015000 182.720000 11.215000 182.920000 ;
        RECT 11.015000 183.125000 11.215000 183.325000 ;
        RECT 11.015000 183.530000 11.215000 183.730000 ;
        RECT 11.015000 183.935000 11.215000 184.135000 ;
        RECT 11.015000 184.340000 11.215000 184.540000 ;
        RECT 11.015000 184.745000 11.215000 184.945000 ;
        RECT 11.015000 185.150000 11.215000 185.350000 ;
        RECT 11.015000 185.555000 11.215000 185.755000 ;
        RECT 11.015000 185.960000 11.215000 186.160000 ;
        RECT 11.015000 186.365000 11.215000 186.565000 ;
        RECT 11.015000 186.770000 11.215000 186.970000 ;
        RECT 11.015000 187.175000 11.215000 187.375000 ;
        RECT 11.015000 187.580000 11.215000 187.780000 ;
        RECT 11.015000 187.985000 11.215000 188.185000 ;
        RECT 11.015000 188.390000 11.215000 188.590000 ;
        RECT 11.015000 188.795000 11.215000 188.995000 ;
        RECT 11.015000 189.200000 11.215000 189.400000 ;
        RECT 11.015000 189.605000 11.215000 189.805000 ;
        RECT 11.015000 190.010000 11.215000 190.210000 ;
        RECT 11.015000 190.415000 11.215000 190.615000 ;
        RECT 11.015000 190.820000 11.215000 191.020000 ;
        RECT 11.015000 191.225000 11.215000 191.425000 ;
        RECT 11.015000 191.630000 11.215000 191.830000 ;
        RECT 11.015000 192.035000 11.215000 192.235000 ;
        RECT 11.015000 192.440000 11.215000 192.640000 ;
        RECT 11.015000 192.845000 11.215000 193.045000 ;
        RECT 11.015000 193.250000 11.215000 193.450000 ;
        RECT 11.015000 193.655000 11.215000 193.855000 ;
        RECT 11.015000 194.060000 11.215000 194.260000 ;
        RECT 11.015000 194.465000 11.215000 194.665000 ;
        RECT 11.015000 194.870000 11.215000 195.070000 ;
        RECT 11.015000 195.275000 11.215000 195.475000 ;
        RECT 11.015000 195.680000 11.215000 195.880000 ;
        RECT 11.015000 196.085000 11.215000 196.285000 ;
        RECT 11.015000 196.490000 11.215000 196.690000 ;
        RECT 11.015000 196.895000 11.215000 197.095000 ;
        RECT 11.015000 197.300000 11.215000 197.500000 ;
        RECT 11.015000 197.705000 11.215000 197.905000 ;
        RECT 11.150000  23.910000 11.350000  24.110000 ;
        RECT 11.150000  24.340000 11.350000  24.540000 ;
        RECT 11.150000  24.770000 11.350000  24.970000 ;
        RECT 11.150000  25.200000 11.350000  25.400000 ;
        RECT 11.150000  25.630000 11.350000  25.830000 ;
        RECT 11.150000  26.060000 11.350000  26.260000 ;
        RECT 11.150000  26.490000 11.350000  26.690000 ;
        RECT 11.150000  26.920000 11.350000  27.120000 ;
        RECT 11.150000  27.350000 11.350000  27.550000 ;
        RECT 11.150000  27.780000 11.350000  27.980000 ;
        RECT 11.150000  28.210000 11.350000  28.410000 ;
        RECT 11.415000 173.900000 11.615000 174.100000 ;
        RECT 11.415000 174.300000 11.615000 174.500000 ;
        RECT 11.415000 174.700000 11.615000 174.900000 ;
        RECT 11.415000 175.100000 11.615000 175.300000 ;
        RECT 11.415000 175.500000 11.615000 175.700000 ;
        RECT 11.415000 175.900000 11.615000 176.100000 ;
        RECT 11.415000 176.300000 11.615000 176.500000 ;
        RECT 11.415000 176.700000 11.615000 176.900000 ;
        RECT 11.415000 177.100000 11.615000 177.300000 ;
        RECT 11.415000 177.500000 11.615000 177.700000 ;
        RECT 11.415000 177.900000 11.615000 178.100000 ;
        RECT 11.415000 178.300000 11.615000 178.500000 ;
        RECT 11.415000 178.700000 11.615000 178.900000 ;
        RECT 11.415000 179.100000 11.615000 179.300000 ;
        RECT 11.415000 179.500000 11.615000 179.700000 ;
        RECT 11.415000 179.900000 11.615000 180.100000 ;
        RECT 11.415000 180.300000 11.615000 180.500000 ;
        RECT 11.415000 180.700000 11.615000 180.900000 ;
        RECT 11.415000 181.100000 11.615000 181.300000 ;
        RECT 11.415000 181.505000 11.615000 181.705000 ;
        RECT 11.415000 181.910000 11.615000 182.110000 ;
        RECT 11.415000 182.315000 11.615000 182.515000 ;
        RECT 11.415000 182.720000 11.615000 182.920000 ;
        RECT 11.415000 183.125000 11.615000 183.325000 ;
        RECT 11.415000 183.530000 11.615000 183.730000 ;
        RECT 11.415000 183.935000 11.615000 184.135000 ;
        RECT 11.415000 184.340000 11.615000 184.540000 ;
        RECT 11.415000 184.745000 11.615000 184.945000 ;
        RECT 11.415000 185.150000 11.615000 185.350000 ;
        RECT 11.415000 185.555000 11.615000 185.755000 ;
        RECT 11.415000 185.960000 11.615000 186.160000 ;
        RECT 11.415000 186.365000 11.615000 186.565000 ;
        RECT 11.415000 186.770000 11.615000 186.970000 ;
        RECT 11.415000 187.175000 11.615000 187.375000 ;
        RECT 11.415000 187.580000 11.615000 187.780000 ;
        RECT 11.415000 187.985000 11.615000 188.185000 ;
        RECT 11.415000 188.390000 11.615000 188.590000 ;
        RECT 11.415000 188.795000 11.615000 188.995000 ;
        RECT 11.415000 189.200000 11.615000 189.400000 ;
        RECT 11.415000 189.605000 11.615000 189.805000 ;
        RECT 11.415000 190.010000 11.615000 190.210000 ;
        RECT 11.415000 190.415000 11.615000 190.615000 ;
        RECT 11.415000 190.820000 11.615000 191.020000 ;
        RECT 11.415000 191.225000 11.615000 191.425000 ;
        RECT 11.415000 191.630000 11.615000 191.830000 ;
        RECT 11.415000 192.035000 11.615000 192.235000 ;
        RECT 11.415000 192.440000 11.615000 192.640000 ;
        RECT 11.415000 192.845000 11.615000 193.045000 ;
        RECT 11.415000 193.250000 11.615000 193.450000 ;
        RECT 11.415000 193.655000 11.615000 193.855000 ;
        RECT 11.415000 194.060000 11.615000 194.260000 ;
        RECT 11.415000 194.465000 11.615000 194.665000 ;
        RECT 11.415000 194.870000 11.615000 195.070000 ;
        RECT 11.415000 195.275000 11.615000 195.475000 ;
        RECT 11.415000 195.680000 11.615000 195.880000 ;
        RECT 11.415000 196.085000 11.615000 196.285000 ;
        RECT 11.415000 196.490000 11.615000 196.690000 ;
        RECT 11.415000 196.895000 11.615000 197.095000 ;
        RECT 11.415000 197.300000 11.615000 197.500000 ;
        RECT 11.415000 197.705000 11.615000 197.905000 ;
        RECT 11.555000  23.910000 11.755000  24.110000 ;
        RECT 11.555000  24.340000 11.755000  24.540000 ;
        RECT 11.555000  24.770000 11.755000  24.970000 ;
        RECT 11.555000  25.200000 11.755000  25.400000 ;
        RECT 11.555000  25.630000 11.755000  25.830000 ;
        RECT 11.555000  26.060000 11.755000  26.260000 ;
        RECT 11.555000  26.490000 11.755000  26.690000 ;
        RECT 11.555000  26.920000 11.755000  27.120000 ;
        RECT 11.555000  27.350000 11.755000  27.550000 ;
        RECT 11.555000  27.780000 11.755000  27.980000 ;
        RECT 11.555000  28.210000 11.755000  28.410000 ;
        RECT 11.815000 173.900000 12.015000 174.100000 ;
        RECT 11.815000 174.300000 12.015000 174.500000 ;
        RECT 11.815000 174.700000 12.015000 174.900000 ;
        RECT 11.815000 175.100000 12.015000 175.300000 ;
        RECT 11.815000 175.500000 12.015000 175.700000 ;
        RECT 11.815000 175.900000 12.015000 176.100000 ;
        RECT 11.815000 176.300000 12.015000 176.500000 ;
        RECT 11.815000 176.700000 12.015000 176.900000 ;
        RECT 11.815000 177.100000 12.015000 177.300000 ;
        RECT 11.815000 177.500000 12.015000 177.700000 ;
        RECT 11.815000 177.900000 12.015000 178.100000 ;
        RECT 11.815000 178.300000 12.015000 178.500000 ;
        RECT 11.815000 178.700000 12.015000 178.900000 ;
        RECT 11.815000 179.100000 12.015000 179.300000 ;
        RECT 11.815000 179.500000 12.015000 179.700000 ;
        RECT 11.815000 179.900000 12.015000 180.100000 ;
        RECT 11.815000 180.300000 12.015000 180.500000 ;
        RECT 11.815000 180.700000 12.015000 180.900000 ;
        RECT 11.815000 181.100000 12.015000 181.300000 ;
        RECT 11.815000 181.505000 12.015000 181.705000 ;
        RECT 11.815000 181.910000 12.015000 182.110000 ;
        RECT 11.815000 182.315000 12.015000 182.515000 ;
        RECT 11.815000 182.720000 12.015000 182.920000 ;
        RECT 11.815000 183.125000 12.015000 183.325000 ;
        RECT 11.815000 183.530000 12.015000 183.730000 ;
        RECT 11.815000 183.935000 12.015000 184.135000 ;
        RECT 11.815000 184.340000 12.015000 184.540000 ;
        RECT 11.815000 184.745000 12.015000 184.945000 ;
        RECT 11.815000 185.150000 12.015000 185.350000 ;
        RECT 11.815000 185.555000 12.015000 185.755000 ;
        RECT 11.815000 185.960000 12.015000 186.160000 ;
        RECT 11.815000 186.365000 12.015000 186.565000 ;
        RECT 11.815000 186.770000 12.015000 186.970000 ;
        RECT 11.815000 187.175000 12.015000 187.375000 ;
        RECT 11.815000 187.580000 12.015000 187.780000 ;
        RECT 11.815000 187.985000 12.015000 188.185000 ;
        RECT 11.815000 188.390000 12.015000 188.590000 ;
        RECT 11.815000 188.795000 12.015000 188.995000 ;
        RECT 11.815000 189.200000 12.015000 189.400000 ;
        RECT 11.815000 189.605000 12.015000 189.805000 ;
        RECT 11.815000 190.010000 12.015000 190.210000 ;
        RECT 11.815000 190.415000 12.015000 190.615000 ;
        RECT 11.815000 190.820000 12.015000 191.020000 ;
        RECT 11.815000 191.225000 12.015000 191.425000 ;
        RECT 11.815000 191.630000 12.015000 191.830000 ;
        RECT 11.815000 192.035000 12.015000 192.235000 ;
        RECT 11.815000 192.440000 12.015000 192.640000 ;
        RECT 11.815000 192.845000 12.015000 193.045000 ;
        RECT 11.815000 193.250000 12.015000 193.450000 ;
        RECT 11.815000 193.655000 12.015000 193.855000 ;
        RECT 11.815000 194.060000 12.015000 194.260000 ;
        RECT 11.815000 194.465000 12.015000 194.665000 ;
        RECT 11.815000 194.870000 12.015000 195.070000 ;
        RECT 11.815000 195.275000 12.015000 195.475000 ;
        RECT 11.815000 195.680000 12.015000 195.880000 ;
        RECT 11.815000 196.085000 12.015000 196.285000 ;
        RECT 11.815000 196.490000 12.015000 196.690000 ;
        RECT 11.815000 196.895000 12.015000 197.095000 ;
        RECT 11.815000 197.300000 12.015000 197.500000 ;
        RECT 11.815000 197.705000 12.015000 197.905000 ;
        RECT 11.960000  23.910000 12.160000  24.110000 ;
        RECT 11.960000  24.340000 12.160000  24.540000 ;
        RECT 11.960000  24.770000 12.160000  24.970000 ;
        RECT 11.960000  25.200000 12.160000  25.400000 ;
        RECT 11.960000  25.630000 12.160000  25.830000 ;
        RECT 11.960000  26.060000 12.160000  26.260000 ;
        RECT 11.960000  26.490000 12.160000  26.690000 ;
        RECT 11.960000  26.920000 12.160000  27.120000 ;
        RECT 11.960000  27.350000 12.160000  27.550000 ;
        RECT 11.960000  27.780000 12.160000  27.980000 ;
        RECT 11.960000  28.210000 12.160000  28.410000 ;
        RECT 12.215000 173.900000 12.415000 174.100000 ;
        RECT 12.215000 174.300000 12.415000 174.500000 ;
        RECT 12.215000 174.700000 12.415000 174.900000 ;
        RECT 12.215000 175.100000 12.415000 175.300000 ;
        RECT 12.215000 175.500000 12.415000 175.700000 ;
        RECT 12.215000 175.900000 12.415000 176.100000 ;
        RECT 12.215000 176.300000 12.415000 176.500000 ;
        RECT 12.215000 176.700000 12.415000 176.900000 ;
        RECT 12.215000 177.100000 12.415000 177.300000 ;
        RECT 12.215000 177.500000 12.415000 177.700000 ;
        RECT 12.215000 177.900000 12.415000 178.100000 ;
        RECT 12.215000 178.300000 12.415000 178.500000 ;
        RECT 12.215000 178.700000 12.415000 178.900000 ;
        RECT 12.215000 179.100000 12.415000 179.300000 ;
        RECT 12.215000 179.500000 12.415000 179.700000 ;
        RECT 12.215000 179.900000 12.415000 180.100000 ;
        RECT 12.215000 180.300000 12.415000 180.500000 ;
        RECT 12.215000 180.700000 12.415000 180.900000 ;
        RECT 12.215000 181.100000 12.415000 181.300000 ;
        RECT 12.215000 181.505000 12.415000 181.705000 ;
        RECT 12.215000 181.910000 12.415000 182.110000 ;
        RECT 12.215000 182.315000 12.415000 182.515000 ;
        RECT 12.215000 182.720000 12.415000 182.920000 ;
        RECT 12.215000 183.125000 12.415000 183.325000 ;
        RECT 12.215000 183.530000 12.415000 183.730000 ;
        RECT 12.215000 183.935000 12.415000 184.135000 ;
        RECT 12.215000 184.340000 12.415000 184.540000 ;
        RECT 12.215000 184.745000 12.415000 184.945000 ;
        RECT 12.215000 185.150000 12.415000 185.350000 ;
        RECT 12.215000 185.555000 12.415000 185.755000 ;
        RECT 12.215000 185.960000 12.415000 186.160000 ;
        RECT 12.215000 186.365000 12.415000 186.565000 ;
        RECT 12.215000 186.770000 12.415000 186.970000 ;
        RECT 12.215000 187.175000 12.415000 187.375000 ;
        RECT 12.215000 187.580000 12.415000 187.780000 ;
        RECT 12.215000 187.985000 12.415000 188.185000 ;
        RECT 12.215000 188.390000 12.415000 188.590000 ;
        RECT 12.215000 188.795000 12.415000 188.995000 ;
        RECT 12.215000 189.200000 12.415000 189.400000 ;
        RECT 12.215000 189.605000 12.415000 189.805000 ;
        RECT 12.215000 190.010000 12.415000 190.210000 ;
        RECT 12.215000 190.415000 12.415000 190.615000 ;
        RECT 12.215000 190.820000 12.415000 191.020000 ;
        RECT 12.215000 191.225000 12.415000 191.425000 ;
        RECT 12.215000 191.630000 12.415000 191.830000 ;
        RECT 12.215000 192.035000 12.415000 192.235000 ;
        RECT 12.215000 192.440000 12.415000 192.640000 ;
        RECT 12.215000 192.845000 12.415000 193.045000 ;
        RECT 12.215000 193.250000 12.415000 193.450000 ;
        RECT 12.215000 193.655000 12.415000 193.855000 ;
        RECT 12.215000 194.060000 12.415000 194.260000 ;
        RECT 12.215000 194.465000 12.415000 194.665000 ;
        RECT 12.215000 194.870000 12.415000 195.070000 ;
        RECT 12.215000 195.275000 12.415000 195.475000 ;
        RECT 12.215000 195.680000 12.415000 195.880000 ;
        RECT 12.215000 196.085000 12.415000 196.285000 ;
        RECT 12.215000 196.490000 12.415000 196.690000 ;
        RECT 12.215000 196.895000 12.415000 197.095000 ;
        RECT 12.215000 197.300000 12.415000 197.500000 ;
        RECT 12.215000 197.705000 12.415000 197.905000 ;
        RECT 12.365000  23.910000 12.565000  24.110000 ;
        RECT 12.365000  24.340000 12.565000  24.540000 ;
        RECT 12.365000  24.770000 12.565000  24.970000 ;
        RECT 12.365000  25.200000 12.565000  25.400000 ;
        RECT 12.365000  25.630000 12.565000  25.830000 ;
        RECT 12.365000  26.060000 12.565000  26.260000 ;
        RECT 12.365000  26.490000 12.565000  26.690000 ;
        RECT 12.365000  26.920000 12.565000  27.120000 ;
        RECT 12.365000  27.350000 12.565000  27.550000 ;
        RECT 12.365000  27.780000 12.565000  27.980000 ;
        RECT 12.365000  28.210000 12.565000  28.410000 ;
        RECT 12.615000 173.900000 12.815000 174.100000 ;
        RECT 12.615000 174.300000 12.815000 174.500000 ;
        RECT 12.615000 174.700000 12.815000 174.900000 ;
        RECT 12.615000 175.100000 12.815000 175.300000 ;
        RECT 12.615000 175.500000 12.815000 175.700000 ;
        RECT 12.615000 175.900000 12.815000 176.100000 ;
        RECT 12.615000 176.300000 12.815000 176.500000 ;
        RECT 12.615000 176.700000 12.815000 176.900000 ;
        RECT 12.615000 177.100000 12.815000 177.300000 ;
        RECT 12.615000 177.500000 12.815000 177.700000 ;
        RECT 12.615000 177.900000 12.815000 178.100000 ;
        RECT 12.615000 178.300000 12.815000 178.500000 ;
        RECT 12.615000 178.700000 12.815000 178.900000 ;
        RECT 12.615000 179.100000 12.815000 179.300000 ;
        RECT 12.615000 179.500000 12.815000 179.700000 ;
        RECT 12.615000 179.900000 12.815000 180.100000 ;
        RECT 12.615000 180.300000 12.815000 180.500000 ;
        RECT 12.615000 180.700000 12.815000 180.900000 ;
        RECT 12.615000 181.100000 12.815000 181.300000 ;
        RECT 12.615000 181.505000 12.815000 181.705000 ;
        RECT 12.615000 181.910000 12.815000 182.110000 ;
        RECT 12.615000 182.315000 12.815000 182.515000 ;
        RECT 12.615000 182.720000 12.815000 182.920000 ;
        RECT 12.615000 183.125000 12.815000 183.325000 ;
        RECT 12.615000 183.530000 12.815000 183.730000 ;
        RECT 12.615000 183.935000 12.815000 184.135000 ;
        RECT 12.615000 184.340000 12.815000 184.540000 ;
        RECT 12.615000 184.745000 12.815000 184.945000 ;
        RECT 12.615000 185.150000 12.815000 185.350000 ;
        RECT 12.615000 185.555000 12.815000 185.755000 ;
        RECT 12.615000 185.960000 12.815000 186.160000 ;
        RECT 12.615000 186.365000 12.815000 186.565000 ;
        RECT 12.615000 186.770000 12.815000 186.970000 ;
        RECT 12.615000 187.175000 12.815000 187.375000 ;
        RECT 12.615000 187.580000 12.815000 187.780000 ;
        RECT 12.615000 187.985000 12.815000 188.185000 ;
        RECT 12.615000 188.390000 12.815000 188.590000 ;
        RECT 12.615000 188.795000 12.815000 188.995000 ;
        RECT 12.615000 189.200000 12.815000 189.400000 ;
        RECT 12.615000 189.605000 12.815000 189.805000 ;
        RECT 12.615000 190.010000 12.815000 190.210000 ;
        RECT 12.615000 190.415000 12.815000 190.615000 ;
        RECT 12.615000 190.820000 12.815000 191.020000 ;
        RECT 12.615000 191.225000 12.815000 191.425000 ;
        RECT 12.615000 191.630000 12.815000 191.830000 ;
        RECT 12.615000 192.035000 12.815000 192.235000 ;
        RECT 12.615000 192.440000 12.815000 192.640000 ;
        RECT 12.615000 192.845000 12.815000 193.045000 ;
        RECT 12.615000 193.250000 12.815000 193.450000 ;
        RECT 12.615000 193.655000 12.815000 193.855000 ;
        RECT 12.615000 194.060000 12.815000 194.260000 ;
        RECT 12.615000 194.465000 12.815000 194.665000 ;
        RECT 12.615000 194.870000 12.815000 195.070000 ;
        RECT 12.615000 195.275000 12.815000 195.475000 ;
        RECT 12.615000 195.680000 12.815000 195.880000 ;
        RECT 12.615000 196.085000 12.815000 196.285000 ;
        RECT 12.615000 196.490000 12.815000 196.690000 ;
        RECT 12.615000 196.895000 12.815000 197.095000 ;
        RECT 12.615000 197.300000 12.815000 197.500000 ;
        RECT 12.615000 197.705000 12.815000 197.905000 ;
        RECT 12.770000  23.910000 12.970000  24.110000 ;
        RECT 12.770000  24.340000 12.970000  24.540000 ;
        RECT 12.770000  24.770000 12.970000  24.970000 ;
        RECT 12.770000  25.200000 12.970000  25.400000 ;
        RECT 12.770000  25.630000 12.970000  25.830000 ;
        RECT 12.770000  26.060000 12.970000  26.260000 ;
        RECT 12.770000  26.490000 12.970000  26.690000 ;
        RECT 12.770000  26.920000 12.970000  27.120000 ;
        RECT 12.770000  27.350000 12.970000  27.550000 ;
        RECT 12.770000  27.780000 12.970000  27.980000 ;
        RECT 12.770000  28.210000 12.970000  28.410000 ;
        RECT 13.175000  23.910000 13.375000  24.110000 ;
        RECT 13.175000  24.340000 13.375000  24.540000 ;
        RECT 13.175000  24.770000 13.375000  24.970000 ;
        RECT 13.175000  25.200000 13.375000  25.400000 ;
        RECT 13.175000  25.630000 13.375000  25.830000 ;
        RECT 13.175000  26.060000 13.375000  26.260000 ;
        RECT 13.175000  26.490000 13.375000  26.690000 ;
        RECT 13.175000  26.920000 13.375000  27.120000 ;
        RECT 13.175000  27.350000 13.375000  27.550000 ;
        RECT 13.175000  27.780000 13.375000  27.980000 ;
        RECT 13.175000  28.210000 13.375000  28.410000 ;
        RECT 13.580000  23.910000 13.780000  24.110000 ;
        RECT 13.580000  24.340000 13.780000  24.540000 ;
        RECT 13.580000  24.770000 13.780000  24.970000 ;
        RECT 13.580000  25.200000 13.780000  25.400000 ;
        RECT 13.580000  25.630000 13.780000  25.830000 ;
        RECT 13.580000  26.060000 13.780000  26.260000 ;
        RECT 13.580000  26.490000 13.780000  26.690000 ;
        RECT 13.580000  26.920000 13.780000  27.120000 ;
        RECT 13.580000  27.350000 13.780000  27.550000 ;
        RECT 13.580000  27.780000 13.780000  27.980000 ;
        RECT 13.580000  28.210000 13.780000  28.410000 ;
        RECT 13.985000  23.910000 14.185000  24.110000 ;
        RECT 13.985000  24.340000 14.185000  24.540000 ;
        RECT 13.985000  24.770000 14.185000  24.970000 ;
        RECT 13.985000  25.200000 14.185000  25.400000 ;
        RECT 13.985000  25.630000 14.185000  25.830000 ;
        RECT 13.985000  26.060000 14.185000  26.260000 ;
        RECT 13.985000  26.490000 14.185000  26.690000 ;
        RECT 13.985000  26.920000 14.185000  27.120000 ;
        RECT 13.985000  27.350000 14.185000  27.550000 ;
        RECT 13.985000  27.780000 14.185000  27.980000 ;
        RECT 13.985000  28.210000 14.185000  28.410000 ;
        RECT 14.390000  23.910000 14.590000  24.110000 ;
        RECT 14.390000  24.340000 14.590000  24.540000 ;
        RECT 14.390000  24.770000 14.590000  24.970000 ;
        RECT 14.390000  25.200000 14.590000  25.400000 ;
        RECT 14.390000  25.630000 14.590000  25.830000 ;
        RECT 14.390000  26.060000 14.590000  26.260000 ;
        RECT 14.390000  26.490000 14.590000  26.690000 ;
        RECT 14.390000  26.920000 14.590000  27.120000 ;
        RECT 14.390000  27.350000 14.590000  27.550000 ;
        RECT 14.390000  27.780000 14.590000  27.980000 ;
        RECT 14.390000  28.210000 14.590000  28.410000 ;
        RECT 14.795000  23.910000 14.995000  24.110000 ;
        RECT 14.795000  24.340000 14.995000  24.540000 ;
        RECT 14.795000  24.770000 14.995000  24.970000 ;
        RECT 14.795000  25.200000 14.995000  25.400000 ;
        RECT 14.795000  25.630000 14.995000  25.830000 ;
        RECT 14.795000  26.060000 14.995000  26.260000 ;
        RECT 14.795000  26.490000 14.995000  26.690000 ;
        RECT 14.795000  26.920000 14.995000  27.120000 ;
        RECT 14.795000  27.350000 14.995000  27.550000 ;
        RECT 14.795000  27.780000 14.995000  27.980000 ;
        RECT 14.795000  28.210000 14.995000  28.410000 ;
        RECT 15.200000  23.910000 15.400000  24.110000 ;
        RECT 15.200000  24.340000 15.400000  24.540000 ;
        RECT 15.200000  24.770000 15.400000  24.970000 ;
        RECT 15.200000  25.200000 15.400000  25.400000 ;
        RECT 15.200000  25.630000 15.400000  25.830000 ;
        RECT 15.200000  26.060000 15.400000  26.260000 ;
        RECT 15.200000  26.490000 15.400000  26.690000 ;
        RECT 15.200000  26.920000 15.400000  27.120000 ;
        RECT 15.200000  27.350000 15.400000  27.550000 ;
        RECT 15.200000  27.780000 15.400000  27.980000 ;
        RECT 15.200000  28.210000 15.400000  28.410000 ;
        RECT 15.605000  23.910000 15.805000  24.110000 ;
        RECT 15.605000  24.340000 15.805000  24.540000 ;
        RECT 15.605000  24.770000 15.805000  24.970000 ;
        RECT 15.605000  25.200000 15.805000  25.400000 ;
        RECT 15.605000  25.630000 15.805000  25.830000 ;
        RECT 15.605000  26.060000 15.805000  26.260000 ;
        RECT 15.605000  26.490000 15.805000  26.690000 ;
        RECT 15.605000  26.920000 15.805000  27.120000 ;
        RECT 15.605000  27.350000 15.805000  27.550000 ;
        RECT 15.605000  27.780000 15.805000  27.980000 ;
        RECT 15.605000  28.210000 15.805000  28.410000 ;
        RECT 16.010000  23.910000 16.210000  24.110000 ;
        RECT 16.010000  24.340000 16.210000  24.540000 ;
        RECT 16.010000  24.770000 16.210000  24.970000 ;
        RECT 16.010000  25.200000 16.210000  25.400000 ;
        RECT 16.010000  25.630000 16.210000  25.830000 ;
        RECT 16.010000  26.060000 16.210000  26.260000 ;
        RECT 16.010000  26.490000 16.210000  26.690000 ;
        RECT 16.010000  26.920000 16.210000  27.120000 ;
        RECT 16.010000  27.350000 16.210000  27.550000 ;
        RECT 16.010000  27.780000 16.210000  27.980000 ;
        RECT 16.010000  28.210000 16.210000  28.410000 ;
        RECT 16.415000  23.910000 16.615000  24.110000 ;
        RECT 16.415000  24.340000 16.615000  24.540000 ;
        RECT 16.415000  24.770000 16.615000  24.970000 ;
        RECT 16.415000  25.200000 16.615000  25.400000 ;
        RECT 16.415000  25.630000 16.615000  25.830000 ;
        RECT 16.415000  26.060000 16.615000  26.260000 ;
        RECT 16.415000  26.490000 16.615000  26.690000 ;
        RECT 16.415000  26.920000 16.615000  27.120000 ;
        RECT 16.415000  27.350000 16.615000  27.550000 ;
        RECT 16.415000  27.780000 16.615000  27.980000 ;
        RECT 16.415000  28.210000 16.615000  28.410000 ;
        RECT 16.820000  23.910000 17.020000  24.110000 ;
        RECT 16.820000  24.340000 17.020000  24.540000 ;
        RECT 16.820000  24.770000 17.020000  24.970000 ;
        RECT 16.820000  25.200000 17.020000  25.400000 ;
        RECT 16.820000  25.630000 17.020000  25.830000 ;
        RECT 16.820000  26.060000 17.020000  26.260000 ;
        RECT 16.820000  26.490000 17.020000  26.690000 ;
        RECT 16.820000  26.920000 17.020000  27.120000 ;
        RECT 16.820000  27.350000 17.020000  27.550000 ;
        RECT 16.820000  27.780000 17.020000  27.980000 ;
        RECT 16.820000  28.210000 17.020000  28.410000 ;
        RECT 17.225000  23.910000 17.425000  24.110000 ;
        RECT 17.225000  24.340000 17.425000  24.540000 ;
        RECT 17.225000  24.770000 17.425000  24.970000 ;
        RECT 17.225000  25.200000 17.425000  25.400000 ;
        RECT 17.225000  25.630000 17.425000  25.830000 ;
        RECT 17.225000  26.060000 17.425000  26.260000 ;
        RECT 17.225000  26.490000 17.425000  26.690000 ;
        RECT 17.225000  26.920000 17.425000  27.120000 ;
        RECT 17.225000  27.350000 17.425000  27.550000 ;
        RECT 17.225000  27.780000 17.425000  27.980000 ;
        RECT 17.225000  28.210000 17.425000  28.410000 ;
        RECT 17.630000  23.910000 17.830000  24.110000 ;
        RECT 17.630000  24.340000 17.830000  24.540000 ;
        RECT 17.630000  24.770000 17.830000  24.970000 ;
        RECT 17.630000  25.200000 17.830000  25.400000 ;
        RECT 17.630000  25.630000 17.830000  25.830000 ;
        RECT 17.630000  26.060000 17.830000  26.260000 ;
        RECT 17.630000  26.490000 17.830000  26.690000 ;
        RECT 17.630000  26.920000 17.830000  27.120000 ;
        RECT 17.630000  27.350000 17.830000  27.550000 ;
        RECT 17.630000  27.780000 17.830000  27.980000 ;
        RECT 17.630000  28.210000 17.830000  28.410000 ;
        RECT 18.035000  23.910000 18.235000  24.110000 ;
        RECT 18.035000  24.340000 18.235000  24.540000 ;
        RECT 18.035000  24.770000 18.235000  24.970000 ;
        RECT 18.035000  25.200000 18.235000  25.400000 ;
        RECT 18.035000  25.630000 18.235000  25.830000 ;
        RECT 18.035000  26.060000 18.235000  26.260000 ;
        RECT 18.035000  26.490000 18.235000  26.690000 ;
        RECT 18.035000  26.920000 18.235000  27.120000 ;
        RECT 18.035000  27.350000 18.235000  27.550000 ;
        RECT 18.035000  27.780000 18.235000  27.980000 ;
        RECT 18.035000  28.210000 18.235000  28.410000 ;
        RECT 18.440000  23.910000 18.640000  24.110000 ;
        RECT 18.440000  24.340000 18.640000  24.540000 ;
        RECT 18.440000  24.770000 18.640000  24.970000 ;
        RECT 18.440000  25.200000 18.640000  25.400000 ;
        RECT 18.440000  25.630000 18.640000  25.830000 ;
        RECT 18.440000  26.060000 18.640000  26.260000 ;
        RECT 18.440000  26.490000 18.640000  26.690000 ;
        RECT 18.440000  26.920000 18.640000  27.120000 ;
        RECT 18.440000  27.350000 18.640000  27.550000 ;
        RECT 18.440000  27.780000 18.640000  27.980000 ;
        RECT 18.440000  28.210000 18.640000  28.410000 ;
        RECT 18.845000  23.910000 19.045000  24.110000 ;
        RECT 18.845000  24.340000 19.045000  24.540000 ;
        RECT 18.845000  24.770000 19.045000  24.970000 ;
        RECT 18.845000  25.200000 19.045000  25.400000 ;
        RECT 18.845000  25.630000 19.045000  25.830000 ;
        RECT 18.845000  26.060000 19.045000  26.260000 ;
        RECT 18.845000  26.490000 19.045000  26.690000 ;
        RECT 18.845000  26.920000 19.045000  27.120000 ;
        RECT 18.845000  27.350000 19.045000  27.550000 ;
        RECT 18.845000  27.780000 19.045000  27.980000 ;
        RECT 18.845000  28.210000 19.045000  28.410000 ;
        RECT 19.250000  23.910000 19.450000  24.110000 ;
        RECT 19.250000  24.340000 19.450000  24.540000 ;
        RECT 19.250000  24.770000 19.450000  24.970000 ;
        RECT 19.250000  25.200000 19.450000  25.400000 ;
        RECT 19.250000  25.630000 19.450000  25.830000 ;
        RECT 19.250000  26.060000 19.450000  26.260000 ;
        RECT 19.250000  26.490000 19.450000  26.690000 ;
        RECT 19.250000  26.920000 19.450000  27.120000 ;
        RECT 19.250000  27.350000 19.450000  27.550000 ;
        RECT 19.250000  27.780000 19.450000  27.980000 ;
        RECT 19.250000  28.210000 19.450000  28.410000 ;
        RECT 19.655000  23.910000 19.855000  24.110000 ;
        RECT 19.655000  24.340000 19.855000  24.540000 ;
        RECT 19.655000  24.770000 19.855000  24.970000 ;
        RECT 19.655000  25.200000 19.855000  25.400000 ;
        RECT 19.655000  25.630000 19.855000  25.830000 ;
        RECT 19.655000  26.060000 19.855000  26.260000 ;
        RECT 19.655000  26.490000 19.855000  26.690000 ;
        RECT 19.655000  26.920000 19.855000  27.120000 ;
        RECT 19.655000  27.350000 19.855000  27.550000 ;
        RECT 19.655000  27.780000 19.855000  27.980000 ;
        RECT 19.655000  28.210000 19.855000  28.410000 ;
        RECT 20.060000  23.910000 20.260000  24.110000 ;
        RECT 20.060000  24.340000 20.260000  24.540000 ;
        RECT 20.060000  24.770000 20.260000  24.970000 ;
        RECT 20.060000  25.200000 20.260000  25.400000 ;
        RECT 20.060000  25.630000 20.260000  25.830000 ;
        RECT 20.060000  26.060000 20.260000  26.260000 ;
        RECT 20.060000  26.490000 20.260000  26.690000 ;
        RECT 20.060000  26.920000 20.260000  27.120000 ;
        RECT 20.060000  27.350000 20.260000  27.550000 ;
        RECT 20.060000  27.780000 20.260000  27.980000 ;
        RECT 20.060000  28.210000 20.260000  28.410000 ;
        RECT 20.465000  23.910000 20.665000  24.110000 ;
        RECT 20.465000  24.340000 20.665000  24.540000 ;
        RECT 20.465000  24.770000 20.665000  24.970000 ;
        RECT 20.465000  25.200000 20.665000  25.400000 ;
        RECT 20.465000  25.630000 20.665000  25.830000 ;
        RECT 20.465000  26.060000 20.665000  26.260000 ;
        RECT 20.465000  26.490000 20.665000  26.690000 ;
        RECT 20.465000  26.920000 20.665000  27.120000 ;
        RECT 20.465000  27.350000 20.665000  27.550000 ;
        RECT 20.465000  27.780000 20.665000  27.980000 ;
        RECT 20.465000  28.210000 20.665000  28.410000 ;
        RECT 20.870000  23.910000 21.070000  24.110000 ;
        RECT 20.870000  24.340000 21.070000  24.540000 ;
        RECT 20.870000  24.770000 21.070000  24.970000 ;
        RECT 20.870000  25.200000 21.070000  25.400000 ;
        RECT 20.870000  25.630000 21.070000  25.830000 ;
        RECT 20.870000  26.060000 21.070000  26.260000 ;
        RECT 20.870000  26.490000 21.070000  26.690000 ;
        RECT 20.870000  26.920000 21.070000  27.120000 ;
        RECT 20.870000  27.350000 21.070000  27.550000 ;
        RECT 20.870000  27.780000 21.070000  27.980000 ;
        RECT 20.870000  28.210000 21.070000  28.410000 ;
        RECT 21.275000  23.910000 21.475000  24.110000 ;
        RECT 21.275000  24.340000 21.475000  24.540000 ;
        RECT 21.275000  24.770000 21.475000  24.970000 ;
        RECT 21.275000  25.200000 21.475000  25.400000 ;
        RECT 21.275000  25.630000 21.475000  25.830000 ;
        RECT 21.275000  26.060000 21.475000  26.260000 ;
        RECT 21.275000  26.490000 21.475000  26.690000 ;
        RECT 21.275000  26.920000 21.475000  27.120000 ;
        RECT 21.275000  27.350000 21.475000  27.550000 ;
        RECT 21.275000  27.780000 21.475000  27.980000 ;
        RECT 21.275000  28.210000 21.475000  28.410000 ;
        RECT 21.680000  23.910000 21.880000  24.110000 ;
        RECT 21.680000  24.340000 21.880000  24.540000 ;
        RECT 21.680000  24.770000 21.880000  24.970000 ;
        RECT 21.680000  25.200000 21.880000  25.400000 ;
        RECT 21.680000  25.630000 21.880000  25.830000 ;
        RECT 21.680000  26.060000 21.880000  26.260000 ;
        RECT 21.680000  26.490000 21.880000  26.690000 ;
        RECT 21.680000  26.920000 21.880000  27.120000 ;
        RECT 21.680000  27.350000 21.880000  27.550000 ;
        RECT 21.680000  27.780000 21.880000  27.980000 ;
        RECT 21.680000  28.210000 21.880000  28.410000 ;
        RECT 22.085000  23.910000 22.285000  24.110000 ;
        RECT 22.085000  24.340000 22.285000  24.540000 ;
        RECT 22.085000  24.770000 22.285000  24.970000 ;
        RECT 22.085000  25.200000 22.285000  25.400000 ;
        RECT 22.085000  25.630000 22.285000  25.830000 ;
        RECT 22.085000  26.060000 22.285000  26.260000 ;
        RECT 22.085000  26.490000 22.285000  26.690000 ;
        RECT 22.085000  26.920000 22.285000  27.120000 ;
        RECT 22.085000  27.350000 22.285000  27.550000 ;
        RECT 22.085000  27.780000 22.285000  27.980000 ;
        RECT 22.085000  28.210000 22.285000  28.410000 ;
        RECT 22.490000  23.910000 22.690000  24.110000 ;
        RECT 22.490000  24.340000 22.690000  24.540000 ;
        RECT 22.490000  24.770000 22.690000  24.970000 ;
        RECT 22.490000  25.200000 22.690000  25.400000 ;
        RECT 22.490000  25.630000 22.690000  25.830000 ;
        RECT 22.490000  26.060000 22.690000  26.260000 ;
        RECT 22.490000  26.490000 22.690000  26.690000 ;
        RECT 22.490000  26.920000 22.690000  27.120000 ;
        RECT 22.490000  27.350000 22.690000  27.550000 ;
        RECT 22.490000  27.780000 22.690000  27.980000 ;
        RECT 22.490000  28.210000 22.690000  28.410000 ;
        RECT 22.895000  23.910000 23.095000  24.110000 ;
        RECT 22.895000  24.340000 23.095000  24.540000 ;
        RECT 22.895000  24.770000 23.095000  24.970000 ;
        RECT 22.895000  25.200000 23.095000  25.400000 ;
        RECT 22.895000  25.630000 23.095000  25.830000 ;
        RECT 22.895000  26.060000 23.095000  26.260000 ;
        RECT 22.895000  26.490000 23.095000  26.690000 ;
        RECT 22.895000  26.920000 23.095000  27.120000 ;
        RECT 22.895000  27.350000 23.095000  27.550000 ;
        RECT 22.895000  27.780000 23.095000  27.980000 ;
        RECT 22.895000  28.210000 23.095000  28.410000 ;
        RECT 23.300000  23.910000 23.500000  24.110000 ;
        RECT 23.300000  24.340000 23.500000  24.540000 ;
        RECT 23.300000  24.770000 23.500000  24.970000 ;
        RECT 23.300000  25.200000 23.500000  25.400000 ;
        RECT 23.300000  25.630000 23.500000  25.830000 ;
        RECT 23.300000  26.060000 23.500000  26.260000 ;
        RECT 23.300000  26.490000 23.500000  26.690000 ;
        RECT 23.300000  26.920000 23.500000  27.120000 ;
        RECT 23.300000  27.350000 23.500000  27.550000 ;
        RECT 23.300000  27.780000 23.500000  27.980000 ;
        RECT 23.300000  28.210000 23.500000  28.410000 ;
        RECT 23.705000  23.910000 23.905000  24.110000 ;
        RECT 23.705000  24.340000 23.905000  24.540000 ;
        RECT 23.705000  24.770000 23.905000  24.970000 ;
        RECT 23.705000  25.200000 23.905000  25.400000 ;
        RECT 23.705000  25.630000 23.905000  25.830000 ;
        RECT 23.705000  26.060000 23.905000  26.260000 ;
        RECT 23.705000  26.490000 23.905000  26.690000 ;
        RECT 23.705000  26.920000 23.905000  27.120000 ;
        RECT 23.705000  27.350000 23.905000  27.550000 ;
        RECT 23.705000  27.780000 23.905000  27.980000 ;
        RECT 23.705000  28.210000 23.905000  28.410000 ;
        RECT 24.110000  23.910000 24.310000  24.110000 ;
        RECT 24.110000  24.340000 24.310000  24.540000 ;
        RECT 24.110000  24.770000 24.310000  24.970000 ;
        RECT 24.110000  25.200000 24.310000  25.400000 ;
        RECT 24.110000  25.630000 24.310000  25.830000 ;
        RECT 24.110000  26.060000 24.310000  26.260000 ;
        RECT 24.110000  26.490000 24.310000  26.690000 ;
        RECT 24.110000  26.920000 24.310000  27.120000 ;
        RECT 24.110000  27.350000 24.310000  27.550000 ;
        RECT 24.110000  27.780000 24.310000  27.980000 ;
        RECT 24.110000  28.210000 24.310000  28.410000 ;
        RECT 50.845000  23.910000 51.045000  24.110000 ;
        RECT 50.845000  24.340000 51.045000  24.540000 ;
        RECT 50.845000  24.770000 51.045000  24.970000 ;
        RECT 50.845000  25.200000 51.045000  25.400000 ;
        RECT 50.845000  25.630000 51.045000  25.830000 ;
        RECT 50.845000  26.060000 51.045000  26.260000 ;
        RECT 50.845000  26.490000 51.045000  26.690000 ;
        RECT 50.845000  26.920000 51.045000  27.120000 ;
        RECT 50.845000  27.350000 51.045000  27.550000 ;
        RECT 50.845000  27.780000 51.045000  27.980000 ;
        RECT 50.845000  28.210000 51.045000  28.410000 ;
        RECT 51.255000  23.910000 51.455000  24.110000 ;
        RECT 51.255000  24.340000 51.455000  24.540000 ;
        RECT 51.255000  24.770000 51.455000  24.970000 ;
        RECT 51.255000  25.200000 51.455000  25.400000 ;
        RECT 51.255000  25.630000 51.455000  25.830000 ;
        RECT 51.255000  26.060000 51.455000  26.260000 ;
        RECT 51.255000  26.490000 51.455000  26.690000 ;
        RECT 51.255000  26.920000 51.455000  27.120000 ;
        RECT 51.255000  27.350000 51.455000  27.550000 ;
        RECT 51.255000  27.780000 51.455000  27.980000 ;
        RECT 51.255000  28.210000 51.455000  28.410000 ;
        RECT 51.665000  23.910000 51.865000  24.110000 ;
        RECT 51.665000  24.340000 51.865000  24.540000 ;
        RECT 51.665000  24.770000 51.865000  24.970000 ;
        RECT 51.665000  25.200000 51.865000  25.400000 ;
        RECT 51.665000  25.630000 51.865000  25.830000 ;
        RECT 51.665000  26.060000 51.865000  26.260000 ;
        RECT 51.665000  26.490000 51.865000  26.690000 ;
        RECT 51.665000  26.920000 51.865000  27.120000 ;
        RECT 51.665000  27.350000 51.865000  27.550000 ;
        RECT 51.665000  27.780000 51.865000  27.980000 ;
        RECT 51.665000  28.210000 51.865000  28.410000 ;
        RECT 52.075000  23.910000 52.275000  24.110000 ;
        RECT 52.075000  24.340000 52.275000  24.540000 ;
        RECT 52.075000  24.770000 52.275000  24.970000 ;
        RECT 52.075000  25.200000 52.275000  25.400000 ;
        RECT 52.075000  25.630000 52.275000  25.830000 ;
        RECT 52.075000  26.060000 52.275000  26.260000 ;
        RECT 52.075000  26.490000 52.275000  26.690000 ;
        RECT 52.075000  26.920000 52.275000  27.120000 ;
        RECT 52.075000  27.350000 52.275000  27.550000 ;
        RECT 52.075000  27.780000 52.275000  27.980000 ;
        RECT 52.075000  28.210000 52.275000  28.410000 ;
        RECT 52.485000  23.910000 52.685000  24.110000 ;
        RECT 52.485000  24.340000 52.685000  24.540000 ;
        RECT 52.485000  24.770000 52.685000  24.970000 ;
        RECT 52.485000  25.200000 52.685000  25.400000 ;
        RECT 52.485000  25.630000 52.685000  25.830000 ;
        RECT 52.485000  26.060000 52.685000  26.260000 ;
        RECT 52.485000  26.490000 52.685000  26.690000 ;
        RECT 52.485000  26.920000 52.685000  27.120000 ;
        RECT 52.485000  27.350000 52.685000  27.550000 ;
        RECT 52.485000  27.780000 52.685000  27.980000 ;
        RECT 52.485000  28.210000 52.685000  28.410000 ;
        RECT 52.895000  23.910000 53.095000  24.110000 ;
        RECT 52.895000  24.340000 53.095000  24.540000 ;
        RECT 52.895000  24.770000 53.095000  24.970000 ;
        RECT 52.895000  25.200000 53.095000  25.400000 ;
        RECT 52.895000  25.630000 53.095000  25.830000 ;
        RECT 52.895000  26.060000 53.095000  26.260000 ;
        RECT 52.895000  26.490000 53.095000  26.690000 ;
        RECT 52.895000  26.920000 53.095000  27.120000 ;
        RECT 52.895000  27.350000 53.095000  27.550000 ;
        RECT 52.895000  27.780000 53.095000  27.980000 ;
        RECT 52.895000  28.210000 53.095000  28.410000 ;
        RECT 53.305000  23.910000 53.505000  24.110000 ;
        RECT 53.305000  24.340000 53.505000  24.540000 ;
        RECT 53.305000  24.770000 53.505000  24.970000 ;
        RECT 53.305000  25.200000 53.505000  25.400000 ;
        RECT 53.305000  25.630000 53.505000  25.830000 ;
        RECT 53.305000  26.060000 53.505000  26.260000 ;
        RECT 53.305000  26.490000 53.505000  26.690000 ;
        RECT 53.305000  26.920000 53.505000  27.120000 ;
        RECT 53.305000  27.350000 53.505000  27.550000 ;
        RECT 53.305000  27.780000 53.505000  27.980000 ;
        RECT 53.305000  28.210000 53.505000  28.410000 ;
        RECT 53.715000  23.910000 53.915000  24.110000 ;
        RECT 53.715000  24.340000 53.915000  24.540000 ;
        RECT 53.715000  24.770000 53.915000  24.970000 ;
        RECT 53.715000  25.200000 53.915000  25.400000 ;
        RECT 53.715000  25.630000 53.915000  25.830000 ;
        RECT 53.715000  26.060000 53.915000  26.260000 ;
        RECT 53.715000  26.490000 53.915000  26.690000 ;
        RECT 53.715000  26.920000 53.915000  27.120000 ;
        RECT 53.715000  27.350000 53.915000  27.550000 ;
        RECT 53.715000  27.780000 53.915000  27.980000 ;
        RECT 53.715000  28.210000 53.915000  28.410000 ;
        RECT 54.125000  23.910000 54.325000  24.110000 ;
        RECT 54.125000  24.340000 54.325000  24.540000 ;
        RECT 54.125000  24.770000 54.325000  24.970000 ;
        RECT 54.125000  25.200000 54.325000  25.400000 ;
        RECT 54.125000  25.630000 54.325000  25.830000 ;
        RECT 54.125000  26.060000 54.325000  26.260000 ;
        RECT 54.125000  26.490000 54.325000  26.690000 ;
        RECT 54.125000  26.920000 54.325000  27.120000 ;
        RECT 54.125000  27.350000 54.325000  27.550000 ;
        RECT 54.125000  27.780000 54.325000  27.980000 ;
        RECT 54.125000  28.210000 54.325000  28.410000 ;
        RECT 54.535000  23.910000 54.735000  24.110000 ;
        RECT 54.535000  24.340000 54.735000  24.540000 ;
        RECT 54.535000  24.770000 54.735000  24.970000 ;
        RECT 54.535000  25.200000 54.735000  25.400000 ;
        RECT 54.535000  25.630000 54.735000  25.830000 ;
        RECT 54.535000  26.060000 54.735000  26.260000 ;
        RECT 54.535000  26.490000 54.735000  26.690000 ;
        RECT 54.535000  26.920000 54.735000  27.120000 ;
        RECT 54.535000  27.350000 54.735000  27.550000 ;
        RECT 54.535000  27.780000 54.735000  27.980000 ;
        RECT 54.535000  28.210000 54.735000  28.410000 ;
        RECT 54.945000  23.910000 55.145000  24.110000 ;
        RECT 54.945000  24.340000 55.145000  24.540000 ;
        RECT 54.945000  24.770000 55.145000  24.970000 ;
        RECT 54.945000  25.200000 55.145000  25.400000 ;
        RECT 54.945000  25.630000 55.145000  25.830000 ;
        RECT 54.945000  26.060000 55.145000  26.260000 ;
        RECT 54.945000  26.490000 55.145000  26.690000 ;
        RECT 54.945000  26.920000 55.145000  27.120000 ;
        RECT 54.945000  27.350000 55.145000  27.550000 ;
        RECT 54.945000  27.780000 55.145000  27.980000 ;
        RECT 54.945000  28.210000 55.145000  28.410000 ;
        RECT 55.355000  23.910000 55.555000  24.110000 ;
        RECT 55.355000  24.340000 55.555000  24.540000 ;
        RECT 55.355000  24.770000 55.555000  24.970000 ;
        RECT 55.355000  25.200000 55.555000  25.400000 ;
        RECT 55.355000  25.630000 55.555000  25.830000 ;
        RECT 55.355000  26.060000 55.555000  26.260000 ;
        RECT 55.355000  26.490000 55.555000  26.690000 ;
        RECT 55.355000  26.920000 55.555000  27.120000 ;
        RECT 55.355000  27.350000 55.555000  27.550000 ;
        RECT 55.355000  27.780000 55.555000  27.980000 ;
        RECT 55.355000  28.210000 55.555000  28.410000 ;
        RECT 55.765000  23.910000 55.965000  24.110000 ;
        RECT 55.765000  24.340000 55.965000  24.540000 ;
        RECT 55.765000  24.770000 55.965000  24.970000 ;
        RECT 55.765000  25.200000 55.965000  25.400000 ;
        RECT 55.765000  25.630000 55.965000  25.830000 ;
        RECT 55.765000  26.060000 55.965000  26.260000 ;
        RECT 55.765000  26.490000 55.965000  26.690000 ;
        RECT 55.765000  26.920000 55.965000  27.120000 ;
        RECT 55.765000  27.350000 55.965000  27.550000 ;
        RECT 55.765000  27.780000 55.965000  27.980000 ;
        RECT 55.765000  28.210000 55.965000  28.410000 ;
        RECT 56.175000  23.910000 56.375000  24.110000 ;
        RECT 56.175000  24.340000 56.375000  24.540000 ;
        RECT 56.175000  24.770000 56.375000  24.970000 ;
        RECT 56.175000  25.200000 56.375000  25.400000 ;
        RECT 56.175000  25.630000 56.375000  25.830000 ;
        RECT 56.175000  26.060000 56.375000  26.260000 ;
        RECT 56.175000  26.490000 56.375000  26.690000 ;
        RECT 56.175000  26.920000 56.375000  27.120000 ;
        RECT 56.175000  27.350000 56.375000  27.550000 ;
        RECT 56.175000  27.780000 56.375000  27.980000 ;
        RECT 56.175000  28.210000 56.375000  28.410000 ;
        RECT 56.585000  23.910000 56.785000  24.110000 ;
        RECT 56.585000  24.340000 56.785000  24.540000 ;
        RECT 56.585000  24.770000 56.785000  24.970000 ;
        RECT 56.585000  25.200000 56.785000  25.400000 ;
        RECT 56.585000  25.630000 56.785000  25.830000 ;
        RECT 56.585000  26.060000 56.785000  26.260000 ;
        RECT 56.585000  26.490000 56.785000  26.690000 ;
        RECT 56.585000  26.920000 56.785000  27.120000 ;
        RECT 56.585000  27.350000 56.785000  27.550000 ;
        RECT 56.585000  27.780000 56.785000  27.980000 ;
        RECT 56.585000  28.210000 56.785000  28.410000 ;
        RECT 56.990000  23.910000 57.190000  24.110000 ;
        RECT 56.990000  24.340000 57.190000  24.540000 ;
        RECT 56.990000  24.770000 57.190000  24.970000 ;
        RECT 56.990000  25.200000 57.190000  25.400000 ;
        RECT 56.990000  25.630000 57.190000  25.830000 ;
        RECT 56.990000  26.060000 57.190000  26.260000 ;
        RECT 56.990000  26.490000 57.190000  26.690000 ;
        RECT 56.990000  26.920000 57.190000  27.120000 ;
        RECT 56.990000  27.350000 57.190000  27.550000 ;
        RECT 56.990000  27.780000 57.190000  27.980000 ;
        RECT 56.990000  28.210000 57.190000  28.410000 ;
        RECT 57.395000  23.910000 57.595000  24.110000 ;
        RECT 57.395000  24.340000 57.595000  24.540000 ;
        RECT 57.395000  24.770000 57.595000  24.970000 ;
        RECT 57.395000  25.200000 57.595000  25.400000 ;
        RECT 57.395000  25.630000 57.595000  25.830000 ;
        RECT 57.395000  26.060000 57.595000  26.260000 ;
        RECT 57.395000  26.490000 57.595000  26.690000 ;
        RECT 57.395000  26.920000 57.595000  27.120000 ;
        RECT 57.395000  27.350000 57.595000  27.550000 ;
        RECT 57.395000  27.780000 57.595000  27.980000 ;
        RECT 57.395000  28.210000 57.595000  28.410000 ;
        RECT 57.800000  23.910000 58.000000  24.110000 ;
        RECT 57.800000  24.340000 58.000000  24.540000 ;
        RECT 57.800000  24.770000 58.000000  24.970000 ;
        RECT 57.800000  25.200000 58.000000  25.400000 ;
        RECT 57.800000  25.630000 58.000000  25.830000 ;
        RECT 57.800000  26.060000 58.000000  26.260000 ;
        RECT 57.800000  26.490000 58.000000  26.690000 ;
        RECT 57.800000  26.920000 58.000000  27.120000 ;
        RECT 57.800000  27.350000 58.000000  27.550000 ;
        RECT 57.800000  27.780000 58.000000  27.980000 ;
        RECT 57.800000  28.210000 58.000000  28.410000 ;
        RECT 58.205000  23.910000 58.405000  24.110000 ;
        RECT 58.205000  24.340000 58.405000  24.540000 ;
        RECT 58.205000  24.770000 58.405000  24.970000 ;
        RECT 58.205000  25.200000 58.405000  25.400000 ;
        RECT 58.205000  25.630000 58.405000  25.830000 ;
        RECT 58.205000  26.060000 58.405000  26.260000 ;
        RECT 58.205000  26.490000 58.405000  26.690000 ;
        RECT 58.205000  26.920000 58.405000  27.120000 ;
        RECT 58.205000  27.350000 58.405000  27.550000 ;
        RECT 58.205000  27.780000 58.405000  27.980000 ;
        RECT 58.205000  28.210000 58.405000  28.410000 ;
        RECT 58.610000  23.910000 58.810000  24.110000 ;
        RECT 58.610000  24.340000 58.810000  24.540000 ;
        RECT 58.610000  24.770000 58.810000  24.970000 ;
        RECT 58.610000  25.200000 58.810000  25.400000 ;
        RECT 58.610000  25.630000 58.810000  25.830000 ;
        RECT 58.610000  26.060000 58.810000  26.260000 ;
        RECT 58.610000  26.490000 58.810000  26.690000 ;
        RECT 58.610000  26.920000 58.810000  27.120000 ;
        RECT 58.610000  27.350000 58.810000  27.550000 ;
        RECT 58.610000  27.780000 58.810000  27.980000 ;
        RECT 58.610000  28.210000 58.810000  28.410000 ;
        RECT 59.015000  23.910000 59.215000  24.110000 ;
        RECT 59.015000  24.340000 59.215000  24.540000 ;
        RECT 59.015000  24.770000 59.215000  24.970000 ;
        RECT 59.015000  25.200000 59.215000  25.400000 ;
        RECT 59.015000  25.630000 59.215000  25.830000 ;
        RECT 59.015000  26.060000 59.215000  26.260000 ;
        RECT 59.015000  26.490000 59.215000  26.690000 ;
        RECT 59.015000  26.920000 59.215000  27.120000 ;
        RECT 59.015000  27.350000 59.215000  27.550000 ;
        RECT 59.015000  27.780000 59.215000  27.980000 ;
        RECT 59.015000  28.210000 59.215000  28.410000 ;
        RECT 59.420000  23.910000 59.620000  24.110000 ;
        RECT 59.420000  24.340000 59.620000  24.540000 ;
        RECT 59.420000  24.770000 59.620000  24.970000 ;
        RECT 59.420000  25.200000 59.620000  25.400000 ;
        RECT 59.420000  25.630000 59.620000  25.830000 ;
        RECT 59.420000  26.060000 59.620000  26.260000 ;
        RECT 59.420000  26.490000 59.620000  26.690000 ;
        RECT 59.420000  26.920000 59.620000  27.120000 ;
        RECT 59.420000  27.350000 59.620000  27.550000 ;
        RECT 59.420000  27.780000 59.620000  27.980000 ;
        RECT 59.420000  28.210000 59.620000  28.410000 ;
        RECT 59.825000  23.910000 60.025000  24.110000 ;
        RECT 59.825000  24.340000 60.025000  24.540000 ;
        RECT 59.825000  24.770000 60.025000  24.970000 ;
        RECT 59.825000  25.200000 60.025000  25.400000 ;
        RECT 59.825000  25.630000 60.025000  25.830000 ;
        RECT 59.825000  26.060000 60.025000  26.260000 ;
        RECT 59.825000  26.490000 60.025000  26.690000 ;
        RECT 59.825000  26.920000 60.025000  27.120000 ;
        RECT 59.825000  27.350000 60.025000  27.550000 ;
        RECT 59.825000  27.780000 60.025000  27.980000 ;
        RECT 59.825000  28.210000 60.025000  28.410000 ;
        RECT 60.230000  23.910000 60.430000  24.110000 ;
        RECT 60.230000  24.340000 60.430000  24.540000 ;
        RECT 60.230000  24.770000 60.430000  24.970000 ;
        RECT 60.230000  25.200000 60.430000  25.400000 ;
        RECT 60.230000  25.630000 60.430000  25.830000 ;
        RECT 60.230000  26.060000 60.430000  26.260000 ;
        RECT 60.230000  26.490000 60.430000  26.690000 ;
        RECT 60.230000  26.920000 60.430000  27.120000 ;
        RECT 60.230000  27.350000 60.430000  27.550000 ;
        RECT 60.230000  27.780000 60.430000  27.980000 ;
        RECT 60.230000  28.210000 60.430000  28.410000 ;
        RECT 60.635000  23.910000 60.835000  24.110000 ;
        RECT 60.635000  24.340000 60.835000  24.540000 ;
        RECT 60.635000  24.770000 60.835000  24.970000 ;
        RECT 60.635000  25.200000 60.835000  25.400000 ;
        RECT 60.635000  25.630000 60.835000  25.830000 ;
        RECT 60.635000  26.060000 60.835000  26.260000 ;
        RECT 60.635000  26.490000 60.835000  26.690000 ;
        RECT 60.635000  26.920000 60.835000  27.120000 ;
        RECT 60.635000  27.350000 60.835000  27.550000 ;
        RECT 60.635000  27.780000 60.835000  27.980000 ;
        RECT 60.635000  28.210000 60.835000  28.410000 ;
        RECT 61.040000  23.910000 61.240000  24.110000 ;
        RECT 61.040000  24.340000 61.240000  24.540000 ;
        RECT 61.040000  24.770000 61.240000  24.970000 ;
        RECT 61.040000  25.200000 61.240000  25.400000 ;
        RECT 61.040000  25.630000 61.240000  25.830000 ;
        RECT 61.040000  26.060000 61.240000  26.260000 ;
        RECT 61.040000  26.490000 61.240000  26.690000 ;
        RECT 61.040000  26.920000 61.240000  27.120000 ;
        RECT 61.040000  27.350000 61.240000  27.550000 ;
        RECT 61.040000  27.780000 61.240000  27.980000 ;
        RECT 61.040000  28.210000 61.240000  28.410000 ;
        RECT 61.445000  23.910000 61.645000  24.110000 ;
        RECT 61.445000  24.340000 61.645000  24.540000 ;
        RECT 61.445000  24.770000 61.645000  24.970000 ;
        RECT 61.445000  25.200000 61.645000  25.400000 ;
        RECT 61.445000  25.630000 61.645000  25.830000 ;
        RECT 61.445000  26.060000 61.645000  26.260000 ;
        RECT 61.445000  26.490000 61.645000  26.690000 ;
        RECT 61.445000  26.920000 61.645000  27.120000 ;
        RECT 61.445000  27.350000 61.645000  27.550000 ;
        RECT 61.445000  27.780000 61.645000  27.980000 ;
        RECT 61.445000  28.210000 61.645000  28.410000 ;
        RECT 61.850000  23.910000 62.050000  24.110000 ;
        RECT 61.850000  24.340000 62.050000  24.540000 ;
        RECT 61.850000  24.770000 62.050000  24.970000 ;
        RECT 61.850000  25.200000 62.050000  25.400000 ;
        RECT 61.850000  25.630000 62.050000  25.830000 ;
        RECT 61.850000  26.060000 62.050000  26.260000 ;
        RECT 61.850000  26.490000 62.050000  26.690000 ;
        RECT 61.850000  26.920000 62.050000  27.120000 ;
        RECT 61.850000  27.350000 62.050000  27.550000 ;
        RECT 61.850000  27.780000 62.050000  27.980000 ;
        RECT 61.850000  28.210000 62.050000  28.410000 ;
        RECT 62.140000 173.900000 62.340000 174.100000 ;
        RECT 62.140000 174.300000 62.340000 174.500000 ;
        RECT 62.140000 174.700000 62.340000 174.900000 ;
        RECT 62.140000 175.100000 62.340000 175.300000 ;
        RECT 62.140000 175.500000 62.340000 175.700000 ;
        RECT 62.140000 175.900000 62.340000 176.100000 ;
        RECT 62.140000 176.300000 62.340000 176.500000 ;
        RECT 62.140000 176.700000 62.340000 176.900000 ;
        RECT 62.140000 177.100000 62.340000 177.300000 ;
        RECT 62.140000 177.500000 62.340000 177.700000 ;
        RECT 62.140000 177.900000 62.340000 178.100000 ;
        RECT 62.140000 178.300000 62.340000 178.500000 ;
        RECT 62.140000 178.700000 62.340000 178.900000 ;
        RECT 62.140000 179.100000 62.340000 179.300000 ;
        RECT 62.140000 179.500000 62.340000 179.700000 ;
        RECT 62.140000 179.900000 62.340000 180.100000 ;
        RECT 62.140000 180.300000 62.340000 180.500000 ;
        RECT 62.140000 180.700000 62.340000 180.900000 ;
        RECT 62.140000 181.100000 62.340000 181.300000 ;
        RECT 62.140000 181.505000 62.340000 181.705000 ;
        RECT 62.140000 181.910000 62.340000 182.110000 ;
        RECT 62.140000 182.315000 62.340000 182.515000 ;
        RECT 62.140000 182.720000 62.340000 182.920000 ;
        RECT 62.140000 183.125000 62.340000 183.325000 ;
        RECT 62.140000 183.530000 62.340000 183.730000 ;
        RECT 62.140000 183.935000 62.340000 184.135000 ;
        RECT 62.140000 184.340000 62.340000 184.540000 ;
        RECT 62.140000 184.745000 62.340000 184.945000 ;
        RECT 62.140000 185.150000 62.340000 185.350000 ;
        RECT 62.140000 185.555000 62.340000 185.755000 ;
        RECT 62.140000 185.960000 62.340000 186.160000 ;
        RECT 62.140000 186.365000 62.340000 186.565000 ;
        RECT 62.140000 186.770000 62.340000 186.970000 ;
        RECT 62.140000 187.175000 62.340000 187.375000 ;
        RECT 62.140000 187.580000 62.340000 187.780000 ;
        RECT 62.140000 187.985000 62.340000 188.185000 ;
        RECT 62.140000 188.390000 62.340000 188.590000 ;
        RECT 62.140000 188.795000 62.340000 188.995000 ;
        RECT 62.140000 189.200000 62.340000 189.400000 ;
        RECT 62.140000 189.605000 62.340000 189.805000 ;
        RECT 62.140000 190.010000 62.340000 190.210000 ;
        RECT 62.140000 190.415000 62.340000 190.615000 ;
        RECT 62.140000 190.820000 62.340000 191.020000 ;
        RECT 62.140000 191.225000 62.340000 191.425000 ;
        RECT 62.140000 191.630000 62.340000 191.830000 ;
        RECT 62.140000 192.035000 62.340000 192.235000 ;
        RECT 62.140000 192.440000 62.340000 192.640000 ;
        RECT 62.140000 192.845000 62.340000 193.045000 ;
        RECT 62.140000 193.250000 62.340000 193.450000 ;
        RECT 62.140000 193.655000 62.340000 193.855000 ;
        RECT 62.140000 194.060000 62.340000 194.260000 ;
        RECT 62.140000 194.465000 62.340000 194.665000 ;
        RECT 62.140000 194.870000 62.340000 195.070000 ;
        RECT 62.140000 195.275000 62.340000 195.475000 ;
        RECT 62.140000 195.680000 62.340000 195.880000 ;
        RECT 62.140000 196.085000 62.340000 196.285000 ;
        RECT 62.140000 196.490000 62.340000 196.690000 ;
        RECT 62.140000 196.895000 62.340000 197.095000 ;
        RECT 62.140000 197.300000 62.340000 197.500000 ;
        RECT 62.140000 197.705000 62.340000 197.905000 ;
        RECT 62.255000  23.910000 62.455000  24.110000 ;
        RECT 62.255000  24.340000 62.455000  24.540000 ;
        RECT 62.255000  24.770000 62.455000  24.970000 ;
        RECT 62.255000  25.200000 62.455000  25.400000 ;
        RECT 62.255000  25.630000 62.455000  25.830000 ;
        RECT 62.255000  26.060000 62.455000  26.260000 ;
        RECT 62.255000  26.490000 62.455000  26.690000 ;
        RECT 62.255000  26.920000 62.455000  27.120000 ;
        RECT 62.255000  27.350000 62.455000  27.550000 ;
        RECT 62.255000  27.780000 62.455000  27.980000 ;
        RECT 62.255000  28.210000 62.455000  28.410000 ;
        RECT 62.550000 173.900000 62.750000 174.100000 ;
        RECT 62.550000 174.300000 62.750000 174.500000 ;
        RECT 62.550000 174.700000 62.750000 174.900000 ;
        RECT 62.550000 175.100000 62.750000 175.300000 ;
        RECT 62.550000 175.500000 62.750000 175.700000 ;
        RECT 62.550000 175.900000 62.750000 176.100000 ;
        RECT 62.550000 176.300000 62.750000 176.500000 ;
        RECT 62.550000 176.700000 62.750000 176.900000 ;
        RECT 62.550000 177.100000 62.750000 177.300000 ;
        RECT 62.550000 177.500000 62.750000 177.700000 ;
        RECT 62.550000 177.900000 62.750000 178.100000 ;
        RECT 62.550000 178.300000 62.750000 178.500000 ;
        RECT 62.550000 178.700000 62.750000 178.900000 ;
        RECT 62.550000 179.100000 62.750000 179.300000 ;
        RECT 62.550000 179.500000 62.750000 179.700000 ;
        RECT 62.550000 179.900000 62.750000 180.100000 ;
        RECT 62.550000 180.300000 62.750000 180.500000 ;
        RECT 62.550000 180.700000 62.750000 180.900000 ;
        RECT 62.550000 181.100000 62.750000 181.300000 ;
        RECT 62.550000 181.505000 62.750000 181.705000 ;
        RECT 62.550000 181.910000 62.750000 182.110000 ;
        RECT 62.550000 182.315000 62.750000 182.515000 ;
        RECT 62.550000 182.720000 62.750000 182.920000 ;
        RECT 62.550000 183.125000 62.750000 183.325000 ;
        RECT 62.550000 183.530000 62.750000 183.730000 ;
        RECT 62.550000 183.935000 62.750000 184.135000 ;
        RECT 62.550000 184.340000 62.750000 184.540000 ;
        RECT 62.550000 184.745000 62.750000 184.945000 ;
        RECT 62.550000 185.150000 62.750000 185.350000 ;
        RECT 62.550000 185.555000 62.750000 185.755000 ;
        RECT 62.550000 185.960000 62.750000 186.160000 ;
        RECT 62.550000 186.365000 62.750000 186.565000 ;
        RECT 62.550000 186.770000 62.750000 186.970000 ;
        RECT 62.550000 187.175000 62.750000 187.375000 ;
        RECT 62.550000 187.580000 62.750000 187.780000 ;
        RECT 62.550000 187.985000 62.750000 188.185000 ;
        RECT 62.550000 188.390000 62.750000 188.590000 ;
        RECT 62.550000 188.795000 62.750000 188.995000 ;
        RECT 62.550000 189.200000 62.750000 189.400000 ;
        RECT 62.550000 189.605000 62.750000 189.805000 ;
        RECT 62.550000 190.010000 62.750000 190.210000 ;
        RECT 62.550000 190.415000 62.750000 190.615000 ;
        RECT 62.550000 190.820000 62.750000 191.020000 ;
        RECT 62.550000 191.225000 62.750000 191.425000 ;
        RECT 62.550000 191.630000 62.750000 191.830000 ;
        RECT 62.550000 192.035000 62.750000 192.235000 ;
        RECT 62.550000 192.440000 62.750000 192.640000 ;
        RECT 62.550000 192.845000 62.750000 193.045000 ;
        RECT 62.550000 193.250000 62.750000 193.450000 ;
        RECT 62.550000 193.655000 62.750000 193.855000 ;
        RECT 62.550000 194.060000 62.750000 194.260000 ;
        RECT 62.550000 194.465000 62.750000 194.665000 ;
        RECT 62.550000 194.870000 62.750000 195.070000 ;
        RECT 62.550000 195.275000 62.750000 195.475000 ;
        RECT 62.550000 195.680000 62.750000 195.880000 ;
        RECT 62.550000 196.085000 62.750000 196.285000 ;
        RECT 62.550000 196.490000 62.750000 196.690000 ;
        RECT 62.550000 196.895000 62.750000 197.095000 ;
        RECT 62.550000 197.300000 62.750000 197.500000 ;
        RECT 62.550000 197.705000 62.750000 197.905000 ;
        RECT 62.660000  23.910000 62.860000  24.110000 ;
        RECT 62.660000  24.340000 62.860000  24.540000 ;
        RECT 62.660000  24.770000 62.860000  24.970000 ;
        RECT 62.660000  25.200000 62.860000  25.400000 ;
        RECT 62.660000  25.630000 62.860000  25.830000 ;
        RECT 62.660000  26.060000 62.860000  26.260000 ;
        RECT 62.660000  26.490000 62.860000  26.690000 ;
        RECT 62.660000  26.920000 62.860000  27.120000 ;
        RECT 62.660000  27.350000 62.860000  27.550000 ;
        RECT 62.660000  27.780000 62.860000  27.980000 ;
        RECT 62.660000  28.210000 62.860000  28.410000 ;
        RECT 62.960000 173.900000 63.160000 174.100000 ;
        RECT 62.960000 174.300000 63.160000 174.500000 ;
        RECT 62.960000 174.700000 63.160000 174.900000 ;
        RECT 62.960000 175.100000 63.160000 175.300000 ;
        RECT 62.960000 175.500000 63.160000 175.700000 ;
        RECT 62.960000 175.900000 63.160000 176.100000 ;
        RECT 62.960000 176.300000 63.160000 176.500000 ;
        RECT 62.960000 176.700000 63.160000 176.900000 ;
        RECT 62.960000 177.100000 63.160000 177.300000 ;
        RECT 62.960000 177.500000 63.160000 177.700000 ;
        RECT 62.960000 177.900000 63.160000 178.100000 ;
        RECT 62.960000 178.300000 63.160000 178.500000 ;
        RECT 62.960000 178.700000 63.160000 178.900000 ;
        RECT 62.960000 179.100000 63.160000 179.300000 ;
        RECT 62.960000 179.500000 63.160000 179.700000 ;
        RECT 62.960000 179.900000 63.160000 180.100000 ;
        RECT 62.960000 180.300000 63.160000 180.500000 ;
        RECT 62.960000 180.700000 63.160000 180.900000 ;
        RECT 62.960000 181.100000 63.160000 181.300000 ;
        RECT 62.960000 181.505000 63.160000 181.705000 ;
        RECT 62.960000 181.910000 63.160000 182.110000 ;
        RECT 62.960000 182.315000 63.160000 182.515000 ;
        RECT 62.960000 182.720000 63.160000 182.920000 ;
        RECT 62.960000 183.125000 63.160000 183.325000 ;
        RECT 62.960000 183.530000 63.160000 183.730000 ;
        RECT 62.960000 183.935000 63.160000 184.135000 ;
        RECT 62.960000 184.340000 63.160000 184.540000 ;
        RECT 62.960000 184.745000 63.160000 184.945000 ;
        RECT 62.960000 185.150000 63.160000 185.350000 ;
        RECT 62.960000 185.555000 63.160000 185.755000 ;
        RECT 62.960000 185.960000 63.160000 186.160000 ;
        RECT 62.960000 186.365000 63.160000 186.565000 ;
        RECT 62.960000 186.770000 63.160000 186.970000 ;
        RECT 62.960000 187.175000 63.160000 187.375000 ;
        RECT 62.960000 187.580000 63.160000 187.780000 ;
        RECT 62.960000 187.985000 63.160000 188.185000 ;
        RECT 62.960000 188.390000 63.160000 188.590000 ;
        RECT 62.960000 188.795000 63.160000 188.995000 ;
        RECT 62.960000 189.200000 63.160000 189.400000 ;
        RECT 62.960000 189.605000 63.160000 189.805000 ;
        RECT 62.960000 190.010000 63.160000 190.210000 ;
        RECT 62.960000 190.415000 63.160000 190.615000 ;
        RECT 62.960000 190.820000 63.160000 191.020000 ;
        RECT 62.960000 191.225000 63.160000 191.425000 ;
        RECT 62.960000 191.630000 63.160000 191.830000 ;
        RECT 62.960000 192.035000 63.160000 192.235000 ;
        RECT 62.960000 192.440000 63.160000 192.640000 ;
        RECT 62.960000 192.845000 63.160000 193.045000 ;
        RECT 62.960000 193.250000 63.160000 193.450000 ;
        RECT 62.960000 193.655000 63.160000 193.855000 ;
        RECT 62.960000 194.060000 63.160000 194.260000 ;
        RECT 62.960000 194.465000 63.160000 194.665000 ;
        RECT 62.960000 194.870000 63.160000 195.070000 ;
        RECT 62.960000 195.275000 63.160000 195.475000 ;
        RECT 62.960000 195.680000 63.160000 195.880000 ;
        RECT 62.960000 196.085000 63.160000 196.285000 ;
        RECT 62.960000 196.490000 63.160000 196.690000 ;
        RECT 62.960000 196.895000 63.160000 197.095000 ;
        RECT 62.960000 197.300000 63.160000 197.500000 ;
        RECT 62.960000 197.705000 63.160000 197.905000 ;
        RECT 63.065000  23.910000 63.265000  24.110000 ;
        RECT 63.065000  24.340000 63.265000  24.540000 ;
        RECT 63.065000  24.770000 63.265000  24.970000 ;
        RECT 63.065000  25.200000 63.265000  25.400000 ;
        RECT 63.065000  25.630000 63.265000  25.830000 ;
        RECT 63.065000  26.060000 63.265000  26.260000 ;
        RECT 63.065000  26.490000 63.265000  26.690000 ;
        RECT 63.065000  26.920000 63.265000  27.120000 ;
        RECT 63.065000  27.350000 63.265000  27.550000 ;
        RECT 63.065000  27.780000 63.265000  27.980000 ;
        RECT 63.065000  28.210000 63.265000  28.410000 ;
        RECT 63.370000 173.900000 63.570000 174.100000 ;
        RECT 63.370000 174.300000 63.570000 174.500000 ;
        RECT 63.370000 174.700000 63.570000 174.900000 ;
        RECT 63.370000 175.100000 63.570000 175.300000 ;
        RECT 63.370000 175.500000 63.570000 175.700000 ;
        RECT 63.370000 175.900000 63.570000 176.100000 ;
        RECT 63.370000 176.300000 63.570000 176.500000 ;
        RECT 63.370000 176.700000 63.570000 176.900000 ;
        RECT 63.370000 177.100000 63.570000 177.300000 ;
        RECT 63.370000 177.500000 63.570000 177.700000 ;
        RECT 63.370000 177.900000 63.570000 178.100000 ;
        RECT 63.370000 178.300000 63.570000 178.500000 ;
        RECT 63.370000 178.700000 63.570000 178.900000 ;
        RECT 63.370000 179.100000 63.570000 179.300000 ;
        RECT 63.370000 179.500000 63.570000 179.700000 ;
        RECT 63.370000 179.900000 63.570000 180.100000 ;
        RECT 63.370000 180.300000 63.570000 180.500000 ;
        RECT 63.370000 180.700000 63.570000 180.900000 ;
        RECT 63.370000 181.100000 63.570000 181.300000 ;
        RECT 63.370000 181.505000 63.570000 181.705000 ;
        RECT 63.370000 181.910000 63.570000 182.110000 ;
        RECT 63.370000 182.315000 63.570000 182.515000 ;
        RECT 63.370000 182.720000 63.570000 182.920000 ;
        RECT 63.370000 183.125000 63.570000 183.325000 ;
        RECT 63.370000 183.530000 63.570000 183.730000 ;
        RECT 63.370000 183.935000 63.570000 184.135000 ;
        RECT 63.370000 184.340000 63.570000 184.540000 ;
        RECT 63.370000 184.745000 63.570000 184.945000 ;
        RECT 63.370000 185.150000 63.570000 185.350000 ;
        RECT 63.370000 185.555000 63.570000 185.755000 ;
        RECT 63.370000 185.960000 63.570000 186.160000 ;
        RECT 63.370000 186.365000 63.570000 186.565000 ;
        RECT 63.370000 186.770000 63.570000 186.970000 ;
        RECT 63.370000 187.175000 63.570000 187.375000 ;
        RECT 63.370000 187.580000 63.570000 187.780000 ;
        RECT 63.370000 187.985000 63.570000 188.185000 ;
        RECT 63.370000 188.390000 63.570000 188.590000 ;
        RECT 63.370000 188.795000 63.570000 188.995000 ;
        RECT 63.370000 189.200000 63.570000 189.400000 ;
        RECT 63.370000 189.605000 63.570000 189.805000 ;
        RECT 63.370000 190.010000 63.570000 190.210000 ;
        RECT 63.370000 190.415000 63.570000 190.615000 ;
        RECT 63.370000 190.820000 63.570000 191.020000 ;
        RECT 63.370000 191.225000 63.570000 191.425000 ;
        RECT 63.370000 191.630000 63.570000 191.830000 ;
        RECT 63.370000 192.035000 63.570000 192.235000 ;
        RECT 63.370000 192.440000 63.570000 192.640000 ;
        RECT 63.370000 192.845000 63.570000 193.045000 ;
        RECT 63.370000 193.250000 63.570000 193.450000 ;
        RECT 63.370000 193.655000 63.570000 193.855000 ;
        RECT 63.370000 194.060000 63.570000 194.260000 ;
        RECT 63.370000 194.465000 63.570000 194.665000 ;
        RECT 63.370000 194.870000 63.570000 195.070000 ;
        RECT 63.370000 195.275000 63.570000 195.475000 ;
        RECT 63.370000 195.680000 63.570000 195.880000 ;
        RECT 63.370000 196.085000 63.570000 196.285000 ;
        RECT 63.370000 196.490000 63.570000 196.690000 ;
        RECT 63.370000 196.895000 63.570000 197.095000 ;
        RECT 63.370000 197.300000 63.570000 197.500000 ;
        RECT 63.370000 197.705000 63.570000 197.905000 ;
        RECT 63.470000  23.910000 63.670000  24.110000 ;
        RECT 63.470000  24.340000 63.670000  24.540000 ;
        RECT 63.470000  24.770000 63.670000  24.970000 ;
        RECT 63.470000  25.200000 63.670000  25.400000 ;
        RECT 63.470000  25.630000 63.670000  25.830000 ;
        RECT 63.470000  26.060000 63.670000  26.260000 ;
        RECT 63.470000  26.490000 63.670000  26.690000 ;
        RECT 63.470000  26.920000 63.670000  27.120000 ;
        RECT 63.470000  27.350000 63.670000  27.550000 ;
        RECT 63.470000  27.780000 63.670000  27.980000 ;
        RECT 63.470000  28.210000 63.670000  28.410000 ;
        RECT 63.780000 173.900000 63.980000 174.100000 ;
        RECT 63.780000 174.300000 63.980000 174.500000 ;
        RECT 63.780000 174.700000 63.980000 174.900000 ;
        RECT 63.780000 175.100000 63.980000 175.300000 ;
        RECT 63.780000 175.500000 63.980000 175.700000 ;
        RECT 63.780000 175.900000 63.980000 176.100000 ;
        RECT 63.780000 176.300000 63.980000 176.500000 ;
        RECT 63.780000 176.700000 63.980000 176.900000 ;
        RECT 63.780000 177.100000 63.980000 177.300000 ;
        RECT 63.780000 177.500000 63.980000 177.700000 ;
        RECT 63.780000 177.900000 63.980000 178.100000 ;
        RECT 63.780000 178.300000 63.980000 178.500000 ;
        RECT 63.780000 178.700000 63.980000 178.900000 ;
        RECT 63.780000 179.100000 63.980000 179.300000 ;
        RECT 63.780000 179.500000 63.980000 179.700000 ;
        RECT 63.780000 179.900000 63.980000 180.100000 ;
        RECT 63.780000 180.300000 63.980000 180.500000 ;
        RECT 63.780000 180.700000 63.980000 180.900000 ;
        RECT 63.780000 181.100000 63.980000 181.300000 ;
        RECT 63.780000 181.505000 63.980000 181.705000 ;
        RECT 63.780000 181.910000 63.980000 182.110000 ;
        RECT 63.780000 182.315000 63.980000 182.515000 ;
        RECT 63.780000 182.720000 63.980000 182.920000 ;
        RECT 63.780000 183.125000 63.980000 183.325000 ;
        RECT 63.780000 183.530000 63.980000 183.730000 ;
        RECT 63.780000 183.935000 63.980000 184.135000 ;
        RECT 63.780000 184.340000 63.980000 184.540000 ;
        RECT 63.780000 184.745000 63.980000 184.945000 ;
        RECT 63.780000 185.150000 63.980000 185.350000 ;
        RECT 63.780000 185.555000 63.980000 185.755000 ;
        RECT 63.780000 185.960000 63.980000 186.160000 ;
        RECT 63.780000 186.365000 63.980000 186.565000 ;
        RECT 63.780000 186.770000 63.980000 186.970000 ;
        RECT 63.780000 187.175000 63.980000 187.375000 ;
        RECT 63.780000 187.580000 63.980000 187.780000 ;
        RECT 63.780000 187.985000 63.980000 188.185000 ;
        RECT 63.780000 188.390000 63.980000 188.590000 ;
        RECT 63.780000 188.795000 63.980000 188.995000 ;
        RECT 63.780000 189.200000 63.980000 189.400000 ;
        RECT 63.780000 189.605000 63.980000 189.805000 ;
        RECT 63.780000 190.010000 63.980000 190.210000 ;
        RECT 63.780000 190.415000 63.980000 190.615000 ;
        RECT 63.780000 190.820000 63.980000 191.020000 ;
        RECT 63.780000 191.225000 63.980000 191.425000 ;
        RECT 63.780000 191.630000 63.980000 191.830000 ;
        RECT 63.780000 192.035000 63.980000 192.235000 ;
        RECT 63.780000 192.440000 63.980000 192.640000 ;
        RECT 63.780000 192.845000 63.980000 193.045000 ;
        RECT 63.780000 193.250000 63.980000 193.450000 ;
        RECT 63.780000 193.655000 63.980000 193.855000 ;
        RECT 63.780000 194.060000 63.980000 194.260000 ;
        RECT 63.780000 194.465000 63.980000 194.665000 ;
        RECT 63.780000 194.870000 63.980000 195.070000 ;
        RECT 63.780000 195.275000 63.980000 195.475000 ;
        RECT 63.780000 195.680000 63.980000 195.880000 ;
        RECT 63.780000 196.085000 63.980000 196.285000 ;
        RECT 63.780000 196.490000 63.980000 196.690000 ;
        RECT 63.780000 196.895000 63.980000 197.095000 ;
        RECT 63.780000 197.300000 63.980000 197.500000 ;
        RECT 63.780000 197.705000 63.980000 197.905000 ;
        RECT 63.875000  23.910000 64.075000  24.110000 ;
        RECT 63.875000  24.340000 64.075000  24.540000 ;
        RECT 63.875000  24.770000 64.075000  24.970000 ;
        RECT 63.875000  25.200000 64.075000  25.400000 ;
        RECT 63.875000  25.630000 64.075000  25.830000 ;
        RECT 63.875000  26.060000 64.075000  26.260000 ;
        RECT 63.875000  26.490000 64.075000  26.690000 ;
        RECT 63.875000  26.920000 64.075000  27.120000 ;
        RECT 63.875000  27.350000 64.075000  27.550000 ;
        RECT 63.875000  27.780000 64.075000  27.980000 ;
        RECT 63.875000  28.210000 64.075000  28.410000 ;
        RECT 64.190000 173.900000 64.390000 174.100000 ;
        RECT 64.190000 174.300000 64.390000 174.500000 ;
        RECT 64.190000 174.700000 64.390000 174.900000 ;
        RECT 64.190000 175.100000 64.390000 175.300000 ;
        RECT 64.190000 175.500000 64.390000 175.700000 ;
        RECT 64.190000 175.900000 64.390000 176.100000 ;
        RECT 64.190000 176.300000 64.390000 176.500000 ;
        RECT 64.190000 176.700000 64.390000 176.900000 ;
        RECT 64.190000 177.100000 64.390000 177.300000 ;
        RECT 64.190000 177.500000 64.390000 177.700000 ;
        RECT 64.190000 177.900000 64.390000 178.100000 ;
        RECT 64.190000 178.300000 64.390000 178.500000 ;
        RECT 64.190000 178.700000 64.390000 178.900000 ;
        RECT 64.190000 179.100000 64.390000 179.300000 ;
        RECT 64.190000 179.500000 64.390000 179.700000 ;
        RECT 64.190000 179.900000 64.390000 180.100000 ;
        RECT 64.190000 180.300000 64.390000 180.500000 ;
        RECT 64.190000 180.700000 64.390000 180.900000 ;
        RECT 64.190000 181.100000 64.390000 181.300000 ;
        RECT 64.190000 181.505000 64.390000 181.705000 ;
        RECT 64.190000 181.910000 64.390000 182.110000 ;
        RECT 64.190000 182.315000 64.390000 182.515000 ;
        RECT 64.190000 182.720000 64.390000 182.920000 ;
        RECT 64.190000 183.125000 64.390000 183.325000 ;
        RECT 64.190000 183.530000 64.390000 183.730000 ;
        RECT 64.190000 183.935000 64.390000 184.135000 ;
        RECT 64.190000 184.340000 64.390000 184.540000 ;
        RECT 64.190000 184.745000 64.390000 184.945000 ;
        RECT 64.190000 185.150000 64.390000 185.350000 ;
        RECT 64.190000 185.555000 64.390000 185.755000 ;
        RECT 64.190000 185.960000 64.390000 186.160000 ;
        RECT 64.190000 186.365000 64.390000 186.565000 ;
        RECT 64.190000 186.770000 64.390000 186.970000 ;
        RECT 64.190000 187.175000 64.390000 187.375000 ;
        RECT 64.190000 187.580000 64.390000 187.780000 ;
        RECT 64.190000 187.985000 64.390000 188.185000 ;
        RECT 64.190000 188.390000 64.390000 188.590000 ;
        RECT 64.190000 188.795000 64.390000 188.995000 ;
        RECT 64.190000 189.200000 64.390000 189.400000 ;
        RECT 64.190000 189.605000 64.390000 189.805000 ;
        RECT 64.190000 190.010000 64.390000 190.210000 ;
        RECT 64.190000 190.415000 64.390000 190.615000 ;
        RECT 64.190000 190.820000 64.390000 191.020000 ;
        RECT 64.190000 191.225000 64.390000 191.425000 ;
        RECT 64.190000 191.630000 64.390000 191.830000 ;
        RECT 64.190000 192.035000 64.390000 192.235000 ;
        RECT 64.190000 192.440000 64.390000 192.640000 ;
        RECT 64.190000 192.845000 64.390000 193.045000 ;
        RECT 64.190000 193.250000 64.390000 193.450000 ;
        RECT 64.190000 193.655000 64.390000 193.855000 ;
        RECT 64.190000 194.060000 64.390000 194.260000 ;
        RECT 64.190000 194.465000 64.390000 194.665000 ;
        RECT 64.190000 194.870000 64.390000 195.070000 ;
        RECT 64.190000 195.275000 64.390000 195.475000 ;
        RECT 64.190000 195.680000 64.390000 195.880000 ;
        RECT 64.190000 196.085000 64.390000 196.285000 ;
        RECT 64.190000 196.490000 64.390000 196.690000 ;
        RECT 64.190000 196.895000 64.390000 197.095000 ;
        RECT 64.190000 197.300000 64.390000 197.500000 ;
        RECT 64.190000 197.705000 64.390000 197.905000 ;
        RECT 64.280000  23.910000 64.480000  24.110000 ;
        RECT 64.280000  24.340000 64.480000  24.540000 ;
        RECT 64.280000  24.770000 64.480000  24.970000 ;
        RECT 64.280000  25.200000 64.480000  25.400000 ;
        RECT 64.280000  25.630000 64.480000  25.830000 ;
        RECT 64.280000  26.060000 64.480000  26.260000 ;
        RECT 64.280000  26.490000 64.480000  26.690000 ;
        RECT 64.280000  26.920000 64.480000  27.120000 ;
        RECT 64.280000  27.350000 64.480000  27.550000 ;
        RECT 64.280000  27.780000 64.480000  27.980000 ;
        RECT 64.280000  28.210000 64.480000  28.410000 ;
        RECT 64.600000 173.900000 64.800000 174.100000 ;
        RECT 64.600000 174.300000 64.800000 174.500000 ;
        RECT 64.600000 174.700000 64.800000 174.900000 ;
        RECT 64.600000 175.100000 64.800000 175.300000 ;
        RECT 64.600000 175.500000 64.800000 175.700000 ;
        RECT 64.600000 175.900000 64.800000 176.100000 ;
        RECT 64.600000 176.300000 64.800000 176.500000 ;
        RECT 64.600000 176.700000 64.800000 176.900000 ;
        RECT 64.600000 177.100000 64.800000 177.300000 ;
        RECT 64.600000 177.500000 64.800000 177.700000 ;
        RECT 64.600000 177.900000 64.800000 178.100000 ;
        RECT 64.600000 178.300000 64.800000 178.500000 ;
        RECT 64.600000 178.700000 64.800000 178.900000 ;
        RECT 64.600000 179.100000 64.800000 179.300000 ;
        RECT 64.600000 179.500000 64.800000 179.700000 ;
        RECT 64.600000 179.900000 64.800000 180.100000 ;
        RECT 64.600000 180.300000 64.800000 180.500000 ;
        RECT 64.600000 180.700000 64.800000 180.900000 ;
        RECT 64.600000 181.100000 64.800000 181.300000 ;
        RECT 64.600000 181.505000 64.800000 181.705000 ;
        RECT 64.600000 181.910000 64.800000 182.110000 ;
        RECT 64.600000 182.315000 64.800000 182.515000 ;
        RECT 64.600000 182.720000 64.800000 182.920000 ;
        RECT 64.600000 183.125000 64.800000 183.325000 ;
        RECT 64.600000 183.530000 64.800000 183.730000 ;
        RECT 64.600000 183.935000 64.800000 184.135000 ;
        RECT 64.600000 184.340000 64.800000 184.540000 ;
        RECT 64.600000 184.745000 64.800000 184.945000 ;
        RECT 64.600000 185.150000 64.800000 185.350000 ;
        RECT 64.600000 185.555000 64.800000 185.755000 ;
        RECT 64.600000 185.960000 64.800000 186.160000 ;
        RECT 64.600000 186.365000 64.800000 186.565000 ;
        RECT 64.600000 186.770000 64.800000 186.970000 ;
        RECT 64.600000 187.175000 64.800000 187.375000 ;
        RECT 64.600000 187.580000 64.800000 187.780000 ;
        RECT 64.600000 187.985000 64.800000 188.185000 ;
        RECT 64.600000 188.390000 64.800000 188.590000 ;
        RECT 64.600000 188.795000 64.800000 188.995000 ;
        RECT 64.600000 189.200000 64.800000 189.400000 ;
        RECT 64.600000 189.605000 64.800000 189.805000 ;
        RECT 64.600000 190.010000 64.800000 190.210000 ;
        RECT 64.600000 190.415000 64.800000 190.615000 ;
        RECT 64.600000 190.820000 64.800000 191.020000 ;
        RECT 64.600000 191.225000 64.800000 191.425000 ;
        RECT 64.600000 191.630000 64.800000 191.830000 ;
        RECT 64.600000 192.035000 64.800000 192.235000 ;
        RECT 64.600000 192.440000 64.800000 192.640000 ;
        RECT 64.600000 192.845000 64.800000 193.045000 ;
        RECT 64.600000 193.250000 64.800000 193.450000 ;
        RECT 64.600000 193.655000 64.800000 193.855000 ;
        RECT 64.600000 194.060000 64.800000 194.260000 ;
        RECT 64.600000 194.465000 64.800000 194.665000 ;
        RECT 64.600000 194.870000 64.800000 195.070000 ;
        RECT 64.600000 195.275000 64.800000 195.475000 ;
        RECT 64.600000 195.680000 64.800000 195.880000 ;
        RECT 64.600000 196.085000 64.800000 196.285000 ;
        RECT 64.600000 196.490000 64.800000 196.690000 ;
        RECT 64.600000 196.895000 64.800000 197.095000 ;
        RECT 64.600000 197.300000 64.800000 197.500000 ;
        RECT 64.600000 197.705000 64.800000 197.905000 ;
        RECT 64.685000  23.910000 64.885000  24.110000 ;
        RECT 64.685000  24.340000 64.885000  24.540000 ;
        RECT 64.685000  24.770000 64.885000  24.970000 ;
        RECT 64.685000  25.200000 64.885000  25.400000 ;
        RECT 64.685000  25.630000 64.885000  25.830000 ;
        RECT 64.685000  26.060000 64.885000  26.260000 ;
        RECT 64.685000  26.490000 64.885000  26.690000 ;
        RECT 64.685000  26.920000 64.885000  27.120000 ;
        RECT 64.685000  27.350000 64.885000  27.550000 ;
        RECT 64.685000  27.780000 64.885000  27.980000 ;
        RECT 64.685000  28.210000 64.885000  28.410000 ;
        RECT 65.010000 173.900000 65.210000 174.100000 ;
        RECT 65.010000 174.300000 65.210000 174.500000 ;
        RECT 65.010000 174.700000 65.210000 174.900000 ;
        RECT 65.010000 175.100000 65.210000 175.300000 ;
        RECT 65.010000 175.500000 65.210000 175.700000 ;
        RECT 65.010000 175.900000 65.210000 176.100000 ;
        RECT 65.010000 176.300000 65.210000 176.500000 ;
        RECT 65.010000 176.700000 65.210000 176.900000 ;
        RECT 65.010000 177.100000 65.210000 177.300000 ;
        RECT 65.010000 177.500000 65.210000 177.700000 ;
        RECT 65.010000 177.900000 65.210000 178.100000 ;
        RECT 65.010000 178.300000 65.210000 178.500000 ;
        RECT 65.010000 178.700000 65.210000 178.900000 ;
        RECT 65.010000 179.100000 65.210000 179.300000 ;
        RECT 65.010000 179.500000 65.210000 179.700000 ;
        RECT 65.010000 179.900000 65.210000 180.100000 ;
        RECT 65.010000 180.300000 65.210000 180.500000 ;
        RECT 65.010000 180.700000 65.210000 180.900000 ;
        RECT 65.010000 181.100000 65.210000 181.300000 ;
        RECT 65.010000 181.505000 65.210000 181.705000 ;
        RECT 65.010000 181.910000 65.210000 182.110000 ;
        RECT 65.010000 182.315000 65.210000 182.515000 ;
        RECT 65.010000 182.720000 65.210000 182.920000 ;
        RECT 65.010000 183.125000 65.210000 183.325000 ;
        RECT 65.010000 183.530000 65.210000 183.730000 ;
        RECT 65.010000 183.935000 65.210000 184.135000 ;
        RECT 65.010000 184.340000 65.210000 184.540000 ;
        RECT 65.010000 184.745000 65.210000 184.945000 ;
        RECT 65.010000 185.150000 65.210000 185.350000 ;
        RECT 65.010000 185.555000 65.210000 185.755000 ;
        RECT 65.010000 185.960000 65.210000 186.160000 ;
        RECT 65.010000 186.365000 65.210000 186.565000 ;
        RECT 65.010000 186.770000 65.210000 186.970000 ;
        RECT 65.010000 187.175000 65.210000 187.375000 ;
        RECT 65.010000 187.580000 65.210000 187.780000 ;
        RECT 65.010000 187.985000 65.210000 188.185000 ;
        RECT 65.010000 188.390000 65.210000 188.590000 ;
        RECT 65.010000 188.795000 65.210000 188.995000 ;
        RECT 65.010000 189.200000 65.210000 189.400000 ;
        RECT 65.010000 189.605000 65.210000 189.805000 ;
        RECT 65.010000 190.010000 65.210000 190.210000 ;
        RECT 65.010000 190.415000 65.210000 190.615000 ;
        RECT 65.010000 190.820000 65.210000 191.020000 ;
        RECT 65.010000 191.225000 65.210000 191.425000 ;
        RECT 65.010000 191.630000 65.210000 191.830000 ;
        RECT 65.010000 192.035000 65.210000 192.235000 ;
        RECT 65.010000 192.440000 65.210000 192.640000 ;
        RECT 65.010000 192.845000 65.210000 193.045000 ;
        RECT 65.010000 193.250000 65.210000 193.450000 ;
        RECT 65.010000 193.655000 65.210000 193.855000 ;
        RECT 65.010000 194.060000 65.210000 194.260000 ;
        RECT 65.010000 194.465000 65.210000 194.665000 ;
        RECT 65.010000 194.870000 65.210000 195.070000 ;
        RECT 65.010000 195.275000 65.210000 195.475000 ;
        RECT 65.010000 195.680000 65.210000 195.880000 ;
        RECT 65.010000 196.085000 65.210000 196.285000 ;
        RECT 65.010000 196.490000 65.210000 196.690000 ;
        RECT 65.010000 196.895000 65.210000 197.095000 ;
        RECT 65.010000 197.300000 65.210000 197.500000 ;
        RECT 65.010000 197.705000 65.210000 197.905000 ;
        RECT 65.090000  23.910000 65.290000  24.110000 ;
        RECT 65.090000  24.340000 65.290000  24.540000 ;
        RECT 65.090000  24.770000 65.290000  24.970000 ;
        RECT 65.090000  25.200000 65.290000  25.400000 ;
        RECT 65.090000  25.630000 65.290000  25.830000 ;
        RECT 65.090000  26.060000 65.290000  26.260000 ;
        RECT 65.090000  26.490000 65.290000  26.690000 ;
        RECT 65.090000  26.920000 65.290000  27.120000 ;
        RECT 65.090000  27.350000 65.290000  27.550000 ;
        RECT 65.090000  27.780000 65.290000  27.980000 ;
        RECT 65.090000  28.210000 65.290000  28.410000 ;
        RECT 65.420000 173.900000 65.620000 174.100000 ;
        RECT 65.420000 174.300000 65.620000 174.500000 ;
        RECT 65.420000 174.700000 65.620000 174.900000 ;
        RECT 65.420000 175.100000 65.620000 175.300000 ;
        RECT 65.420000 175.500000 65.620000 175.700000 ;
        RECT 65.420000 175.900000 65.620000 176.100000 ;
        RECT 65.420000 176.300000 65.620000 176.500000 ;
        RECT 65.420000 176.700000 65.620000 176.900000 ;
        RECT 65.420000 177.100000 65.620000 177.300000 ;
        RECT 65.420000 177.500000 65.620000 177.700000 ;
        RECT 65.420000 177.900000 65.620000 178.100000 ;
        RECT 65.420000 178.300000 65.620000 178.500000 ;
        RECT 65.420000 178.700000 65.620000 178.900000 ;
        RECT 65.420000 179.100000 65.620000 179.300000 ;
        RECT 65.420000 179.500000 65.620000 179.700000 ;
        RECT 65.420000 179.900000 65.620000 180.100000 ;
        RECT 65.420000 180.300000 65.620000 180.500000 ;
        RECT 65.420000 180.700000 65.620000 180.900000 ;
        RECT 65.420000 181.100000 65.620000 181.300000 ;
        RECT 65.420000 181.505000 65.620000 181.705000 ;
        RECT 65.420000 181.910000 65.620000 182.110000 ;
        RECT 65.420000 182.315000 65.620000 182.515000 ;
        RECT 65.420000 182.720000 65.620000 182.920000 ;
        RECT 65.420000 183.125000 65.620000 183.325000 ;
        RECT 65.420000 183.530000 65.620000 183.730000 ;
        RECT 65.420000 183.935000 65.620000 184.135000 ;
        RECT 65.420000 184.340000 65.620000 184.540000 ;
        RECT 65.420000 184.745000 65.620000 184.945000 ;
        RECT 65.420000 185.150000 65.620000 185.350000 ;
        RECT 65.420000 185.555000 65.620000 185.755000 ;
        RECT 65.420000 185.960000 65.620000 186.160000 ;
        RECT 65.420000 186.365000 65.620000 186.565000 ;
        RECT 65.420000 186.770000 65.620000 186.970000 ;
        RECT 65.420000 187.175000 65.620000 187.375000 ;
        RECT 65.420000 187.580000 65.620000 187.780000 ;
        RECT 65.420000 187.985000 65.620000 188.185000 ;
        RECT 65.420000 188.390000 65.620000 188.590000 ;
        RECT 65.420000 188.795000 65.620000 188.995000 ;
        RECT 65.420000 189.200000 65.620000 189.400000 ;
        RECT 65.420000 189.605000 65.620000 189.805000 ;
        RECT 65.420000 190.010000 65.620000 190.210000 ;
        RECT 65.420000 190.415000 65.620000 190.615000 ;
        RECT 65.420000 190.820000 65.620000 191.020000 ;
        RECT 65.420000 191.225000 65.620000 191.425000 ;
        RECT 65.420000 191.630000 65.620000 191.830000 ;
        RECT 65.420000 192.035000 65.620000 192.235000 ;
        RECT 65.420000 192.440000 65.620000 192.640000 ;
        RECT 65.420000 192.845000 65.620000 193.045000 ;
        RECT 65.420000 193.250000 65.620000 193.450000 ;
        RECT 65.420000 193.655000 65.620000 193.855000 ;
        RECT 65.420000 194.060000 65.620000 194.260000 ;
        RECT 65.420000 194.465000 65.620000 194.665000 ;
        RECT 65.420000 194.870000 65.620000 195.070000 ;
        RECT 65.420000 195.275000 65.620000 195.475000 ;
        RECT 65.420000 195.680000 65.620000 195.880000 ;
        RECT 65.420000 196.085000 65.620000 196.285000 ;
        RECT 65.420000 196.490000 65.620000 196.690000 ;
        RECT 65.420000 196.895000 65.620000 197.095000 ;
        RECT 65.420000 197.300000 65.620000 197.500000 ;
        RECT 65.420000 197.705000 65.620000 197.905000 ;
        RECT 65.495000  23.910000 65.695000  24.110000 ;
        RECT 65.495000  24.340000 65.695000  24.540000 ;
        RECT 65.495000  24.770000 65.695000  24.970000 ;
        RECT 65.495000  25.200000 65.695000  25.400000 ;
        RECT 65.495000  25.630000 65.695000  25.830000 ;
        RECT 65.495000  26.060000 65.695000  26.260000 ;
        RECT 65.495000  26.490000 65.695000  26.690000 ;
        RECT 65.495000  26.920000 65.695000  27.120000 ;
        RECT 65.495000  27.350000 65.695000  27.550000 ;
        RECT 65.495000  27.780000 65.695000  27.980000 ;
        RECT 65.495000  28.210000 65.695000  28.410000 ;
        RECT 65.830000 173.900000 66.030000 174.100000 ;
        RECT 65.830000 174.300000 66.030000 174.500000 ;
        RECT 65.830000 174.700000 66.030000 174.900000 ;
        RECT 65.830000 175.100000 66.030000 175.300000 ;
        RECT 65.830000 175.500000 66.030000 175.700000 ;
        RECT 65.830000 175.900000 66.030000 176.100000 ;
        RECT 65.830000 176.300000 66.030000 176.500000 ;
        RECT 65.830000 176.700000 66.030000 176.900000 ;
        RECT 65.830000 177.100000 66.030000 177.300000 ;
        RECT 65.830000 177.500000 66.030000 177.700000 ;
        RECT 65.830000 177.900000 66.030000 178.100000 ;
        RECT 65.830000 178.300000 66.030000 178.500000 ;
        RECT 65.830000 178.700000 66.030000 178.900000 ;
        RECT 65.830000 179.100000 66.030000 179.300000 ;
        RECT 65.830000 179.500000 66.030000 179.700000 ;
        RECT 65.830000 179.900000 66.030000 180.100000 ;
        RECT 65.830000 180.300000 66.030000 180.500000 ;
        RECT 65.830000 180.700000 66.030000 180.900000 ;
        RECT 65.830000 181.100000 66.030000 181.300000 ;
        RECT 65.830000 181.505000 66.030000 181.705000 ;
        RECT 65.830000 181.910000 66.030000 182.110000 ;
        RECT 65.830000 182.315000 66.030000 182.515000 ;
        RECT 65.830000 182.720000 66.030000 182.920000 ;
        RECT 65.830000 183.125000 66.030000 183.325000 ;
        RECT 65.830000 183.530000 66.030000 183.730000 ;
        RECT 65.830000 183.935000 66.030000 184.135000 ;
        RECT 65.830000 184.340000 66.030000 184.540000 ;
        RECT 65.830000 184.745000 66.030000 184.945000 ;
        RECT 65.830000 185.150000 66.030000 185.350000 ;
        RECT 65.830000 185.555000 66.030000 185.755000 ;
        RECT 65.830000 185.960000 66.030000 186.160000 ;
        RECT 65.830000 186.365000 66.030000 186.565000 ;
        RECT 65.830000 186.770000 66.030000 186.970000 ;
        RECT 65.830000 187.175000 66.030000 187.375000 ;
        RECT 65.830000 187.580000 66.030000 187.780000 ;
        RECT 65.830000 187.985000 66.030000 188.185000 ;
        RECT 65.830000 188.390000 66.030000 188.590000 ;
        RECT 65.830000 188.795000 66.030000 188.995000 ;
        RECT 65.830000 189.200000 66.030000 189.400000 ;
        RECT 65.830000 189.605000 66.030000 189.805000 ;
        RECT 65.830000 190.010000 66.030000 190.210000 ;
        RECT 65.830000 190.415000 66.030000 190.615000 ;
        RECT 65.830000 190.820000 66.030000 191.020000 ;
        RECT 65.830000 191.225000 66.030000 191.425000 ;
        RECT 65.830000 191.630000 66.030000 191.830000 ;
        RECT 65.830000 192.035000 66.030000 192.235000 ;
        RECT 65.830000 192.440000 66.030000 192.640000 ;
        RECT 65.830000 192.845000 66.030000 193.045000 ;
        RECT 65.830000 193.250000 66.030000 193.450000 ;
        RECT 65.830000 193.655000 66.030000 193.855000 ;
        RECT 65.830000 194.060000 66.030000 194.260000 ;
        RECT 65.830000 194.465000 66.030000 194.665000 ;
        RECT 65.830000 194.870000 66.030000 195.070000 ;
        RECT 65.830000 195.275000 66.030000 195.475000 ;
        RECT 65.830000 195.680000 66.030000 195.880000 ;
        RECT 65.830000 196.085000 66.030000 196.285000 ;
        RECT 65.830000 196.490000 66.030000 196.690000 ;
        RECT 65.830000 196.895000 66.030000 197.095000 ;
        RECT 65.830000 197.300000 66.030000 197.500000 ;
        RECT 65.830000 197.705000 66.030000 197.905000 ;
        RECT 65.900000  23.910000 66.100000  24.110000 ;
        RECT 65.900000  24.340000 66.100000  24.540000 ;
        RECT 65.900000  24.770000 66.100000  24.970000 ;
        RECT 65.900000  25.200000 66.100000  25.400000 ;
        RECT 65.900000  25.630000 66.100000  25.830000 ;
        RECT 65.900000  26.060000 66.100000  26.260000 ;
        RECT 65.900000  26.490000 66.100000  26.690000 ;
        RECT 65.900000  26.920000 66.100000  27.120000 ;
        RECT 65.900000  27.350000 66.100000  27.550000 ;
        RECT 65.900000  27.780000 66.100000  27.980000 ;
        RECT 65.900000  28.210000 66.100000  28.410000 ;
        RECT 66.240000 173.900000 66.440000 174.100000 ;
        RECT 66.240000 174.300000 66.440000 174.500000 ;
        RECT 66.240000 174.700000 66.440000 174.900000 ;
        RECT 66.240000 175.100000 66.440000 175.300000 ;
        RECT 66.240000 175.500000 66.440000 175.700000 ;
        RECT 66.240000 175.900000 66.440000 176.100000 ;
        RECT 66.240000 176.300000 66.440000 176.500000 ;
        RECT 66.240000 176.700000 66.440000 176.900000 ;
        RECT 66.240000 177.100000 66.440000 177.300000 ;
        RECT 66.240000 177.500000 66.440000 177.700000 ;
        RECT 66.240000 177.900000 66.440000 178.100000 ;
        RECT 66.240000 178.300000 66.440000 178.500000 ;
        RECT 66.240000 178.700000 66.440000 178.900000 ;
        RECT 66.240000 179.100000 66.440000 179.300000 ;
        RECT 66.240000 179.500000 66.440000 179.700000 ;
        RECT 66.240000 179.900000 66.440000 180.100000 ;
        RECT 66.240000 180.300000 66.440000 180.500000 ;
        RECT 66.240000 180.700000 66.440000 180.900000 ;
        RECT 66.240000 181.100000 66.440000 181.300000 ;
        RECT 66.240000 181.505000 66.440000 181.705000 ;
        RECT 66.240000 181.910000 66.440000 182.110000 ;
        RECT 66.240000 182.315000 66.440000 182.515000 ;
        RECT 66.240000 182.720000 66.440000 182.920000 ;
        RECT 66.240000 183.125000 66.440000 183.325000 ;
        RECT 66.240000 183.530000 66.440000 183.730000 ;
        RECT 66.240000 183.935000 66.440000 184.135000 ;
        RECT 66.240000 184.340000 66.440000 184.540000 ;
        RECT 66.240000 184.745000 66.440000 184.945000 ;
        RECT 66.240000 185.150000 66.440000 185.350000 ;
        RECT 66.240000 185.555000 66.440000 185.755000 ;
        RECT 66.240000 185.960000 66.440000 186.160000 ;
        RECT 66.240000 186.365000 66.440000 186.565000 ;
        RECT 66.240000 186.770000 66.440000 186.970000 ;
        RECT 66.240000 187.175000 66.440000 187.375000 ;
        RECT 66.240000 187.580000 66.440000 187.780000 ;
        RECT 66.240000 187.985000 66.440000 188.185000 ;
        RECT 66.240000 188.390000 66.440000 188.590000 ;
        RECT 66.240000 188.795000 66.440000 188.995000 ;
        RECT 66.240000 189.200000 66.440000 189.400000 ;
        RECT 66.240000 189.605000 66.440000 189.805000 ;
        RECT 66.240000 190.010000 66.440000 190.210000 ;
        RECT 66.240000 190.415000 66.440000 190.615000 ;
        RECT 66.240000 190.820000 66.440000 191.020000 ;
        RECT 66.240000 191.225000 66.440000 191.425000 ;
        RECT 66.240000 191.630000 66.440000 191.830000 ;
        RECT 66.240000 192.035000 66.440000 192.235000 ;
        RECT 66.240000 192.440000 66.440000 192.640000 ;
        RECT 66.240000 192.845000 66.440000 193.045000 ;
        RECT 66.240000 193.250000 66.440000 193.450000 ;
        RECT 66.240000 193.655000 66.440000 193.855000 ;
        RECT 66.240000 194.060000 66.440000 194.260000 ;
        RECT 66.240000 194.465000 66.440000 194.665000 ;
        RECT 66.240000 194.870000 66.440000 195.070000 ;
        RECT 66.240000 195.275000 66.440000 195.475000 ;
        RECT 66.240000 195.680000 66.440000 195.880000 ;
        RECT 66.240000 196.085000 66.440000 196.285000 ;
        RECT 66.240000 196.490000 66.440000 196.690000 ;
        RECT 66.240000 196.895000 66.440000 197.095000 ;
        RECT 66.240000 197.300000 66.440000 197.500000 ;
        RECT 66.240000 197.705000 66.440000 197.905000 ;
        RECT 66.305000  23.910000 66.505000  24.110000 ;
        RECT 66.305000  24.340000 66.505000  24.540000 ;
        RECT 66.305000  24.770000 66.505000  24.970000 ;
        RECT 66.305000  25.200000 66.505000  25.400000 ;
        RECT 66.305000  25.630000 66.505000  25.830000 ;
        RECT 66.305000  26.060000 66.505000  26.260000 ;
        RECT 66.305000  26.490000 66.505000  26.690000 ;
        RECT 66.305000  26.920000 66.505000  27.120000 ;
        RECT 66.305000  27.350000 66.505000  27.550000 ;
        RECT 66.305000  27.780000 66.505000  27.980000 ;
        RECT 66.305000  28.210000 66.505000  28.410000 ;
        RECT 66.650000 173.900000 66.850000 174.100000 ;
        RECT 66.650000 174.300000 66.850000 174.500000 ;
        RECT 66.650000 174.700000 66.850000 174.900000 ;
        RECT 66.650000 175.100000 66.850000 175.300000 ;
        RECT 66.650000 175.500000 66.850000 175.700000 ;
        RECT 66.650000 175.900000 66.850000 176.100000 ;
        RECT 66.650000 176.300000 66.850000 176.500000 ;
        RECT 66.650000 176.700000 66.850000 176.900000 ;
        RECT 66.650000 177.100000 66.850000 177.300000 ;
        RECT 66.650000 177.500000 66.850000 177.700000 ;
        RECT 66.650000 177.900000 66.850000 178.100000 ;
        RECT 66.650000 178.300000 66.850000 178.500000 ;
        RECT 66.650000 178.700000 66.850000 178.900000 ;
        RECT 66.650000 179.100000 66.850000 179.300000 ;
        RECT 66.650000 179.500000 66.850000 179.700000 ;
        RECT 66.650000 179.900000 66.850000 180.100000 ;
        RECT 66.650000 180.300000 66.850000 180.500000 ;
        RECT 66.650000 180.700000 66.850000 180.900000 ;
        RECT 66.650000 181.100000 66.850000 181.300000 ;
        RECT 66.650000 181.505000 66.850000 181.705000 ;
        RECT 66.650000 181.910000 66.850000 182.110000 ;
        RECT 66.650000 182.315000 66.850000 182.515000 ;
        RECT 66.650000 182.720000 66.850000 182.920000 ;
        RECT 66.650000 183.125000 66.850000 183.325000 ;
        RECT 66.650000 183.530000 66.850000 183.730000 ;
        RECT 66.650000 183.935000 66.850000 184.135000 ;
        RECT 66.650000 184.340000 66.850000 184.540000 ;
        RECT 66.650000 184.745000 66.850000 184.945000 ;
        RECT 66.650000 185.150000 66.850000 185.350000 ;
        RECT 66.650000 185.555000 66.850000 185.755000 ;
        RECT 66.650000 185.960000 66.850000 186.160000 ;
        RECT 66.650000 186.365000 66.850000 186.565000 ;
        RECT 66.650000 186.770000 66.850000 186.970000 ;
        RECT 66.650000 187.175000 66.850000 187.375000 ;
        RECT 66.650000 187.580000 66.850000 187.780000 ;
        RECT 66.650000 187.985000 66.850000 188.185000 ;
        RECT 66.650000 188.390000 66.850000 188.590000 ;
        RECT 66.650000 188.795000 66.850000 188.995000 ;
        RECT 66.650000 189.200000 66.850000 189.400000 ;
        RECT 66.650000 189.605000 66.850000 189.805000 ;
        RECT 66.650000 190.010000 66.850000 190.210000 ;
        RECT 66.650000 190.415000 66.850000 190.615000 ;
        RECT 66.650000 190.820000 66.850000 191.020000 ;
        RECT 66.650000 191.225000 66.850000 191.425000 ;
        RECT 66.650000 191.630000 66.850000 191.830000 ;
        RECT 66.650000 192.035000 66.850000 192.235000 ;
        RECT 66.650000 192.440000 66.850000 192.640000 ;
        RECT 66.650000 192.845000 66.850000 193.045000 ;
        RECT 66.650000 193.250000 66.850000 193.450000 ;
        RECT 66.650000 193.655000 66.850000 193.855000 ;
        RECT 66.650000 194.060000 66.850000 194.260000 ;
        RECT 66.650000 194.465000 66.850000 194.665000 ;
        RECT 66.650000 194.870000 66.850000 195.070000 ;
        RECT 66.650000 195.275000 66.850000 195.475000 ;
        RECT 66.650000 195.680000 66.850000 195.880000 ;
        RECT 66.650000 196.085000 66.850000 196.285000 ;
        RECT 66.650000 196.490000 66.850000 196.690000 ;
        RECT 66.650000 196.895000 66.850000 197.095000 ;
        RECT 66.650000 197.300000 66.850000 197.500000 ;
        RECT 66.650000 197.705000 66.850000 197.905000 ;
        RECT 66.710000  23.910000 66.910000  24.110000 ;
        RECT 66.710000  24.340000 66.910000  24.540000 ;
        RECT 66.710000  24.770000 66.910000  24.970000 ;
        RECT 66.710000  25.200000 66.910000  25.400000 ;
        RECT 66.710000  25.630000 66.910000  25.830000 ;
        RECT 66.710000  26.060000 66.910000  26.260000 ;
        RECT 66.710000  26.490000 66.910000  26.690000 ;
        RECT 66.710000  26.920000 66.910000  27.120000 ;
        RECT 66.710000  27.350000 66.910000  27.550000 ;
        RECT 66.710000  27.780000 66.910000  27.980000 ;
        RECT 66.710000  28.210000 66.910000  28.410000 ;
        RECT 67.060000 173.900000 67.260000 174.100000 ;
        RECT 67.060000 174.300000 67.260000 174.500000 ;
        RECT 67.060000 174.700000 67.260000 174.900000 ;
        RECT 67.060000 175.100000 67.260000 175.300000 ;
        RECT 67.060000 175.500000 67.260000 175.700000 ;
        RECT 67.060000 175.900000 67.260000 176.100000 ;
        RECT 67.060000 176.300000 67.260000 176.500000 ;
        RECT 67.060000 176.700000 67.260000 176.900000 ;
        RECT 67.060000 177.100000 67.260000 177.300000 ;
        RECT 67.060000 177.500000 67.260000 177.700000 ;
        RECT 67.060000 177.900000 67.260000 178.100000 ;
        RECT 67.060000 178.300000 67.260000 178.500000 ;
        RECT 67.060000 178.700000 67.260000 178.900000 ;
        RECT 67.060000 179.100000 67.260000 179.300000 ;
        RECT 67.060000 179.500000 67.260000 179.700000 ;
        RECT 67.060000 179.900000 67.260000 180.100000 ;
        RECT 67.060000 180.300000 67.260000 180.500000 ;
        RECT 67.060000 180.700000 67.260000 180.900000 ;
        RECT 67.060000 181.100000 67.260000 181.300000 ;
        RECT 67.060000 181.505000 67.260000 181.705000 ;
        RECT 67.060000 181.910000 67.260000 182.110000 ;
        RECT 67.060000 182.315000 67.260000 182.515000 ;
        RECT 67.060000 182.720000 67.260000 182.920000 ;
        RECT 67.060000 183.125000 67.260000 183.325000 ;
        RECT 67.060000 183.530000 67.260000 183.730000 ;
        RECT 67.060000 183.935000 67.260000 184.135000 ;
        RECT 67.060000 184.340000 67.260000 184.540000 ;
        RECT 67.060000 184.745000 67.260000 184.945000 ;
        RECT 67.060000 185.150000 67.260000 185.350000 ;
        RECT 67.060000 185.555000 67.260000 185.755000 ;
        RECT 67.060000 185.960000 67.260000 186.160000 ;
        RECT 67.060000 186.365000 67.260000 186.565000 ;
        RECT 67.060000 186.770000 67.260000 186.970000 ;
        RECT 67.060000 187.175000 67.260000 187.375000 ;
        RECT 67.060000 187.580000 67.260000 187.780000 ;
        RECT 67.060000 187.985000 67.260000 188.185000 ;
        RECT 67.060000 188.390000 67.260000 188.590000 ;
        RECT 67.060000 188.795000 67.260000 188.995000 ;
        RECT 67.060000 189.200000 67.260000 189.400000 ;
        RECT 67.060000 189.605000 67.260000 189.805000 ;
        RECT 67.060000 190.010000 67.260000 190.210000 ;
        RECT 67.060000 190.415000 67.260000 190.615000 ;
        RECT 67.060000 190.820000 67.260000 191.020000 ;
        RECT 67.060000 191.225000 67.260000 191.425000 ;
        RECT 67.060000 191.630000 67.260000 191.830000 ;
        RECT 67.060000 192.035000 67.260000 192.235000 ;
        RECT 67.060000 192.440000 67.260000 192.640000 ;
        RECT 67.060000 192.845000 67.260000 193.045000 ;
        RECT 67.060000 193.250000 67.260000 193.450000 ;
        RECT 67.060000 193.655000 67.260000 193.855000 ;
        RECT 67.060000 194.060000 67.260000 194.260000 ;
        RECT 67.060000 194.465000 67.260000 194.665000 ;
        RECT 67.060000 194.870000 67.260000 195.070000 ;
        RECT 67.060000 195.275000 67.260000 195.475000 ;
        RECT 67.060000 195.680000 67.260000 195.880000 ;
        RECT 67.060000 196.085000 67.260000 196.285000 ;
        RECT 67.060000 196.490000 67.260000 196.690000 ;
        RECT 67.060000 196.895000 67.260000 197.095000 ;
        RECT 67.060000 197.300000 67.260000 197.500000 ;
        RECT 67.060000 197.705000 67.260000 197.905000 ;
        RECT 67.115000  23.910000 67.315000  24.110000 ;
        RECT 67.115000  24.340000 67.315000  24.540000 ;
        RECT 67.115000  24.770000 67.315000  24.970000 ;
        RECT 67.115000  25.200000 67.315000  25.400000 ;
        RECT 67.115000  25.630000 67.315000  25.830000 ;
        RECT 67.115000  26.060000 67.315000  26.260000 ;
        RECT 67.115000  26.490000 67.315000  26.690000 ;
        RECT 67.115000  26.920000 67.315000  27.120000 ;
        RECT 67.115000  27.350000 67.315000  27.550000 ;
        RECT 67.115000  27.780000 67.315000  27.980000 ;
        RECT 67.115000  28.210000 67.315000  28.410000 ;
        RECT 67.470000 173.900000 67.670000 174.100000 ;
        RECT 67.470000 174.300000 67.670000 174.500000 ;
        RECT 67.470000 174.700000 67.670000 174.900000 ;
        RECT 67.470000 175.100000 67.670000 175.300000 ;
        RECT 67.470000 175.500000 67.670000 175.700000 ;
        RECT 67.470000 175.900000 67.670000 176.100000 ;
        RECT 67.470000 176.300000 67.670000 176.500000 ;
        RECT 67.470000 176.700000 67.670000 176.900000 ;
        RECT 67.470000 177.100000 67.670000 177.300000 ;
        RECT 67.470000 177.500000 67.670000 177.700000 ;
        RECT 67.470000 177.900000 67.670000 178.100000 ;
        RECT 67.470000 178.300000 67.670000 178.500000 ;
        RECT 67.470000 178.700000 67.670000 178.900000 ;
        RECT 67.470000 179.100000 67.670000 179.300000 ;
        RECT 67.470000 179.500000 67.670000 179.700000 ;
        RECT 67.470000 179.900000 67.670000 180.100000 ;
        RECT 67.470000 180.300000 67.670000 180.500000 ;
        RECT 67.470000 180.700000 67.670000 180.900000 ;
        RECT 67.470000 181.100000 67.670000 181.300000 ;
        RECT 67.470000 181.505000 67.670000 181.705000 ;
        RECT 67.470000 181.910000 67.670000 182.110000 ;
        RECT 67.470000 182.315000 67.670000 182.515000 ;
        RECT 67.470000 182.720000 67.670000 182.920000 ;
        RECT 67.470000 183.125000 67.670000 183.325000 ;
        RECT 67.470000 183.530000 67.670000 183.730000 ;
        RECT 67.470000 183.935000 67.670000 184.135000 ;
        RECT 67.470000 184.340000 67.670000 184.540000 ;
        RECT 67.470000 184.745000 67.670000 184.945000 ;
        RECT 67.470000 185.150000 67.670000 185.350000 ;
        RECT 67.470000 185.555000 67.670000 185.755000 ;
        RECT 67.470000 185.960000 67.670000 186.160000 ;
        RECT 67.470000 186.365000 67.670000 186.565000 ;
        RECT 67.470000 186.770000 67.670000 186.970000 ;
        RECT 67.470000 187.175000 67.670000 187.375000 ;
        RECT 67.470000 187.580000 67.670000 187.780000 ;
        RECT 67.470000 187.985000 67.670000 188.185000 ;
        RECT 67.470000 188.390000 67.670000 188.590000 ;
        RECT 67.470000 188.795000 67.670000 188.995000 ;
        RECT 67.470000 189.200000 67.670000 189.400000 ;
        RECT 67.470000 189.605000 67.670000 189.805000 ;
        RECT 67.470000 190.010000 67.670000 190.210000 ;
        RECT 67.470000 190.415000 67.670000 190.615000 ;
        RECT 67.470000 190.820000 67.670000 191.020000 ;
        RECT 67.470000 191.225000 67.670000 191.425000 ;
        RECT 67.470000 191.630000 67.670000 191.830000 ;
        RECT 67.470000 192.035000 67.670000 192.235000 ;
        RECT 67.470000 192.440000 67.670000 192.640000 ;
        RECT 67.470000 192.845000 67.670000 193.045000 ;
        RECT 67.470000 193.250000 67.670000 193.450000 ;
        RECT 67.470000 193.655000 67.670000 193.855000 ;
        RECT 67.470000 194.060000 67.670000 194.260000 ;
        RECT 67.470000 194.465000 67.670000 194.665000 ;
        RECT 67.470000 194.870000 67.670000 195.070000 ;
        RECT 67.470000 195.275000 67.670000 195.475000 ;
        RECT 67.470000 195.680000 67.670000 195.880000 ;
        RECT 67.470000 196.085000 67.670000 196.285000 ;
        RECT 67.470000 196.490000 67.670000 196.690000 ;
        RECT 67.470000 196.895000 67.670000 197.095000 ;
        RECT 67.470000 197.300000 67.670000 197.500000 ;
        RECT 67.470000 197.705000 67.670000 197.905000 ;
        RECT 67.520000  23.910000 67.720000  24.110000 ;
        RECT 67.520000  24.340000 67.720000  24.540000 ;
        RECT 67.520000  24.770000 67.720000  24.970000 ;
        RECT 67.520000  25.200000 67.720000  25.400000 ;
        RECT 67.520000  25.630000 67.720000  25.830000 ;
        RECT 67.520000  26.060000 67.720000  26.260000 ;
        RECT 67.520000  26.490000 67.720000  26.690000 ;
        RECT 67.520000  26.920000 67.720000  27.120000 ;
        RECT 67.520000  27.350000 67.720000  27.550000 ;
        RECT 67.520000  27.780000 67.720000  27.980000 ;
        RECT 67.520000  28.210000 67.720000  28.410000 ;
        RECT 67.880000 173.900000 68.080000 174.100000 ;
        RECT 67.880000 174.300000 68.080000 174.500000 ;
        RECT 67.880000 174.700000 68.080000 174.900000 ;
        RECT 67.880000 175.100000 68.080000 175.300000 ;
        RECT 67.880000 175.500000 68.080000 175.700000 ;
        RECT 67.880000 175.900000 68.080000 176.100000 ;
        RECT 67.880000 176.300000 68.080000 176.500000 ;
        RECT 67.880000 176.700000 68.080000 176.900000 ;
        RECT 67.880000 177.100000 68.080000 177.300000 ;
        RECT 67.880000 177.500000 68.080000 177.700000 ;
        RECT 67.880000 177.900000 68.080000 178.100000 ;
        RECT 67.880000 178.300000 68.080000 178.500000 ;
        RECT 67.880000 178.700000 68.080000 178.900000 ;
        RECT 67.880000 179.100000 68.080000 179.300000 ;
        RECT 67.880000 179.500000 68.080000 179.700000 ;
        RECT 67.880000 179.900000 68.080000 180.100000 ;
        RECT 67.880000 180.300000 68.080000 180.500000 ;
        RECT 67.880000 180.700000 68.080000 180.900000 ;
        RECT 67.880000 181.100000 68.080000 181.300000 ;
        RECT 67.880000 181.505000 68.080000 181.705000 ;
        RECT 67.880000 181.910000 68.080000 182.110000 ;
        RECT 67.880000 182.315000 68.080000 182.515000 ;
        RECT 67.880000 182.720000 68.080000 182.920000 ;
        RECT 67.880000 183.125000 68.080000 183.325000 ;
        RECT 67.880000 183.530000 68.080000 183.730000 ;
        RECT 67.880000 183.935000 68.080000 184.135000 ;
        RECT 67.880000 184.340000 68.080000 184.540000 ;
        RECT 67.880000 184.745000 68.080000 184.945000 ;
        RECT 67.880000 185.150000 68.080000 185.350000 ;
        RECT 67.880000 185.555000 68.080000 185.755000 ;
        RECT 67.880000 185.960000 68.080000 186.160000 ;
        RECT 67.880000 186.365000 68.080000 186.565000 ;
        RECT 67.880000 186.770000 68.080000 186.970000 ;
        RECT 67.880000 187.175000 68.080000 187.375000 ;
        RECT 67.880000 187.580000 68.080000 187.780000 ;
        RECT 67.880000 187.985000 68.080000 188.185000 ;
        RECT 67.880000 188.390000 68.080000 188.590000 ;
        RECT 67.880000 188.795000 68.080000 188.995000 ;
        RECT 67.880000 189.200000 68.080000 189.400000 ;
        RECT 67.880000 189.605000 68.080000 189.805000 ;
        RECT 67.880000 190.010000 68.080000 190.210000 ;
        RECT 67.880000 190.415000 68.080000 190.615000 ;
        RECT 67.880000 190.820000 68.080000 191.020000 ;
        RECT 67.880000 191.225000 68.080000 191.425000 ;
        RECT 67.880000 191.630000 68.080000 191.830000 ;
        RECT 67.880000 192.035000 68.080000 192.235000 ;
        RECT 67.880000 192.440000 68.080000 192.640000 ;
        RECT 67.880000 192.845000 68.080000 193.045000 ;
        RECT 67.880000 193.250000 68.080000 193.450000 ;
        RECT 67.880000 193.655000 68.080000 193.855000 ;
        RECT 67.880000 194.060000 68.080000 194.260000 ;
        RECT 67.880000 194.465000 68.080000 194.665000 ;
        RECT 67.880000 194.870000 68.080000 195.070000 ;
        RECT 67.880000 195.275000 68.080000 195.475000 ;
        RECT 67.880000 195.680000 68.080000 195.880000 ;
        RECT 67.880000 196.085000 68.080000 196.285000 ;
        RECT 67.880000 196.490000 68.080000 196.690000 ;
        RECT 67.880000 196.895000 68.080000 197.095000 ;
        RECT 67.880000 197.300000 68.080000 197.500000 ;
        RECT 67.880000 197.705000 68.080000 197.905000 ;
        RECT 67.925000  23.910000 68.125000  24.110000 ;
        RECT 67.925000  24.340000 68.125000  24.540000 ;
        RECT 67.925000  24.770000 68.125000  24.970000 ;
        RECT 67.925000  25.200000 68.125000  25.400000 ;
        RECT 67.925000  25.630000 68.125000  25.830000 ;
        RECT 67.925000  26.060000 68.125000  26.260000 ;
        RECT 67.925000  26.490000 68.125000  26.690000 ;
        RECT 67.925000  26.920000 68.125000  27.120000 ;
        RECT 67.925000  27.350000 68.125000  27.550000 ;
        RECT 67.925000  27.780000 68.125000  27.980000 ;
        RECT 67.925000  28.210000 68.125000  28.410000 ;
        RECT 68.290000 173.900000 68.490000 174.100000 ;
        RECT 68.290000 174.300000 68.490000 174.500000 ;
        RECT 68.290000 174.700000 68.490000 174.900000 ;
        RECT 68.290000 175.100000 68.490000 175.300000 ;
        RECT 68.290000 175.500000 68.490000 175.700000 ;
        RECT 68.290000 175.900000 68.490000 176.100000 ;
        RECT 68.290000 176.300000 68.490000 176.500000 ;
        RECT 68.290000 176.700000 68.490000 176.900000 ;
        RECT 68.290000 177.100000 68.490000 177.300000 ;
        RECT 68.290000 177.500000 68.490000 177.700000 ;
        RECT 68.290000 177.900000 68.490000 178.100000 ;
        RECT 68.290000 178.300000 68.490000 178.500000 ;
        RECT 68.290000 178.700000 68.490000 178.900000 ;
        RECT 68.290000 179.100000 68.490000 179.300000 ;
        RECT 68.290000 179.500000 68.490000 179.700000 ;
        RECT 68.290000 179.900000 68.490000 180.100000 ;
        RECT 68.290000 180.300000 68.490000 180.500000 ;
        RECT 68.290000 180.700000 68.490000 180.900000 ;
        RECT 68.290000 181.100000 68.490000 181.300000 ;
        RECT 68.290000 181.505000 68.490000 181.705000 ;
        RECT 68.290000 181.910000 68.490000 182.110000 ;
        RECT 68.290000 182.315000 68.490000 182.515000 ;
        RECT 68.290000 182.720000 68.490000 182.920000 ;
        RECT 68.290000 183.125000 68.490000 183.325000 ;
        RECT 68.290000 183.530000 68.490000 183.730000 ;
        RECT 68.290000 183.935000 68.490000 184.135000 ;
        RECT 68.290000 184.340000 68.490000 184.540000 ;
        RECT 68.290000 184.745000 68.490000 184.945000 ;
        RECT 68.290000 185.150000 68.490000 185.350000 ;
        RECT 68.290000 185.555000 68.490000 185.755000 ;
        RECT 68.290000 185.960000 68.490000 186.160000 ;
        RECT 68.290000 186.365000 68.490000 186.565000 ;
        RECT 68.290000 186.770000 68.490000 186.970000 ;
        RECT 68.290000 187.175000 68.490000 187.375000 ;
        RECT 68.290000 187.580000 68.490000 187.780000 ;
        RECT 68.290000 187.985000 68.490000 188.185000 ;
        RECT 68.290000 188.390000 68.490000 188.590000 ;
        RECT 68.290000 188.795000 68.490000 188.995000 ;
        RECT 68.290000 189.200000 68.490000 189.400000 ;
        RECT 68.290000 189.605000 68.490000 189.805000 ;
        RECT 68.290000 190.010000 68.490000 190.210000 ;
        RECT 68.290000 190.415000 68.490000 190.615000 ;
        RECT 68.290000 190.820000 68.490000 191.020000 ;
        RECT 68.290000 191.225000 68.490000 191.425000 ;
        RECT 68.290000 191.630000 68.490000 191.830000 ;
        RECT 68.290000 192.035000 68.490000 192.235000 ;
        RECT 68.290000 192.440000 68.490000 192.640000 ;
        RECT 68.290000 192.845000 68.490000 193.045000 ;
        RECT 68.290000 193.250000 68.490000 193.450000 ;
        RECT 68.290000 193.655000 68.490000 193.855000 ;
        RECT 68.290000 194.060000 68.490000 194.260000 ;
        RECT 68.290000 194.465000 68.490000 194.665000 ;
        RECT 68.290000 194.870000 68.490000 195.070000 ;
        RECT 68.290000 195.275000 68.490000 195.475000 ;
        RECT 68.290000 195.680000 68.490000 195.880000 ;
        RECT 68.290000 196.085000 68.490000 196.285000 ;
        RECT 68.290000 196.490000 68.490000 196.690000 ;
        RECT 68.290000 196.895000 68.490000 197.095000 ;
        RECT 68.290000 197.300000 68.490000 197.500000 ;
        RECT 68.290000 197.705000 68.490000 197.905000 ;
        RECT 68.330000  23.910000 68.530000  24.110000 ;
        RECT 68.330000  24.340000 68.530000  24.540000 ;
        RECT 68.330000  24.770000 68.530000  24.970000 ;
        RECT 68.330000  25.200000 68.530000  25.400000 ;
        RECT 68.330000  25.630000 68.530000  25.830000 ;
        RECT 68.330000  26.060000 68.530000  26.260000 ;
        RECT 68.330000  26.490000 68.530000  26.690000 ;
        RECT 68.330000  26.920000 68.530000  27.120000 ;
        RECT 68.330000  27.350000 68.530000  27.550000 ;
        RECT 68.330000  27.780000 68.530000  27.980000 ;
        RECT 68.330000  28.210000 68.530000  28.410000 ;
        RECT 68.700000 173.900000 68.900000 174.100000 ;
        RECT 68.700000 174.300000 68.900000 174.500000 ;
        RECT 68.700000 174.700000 68.900000 174.900000 ;
        RECT 68.700000 175.100000 68.900000 175.300000 ;
        RECT 68.700000 175.500000 68.900000 175.700000 ;
        RECT 68.700000 175.900000 68.900000 176.100000 ;
        RECT 68.700000 176.300000 68.900000 176.500000 ;
        RECT 68.700000 176.700000 68.900000 176.900000 ;
        RECT 68.700000 177.100000 68.900000 177.300000 ;
        RECT 68.700000 177.500000 68.900000 177.700000 ;
        RECT 68.700000 177.900000 68.900000 178.100000 ;
        RECT 68.700000 178.300000 68.900000 178.500000 ;
        RECT 68.700000 178.700000 68.900000 178.900000 ;
        RECT 68.700000 179.100000 68.900000 179.300000 ;
        RECT 68.700000 179.500000 68.900000 179.700000 ;
        RECT 68.700000 179.900000 68.900000 180.100000 ;
        RECT 68.700000 180.300000 68.900000 180.500000 ;
        RECT 68.700000 180.700000 68.900000 180.900000 ;
        RECT 68.700000 181.100000 68.900000 181.300000 ;
        RECT 68.700000 181.505000 68.900000 181.705000 ;
        RECT 68.700000 181.910000 68.900000 182.110000 ;
        RECT 68.700000 182.315000 68.900000 182.515000 ;
        RECT 68.700000 182.720000 68.900000 182.920000 ;
        RECT 68.700000 183.125000 68.900000 183.325000 ;
        RECT 68.700000 183.530000 68.900000 183.730000 ;
        RECT 68.700000 183.935000 68.900000 184.135000 ;
        RECT 68.700000 184.340000 68.900000 184.540000 ;
        RECT 68.700000 184.745000 68.900000 184.945000 ;
        RECT 68.700000 185.150000 68.900000 185.350000 ;
        RECT 68.700000 185.555000 68.900000 185.755000 ;
        RECT 68.700000 185.960000 68.900000 186.160000 ;
        RECT 68.700000 186.365000 68.900000 186.565000 ;
        RECT 68.700000 186.770000 68.900000 186.970000 ;
        RECT 68.700000 187.175000 68.900000 187.375000 ;
        RECT 68.700000 187.580000 68.900000 187.780000 ;
        RECT 68.700000 187.985000 68.900000 188.185000 ;
        RECT 68.700000 188.390000 68.900000 188.590000 ;
        RECT 68.700000 188.795000 68.900000 188.995000 ;
        RECT 68.700000 189.200000 68.900000 189.400000 ;
        RECT 68.700000 189.605000 68.900000 189.805000 ;
        RECT 68.700000 190.010000 68.900000 190.210000 ;
        RECT 68.700000 190.415000 68.900000 190.615000 ;
        RECT 68.700000 190.820000 68.900000 191.020000 ;
        RECT 68.700000 191.225000 68.900000 191.425000 ;
        RECT 68.700000 191.630000 68.900000 191.830000 ;
        RECT 68.700000 192.035000 68.900000 192.235000 ;
        RECT 68.700000 192.440000 68.900000 192.640000 ;
        RECT 68.700000 192.845000 68.900000 193.045000 ;
        RECT 68.700000 193.250000 68.900000 193.450000 ;
        RECT 68.700000 193.655000 68.900000 193.855000 ;
        RECT 68.700000 194.060000 68.900000 194.260000 ;
        RECT 68.700000 194.465000 68.900000 194.665000 ;
        RECT 68.700000 194.870000 68.900000 195.070000 ;
        RECT 68.700000 195.275000 68.900000 195.475000 ;
        RECT 68.700000 195.680000 68.900000 195.880000 ;
        RECT 68.700000 196.085000 68.900000 196.285000 ;
        RECT 68.700000 196.490000 68.900000 196.690000 ;
        RECT 68.700000 196.895000 68.900000 197.095000 ;
        RECT 68.700000 197.300000 68.900000 197.500000 ;
        RECT 68.700000 197.705000 68.900000 197.905000 ;
        RECT 68.735000  23.910000 68.935000  24.110000 ;
        RECT 68.735000  24.340000 68.935000  24.540000 ;
        RECT 68.735000  24.770000 68.935000  24.970000 ;
        RECT 68.735000  25.200000 68.935000  25.400000 ;
        RECT 68.735000  25.630000 68.935000  25.830000 ;
        RECT 68.735000  26.060000 68.935000  26.260000 ;
        RECT 68.735000  26.490000 68.935000  26.690000 ;
        RECT 68.735000  26.920000 68.935000  27.120000 ;
        RECT 68.735000  27.350000 68.935000  27.550000 ;
        RECT 68.735000  27.780000 68.935000  27.980000 ;
        RECT 68.735000  28.210000 68.935000  28.410000 ;
        RECT 69.110000 173.900000 69.310000 174.100000 ;
        RECT 69.110000 174.300000 69.310000 174.500000 ;
        RECT 69.110000 174.700000 69.310000 174.900000 ;
        RECT 69.110000 175.100000 69.310000 175.300000 ;
        RECT 69.110000 175.500000 69.310000 175.700000 ;
        RECT 69.110000 175.900000 69.310000 176.100000 ;
        RECT 69.110000 176.300000 69.310000 176.500000 ;
        RECT 69.110000 176.700000 69.310000 176.900000 ;
        RECT 69.110000 177.100000 69.310000 177.300000 ;
        RECT 69.110000 177.500000 69.310000 177.700000 ;
        RECT 69.110000 177.900000 69.310000 178.100000 ;
        RECT 69.110000 178.300000 69.310000 178.500000 ;
        RECT 69.110000 178.700000 69.310000 178.900000 ;
        RECT 69.110000 179.100000 69.310000 179.300000 ;
        RECT 69.110000 179.500000 69.310000 179.700000 ;
        RECT 69.110000 179.900000 69.310000 180.100000 ;
        RECT 69.110000 180.300000 69.310000 180.500000 ;
        RECT 69.110000 180.700000 69.310000 180.900000 ;
        RECT 69.110000 181.100000 69.310000 181.300000 ;
        RECT 69.110000 181.505000 69.310000 181.705000 ;
        RECT 69.110000 181.910000 69.310000 182.110000 ;
        RECT 69.110000 182.315000 69.310000 182.515000 ;
        RECT 69.110000 182.720000 69.310000 182.920000 ;
        RECT 69.110000 183.125000 69.310000 183.325000 ;
        RECT 69.110000 183.530000 69.310000 183.730000 ;
        RECT 69.110000 183.935000 69.310000 184.135000 ;
        RECT 69.110000 184.340000 69.310000 184.540000 ;
        RECT 69.110000 184.745000 69.310000 184.945000 ;
        RECT 69.110000 185.150000 69.310000 185.350000 ;
        RECT 69.110000 185.555000 69.310000 185.755000 ;
        RECT 69.110000 185.960000 69.310000 186.160000 ;
        RECT 69.110000 186.365000 69.310000 186.565000 ;
        RECT 69.110000 186.770000 69.310000 186.970000 ;
        RECT 69.110000 187.175000 69.310000 187.375000 ;
        RECT 69.110000 187.580000 69.310000 187.780000 ;
        RECT 69.110000 187.985000 69.310000 188.185000 ;
        RECT 69.110000 188.390000 69.310000 188.590000 ;
        RECT 69.110000 188.795000 69.310000 188.995000 ;
        RECT 69.110000 189.200000 69.310000 189.400000 ;
        RECT 69.110000 189.605000 69.310000 189.805000 ;
        RECT 69.110000 190.010000 69.310000 190.210000 ;
        RECT 69.110000 190.415000 69.310000 190.615000 ;
        RECT 69.110000 190.820000 69.310000 191.020000 ;
        RECT 69.110000 191.225000 69.310000 191.425000 ;
        RECT 69.110000 191.630000 69.310000 191.830000 ;
        RECT 69.110000 192.035000 69.310000 192.235000 ;
        RECT 69.110000 192.440000 69.310000 192.640000 ;
        RECT 69.110000 192.845000 69.310000 193.045000 ;
        RECT 69.110000 193.250000 69.310000 193.450000 ;
        RECT 69.110000 193.655000 69.310000 193.855000 ;
        RECT 69.110000 194.060000 69.310000 194.260000 ;
        RECT 69.110000 194.465000 69.310000 194.665000 ;
        RECT 69.110000 194.870000 69.310000 195.070000 ;
        RECT 69.110000 195.275000 69.310000 195.475000 ;
        RECT 69.110000 195.680000 69.310000 195.880000 ;
        RECT 69.110000 196.085000 69.310000 196.285000 ;
        RECT 69.110000 196.490000 69.310000 196.690000 ;
        RECT 69.110000 196.895000 69.310000 197.095000 ;
        RECT 69.110000 197.300000 69.310000 197.500000 ;
        RECT 69.110000 197.705000 69.310000 197.905000 ;
        RECT 69.140000  23.910000 69.340000  24.110000 ;
        RECT 69.140000  24.340000 69.340000  24.540000 ;
        RECT 69.140000  24.770000 69.340000  24.970000 ;
        RECT 69.140000  25.200000 69.340000  25.400000 ;
        RECT 69.140000  25.630000 69.340000  25.830000 ;
        RECT 69.140000  26.060000 69.340000  26.260000 ;
        RECT 69.140000  26.490000 69.340000  26.690000 ;
        RECT 69.140000  26.920000 69.340000  27.120000 ;
        RECT 69.140000  27.350000 69.340000  27.550000 ;
        RECT 69.140000  27.780000 69.340000  27.980000 ;
        RECT 69.140000  28.210000 69.340000  28.410000 ;
        RECT 69.520000 173.900000 69.720000 174.100000 ;
        RECT 69.520000 174.300000 69.720000 174.500000 ;
        RECT 69.520000 174.700000 69.720000 174.900000 ;
        RECT 69.520000 175.100000 69.720000 175.300000 ;
        RECT 69.520000 175.500000 69.720000 175.700000 ;
        RECT 69.520000 175.900000 69.720000 176.100000 ;
        RECT 69.520000 176.300000 69.720000 176.500000 ;
        RECT 69.520000 176.700000 69.720000 176.900000 ;
        RECT 69.520000 177.100000 69.720000 177.300000 ;
        RECT 69.520000 177.500000 69.720000 177.700000 ;
        RECT 69.520000 177.900000 69.720000 178.100000 ;
        RECT 69.520000 178.300000 69.720000 178.500000 ;
        RECT 69.520000 178.700000 69.720000 178.900000 ;
        RECT 69.520000 179.100000 69.720000 179.300000 ;
        RECT 69.520000 179.500000 69.720000 179.700000 ;
        RECT 69.520000 179.900000 69.720000 180.100000 ;
        RECT 69.520000 180.300000 69.720000 180.500000 ;
        RECT 69.520000 180.700000 69.720000 180.900000 ;
        RECT 69.520000 181.100000 69.720000 181.300000 ;
        RECT 69.520000 181.505000 69.720000 181.705000 ;
        RECT 69.520000 181.910000 69.720000 182.110000 ;
        RECT 69.520000 182.315000 69.720000 182.515000 ;
        RECT 69.520000 182.720000 69.720000 182.920000 ;
        RECT 69.520000 183.125000 69.720000 183.325000 ;
        RECT 69.520000 183.530000 69.720000 183.730000 ;
        RECT 69.520000 183.935000 69.720000 184.135000 ;
        RECT 69.520000 184.340000 69.720000 184.540000 ;
        RECT 69.520000 184.745000 69.720000 184.945000 ;
        RECT 69.520000 185.150000 69.720000 185.350000 ;
        RECT 69.520000 185.555000 69.720000 185.755000 ;
        RECT 69.520000 185.960000 69.720000 186.160000 ;
        RECT 69.520000 186.365000 69.720000 186.565000 ;
        RECT 69.520000 186.770000 69.720000 186.970000 ;
        RECT 69.520000 187.175000 69.720000 187.375000 ;
        RECT 69.520000 187.580000 69.720000 187.780000 ;
        RECT 69.520000 187.985000 69.720000 188.185000 ;
        RECT 69.520000 188.390000 69.720000 188.590000 ;
        RECT 69.520000 188.795000 69.720000 188.995000 ;
        RECT 69.520000 189.200000 69.720000 189.400000 ;
        RECT 69.520000 189.605000 69.720000 189.805000 ;
        RECT 69.520000 190.010000 69.720000 190.210000 ;
        RECT 69.520000 190.415000 69.720000 190.615000 ;
        RECT 69.520000 190.820000 69.720000 191.020000 ;
        RECT 69.520000 191.225000 69.720000 191.425000 ;
        RECT 69.520000 191.630000 69.720000 191.830000 ;
        RECT 69.520000 192.035000 69.720000 192.235000 ;
        RECT 69.520000 192.440000 69.720000 192.640000 ;
        RECT 69.520000 192.845000 69.720000 193.045000 ;
        RECT 69.520000 193.250000 69.720000 193.450000 ;
        RECT 69.520000 193.655000 69.720000 193.855000 ;
        RECT 69.520000 194.060000 69.720000 194.260000 ;
        RECT 69.520000 194.465000 69.720000 194.665000 ;
        RECT 69.520000 194.870000 69.720000 195.070000 ;
        RECT 69.520000 195.275000 69.720000 195.475000 ;
        RECT 69.520000 195.680000 69.720000 195.880000 ;
        RECT 69.520000 196.085000 69.720000 196.285000 ;
        RECT 69.520000 196.490000 69.720000 196.690000 ;
        RECT 69.520000 196.895000 69.720000 197.095000 ;
        RECT 69.520000 197.300000 69.720000 197.500000 ;
        RECT 69.520000 197.705000 69.720000 197.905000 ;
        RECT 69.545000  23.910000 69.745000  24.110000 ;
        RECT 69.545000  24.340000 69.745000  24.540000 ;
        RECT 69.545000  24.770000 69.745000  24.970000 ;
        RECT 69.545000  25.200000 69.745000  25.400000 ;
        RECT 69.545000  25.630000 69.745000  25.830000 ;
        RECT 69.545000  26.060000 69.745000  26.260000 ;
        RECT 69.545000  26.490000 69.745000  26.690000 ;
        RECT 69.545000  26.920000 69.745000  27.120000 ;
        RECT 69.545000  27.350000 69.745000  27.550000 ;
        RECT 69.545000  27.780000 69.745000  27.980000 ;
        RECT 69.545000  28.210000 69.745000  28.410000 ;
        RECT 69.930000 173.900000 70.130000 174.100000 ;
        RECT 69.930000 174.300000 70.130000 174.500000 ;
        RECT 69.930000 174.700000 70.130000 174.900000 ;
        RECT 69.930000 175.100000 70.130000 175.300000 ;
        RECT 69.930000 175.500000 70.130000 175.700000 ;
        RECT 69.930000 175.900000 70.130000 176.100000 ;
        RECT 69.930000 176.300000 70.130000 176.500000 ;
        RECT 69.930000 176.700000 70.130000 176.900000 ;
        RECT 69.930000 177.100000 70.130000 177.300000 ;
        RECT 69.930000 177.500000 70.130000 177.700000 ;
        RECT 69.930000 177.900000 70.130000 178.100000 ;
        RECT 69.930000 178.300000 70.130000 178.500000 ;
        RECT 69.930000 178.700000 70.130000 178.900000 ;
        RECT 69.930000 179.100000 70.130000 179.300000 ;
        RECT 69.930000 179.500000 70.130000 179.700000 ;
        RECT 69.930000 179.900000 70.130000 180.100000 ;
        RECT 69.930000 180.300000 70.130000 180.500000 ;
        RECT 69.930000 180.700000 70.130000 180.900000 ;
        RECT 69.930000 181.100000 70.130000 181.300000 ;
        RECT 69.930000 181.505000 70.130000 181.705000 ;
        RECT 69.930000 181.910000 70.130000 182.110000 ;
        RECT 69.930000 182.315000 70.130000 182.515000 ;
        RECT 69.930000 182.720000 70.130000 182.920000 ;
        RECT 69.930000 183.125000 70.130000 183.325000 ;
        RECT 69.930000 183.530000 70.130000 183.730000 ;
        RECT 69.930000 183.935000 70.130000 184.135000 ;
        RECT 69.930000 184.340000 70.130000 184.540000 ;
        RECT 69.930000 184.745000 70.130000 184.945000 ;
        RECT 69.930000 185.150000 70.130000 185.350000 ;
        RECT 69.930000 185.555000 70.130000 185.755000 ;
        RECT 69.930000 185.960000 70.130000 186.160000 ;
        RECT 69.930000 186.365000 70.130000 186.565000 ;
        RECT 69.930000 186.770000 70.130000 186.970000 ;
        RECT 69.930000 187.175000 70.130000 187.375000 ;
        RECT 69.930000 187.580000 70.130000 187.780000 ;
        RECT 69.930000 187.985000 70.130000 188.185000 ;
        RECT 69.930000 188.390000 70.130000 188.590000 ;
        RECT 69.930000 188.795000 70.130000 188.995000 ;
        RECT 69.930000 189.200000 70.130000 189.400000 ;
        RECT 69.930000 189.605000 70.130000 189.805000 ;
        RECT 69.930000 190.010000 70.130000 190.210000 ;
        RECT 69.930000 190.415000 70.130000 190.615000 ;
        RECT 69.930000 190.820000 70.130000 191.020000 ;
        RECT 69.930000 191.225000 70.130000 191.425000 ;
        RECT 69.930000 191.630000 70.130000 191.830000 ;
        RECT 69.930000 192.035000 70.130000 192.235000 ;
        RECT 69.930000 192.440000 70.130000 192.640000 ;
        RECT 69.930000 192.845000 70.130000 193.045000 ;
        RECT 69.930000 193.250000 70.130000 193.450000 ;
        RECT 69.930000 193.655000 70.130000 193.855000 ;
        RECT 69.930000 194.060000 70.130000 194.260000 ;
        RECT 69.930000 194.465000 70.130000 194.665000 ;
        RECT 69.930000 194.870000 70.130000 195.070000 ;
        RECT 69.930000 195.275000 70.130000 195.475000 ;
        RECT 69.930000 195.680000 70.130000 195.880000 ;
        RECT 69.930000 196.085000 70.130000 196.285000 ;
        RECT 69.930000 196.490000 70.130000 196.690000 ;
        RECT 69.930000 196.895000 70.130000 197.095000 ;
        RECT 69.930000 197.300000 70.130000 197.500000 ;
        RECT 69.930000 197.705000 70.130000 197.905000 ;
        RECT 69.950000  23.910000 70.150000  24.110000 ;
        RECT 69.950000  24.340000 70.150000  24.540000 ;
        RECT 69.950000  24.770000 70.150000  24.970000 ;
        RECT 69.950000  25.200000 70.150000  25.400000 ;
        RECT 69.950000  25.630000 70.150000  25.830000 ;
        RECT 69.950000  26.060000 70.150000  26.260000 ;
        RECT 69.950000  26.490000 70.150000  26.690000 ;
        RECT 69.950000  26.920000 70.150000  27.120000 ;
        RECT 69.950000  27.350000 70.150000  27.550000 ;
        RECT 69.950000  27.780000 70.150000  27.980000 ;
        RECT 69.950000  28.210000 70.150000  28.410000 ;
        RECT 70.340000 173.900000 70.540000 174.100000 ;
        RECT 70.340000 174.300000 70.540000 174.500000 ;
        RECT 70.340000 174.700000 70.540000 174.900000 ;
        RECT 70.340000 175.100000 70.540000 175.300000 ;
        RECT 70.340000 175.500000 70.540000 175.700000 ;
        RECT 70.340000 175.900000 70.540000 176.100000 ;
        RECT 70.340000 176.300000 70.540000 176.500000 ;
        RECT 70.340000 176.700000 70.540000 176.900000 ;
        RECT 70.340000 177.100000 70.540000 177.300000 ;
        RECT 70.340000 177.500000 70.540000 177.700000 ;
        RECT 70.340000 177.900000 70.540000 178.100000 ;
        RECT 70.340000 178.300000 70.540000 178.500000 ;
        RECT 70.340000 178.700000 70.540000 178.900000 ;
        RECT 70.340000 179.100000 70.540000 179.300000 ;
        RECT 70.340000 179.500000 70.540000 179.700000 ;
        RECT 70.340000 179.900000 70.540000 180.100000 ;
        RECT 70.340000 180.300000 70.540000 180.500000 ;
        RECT 70.340000 180.700000 70.540000 180.900000 ;
        RECT 70.340000 181.100000 70.540000 181.300000 ;
        RECT 70.340000 181.505000 70.540000 181.705000 ;
        RECT 70.340000 181.910000 70.540000 182.110000 ;
        RECT 70.340000 182.315000 70.540000 182.515000 ;
        RECT 70.340000 182.720000 70.540000 182.920000 ;
        RECT 70.340000 183.125000 70.540000 183.325000 ;
        RECT 70.340000 183.530000 70.540000 183.730000 ;
        RECT 70.340000 183.935000 70.540000 184.135000 ;
        RECT 70.340000 184.340000 70.540000 184.540000 ;
        RECT 70.340000 184.745000 70.540000 184.945000 ;
        RECT 70.340000 185.150000 70.540000 185.350000 ;
        RECT 70.340000 185.555000 70.540000 185.755000 ;
        RECT 70.340000 185.960000 70.540000 186.160000 ;
        RECT 70.340000 186.365000 70.540000 186.565000 ;
        RECT 70.340000 186.770000 70.540000 186.970000 ;
        RECT 70.340000 187.175000 70.540000 187.375000 ;
        RECT 70.340000 187.580000 70.540000 187.780000 ;
        RECT 70.340000 187.985000 70.540000 188.185000 ;
        RECT 70.340000 188.390000 70.540000 188.590000 ;
        RECT 70.340000 188.795000 70.540000 188.995000 ;
        RECT 70.340000 189.200000 70.540000 189.400000 ;
        RECT 70.340000 189.605000 70.540000 189.805000 ;
        RECT 70.340000 190.010000 70.540000 190.210000 ;
        RECT 70.340000 190.415000 70.540000 190.615000 ;
        RECT 70.340000 190.820000 70.540000 191.020000 ;
        RECT 70.340000 191.225000 70.540000 191.425000 ;
        RECT 70.340000 191.630000 70.540000 191.830000 ;
        RECT 70.340000 192.035000 70.540000 192.235000 ;
        RECT 70.340000 192.440000 70.540000 192.640000 ;
        RECT 70.340000 192.845000 70.540000 193.045000 ;
        RECT 70.340000 193.250000 70.540000 193.450000 ;
        RECT 70.340000 193.655000 70.540000 193.855000 ;
        RECT 70.340000 194.060000 70.540000 194.260000 ;
        RECT 70.340000 194.465000 70.540000 194.665000 ;
        RECT 70.340000 194.870000 70.540000 195.070000 ;
        RECT 70.340000 195.275000 70.540000 195.475000 ;
        RECT 70.340000 195.680000 70.540000 195.880000 ;
        RECT 70.340000 196.085000 70.540000 196.285000 ;
        RECT 70.340000 196.490000 70.540000 196.690000 ;
        RECT 70.340000 196.895000 70.540000 197.095000 ;
        RECT 70.340000 197.300000 70.540000 197.500000 ;
        RECT 70.340000 197.705000 70.540000 197.905000 ;
        RECT 70.355000  23.910000 70.555000  24.110000 ;
        RECT 70.355000  24.340000 70.555000  24.540000 ;
        RECT 70.355000  24.770000 70.555000  24.970000 ;
        RECT 70.355000  25.200000 70.555000  25.400000 ;
        RECT 70.355000  25.630000 70.555000  25.830000 ;
        RECT 70.355000  26.060000 70.555000  26.260000 ;
        RECT 70.355000  26.490000 70.555000  26.690000 ;
        RECT 70.355000  26.920000 70.555000  27.120000 ;
        RECT 70.355000  27.350000 70.555000  27.550000 ;
        RECT 70.355000  27.780000 70.555000  27.980000 ;
        RECT 70.355000  28.210000 70.555000  28.410000 ;
        RECT 70.750000 173.900000 70.950000 174.100000 ;
        RECT 70.750000 174.300000 70.950000 174.500000 ;
        RECT 70.750000 174.700000 70.950000 174.900000 ;
        RECT 70.750000 175.100000 70.950000 175.300000 ;
        RECT 70.750000 175.500000 70.950000 175.700000 ;
        RECT 70.750000 175.900000 70.950000 176.100000 ;
        RECT 70.750000 176.300000 70.950000 176.500000 ;
        RECT 70.750000 176.700000 70.950000 176.900000 ;
        RECT 70.750000 177.100000 70.950000 177.300000 ;
        RECT 70.750000 177.500000 70.950000 177.700000 ;
        RECT 70.750000 177.900000 70.950000 178.100000 ;
        RECT 70.750000 178.300000 70.950000 178.500000 ;
        RECT 70.750000 178.700000 70.950000 178.900000 ;
        RECT 70.750000 179.100000 70.950000 179.300000 ;
        RECT 70.750000 179.500000 70.950000 179.700000 ;
        RECT 70.750000 179.900000 70.950000 180.100000 ;
        RECT 70.750000 180.300000 70.950000 180.500000 ;
        RECT 70.750000 180.700000 70.950000 180.900000 ;
        RECT 70.750000 181.100000 70.950000 181.300000 ;
        RECT 70.750000 181.505000 70.950000 181.705000 ;
        RECT 70.750000 181.910000 70.950000 182.110000 ;
        RECT 70.750000 182.315000 70.950000 182.515000 ;
        RECT 70.750000 182.720000 70.950000 182.920000 ;
        RECT 70.750000 183.125000 70.950000 183.325000 ;
        RECT 70.750000 183.530000 70.950000 183.730000 ;
        RECT 70.750000 183.935000 70.950000 184.135000 ;
        RECT 70.750000 184.340000 70.950000 184.540000 ;
        RECT 70.750000 184.745000 70.950000 184.945000 ;
        RECT 70.750000 185.150000 70.950000 185.350000 ;
        RECT 70.750000 185.555000 70.950000 185.755000 ;
        RECT 70.750000 185.960000 70.950000 186.160000 ;
        RECT 70.750000 186.365000 70.950000 186.565000 ;
        RECT 70.750000 186.770000 70.950000 186.970000 ;
        RECT 70.750000 187.175000 70.950000 187.375000 ;
        RECT 70.750000 187.580000 70.950000 187.780000 ;
        RECT 70.750000 187.985000 70.950000 188.185000 ;
        RECT 70.750000 188.390000 70.950000 188.590000 ;
        RECT 70.750000 188.795000 70.950000 188.995000 ;
        RECT 70.750000 189.200000 70.950000 189.400000 ;
        RECT 70.750000 189.605000 70.950000 189.805000 ;
        RECT 70.750000 190.010000 70.950000 190.210000 ;
        RECT 70.750000 190.415000 70.950000 190.615000 ;
        RECT 70.750000 190.820000 70.950000 191.020000 ;
        RECT 70.750000 191.225000 70.950000 191.425000 ;
        RECT 70.750000 191.630000 70.950000 191.830000 ;
        RECT 70.750000 192.035000 70.950000 192.235000 ;
        RECT 70.750000 192.440000 70.950000 192.640000 ;
        RECT 70.750000 192.845000 70.950000 193.045000 ;
        RECT 70.750000 193.250000 70.950000 193.450000 ;
        RECT 70.750000 193.655000 70.950000 193.855000 ;
        RECT 70.750000 194.060000 70.950000 194.260000 ;
        RECT 70.750000 194.465000 70.950000 194.665000 ;
        RECT 70.750000 194.870000 70.950000 195.070000 ;
        RECT 70.750000 195.275000 70.950000 195.475000 ;
        RECT 70.750000 195.680000 70.950000 195.880000 ;
        RECT 70.750000 196.085000 70.950000 196.285000 ;
        RECT 70.750000 196.490000 70.950000 196.690000 ;
        RECT 70.750000 196.895000 70.950000 197.095000 ;
        RECT 70.750000 197.300000 70.950000 197.500000 ;
        RECT 70.750000 197.705000 70.950000 197.905000 ;
        RECT 70.760000  23.910000 70.960000  24.110000 ;
        RECT 70.760000  24.340000 70.960000  24.540000 ;
        RECT 70.760000  24.770000 70.960000  24.970000 ;
        RECT 70.760000  25.200000 70.960000  25.400000 ;
        RECT 70.760000  25.630000 70.960000  25.830000 ;
        RECT 70.760000  26.060000 70.960000  26.260000 ;
        RECT 70.760000  26.490000 70.960000  26.690000 ;
        RECT 70.760000  26.920000 70.960000  27.120000 ;
        RECT 70.760000  27.350000 70.960000  27.550000 ;
        RECT 70.760000  27.780000 70.960000  27.980000 ;
        RECT 70.760000  28.210000 70.960000  28.410000 ;
        RECT 71.160000 173.900000 71.360000 174.100000 ;
        RECT 71.160000 174.300000 71.360000 174.500000 ;
        RECT 71.160000 174.700000 71.360000 174.900000 ;
        RECT 71.160000 175.100000 71.360000 175.300000 ;
        RECT 71.160000 175.500000 71.360000 175.700000 ;
        RECT 71.160000 175.900000 71.360000 176.100000 ;
        RECT 71.160000 176.300000 71.360000 176.500000 ;
        RECT 71.160000 176.700000 71.360000 176.900000 ;
        RECT 71.160000 177.100000 71.360000 177.300000 ;
        RECT 71.160000 177.500000 71.360000 177.700000 ;
        RECT 71.160000 177.900000 71.360000 178.100000 ;
        RECT 71.160000 178.300000 71.360000 178.500000 ;
        RECT 71.160000 178.700000 71.360000 178.900000 ;
        RECT 71.160000 179.100000 71.360000 179.300000 ;
        RECT 71.160000 179.500000 71.360000 179.700000 ;
        RECT 71.160000 179.900000 71.360000 180.100000 ;
        RECT 71.160000 180.300000 71.360000 180.500000 ;
        RECT 71.160000 180.700000 71.360000 180.900000 ;
        RECT 71.160000 181.100000 71.360000 181.300000 ;
        RECT 71.160000 181.505000 71.360000 181.705000 ;
        RECT 71.160000 181.910000 71.360000 182.110000 ;
        RECT 71.160000 182.315000 71.360000 182.515000 ;
        RECT 71.160000 182.720000 71.360000 182.920000 ;
        RECT 71.160000 183.125000 71.360000 183.325000 ;
        RECT 71.160000 183.530000 71.360000 183.730000 ;
        RECT 71.160000 183.935000 71.360000 184.135000 ;
        RECT 71.160000 184.340000 71.360000 184.540000 ;
        RECT 71.160000 184.745000 71.360000 184.945000 ;
        RECT 71.160000 185.150000 71.360000 185.350000 ;
        RECT 71.160000 185.555000 71.360000 185.755000 ;
        RECT 71.160000 185.960000 71.360000 186.160000 ;
        RECT 71.160000 186.365000 71.360000 186.565000 ;
        RECT 71.160000 186.770000 71.360000 186.970000 ;
        RECT 71.160000 187.175000 71.360000 187.375000 ;
        RECT 71.160000 187.580000 71.360000 187.780000 ;
        RECT 71.160000 187.985000 71.360000 188.185000 ;
        RECT 71.160000 188.390000 71.360000 188.590000 ;
        RECT 71.160000 188.795000 71.360000 188.995000 ;
        RECT 71.160000 189.200000 71.360000 189.400000 ;
        RECT 71.160000 189.605000 71.360000 189.805000 ;
        RECT 71.160000 190.010000 71.360000 190.210000 ;
        RECT 71.160000 190.415000 71.360000 190.615000 ;
        RECT 71.160000 190.820000 71.360000 191.020000 ;
        RECT 71.160000 191.225000 71.360000 191.425000 ;
        RECT 71.160000 191.630000 71.360000 191.830000 ;
        RECT 71.160000 192.035000 71.360000 192.235000 ;
        RECT 71.160000 192.440000 71.360000 192.640000 ;
        RECT 71.160000 192.845000 71.360000 193.045000 ;
        RECT 71.160000 193.250000 71.360000 193.450000 ;
        RECT 71.160000 193.655000 71.360000 193.855000 ;
        RECT 71.160000 194.060000 71.360000 194.260000 ;
        RECT 71.160000 194.465000 71.360000 194.665000 ;
        RECT 71.160000 194.870000 71.360000 195.070000 ;
        RECT 71.160000 195.275000 71.360000 195.475000 ;
        RECT 71.160000 195.680000 71.360000 195.880000 ;
        RECT 71.160000 196.085000 71.360000 196.285000 ;
        RECT 71.160000 196.490000 71.360000 196.690000 ;
        RECT 71.160000 196.895000 71.360000 197.095000 ;
        RECT 71.160000 197.300000 71.360000 197.500000 ;
        RECT 71.160000 197.705000 71.360000 197.905000 ;
        RECT 71.165000  23.910000 71.365000  24.110000 ;
        RECT 71.165000  24.340000 71.365000  24.540000 ;
        RECT 71.165000  24.770000 71.365000  24.970000 ;
        RECT 71.165000  25.200000 71.365000  25.400000 ;
        RECT 71.165000  25.630000 71.365000  25.830000 ;
        RECT 71.165000  26.060000 71.365000  26.260000 ;
        RECT 71.165000  26.490000 71.365000  26.690000 ;
        RECT 71.165000  26.920000 71.365000  27.120000 ;
        RECT 71.165000  27.350000 71.365000  27.550000 ;
        RECT 71.165000  27.780000 71.365000  27.980000 ;
        RECT 71.165000  28.210000 71.365000  28.410000 ;
        RECT 71.570000  23.910000 71.770000  24.110000 ;
        RECT 71.570000  24.340000 71.770000  24.540000 ;
        RECT 71.570000  24.770000 71.770000  24.970000 ;
        RECT 71.570000  25.200000 71.770000  25.400000 ;
        RECT 71.570000  25.630000 71.770000  25.830000 ;
        RECT 71.570000  26.060000 71.770000  26.260000 ;
        RECT 71.570000  26.490000 71.770000  26.690000 ;
        RECT 71.570000  26.920000 71.770000  27.120000 ;
        RECT 71.570000  27.350000 71.770000  27.550000 ;
        RECT 71.570000  27.780000 71.770000  27.980000 ;
        RECT 71.570000  28.210000 71.770000  28.410000 ;
        RECT 71.570000 173.900000 71.770000 174.100000 ;
        RECT 71.570000 174.300000 71.770000 174.500000 ;
        RECT 71.570000 174.700000 71.770000 174.900000 ;
        RECT 71.570000 175.100000 71.770000 175.300000 ;
        RECT 71.570000 175.500000 71.770000 175.700000 ;
        RECT 71.570000 175.900000 71.770000 176.100000 ;
        RECT 71.570000 176.300000 71.770000 176.500000 ;
        RECT 71.570000 176.700000 71.770000 176.900000 ;
        RECT 71.570000 177.100000 71.770000 177.300000 ;
        RECT 71.570000 177.500000 71.770000 177.700000 ;
        RECT 71.570000 177.900000 71.770000 178.100000 ;
        RECT 71.570000 178.300000 71.770000 178.500000 ;
        RECT 71.570000 178.700000 71.770000 178.900000 ;
        RECT 71.570000 179.100000 71.770000 179.300000 ;
        RECT 71.570000 179.500000 71.770000 179.700000 ;
        RECT 71.570000 179.900000 71.770000 180.100000 ;
        RECT 71.570000 180.300000 71.770000 180.500000 ;
        RECT 71.570000 180.700000 71.770000 180.900000 ;
        RECT 71.570000 181.100000 71.770000 181.300000 ;
        RECT 71.570000 181.505000 71.770000 181.705000 ;
        RECT 71.570000 181.910000 71.770000 182.110000 ;
        RECT 71.570000 182.315000 71.770000 182.515000 ;
        RECT 71.570000 182.720000 71.770000 182.920000 ;
        RECT 71.570000 183.125000 71.770000 183.325000 ;
        RECT 71.570000 183.530000 71.770000 183.730000 ;
        RECT 71.570000 183.935000 71.770000 184.135000 ;
        RECT 71.570000 184.340000 71.770000 184.540000 ;
        RECT 71.570000 184.745000 71.770000 184.945000 ;
        RECT 71.570000 185.150000 71.770000 185.350000 ;
        RECT 71.570000 185.555000 71.770000 185.755000 ;
        RECT 71.570000 185.960000 71.770000 186.160000 ;
        RECT 71.570000 186.365000 71.770000 186.565000 ;
        RECT 71.570000 186.770000 71.770000 186.970000 ;
        RECT 71.570000 187.175000 71.770000 187.375000 ;
        RECT 71.570000 187.580000 71.770000 187.780000 ;
        RECT 71.570000 187.985000 71.770000 188.185000 ;
        RECT 71.570000 188.390000 71.770000 188.590000 ;
        RECT 71.570000 188.795000 71.770000 188.995000 ;
        RECT 71.570000 189.200000 71.770000 189.400000 ;
        RECT 71.570000 189.605000 71.770000 189.805000 ;
        RECT 71.570000 190.010000 71.770000 190.210000 ;
        RECT 71.570000 190.415000 71.770000 190.615000 ;
        RECT 71.570000 190.820000 71.770000 191.020000 ;
        RECT 71.570000 191.225000 71.770000 191.425000 ;
        RECT 71.570000 191.630000 71.770000 191.830000 ;
        RECT 71.570000 192.035000 71.770000 192.235000 ;
        RECT 71.570000 192.440000 71.770000 192.640000 ;
        RECT 71.570000 192.845000 71.770000 193.045000 ;
        RECT 71.570000 193.250000 71.770000 193.450000 ;
        RECT 71.570000 193.655000 71.770000 193.855000 ;
        RECT 71.570000 194.060000 71.770000 194.260000 ;
        RECT 71.570000 194.465000 71.770000 194.665000 ;
        RECT 71.570000 194.870000 71.770000 195.070000 ;
        RECT 71.570000 195.275000 71.770000 195.475000 ;
        RECT 71.570000 195.680000 71.770000 195.880000 ;
        RECT 71.570000 196.085000 71.770000 196.285000 ;
        RECT 71.570000 196.490000 71.770000 196.690000 ;
        RECT 71.570000 196.895000 71.770000 197.095000 ;
        RECT 71.570000 197.300000 71.770000 197.500000 ;
        RECT 71.570000 197.705000 71.770000 197.905000 ;
        RECT 71.975000  23.910000 72.175000  24.110000 ;
        RECT 71.975000  24.340000 72.175000  24.540000 ;
        RECT 71.975000  24.770000 72.175000  24.970000 ;
        RECT 71.975000  25.200000 72.175000  25.400000 ;
        RECT 71.975000  25.630000 72.175000  25.830000 ;
        RECT 71.975000  26.060000 72.175000  26.260000 ;
        RECT 71.975000  26.490000 72.175000  26.690000 ;
        RECT 71.975000  26.920000 72.175000  27.120000 ;
        RECT 71.975000  27.350000 72.175000  27.550000 ;
        RECT 71.975000  27.780000 72.175000  27.980000 ;
        RECT 71.975000  28.210000 72.175000  28.410000 ;
        RECT 71.980000 173.900000 72.180000 174.100000 ;
        RECT 71.980000 174.300000 72.180000 174.500000 ;
        RECT 71.980000 174.700000 72.180000 174.900000 ;
        RECT 71.980000 175.100000 72.180000 175.300000 ;
        RECT 71.980000 175.500000 72.180000 175.700000 ;
        RECT 71.980000 175.900000 72.180000 176.100000 ;
        RECT 71.980000 176.300000 72.180000 176.500000 ;
        RECT 71.980000 176.700000 72.180000 176.900000 ;
        RECT 71.980000 177.100000 72.180000 177.300000 ;
        RECT 71.980000 177.500000 72.180000 177.700000 ;
        RECT 71.980000 177.900000 72.180000 178.100000 ;
        RECT 71.980000 178.300000 72.180000 178.500000 ;
        RECT 71.980000 178.700000 72.180000 178.900000 ;
        RECT 71.980000 179.100000 72.180000 179.300000 ;
        RECT 71.980000 179.500000 72.180000 179.700000 ;
        RECT 71.980000 179.900000 72.180000 180.100000 ;
        RECT 71.980000 180.300000 72.180000 180.500000 ;
        RECT 71.980000 180.700000 72.180000 180.900000 ;
        RECT 71.980000 181.100000 72.180000 181.300000 ;
        RECT 71.980000 181.505000 72.180000 181.705000 ;
        RECT 71.980000 181.910000 72.180000 182.110000 ;
        RECT 71.980000 182.315000 72.180000 182.515000 ;
        RECT 71.980000 182.720000 72.180000 182.920000 ;
        RECT 71.980000 183.125000 72.180000 183.325000 ;
        RECT 71.980000 183.530000 72.180000 183.730000 ;
        RECT 71.980000 183.935000 72.180000 184.135000 ;
        RECT 71.980000 184.340000 72.180000 184.540000 ;
        RECT 71.980000 184.745000 72.180000 184.945000 ;
        RECT 71.980000 185.150000 72.180000 185.350000 ;
        RECT 71.980000 185.555000 72.180000 185.755000 ;
        RECT 71.980000 185.960000 72.180000 186.160000 ;
        RECT 71.980000 186.365000 72.180000 186.565000 ;
        RECT 71.980000 186.770000 72.180000 186.970000 ;
        RECT 71.980000 187.175000 72.180000 187.375000 ;
        RECT 71.980000 187.580000 72.180000 187.780000 ;
        RECT 71.980000 187.985000 72.180000 188.185000 ;
        RECT 71.980000 188.390000 72.180000 188.590000 ;
        RECT 71.980000 188.795000 72.180000 188.995000 ;
        RECT 71.980000 189.200000 72.180000 189.400000 ;
        RECT 71.980000 189.605000 72.180000 189.805000 ;
        RECT 71.980000 190.010000 72.180000 190.210000 ;
        RECT 71.980000 190.415000 72.180000 190.615000 ;
        RECT 71.980000 190.820000 72.180000 191.020000 ;
        RECT 71.980000 191.225000 72.180000 191.425000 ;
        RECT 71.980000 191.630000 72.180000 191.830000 ;
        RECT 71.980000 192.035000 72.180000 192.235000 ;
        RECT 71.980000 192.440000 72.180000 192.640000 ;
        RECT 71.980000 192.845000 72.180000 193.045000 ;
        RECT 71.980000 193.250000 72.180000 193.450000 ;
        RECT 71.980000 193.655000 72.180000 193.855000 ;
        RECT 71.980000 194.060000 72.180000 194.260000 ;
        RECT 71.980000 194.465000 72.180000 194.665000 ;
        RECT 71.980000 194.870000 72.180000 195.070000 ;
        RECT 71.980000 195.275000 72.180000 195.475000 ;
        RECT 71.980000 195.680000 72.180000 195.880000 ;
        RECT 71.980000 196.085000 72.180000 196.285000 ;
        RECT 71.980000 196.490000 72.180000 196.690000 ;
        RECT 71.980000 196.895000 72.180000 197.095000 ;
        RECT 71.980000 197.300000 72.180000 197.500000 ;
        RECT 71.980000 197.705000 72.180000 197.905000 ;
        RECT 72.380000  23.910000 72.580000  24.110000 ;
        RECT 72.380000  24.340000 72.580000  24.540000 ;
        RECT 72.380000  24.770000 72.580000  24.970000 ;
        RECT 72.380000  25.200000 72.580000  25.400000 ;
        RECT 72.380000  25.630000 72.580000  25.830000 ;
        RECT 72.380000  26.060000 72.580000  26.260000 ;
        RECT 72.380000  26.490000 72.580000  26.690000 ;
        RECT 72.380000  26.920000 72.580000  27.120000 ;
        RECT 72.380000  27.350000 72.580000  27.550000 ;
        RECT 72.380000  27.780000 72.580000  27.980000 ;
        RECT 72.380000  28.210000 72.580000  28.410000 ;
        RECT 72.390000 173.900000 72.590000 174.100000 ;
        RECT 72.390000 174.300000 72.590000 174.500000 ;
        RECT 72.390000 174.700000 72.590000 174.900000 ;
        RECT 72.390000 175.100000 72.590000 175.300000 ;
        RECT 72.390000 175.500000 72.590000 175.700000 ;
        RECT 72.390000 175.900000 72.590000 176.100000 ;
        RECT 72.390000 176.300000 72.590000 176.500000 ;
        RECT 72.390000 176.700000 72.590000 176.900000 ;
        RECT 72.390000 177.100000 72.590000 177.300000 ;
        RECT 72.390000 177.500000 72.590000 177.700000 ;
        RECT 72.390000 177.900000 72.590000 178.100000 ;
        RECT 72.390000 178.300000 72.590000 178.500000 ;
        RECT 72.390000 178.700000 72.590000 178.900000 ;
        RECT 72.390000 179.100000 72.590000 179.300000 ;
        RECT 72.390000 179.500000 72.590000 179.700000 ;
        RECT 72.390000 179.900000 72.590000 180.100000 ;
        RECT 72.390000 180.300000 72.590000 180.500000 ;
        RECT 72.390000 180.700000 72.590000 180.900000 ;
        RECT 72.390000 181.100000 72.590000 181.300000 ;
        RECT 72.390000 181.505000 72.590000 181.705000 ;
        RECT 72.390000 181.910000 72.590000 182.110000 ;
        RECT 72.390000 182.315000 72.590000 182.515000 ;
        RECT 72.390000 182.720000 72.590000 182.920000 ;
        RECT 72.390000 183.125000 72.590000 183.325000 ;
        RECT 72.390000 183.530000 72.590000 183.730000 ;
        RECT 72.390000 183.935000 72.590000 184.135000 ;
        RECT 72.390000 184.340000 72.590000 184.540000 ;
        RECT 72.390000 184.745000 72.590000 184.945000 ;
        RECT 72.390000 185.150000 72.590000 185.350000 ;
        RECT 72.390000 185.555000 72.590000 185.755000 ;
        RECT 72.390000 185.960000 72.590000 186.160000 ;
        RECT 72.390000 186.365000 72.590000 186.565000 ;
        RECT 72.390000 186.770000 72.590000 186.970000 ;
        RECT 72.390000 187.175000 72.590000 187.375000 ;
        RECT 72.390000 187.580000 72.590000 187.780000 ;
        RECT 72.390000 187.985000 72.590000 188.185000 ;
        RECT 72.390000 188.390000 72.590000 188.590000 ;
        RECT 72.390000 188.795000 72.590000 188.995000 ;
        RECT 72.390000 189.200000 72.590000 189.400000 ;
        RECT 72.390000 189.605000 72.590000 189.805000 ;
        RECT 72.390000 190.010000 72.590000 190.210000 ;
        RECT 72.390000 190.415000 72.590000 190.615000 ;
        RECT 72.390000 190.820000 72.590000 191.020000 ;
        RECT 72.390000 191.225000 72.590000 191.425000 ;
        RECT 72.390000 191.630000 72.590000 191.830000 ;
        RECT 72.390000 192.035000 72.590000 192.235000 ;
        RECT 72.390000 192.440000 72.590000 192.640000 ;
        RECT 72.390000 192.845000 72.590000 193.045000 ;
        RECT 72.390000 193.250000 72.590000 193.450000 ;
        RECT 72.390000 193.655000 72.590000 193.855000 ;
        RECT 72.390000 194.060000 72.590000 194.260000 ;
        RECT 72.390000 194.465000 72.590000 194.665000 ;
        RECT 72.390000 194.870000 72.590000 195.070000 ;
        RECT 72.390000 195.275000 72.590000 195.475000 ;
        RECT 72.390000 195.680000 72.590000 195.880000 ;
        RECT 72.390000 196.085000 72.590000 196.285000 ;
        RECT 72.390000 196.490000 72.590000 196.690000 ;
        RECT 72.390000 196.895000 72.590000 197.095000 ;
        RECT 72.390000 197.300000 72.590000 197.500000 ;
        RECT 72.390000 197.705000 72.590000 197.905000 ;
        RECT 72.785000  23.910000 72.985000  24.110000 ;
        RECT 72.785000  24.340000 72.985000  24.540000 ;
        RECT 72.785000  24.770000 72.985000  24.970000 ;
        RECT 72.785000  25.200000 72.985000  25.400000 ;
        RECT 72.785000  25.630000 72.985000  25.830000 ;
        RECT 72.785000  26.060000 72.985000  26.260000 ;
        RECT 72.785000  26.490000 72.985000  26.690000 ;
        RECT 72.785000  26.920000 72.985000  27.120000 ;
        RECT 72.785000  27.350000 72.985000  27.550000 ;
        RECT 72.785000  27.780000 72.985000  27.980000 ;
        RECT 72.785000  28.210000 72.985000  28.410000 ;
        RECT 72.800000 173.900000 73.000000 174.100000 ;
        RECT 72.800000 174.300000 73.000000 174.500000 ;
        RECT 72.800000 174.700000 73.000000 174.900000 ;
        RECT 72.800000 175.100000 73.000000 175.300000 ;
        RECT 72.800000 175.500000 73.000000 175.700000 ;
        RECT 72.800000 175.900000 73.000000 176.100000 ;
        RECT 72.800000 176.300000 73.000000 176.500000 ;
        RECT 72.800000 176.700000 73.000000 176.900000 ;
        RECT 72.800000 177.100000 73.000000 177.300000 ;
        RECT 72.800000 177.500000 73.000000 177.700000 ;
        RECT 72.800000 177.900000 73.000000 178.100000 ;
        RECT 72.800000 178.300000 73.000000 178.500000 ;
        RECT 72.800000 178.700000 73.000000 178.900000 ;
        RECT 72.800000 179.100000 73.000000 179.300000 ;
        RECT 72.800000 179.500000 73.000000 179.700000 ;
        RECT 72.800000 179.900000 73.000000 180.100000 ;
        RECT 72.800000 180.300000 73.000000 180.500000 ;
        RECT 72.800000 180.700000 73.000000 180.900000 ;
        RECT 72.800000 181.100000 73.000000 181.300000 ;
        RECT 72.800000 181.505000 73.000000 181.705000 ;
        RECT 72.800000 181.910000 73.000000 182.110000 ;
        RECT 72.800000 182.315000 73.000000 182.515000 ;
        RECT 72.800000 182.720000 73.000000 182.920000 ;
        RECT 72.800000 183.125000 73.000000 183.325000 ;
        RECT 72.800000 183.530000 73.000000 183.730000 ;
        RECT 72.800000 183.935000 73.000000 184.135000 ;
        RECT 72.800000 184.340000 73.000000 184.540000 ;
        RECT 72.800000 184.745000 73.000000 184.945000 ;
        RECT 72.800000 185.150000 73.000000 185.350000 ;
        RECT 72.800000 185.555000 73.000000 185.755000 ;
        RECT 72.800000 185.960000 73.000000 186.160000 ;
        RECT 72.800000 186.365000 73.000000 186.565000 ;
        RECT 72.800000 186.770000 73.000000 186.970000 ;
        RECT 72.800000 187.175000 73.000000 187.375000 ;
        RECT 72.800000 187.580000 73.000000 187.780000 ;
        RECT 72.800000 187.985000 73.000000 188.185000 ;
        RECT 72.800000 188.390000 73.000000 188.590000 ;
        RECT 72.800000 188.795000 73.000000 188.995000 ;
        RECT 72.800000 189.200000 73.000000 189.400000 ;
        RECT 72.800000 189.605000 73.000000 189.805000 ;
        RECT 72.800000 190.010000 73.000000 190.210000 ;
        RECT 72.800000 190.415000 73.000000 190.615000 ;
        RECT 72.800000 190.820000 73.000000 191.020000 ;
        RECT 72.800000 191.225000 73.000000 191.425000 ;
        RECT 72.800000 191.630000 73.000000 191.830000 ;
        RECT 72.800000 192.035000 73.000000 192.235000 ;
        RECT 72.800000 192.440000 73.000000 192.640000 ;
        RECT 72.800000 192.845000 73.000000 193.045000 ;
        RECT 72.800000 193.250000 73.000000 193.450000 ;
        RECT 72.800000 193.655000 73.000000 193.855000 ;
        RECT 72.800000 194.060000 73.000000 194.260000 ;
        RECT 72.800000 194.465000 73.000000 194.665000 ;
        RECT 72.800000 194.870000 73.000000 195.070000 ;
        RECT 72.800000 195.275000 73.000000 195.475000 ;
        RECT 72.800000 195.680000 73.000000 195.880000 ;
        RECT 72.800000 196.085000 73.000000 196.285000 ;
        RECT 72.800000 196.490000 73.000000 196.690000 ;
        RECT 72.800000 196.895000 73.000000 197.095000 ;
        RECT 72.800000 197.300000 73.000000 197.500000 ;
        RECT 72.800000 197.705000 73.000000 197.905000 ;
        RECT 73.190000  23.910000 73.390000  24.110000 ;
        RECT 73.190000  24.340000 73.390000  24.540000 ;
        RECT 73.190000  24.770000 73.390000  24.970000 ;
        RECT 73.190000  25.200000 73.390000  25.400000 ;
        RECT 73.190000  25.630000 73.390000  25.830000 ;
        RECT 73.190000  26.060000 73.390000  26.260000 ;
        RECT 73.190000  26.490000 73.390000  26.690000 ;
        RECT 73.190000  26.920000 73.390000  27.120000 ;
        RECT 73.190000  27.350000 73.390000  27.550000 ;
        RECT 73.190000  27.780000 73.390000  27.980000 ;
        RECT 73.190000  28.210000 73.390000  28.410000 ;
        RECT 73.210000 173.900000 73.410000 174.100000 ;
        RECT 73.210000 174.300000 73.410000 174.500000 ;
        RECT 73.210000 174.700000 73.410000 174.900000 ;
        RECT 73.210000 175.100000 73.410000 175.300000 ;
        RECT 73.210000 175.500000 73.410000 175.700000 ;
        RECT 73.210000 175.900000 73.410000 176.100000 ;
        RECT 73.210000 176.300000 73.410000 176.500000 ;
        RECT 73.210000 176.700000 73.410000 176.900000 ;
        RECT 73.210000 177.100000 73.410000 177.300000 ;
        RECT 73.210000 177.500000 73.410000 177.700000 ;
        RECT 73.210000 177.900000 73.410000 178.100000 ;
        RECT 73.210000 178.300000 73.410000 178.500000 ;
        RECT 73.210000 178.700000 73.410000 178.900000 ;
        RECT 73.210000 179.100000 73.410000 179.300000 ;
        RECT 73.210000 179.500000 73.410000 179.700000 ;
        RECT 73.210000 179.900000 73.410000 180.100000 ;
        RECT 73.210000 180.300000 73.410000 180.500000 ;
        RECT 73.210000 180.700000 73.410000 180.900000 ;
        RECT 73.210000 181.100000 73.410000 181.300000 ;
        RECT 73.210000 181.505000 73.410000 181.705000 ;
        RECT 73.210000 181.910000 73.410000 182.110000 ;
        RECT 73.210000 182.315000 73.410000 182.515000 ;
        RECT 73.210000 182.720000 73.410000 182.920000 ;
        RECT 73.210000 183.125000 73.410000 183.325000 ;
        RECT 73.210000 183.530000 73.410000 183.730000 ;
        RECT 73.210000 183.935000 73.410000 184.135000 ;
        RECT 73.210000 184.340000 73.410000 184.540000 ;
        RECT 73.210000 184.745000 73.410000 184.945000 ;
        RECT 73.210000 185.150000 73.410000 185.350000 ;
        RECT 73.210000 185.555000 73.410000 185.755000 ;
        RECT 73.210000 185.960000 73.410000 186.160000 ;
        RECT 73.210000 186.365000 73.410000 186.565000 ;
        RECT 73.210000 186.770000 73.410000 186.970000 ;
        RECT 73.210000 187.175000 73.410000 187.375000 ;
        RECT 73.210000 187.580000 73.410000 187.780000 ;
        RECT 73.210000 187.985000 73.410000 188.185000 ;
        RECT 73.210000 188.390000 73.410000 188.590000 ;
        RECT 73.210000 188.795000 73.410000 188.995000 ;
        RECT 73.210000 189.200000 73.410000 189.400000 ;
        RECT 73.210000 189.605000 73.410000 189.805000 ;
        RECT 73.210000 190.010000 73.410000 190.210000 ;
        RECT 73.210000 190.415000 73.410000 190.615000 ;
        RECT 73.210000 190.820000 73.410000 191.020000 ;
        RECT 73.210000 191.225000 73.410000 191.425000 ;
        RECT 73.210000 191.630000 73.410000 191.830000 ;
        RECT 73.210000 192.035000 73.410000 192.235000 ;
        RECT 73.210000 192.440000 73.410000 192.640000 ;
        RECT 73.210000 192.845000 73.410000 193.045000 ;
        RECT 73.210000 193.250000 73.410000 193.450000 ;
        RECT 73.210000 193.655000 73.410000 193.855000 ;
        RECT 73.210000 194.060000 73.410000 194.260000 ;
        RECT 73.210000 194.465000 73.410000 194.665000 ;
        RECT 73.210000 194.870000 73.410000 195.070000 ;
        RECT 73.210000 195.275000 73.410000 195.475000 ;
        RECT 73.210000 195.680000 73.410000 195.880000 ;
        RECT 73.210000 196.085000 73.410000 196.285000 ;
        RECT 73.210000 196.490000 73.410000 196.690000 ;
        RECT 73.210000 196.895000 73.410000 197.095000 ;
        RECT 73.210000 197.300000 73.410000 197.500000 ;
        RECT 73.210000 197.705000 73.410000 197.905000 ;
        RECT 73.595000  23.910000 73.795000  24.110000 ;
        RECT 73.595000  24.340000 73.795000  24.540000 ;
        RECT 73.595000  24.770000 73.795000  24.970000 ;
        RECT 73.595000  25.200000 73.795000  25.400000 ;
        RECT 73.595000  25.630000 73.795000  25.830000 ;
        RECT 73.595000  26.060000 73.795000  26.260000 ;
        RECT 73.595000  26.490000 73.795000  26.690000 ;
        RECT 73.595000  26.920000 73.795000  27.120000 ;
        RECT 73.595000  27.350000 73.795000  27.550000 ;
        RECT 73.595000  27.780000 73.795000  27.980000 ;
        RECT 73.595000  28.210000 73.795000  28.410000 ;
        RECT 73.620000 173.900000 73.820000 174.100000 ;
        RECT 73.620000 174.300000 73.820000 174.500000 ;
        RECT 73.620000 174.700000 73.820000 174.900000 ;
        RECT 73.620000 175.100000 73.820000 175.300000 ;
        RECT 73.620000 175.500000 73.820000 175.700000 ;
        RECT 73.620000 175.900000 73.820000 176.100000 ;
        RECT 73.620000 176.300000 73.820000 176.500000 ;
        RECT 73.620000 176.700000 73.820000 176.900000 ;
        RECT 73.620000 177.100000 73.820000 177.300000 ;
        RECT 73.620000 177.500000 73.820000 177.700000 ;
        RECT 73.620000 177.900000 73.820000 178.100000 ;
        RECT 73.620000 178.300000 73.820000 178.500000 ;
        RECT 73.620000 178.700000 73.820000 178.900000 ;
        RECT 73.620000 179.100000 73.820000 179.300000 ;
        RECT 73.620000 179.500000 73.820000 179.700000 ;
        RECT 73.620000 179.900000 73.820000 180.100000 ;
        RECT 73.620000 180.300000 73.820000 180.500000 ;
        RECT 73.620000 180.700000 73.820000 180.900000 ;
        RECT 73.620000 181.100000 73.820000 181.300000 ;
        RECT 73.620000 181.505000 73.820000 181.705000 ;
        RECT 73.620000 181.910000 73.820000 182.110000 ;
        RECT 73.620000 182.315000 73.820000 182.515000 ;
        RECT 73.620000 182.720000 73.820000 182.920000 ;
        RECT 73.620000 183.125000 73.820000 183.325000 ;
        RECT 73.620000 183.530000 73.820000 183.730000 ;
        RECT 73.620000 183.935000 73.820000 184.135000 ;
        RECT 73.620000 184.340000 73.820000 184.540000 ;
        RECT 73.620000 184.745000 73.820000 184.945000 ;
        RECT 73.620000 185.150000 73.820000 185.350000 ;
        RECT 73.620000 185.555000 73.820000 185.755000 ;
        RECT 73.620000 185.960000 73.820000 186.160000 ;
        RECT 73.620000 186.365000 73.820000 186.565000 ;
        RECT 73.620000 186.770000 73.820000 186.970000 ;
        RECT 73.620000 187.175000 73.820000 187.375000 ;
        RECT 73.620000 187.580000 73.820000 187.780000 ;
        RECT 73.620000 187.985000 73.820000 188.185000 ;
        RECT 73.620000 188.390000 73.820000 188.590000 ;
        RECT 73.620000 188.795000 73.820000 188.995000 ;
        RECT 73.620000 189.200000 73.820000 189.400000 ;
        RECT 73.620000 189.605000 73.820000 189.805000 ;
        RECT 73.620000 190.010000 73.820000 190.210000 ;
        RECT 73.620000 190.415000 73.820000 190.615000 ;
        RECT 73.620000 190.820000 73.820000 191.020000 ;
        RECT 73.620000 191.225000 73.820000 191.425000 ;
        RECT 73.620000 191.630000 73.820000 191.830000 ;
        RECT 73.620000 192.035000 73.820000 192.235000 ;
        RECT 73.620000 192.440000 73.820000 192.640000 ;
        RECT 73.620000 192.845000 73.820000 193.045000 ;
        RECT 73.620000 193.250000 73.820000 193.450000 ;
        RECT 73.620000 193.655000 73.820000 193.855000 ;
        RECT 73.620000 194.060000 73.820000 194.260000 ;
        RECT 73.620000 194.465000 73.820000 194.665000 ;
        RECT 73.620000 194.870000 73.820000 195.070000 ;
        RECT 73.620000 195.275000 73.820000 195.475000 ;
        RECT 73.620000 195.680000 73.820000 195.880000 ;
        RECT 73.620000 196.085000 73.820000 196.285000 ;
        RECT 73.620000 196.490000 73.820000 196.690000 ;
        RECT 73.620000 196.895000 73.820000 197.095000 ;
        RECT 73.620000 197.300000 73.820000 197.500000 ;
        RECT 73.620000 197.705000 73.820000 197.905000 ;
        RECT 74.000000  23.910000 74.200000  24.110000 ;
        RECT 74.000000  24.340000 74.200000  24.540000 ;
        RECT 74.000000  24.770000 74.200000  24.970000 ;
        RECT 74.000000  25.200000 74.200000  25.400000 ;
        RECT 74.000000  25.630000 74.200000  25.830000 ;
        RECT 74.000000  26.060000 74.200000  26.260000 ;
        RECT 74.000000  26.490000 74.200000  26.690000 ;
        RECT 74.000000  26.920000 74.200000  27.120000 ;
        RECT 74.000000  27.350000 74.200000  27.550000 ;
        RECT 74.000000  27.780000 74.200000  27.980000 ;
        RECT 74.000000  28.210000 74.200000  28.410000 ;
        RECT 74.030000 173.900000 74.230000 174.100000 ;
        RECT 74.030000 174.300000 74.230000 174.500000 ;
        RECT 74.030000 174.700000 74.230000 174.900000 ;
        RECT 74.030000 175.100000 74.230000 175.300000 ;
        RECT 74.030000 175.500000 74.230000 175.700000 ;
        RECT 74.030000 175.900000 74.230000 176.100000 ;
        RECT 74.030000 176.300000 74.230000 176.500000 ;
        RECT 74.030000 176.700000 74.230000 176.900000 ;
        RECT 74.030000 177.100000 74.230000 177.300000 ;
        RECT 74.030000 177.500000 74.230000 177.700000 ;
        RECT 74.030000 177.900000 74.230000 178.100000 ;
        RECT 74.030000 178.300000 74.230000 178.500000 ;
        RECT 74.030000 178.700000 74.230000 178.900000 ;
        RECT 74.030000 179.100000 74.230000 179.300000 ;
        RECT 74.030000 179.500000 74.230000 179.700000 ;
        RECT 74.030000 179.900000 74.230000 180.100000 ;
        RECT 74.030000 180.300000 74.230000 180.500000 ;
        RECT 74.030000 180.700000 74.230000 180.900000 ;
        RECT 74.030000 181.100000 74.230000 181.300000 ;
        RECT 74.030000 181.505000 74.230000 181.705000 ;
        RECT 74.030000 181.910000 74.230000 182.110000 ;
        RECT 74.030000 182.315000 74.230000 182.515000 ;
        RECT 74.030000 182.720000 74.230000 182.920000 ;
        RECT 74.030000 183.125000 74.230000 183.325000 ;
        RECT 74.030000 183.530000 74.230000 183.730000 ;
        RECT 74.030000 183.935000 74.230000 184.135000 ;
        RECT 74.030000 184.340000 74.230000 184.540000 ;
        RECT 74.030000 184.745000 74.230000 184.945000 ;
        RECT 74.030000 185.150000 74.230000 185.350000 ;
        RECT 74.030000 185.555000 74.230000 185.755000 ;
        RECT 74.030000 185.960000 74.230000 186.160000 ;
        RECT 74.030000 186.365000 74.230000 186.565000 ;
        RECT 74.030000 186.770000 74.230000 186.970000 ;
        RECT 74.030000 187.175000 74.230000 187.375000 ;
        RECT 74.030000 187.580000 74.230000 187.780000 ;
        RECT 74.030000 187.985000 74.230000 188.185000 ;
        RECT 74.030000 188.390000 74.230000 188.590000 ;
        RECT 74.030000 188.795000 74.230000 188.995000 ;
        RECT 74.030000 189.200000 74.230000 189.400000 ;
        RECT 74.030000 189.605000 74.230000 189.805000 ;
        RECT 74.030000 190.010000 74.230000 190.210000 ;
        RECT 74.030000 190.415000 74.230000 190.615000 ;
        RECT 74.030000 190.820000 74.230000 191.020000 ;
        RECT 74.030000 191.225000 74.230000 191.425000 ;
        RECT 74.030000 191.630000 74.230000 191.830000 ;
        RECT 74.030000 192.035000 74.230000 192.235000 ;
        RECT 74.030000 192.440000 74.230000 192.640000 ;
        RECT 74.030000 192.845000 74.230000 193.045000 ;
        RECT 74.030000 193.250000 74.230000 193.450000 ;
        RECT 74.030000 193.655000 74.230000 193.855000 ;
        RECT 74.030000 194.060000 74.230000 194.260000 ;
        RECT 74.030000 194.465000 74.230000 194.665000 ;
        RECT 74.030000 194.870000 74.230000 195.070000 ;
        RECT 74.030000 195.275000 74.230000 195.475000 ;
        RECT 74.030000 195.680000 74.230000 195.880000 ;
        RECT 74.030000 196.085000 74.230000 196.285000 ;
        RECT 74.030000 196.490000 74.230000 196.690000 ;
        RECT 74.030000 196.895000 74.230000 197.095000 ;
        RECT 74.030000 197.300000 74.230000 197.500000 ;
        RECT 74.030000 197.705000 74.230000 197.905000 ;
        RECT 74.440000 173.900000 74.640000 174.100000 ;
        RECT 74.440000 174.300000 74.640000 174.500000 ;
        RECT 74.440000 174.700000 74.640000 174.900000 ;
        RECT 74.440000 175.100000 74.640000 175.300000 ;
        RECT 74.440000 175.500000 74.640000 175.700000 ;
        RECT 74.440000 175.900000 74.640000 176.100000 ;
        RECT 74.440000 176.300000 74.640000 176.500000 ;
        RECT 74.440000 176.700000 74.640000 176.900000 ;
        RECT 74.440000 177.100000 74.640000 177.300000 ;
        RECT 74.440000 177.500000 74.640000 177.700000 ;
        RECT 74.440000 177.900000 74.640000 178.100000 ;
        RECT 74.440000 178.300000 74.640000 178.500000 ;
        RECT 74.440000 178.700000 74.640000 178.900000 ;
        RECT 74.440000 179.100000 74.640000 179.300000 ;
        RECT 74.440000 179.500000 74.640000 179.700000 ;
        RECT 74.440000 179.900000 74.640000 180.100000 ;
        RECT 74.440000 180.300000 74.640000 180.500000 ;
        RECT 74.440000 180.700000 74.640000 180.900000 ;
        RECT 74.440000 181.100000 74.640000 181.300000 ;
        RECT 74.440000 181.505000 74.640000 181.705000 ;
        RECT 74.440000 181.910000 74.640000 182.110000 ;
        RECT 74.440000 182.315000 74.640000 182.515000 ;
        RECT 74.440000 182.720000 74.640000 182.920000 ;
        RECT 74.440000 183.125000 74.640000 183.325000 ;
        RECT 74.440000 183.530000 74.640000 183.730000 ;
        RECT 74.440000 183.935000 74.640000 184.135000 ;
        RECT 74.440000 184.340000 74.640000 184.540000 ;
        RECT 74.440000 184.745000 74.640000 184.945000 ;
        RECT 74.440000 185.150000 74.640000 185.350000 ;
        RECT 74.440000 185.555000 74.640000 185.755000 ;
        RECT 74.440000 185.960000 74.640000 186.160000 ;
        RECT 74.440000 186.365000 74.640000 186.565000 ;
        RECT 74.440000 186.770000 74.640000 186.970000 ;
        RECT 74.440000 187.175000 74.640000 187.375000 ;
        RECT 74.440000 187.580000 74.640000 187.780000 ;
        RECT 74.440000 187.985000 74.640000 188.185000 ;
        RECT 74.440000 188.390000 74.640000 188.590000 ;
        RECT 74.440000 188.795000 74.640000 188.995000 ;
        RECT 74.440000 189.200000 74.640000 189.400000 ;
        RECT 74.440000 189.605000 74.640000 189.805000 ;
        RECT 74.440000 190.010000 74.640000 190.210000 ;
        RECT 74.440000 190.415000 74.640000 190.615000 ;
        RECT 74.440000 190.820000 74.640000 191.020000 ;
        RECT 74.440000 191.225000 74.640000 191.425000 ;
        RECT 74.440000 191.630000 74.640000 191.830000 ;
        RECT 74.440000 192.035000 74.640000 192.235000 ;
        RECT 74.440000 192.440000 74.640000 192.640000 ;
        RECT 74.440000 192.845000 74.640000 193.045000 ;
        RECT 74.440000 193.250000 74.640000 193.450000 ;
        RECT 74.440000 193.655000 74.640000 193.855000 ;
        RECT 74.440000 194.060000 74.640000 194.260000 ;
        RECT 74.440000 194.465000 74.640000 194.665000 ;
        RECT 74.440000 194.870000 74.640000 195.070000 ;
        RECT 74.440000 195.275000 74.640000 195.475000 ;
        RECT 74.440000 195.680000 74.640000 195.880000 ;
        RECT 74.440000 196.085000 74.640000 196.285000 ;
        RECT 74.440000 196.490000 74.640000 196.690000 ;
        RECT 74.440000 196.895000 74.640000 197.095000 ;
        RECT 74.440000 197.300000 74.640000 197.500000 ;
        RECT 74.440000 197.705000 74.640000 197.905000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.500000 56.240000 24.400000 60.680000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755000 56.240000 74.290000 60.680000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 56.235000 24.375000 60.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.780000 56.235000 75.000000 60.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 56.335000 1.270000 60.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 56.335000 75.000000 60.585000 ;
    END
    PORT
      LAYER via3 ;
        RECT  0.590000 56.310000  0.790000 56.510000 ;
        RECT  0.590000 56.720000  0.790000 56.920000 ;
        RECT  0.590000 57.130000  0.790000 57.330000 ;
        RECT  0.590000 57.540000  0.790000 57.740000 ;
        RECT  0.590000 57.950000  0.790000 58.150000 ;
        RECT  0.590000 58.360000  0.790000 58.560000 ;
        RECT  0.590000 58.770000  0.790000 58.970000 ;
        RECT  0.590000 59.180000  0.790000 59.380000 ;
        RECT  0.590000 59.590000  0.790000 59.790000 ;
        RECT  0.590000 60.000000  0.790000 60.200000 ;
        RECT  0.590000 60.410000  0.790000 60.610000 ;
        RECT  1.000000 56.310000  1.200000 56.510000 ;
        RECT  1.000000 56.720000  1.200000 56.920000 ;
        RECT  1.000000 57.130000  1.200000 57.330000 ;
        RECT  1.000000 57.540000  1.200000 57.740000 ;
        RECT  1.000000 57.950000  1.200000 58.150000 ;
        RECT  1.000000 58.360000  1.200000 58.560000 ;
        RECT  1.000000 58.770000  1.200000 58.970000 ;
        RECT  1.000000 59.180000  1.200000 59.380000 ;
        RECT  1.000000 59.590000  1.200000 59.790000 ;
        RECT  1.000000 60.000000  1.200000 60.200000 ;
        RECT  1.000000 60.410000  1.200000 60.610000 ;
        RECT  1.410000 56.310000  1.610000 56.510000 ;
        RECT  1.410000 56.720000  1.610000 56.920000 ;
        RECT  1.410000 57.130000  1.610000 57.330000 ;
        RECT  1.410000 57.540000  1.610000 57.740000 ;
        RECT  1.410000 57.950000  1.610000 58.150000 ;
        RECT  1.410000 58.360000  1.610000 58.560000 ;
        RECT  1.410000 58.770000  1.610000 58.970000 ;
        RECT  1.410000 59.180000  1.610000 59.380000 ;
        RECT  1.410000 59.590000  1.610000 59.790000 ;
        RECT  1.410000 60.000000  1.610000 60.200000 ;
        RECT  1.410000 60.410000  1.610000 60.610000 ;
        RECT  1.820000 56.310000  2.020000 56.510000 ;
        RECT  1.820000 56.720000  2.020000 56.920000 ;
        RECT  1.820000 57.130000  2.020000 57.330000 ;
        RECT  1.820000 57.540000  2.020000 57.740000 ;
        RECT  1.820000 57.950000  2.020000 58.150000 ;
        RECT  1.820000 58.360000  2.020000 58.560000 ;
        RECT  1.820000 58.770000  2.020000 58.970000 ;
        RECT  1.820000 59.180000  2.020000 59.380000 ;
        RECT  1.820000 59.590000  2.020000 59.790000 ;
        RECT  1.820000 60.000000  2.020000 60.200000 ;
        RECT  1.820000 60.410000  2.020000 60.610000 ;
        RECT  2.230000 56.310000  2.430000 56.510000 ;
        RECT  2.230000 56.720000  2.430000 56.920000 ;
        RECT  2.230000 57.130000  2.430000 57.330000 ;
        RECT  2.230000 57.540000  2.430000 57.740000 ;
        RECT  2.230000 57.950000  2.430000 58.150000 ;
        RECT  2.230000 58.360000  2.430000 58.560000 ;
        RECT  2.230000 58.770000  2.430000 58.970000 ;
        RECT  2.230000 59.180000  2.430000 59.380000 ;
        RECT  2.230000 59.590000  2.430000 59.790000 ;
        RECT  2.230000 60.000000  2.430000 60.200000 ;
        RECT  2.230000 60.410000  2.430000 60.610000 ;
        RECT  2.640000 56.310000  2.840000 56.510000 ;
        RECT  2.640000 56.720000  2.840000 56.920000 ;
        RECT  2.640000 57.130000  2.840000 57.330000 ;
        RECT  2.640000 57.540000  2.840000 57.740000 ;
        RECT  2.640000 57.950000  2.840000 58.150000 ;
        RECT  2.640000 58.360000  2.840000 58.560000 ;
        RECT  2.640000 58.770000  2.840000 58.970000 ;
        RECT  2.640000 59.180000  2.840000 59.380000 ;
        RECT  2.640000 59.590000  2.840000 59.790000 ;
        RECT  2.640000 60.000000  2.840000 60.200000 ;
        RECT  2.640000 60.410000  2.840000 60.610000 ;
        RECT  3.050000 56.310000  3.250000 56.510000 ;
        RECT  3.050000 56.720000  3.250000 56.920000 ;
        RECT  3.050000 57.130000  3.250000 57.330000 ;
        RECT  3.050000 57.540000  3.250000 57.740000 ;
        RECT  3.050000 57.950000  3.250000 58.150000 ;
        RECT  3.050000 58.360000  3.250000 58.560000 ;
        RECT  3.050000 58.770000  3.250000 58.970000 ;
        RECT  3.050000 59.180000  3.250000 59.380000 ;
        RECT  3.050000 59.590000  3.250000 59.790000 ;
        RECT  3.050000 60.000000  3.250000 60.200000 ;
        RECT  3.050000 60.410000  3.250000 60.610000 ;
        RECT  3.455000 56.310000  3.655000 56.510000 ;
        RECT  3.455000 56.720000  3.655000 56.920000 ;
        RECT  3.455000 57.130000  3.655000 57.330000 ;
        RECT  3.455000 57.540000  3.655000 57.740000 ;
        RECT  3.455000 57.950000  3.655000 58.150000 ;
        RECT  3.455000 58.360000  3.655000 58.560000 ;
        RECT  3.455000 58.770000  3.655000 58.970000 ;
        RECT  3.455000 59.180000  3.655000 59.380000 ;
        RECT  3.455000 59.590000  3.655000 59.790000 ;
        RECT  3.455000 60.000000  3.655000 60.200000 ;
        RECT  3.455000 60.410000  3.655000 60.610000 ;
        RECT  3.860000 56.310000  4.060000 56.510000 ;
        RECT  3.860000 56.720000  4.060000 56.920000 ;
        RECT  3.860000 57.130000  4.060000 57.330000 ;
        RECT  3.860000 57.540000  4.060000 57.740000 ;
        RECT  3.860000 57.950000  4.060000 58.150000 ;
        RECT  3.860000 58.360000  4.060000 58.560000 ;
        RECT  3.860000 58.770000  4.060000 58.970000 ;
        RECT  3.860000 59.180000  4.060000 59.380000 ;
        RECT  3.860000 59.590000  4.060000 59.790000 ;
        RECT  3.860000 60.000000  4.060000 60.200000 ;
        RECT  3.860000 60.410000  4.060000 60.610000 ;
        RECT  4.265000 56.310000  4.465000 56.510000 ;
        RECT  4.265000 56.720000  4.465000 56.920000 ;
        RECT  4.265000 57.130000  4.465000 57.330000 ;
        RECT  4.265000 57.540000  4.465000 57.740000 ;
        RECT  4.265000 57.950000  4.465000 58.150000 ;
        RECT  4.265000 58.360000  4.465000 58.560000 ;
        RECT  4.265000 58.770000  4.465000 58.970000 ;
        RECT  4.265000 59.180000  4.465000 59.380000 ;
        RECT  4.265000 59.590000  4.465000 59.790000 ;
        RECT  4.265000 60.000000  4.465000 60.200000 ;
        RECT  4.265000 60.410000  4.465000 60.610000 ;
        RECT  4.670000 56.310000  4.870000 56.510000 ;
        RECT  4.670000 56.720000  4.870000 56.920000 ;
        RECT  4.670000 57.130000  4.870000 57.330000 ;
        RECT  4.670000 57.540000  4.870000 57.740000 ;
        RECT  4.670000 57.950000  4.870000 58.150000 ;
        RECT  4.670000 58.360000  4.870000 58.560000 ;
        RECT  4.670000 58.770000  4.870000 58.970000 ;
        RECT  4.670000 59.180000  4.870000 59.380000 ;
        RECT  4.670000 59.590000  4.870000 59.790000 ;
        RECT  4.670000 60.000000  4.870000 60.200000 ;
        RECT  4.670000 60.410000  4.870000 60.610000 ;
        RECT  5.075000 56.310000  5.275000 56.510000 ;
        RECT  5.075000 56.720000  5.275000 56.920000 ;
        RECT  5.075000 57.130000  5.275000 57.330000 ;
        RECT  5.075000 57.540000  5.275000 57.740000 ;
        RECT  5.075000 57.950000  5.275000 58.150000 ;
        RECT  5.075000 58.360000  5.275000 58.560000 ;
        RECT  5.075000 58.770000  5.275000 58.970000 ;
        RECT  5.075000 59.180000  5.275000 59.380000 ;
        RECT  5.075000 59.590000  5.275000 59.790000 ;
        RECT  5.075000 60.000000  5.275000 60.200000 ;
        RECT  5.075000 60.410000  5.275000 60.610000 ;
        RECT  5.480000 56.310000  5.680000 56.510000 ;
        RECT  5.480000 56.720000  5.680000 56.920000 ;
        RECT  5.480000 57.130000  5.680000 57.330000 ;
        RECT  5.480000 57.540000  5.680000 57.740000 ;
        RECT  5.480000 57.950000  5.680000 58.150000 ;
        RECT  5.480000 58.360000  5.680000 58.560000 ;
        RECT  5.480000 58.770000  5.680000 58.970000 ;
        RECT  5.480000 59.180000  5.680000 59.380000 ;
        RECT  5.480000 59.590000  5.680000 59.790000 ;
        RECT  5.480000 60.000000  5.680000 60.200000 ;
        RECT  5.480000 60.410000  5.680000 60.610000 ;
        RECT  5.885000 56.310000  6.085000 56.510000 ;
        RECT  5.885000 56.720000  6.085000 56.920000 ;
        RECT  5.885000 57.130000  6.085000 57.330000 ;
        RECT  5.885000 57.540000  6.085000 57.740000 ;
        RECT  5.885000 57.950000  6.085000 58.150000 ;
        RECT  5.885000 58.360000  6.085000 58.560000 ;
        RECT  5.885000 58.770000  6.085000 58.970000 ;
        RECT  5.885000 59.180000  6.085000 59.380000 ;
        RECT  5.885000 59.590000  6.085000 59.790000 ;
        RECT  5.885000 60.000000  6.085000 60.200000 ;
        RECT  5.885000 60.410000  6.085000 60.610000 ;
        RECT  6.290000 56.310000  6.490000 56.510000 ;
        RECT  6.290000 56.720000  6.490000 56.920000 ;
        RECT  6.290000 57.130000  6.490000 57.330000 ;
        RECT  6.290000 57.540000  6.490000 57.740000 ;
        RECT  6.290000 57.950000  6.490000 58.150000 ;
        RECT  6.290000 58.360000  6.490000 58.560000 ;
        RECT  6.290000 58.770000  6.490000 58.970000 ;
        RECT  6.290000 59.180000  6.490000 59.380000 ;
        RECT  6.290000 59.590000  6.490000 59.790000 ;
        RECT  6.290000 60.000000  6.490000 60.200000 ;
        RECT  6.290000 60.410000  6.490000 60.610000 ;
        RECT  6.695000 56.310000  6.895000 56.510000 ;
        RECT  6.695000 56.720000  6.895000 56.920000 ;
        RECT  6.695000 57.130000  6.895000 57.330000 ;
        RECT  6.695000 57.540000  6.895000 57.740000 ;
        RECT  6.695000 57.950000  6.895000 58.150000 ;
        RECT  6.695000 58.360000  6.895000 58.560000 ;
        RECT  6.695000 58.770000  6.895000 58.970000 ;
        RECT  6.695000 59.180000  6.895000 59.380000 ;
        RECT  6.695000 59.590000  6.895000 59.790000 ;
        RECT  6.695000 60.000000  6.895000 60.200000 ;
        RECT  6.695000 60.410000  6.895000 60.610000 ;
        RECT  7.100000 56.310000  7.300000 56.510000 ;
        RECT  7.100000 56.720000  7.300000 56.920000 ;
        RECT  7.100000 57.130000  7.300000 57.330000 ;
        RECT  7.100000 57.540000  7.300000 57.740000 ;
        RECT  7.100000 57.950000  7.300000 58.150000 ;
        RECT  7.100000 58.360000  7.300000 58.560000 ;
        RECT  7.100000 58.770000  7.300000 58.970000 ;
        RECT  7.100000 59.180000  7.300000 59.380000 ;
        RECT  7.100000 59.590000  7.300000 59.790000 ;
        RECT  7.100000 60.000000  7.300000 60.200000 ;
        RECT  7.100000 60.410000  7.300000 60.610000 ;
        RECT  7.505000 56.310000  7.705000 56.510000 ;
        RECT  7.505000 56.720000  7.705000 56.920000 ;
        RECT  7.505000 57.130000  7.705000 57.330000 ;
        RECT  7.505000 57.540000  7.705000 57.740000 ;
        RECT  7.505000 57.950000  7.705000 58.150000 ;
        RECT  7.505000 58.360000  7.705000 58.560000 ;
        RECT  7.505000 58.770000  7.705000 58.970000 ;
        RECT  7.505000 59.180000  7.705000 59.380000 ;
        RECT  7.505000 59.590000  7.705000 59.790000 ;
        RECT  7.505000 60.000000  7.705000 60.200000 ;
        RECT  7.505000 60.410000  7.705000 60.610000 ;
        RECT  7.910000 56.310000  8.110000 56.510000 ;
        RECT  7.910000 56.720000  8.110000 56.920000 ;
        RECT  7.910000 57.130000  8.110000 57.330000 ;
        RECT  7.910000 57.540000  8.110000 57.740000 ;
        RECT  7.910000 57.950000  8.110000 58.150000 ;
        RECT  7.910000 58.360000  8.110000 58.560000 ;
        RECT  7.910000 58.770000  8.110000 58.970000 ;
        RECT  7.910000 59.180000  8.110000 59.380000 ;
        RECT  7.910000 59.590000  8.110000 59.790000 ;
        RECT  7.910000 60.000000  8.110000 60.200000 ;
        RECT  7.910000 60.410000  8.110000 60.610000 ;
        RECT  8.315000 56.310000  8.515000 56.510000 ;
        RECT  8.315000 56.720000  8.515000 56.920000 ;
        RECT  8.315000 57.130000  8.515000 57.330000 ;
        RECT  8.315000 57.540000  8.515000 57.740000 ;
        RECT  8.315000 57.950000  8.515000 58.150000 ;
        RECT  8.315000 58.360000  8.515000 58.560000 ;
        RECT  8.315000 58.770000  8.515000 58.970000 ;
        RECT  8.315000 59.180000  8.515000 59.380000 ;
        RECT  8.315000 59.590000  8.515000 59.790000 ;
        RECT  8.315000 60.000000  8.515000 60.200000 ;
        RECT  8.315000 60.410000  8.515000 60.610000 ;
        RECT  8.720000 56.310000  8.920000 56.510000 ;
        RECT  8.720000 56.720000  8.920000 56.920000 ;
        RECT  8.720000 57.130000  8.920000 57.330000 ;
        RECT  8.720000 57.540000  8.920000 57.740000 ;
        RECT  8.720000 57.950000  8.920000 58.150000 ;
        RECT  8.720000 58.360000  8.920000 58.560000 ;
        RECT  8.720000 58.770000  8.920000 58.970000 ;
        RECT  8.720000 59.180000  8.920000 59.380000 ;
        RECT  8.720000 59.590000  8.920000 59.790000 ;
        RECT  8.720000 60.000000  8.920000 60.200000 ;
        RECT  8.720000 60.410000  8.920000 60.610000 ;
        RECT  9.125000 56.310000  9.325000 56.510000 ;
        RECT  9.125000 56.720000  9.325000 56.920000 ;
        RECT  9.125000 57.130000  9.325000 57.330000 ;
        RECT  9.125000 57.540000  9.325000 57.740000 ;
        RECT  9.125000 57.950000  9.325000 58.150000 ;
        RECT  9.125000 58.360000  9.325000 58.560000 ;
        RECT  9.125000 58.770000  9.325000 58.970000 ;
        RECT  9.125000 59.180000  9.325000 59.380000 ;
        RECT  9.125000 59.590000  9.325000 59.790000 ;
        RECT  9.125000 60.000000  9.325000 60.200000 ;
        RECT  9.125000 60.410000  9.325000 60.610000 ;
        RECT  9.530000 56.310000  9.730000 56.510000 ;
        RECT  9.530000 56.720000  9.730000 56.920000 ;
        RECT  9.530000 57.130000  9.730000 57.330000 ;
        RECT  9.530000 57.540000  9.730000 57.740000 ;
        RECT  9.530000 57.950000  9.730000 58.150000 ;
        RECT  9.530000 58.360000  9.730000 58.560000 ;
        RECT  9.530000 58.770000  9.730000 58.970000 ;
        RECT  9.530000 59.180000  9.730000 59.380000 ;
        RECT  9.530000 59.590000  9.730000 59.790000 ;
        RECT  9.530000 60.000000  9.730000 60.200000 ;
        RECT  9.530000 60.410000  9.730000 60.610000 ;
        RECT  9.935000 56.310000 10.135000 56.510000 ;
        RECT  9.935000 56.720000 10.135000 56.920000 ;
        RECT  9.935000 57.130000 10.135000 57.330000 ;
        RECT  9.935000 57.540000 10.135000 57.740000 ;
        RECT  9.935000 57.950000 10.135000 58.150000 ;
        RECT  9.935000 58.360000 10.135000 58.560000 ;
        RECT  9.935000 58.770000 10.135000 58.970000 ;
        RECT  9.935000 59.180000 10.135000 59.380000 ;
        RECT  9.935000 59.590000 10.135000 59.790000 ;
        RECT  9.935000 60.000000 10.135000 60.200000 ;
        RECT  9.935000 60.410000 10.135000 60.610000 ;
        RECT 10.340000 56.310000 10.540000 56.510000 ;
        RECT 10.340000 56.720000 10.540000 56.920000 ;
        RECT 10.340000 57.130000 10.540000 57.330000 ;
        RECT 10.340000 57.540000 10.540000 57.740000 ;
        RECT 10.340000 57.950000 10.540000 58.150000 ;
        RECT 10.340000 58.360000 10.540000 58.560000 ;
        RECT 10.340000 58.770000 10.540000 58.970000 ;
        RECT 10.340000 59.180000 10.540000 59.380000 ;
        RECT 10.340000 59.590000 10.540000 59.790000 ;
        RECT 10.340000 60.000000 10.540000 60.200000 ;
        RECT 10.340000 60.410000 10.540000 60.610000 ;
        RECT 10.745000 56.310000 10.945000 56.510000 ;
        RECT 10.745000 56.720000 10.945000 56.920000 ;
        RECT 10.745000 57.130000 10.945000 57.330000 ;
        RECT 10.745000 57.540000 10.945000 57.740000 ;
        RECT 10.745000 57.950000 10.945000 58.150000 ;
        RECT 10.745000 58.360000 10.945000 58.560000 ;
        RECT 10.745000 58.770000 10.945000 58.970000 ;
        RECT 10.745000 59.180000 10.945000 59.380000 ;
        RECT 10.745000 59.590000 10.945000 59.790000 ;
        RECT 10.745000 60.000000 10.945000 60.200000 ;
        RECT 10.745000 60.410000 10.945000 60.610000 ;
        RECT 11.150000 56.310000 11.350000 56.510000 ;
        RECT 11.150000 56.720000 11.350000 56.920000 ;
        RECT 11.150000 57.130000 11.350000 57.330000 ;
        RECT 11.150000 57.540000 11.350000 57.740000 ;
        RECT 11.150000 57.950000 11.350000 58.150000 ;
        RECT 11.150000 58.360000 11.350000 58.560000 ;
        RECT 11.150000 58.770000 11.350000 58.970000 ;
        RECT 11.150000 59.180000 11.350000 59.380000 ;
        RECT 11.150000 59.590000 11.350000 59.790000 ;
        RECT 11.150000 60.000000 11.350000 60.200000 ;
        RECT 11.150000 60.410000 11.350000 60.610000 ;
        RECT 11.555000 56.310000 11.755000 56.510000 ;
        RECT 11.555000 56.720000 11.755000 56.920000 ;
        RECT 11.555000 57.130000 11.755000 57.330000 ;
        RECT 11.555000 57.540000 11.755000 57.740000 ;
        RECT 11.555000 57.950000 11.755000 58.150000 ;
        RECT 11.555000 58.360000 11.755000 58.560000 ;
        RECT 11.555000 58.770000 11.755000 58.970000 ;
        RECT 11.555000 59.180000 11.755000 59.380000 ;
        RECT 11.555000 59.590000 11.755000 59.790000 ;
        RECT 11.555000 60.000000 11.755000 60.200000 ;
        RECT 11.555000 60.410000 11.755000 60.610000 ;
        RECT 11.960000 56.310000 12.160000 56.510000 ;
        RECT 11.960000 56.720000 12.160000 56.920000 ;
        RECT 11.960000 57.130000 12.160000 57.330000 ;
        RECT 11.960000 57.540000 12.160000 57.740000 ;
        RECT 11.960000 57.950000 12.160000 58.150000 ;
        RECT 11.960000 58.360000 12.160000 58.560000 ;
        RECT 11.960000 58.770000 12.160000 58.970000 ;
        RECT 11.960000 59.180000 12.160000 59.380000 ;
        RECT 11.960000 59.590000 12.160000 59.790000 ;
        RECT 11.960000 60.000000 12.160000 60.200000 ;
        RECT 11.960000 60.410000 12.160000 60.610000 ;
        RECT 12.365000 56.310000 12.565000 56.510000 ;
        RECT 12.365000 56.720000 12.565000 56.920000 ;
        RECT 12.365000 57.130000 12.565000 57.330000 ;
        RECT 12.365000 57.540000 12.565000 57.740000 ;
        RECT 12.365000 57.950000 12.565000 58.150000 ;
        RECT 12.365000 58.360000 12.565000 58.560000 ;
        RECT 12.365000 58.770000 12.565000 58.970000 ;
        RECT 12.365000 59.180000 12.565000 59.380000 ;
        RECT 12.365000 59.590000 12.565000 59.790000 ;
        RECT 12.365000 60.000000 12.565000 60.200000 ;
        RECT 12.365000 60.410000 12.565000 60.610000 ;
        RECT 12.770000 56.310000 12.970000 56.510000 ;
        RECT 12.770000 56.720000 12.970000 56.920000 ;
        RECT 12.770000 57.130000 12.970000 57.330000 ;
        RECT 12.770000 57.540000 12.970000 57.740000 ;
        RECT 12.770000 57.950000 12.970000 58.150000 ;
        RECT 12.770000 58.360000 12.970000 58.560000 ;
        RECT 12.770000 58.770000 12.970000 58.970000 ;
        RECT 12.770000 59.180000 12.970000 59.380000 ;
        RECT 12.770000 59.590000 12.970000 59.790000 ;
        RECT 12.770000 60.000000 12.970000 60.200000 ;
        RECT 12.770000 60.410000 12.970000 60.610000 ;
        RECT 13.175000 56.310000 13.375000 56.510000 ;
        RECT 13.175000 56.720000 13.375000 56.920000 ;
        RECT 13.175000 57.130000 13.375000 57.330000 ;
        RECT 13.175000 57.540000 13.375000 57.740000 ;
        RECT 13.175000 57.950000 13.375000 58.150000 ;
        RECT 13.175000 58.360000 13.375000 58.560000 ;
        RECT 13.175000 58.770000 13.375000 58.970000 ;
        RECT 13.175000 59.180000 13.375000 59.380000 ;
        RECT 13.175000 59.590000 13.375000 59.790000 ;
        RECT 13.175000 60.000000 13.375000 60.200000 ;
        RECT 13.175000 60.410000 13.375000 60.610000 ;
        RECT 13.580000 56.310000 13.780000 56.510000 ;
        RECT 13.580000 56.720000 13.780000 56.920000 ;
        RECT 13.580000 57.130000 13.780000 57.330000 ;
        RECT 13.580000 57.540000 13.780000 57.740000 ;
        RECT 13.580000 57.950000 13.780000 58.150000 ;
        RECT 13.580000 58.360000 13.780000 58.560000 ;
        RECT 13.580000 58.770000 13.780000 58.970000 ;
        RECT 13.580000 59.180000 13.780000 59.380000 ;
        RECT 13.580000 59.590000 13.780000 59.790000 ;
        RECT 13.580000 60.000000 13.780000 60.200000 ;
        RECT 13.580000 60.410000 13.780000 60.610000 ;
        RECT 13.985000 56.310000 14.185000 56.510000 ;
        RECT 13.985000 56.720000 14.185000 56.920000 ;
        RECT 13.985000 57.130000 14.185000 57.330000 ;
        RECT 13.985000 57.540000 14.185000 57.740000 ;
        RECT 13.985000 57.950000 14.185000 58.150000 ;
        RECT 13.985000 58.360000 14.185000 58.560000 ;
        RECT 13.985000 58.770000 14.185000 58.970000 ;
        RECT 13.985000 59.180000 14.185000 59.380000 ;
        RECT 13.985000 59.590000 14.185000 59.790000 ;
        RECT 13.985000 60.000000 14.185000 60.200000 ;
        RECT 13.985000 60.410000 14.185000 60.610000 ;
        RECT 14.390000 56.310000 14.590000 56.510000 ;
        RECT 14.390000 56.720000 14.590000 56.920000 ;
        RECT 14.390000 57.130000 14.590000 57.330000 ;
        RECT 14.390000 57.540000 14.590000 57.740000 ;
        RECT 14.390000 57.950000 14.590000 58.150000 ;
        RECT 14.390000 58.360000 14.590000 58.560000 ;
        RECT 14.390000 58.770000 14.590000 58.970000 ;
        RECT 14.390000 59.180000 14.590000 59.380000 ;
        RECT 14.390000 59.590000 14.590000 59.790000 ;
        RECT 14.390000 60.000000 14.590000 60.200000 ;
        RECT 14.390000 60.410000 14.590000 60.610000 ;
        RECT 14.795000 56.310000 14.995000 56.510000 ;
        RECT 14.795000 56.720000 14.995000 56.920000 ;
        RECT 14.795000 57.130000 14.995000 57.330000 ;
        RECT 14.795000 57.540000 14.995000 57.740000 ;
        RECT 14.795000 57.950000 14.995000 58.150000 ;
        RECT 14.795000 58.360000 14.995000 58.560000 ;
        RECT 14.795000 58.770000 14.995000 58.970000 ;
        RECT 14.795000 59.180000 14.995000 59.380000 ;
        RECT 14.795000 59.590000 14.995000 59.790000 ;
        RECT 14.795000 60.000000 14.995000 60.200000 ;
        RECT 14.795000 60.410000 14.995000 60.610000 ;
        RECT 15.200000 56.310000 15.400000 56.510000 ;
        RECT 15.200000 56.720000 15.400000 56.920000 ;
        RECT 15.200000 57.130000 15.400000 57.330000 ;
        RECT 15.200000 57.540000 15.400000 57.740000 ;
        RECT 15.200000 57.950000 15.400000 58.150000 ;
        RECT 15.200000 58.360000 15.400000 58.560000 ;
        RECT 15.200000 58.770000 15.400000 58.970000 ;
        RECT 15.200000 59.180000 15.400000 59.380000 ;
        RECT 15.200000 59.590000 15.400000 59.790000 ;
        RECT 15.200000 60.000000 15.400000 60.200000 ;
        RECT 15.200000 60.410000 15.400000 60.610000 ;
        RECT 15.605000 56.310000 15.805000 56.510000 ;
        RECT 15.605000 56.720000 15.805000 56.920000 ;
        RECT 15.605000 57.130000 15.805000 57.330000 ;
        RECT 15.605000 57.540000 15.805000 57.740000 ;
        RECT 15.605000 57.950000 15.805000 58.150000 ;
        RECT 15.605000 58.360000 15.805000 58.560000 ;
        RECT 15.605000 58.770000 15.805000 58.970000 ;
        RECT 15.605000 59.180000 15.805000 59.380000 ;
        RECT 15.605000 59.590000 15.805000 59.790000 ;
        RECT 15.605000 60.000000 15.805000 60.200000 ;
        RECT 15.605000 60.410000 15.805000 60.610000 ;
        RECT 16.010000 56.310000 16.210000 56.510000 ;
        RECT 16.010000 56.720000 16.210000 56.920000 ;
        RECT 16.010000 57.130000 16.210000 57.330000 ;
        RECT 16.010000 57.540000 16.210000 57.740000 ;
        RECT 16.010000 57.950000 16.210000 58.150000 ;
        RECT 16.010000 58.360000 16.210000 58.560000 ;
        RECT 16.010000 58.770000 16.210000 58.970000 ;
        RECT 16.010000 59.180000 16.210000 59.380000 ;
        RECT 16.010000 59.590000 16.210000 59.790000 ;
        RECT 16.010000 60.000000 16.210000 60.200000 ;
        RECT 16.010000 60.410000 16.210000 60.610000 ;
        RECT 16.415000 56.310000 16.615000 56.510000 ;
        RECT 16.415000 56.720000 16.615000 56.920000 ;
        RECT 16.415000 57.130000 16.615000 57.330000 ;
        RECT 16.415000 57.540000 16.615000 57.740000 ;
        RECT 16.415000 57.950000 16.615000 58.150000 ;
        RECT 16.415000 58.360000 16.615000 58.560000 ;
        RECT 16.415000 58.770000 16.615000 58.970000 ;
        RECT 16.415000 59.180000 16.615000 59.380000 ;
        RECT 16.415000 59.590000 16.615000 59.790000 ;
        RECT 16.415000 60.000000 16.615000 60.200000 ;
        RECT 16.415000 60.410000 16.615000 60.610000 ;
        RECT 16.820000 56.310000 17.020000 56.510000 ;
        RECT 16.820000 56.720000 17.020000 56.920000 ;
        RECT 16.820000 57.130000 17.020000 57.330000 ;
        RECT 16.820000 57.540000 17.020000 57.740000 ;
        RECT 16.820000 57.950000 17.020000 58.150000 ;
        RECT 16.820000 58.360000 17.020000 58.560000 ;
        RECT 16.820000 58.770000 17.020000 58.970000 ;
        RECT 16.820000 59.180000 17.020000 59.380000 ;
        RECT 16.820000 59.590000 17.020000 59.790000 ;
        RECT 16.820000 60.000000 17.020000 60.200000 ;
        RECT 16.820000 60.410000 17.020000 60.610000 ;
        RECT 17.225000 56.310000 17.425000 56.510000 ;
        RECT 17.225000 56.720000 17.425000 56.920000 ;
        RECT 17.225000 57.130000 17.425000 57.330000 ;
        RECT 17.225000 57.540000 17.425000 57.740000 ;
        RECT 17.225000 57.950000 17.425000 58.150000 ;
        RECT 17.225000 58.360000 17.425000 58.560000 ;
        RECT 17.225000 58.770000 17.425000 58.970000 ;
        RECT 17.225000 59.180000 17.425000 59.380000 ;
        RECT 17.225000 59.590000 17.425000 59.790000 ;
        RECT 17.225000 60.000000 17.425000 60.200000 ;
        RECT 17.225000 60.410000 17.425000 60.610000 ;
        RECT 17.630000 56.310000 17.830000 56.510000 ;
        RECT 17.630000 56.720000 17.830000 56.920000 ;
        RECT 17.630000 57.130000 17.830000 57.330000 ;
        RECT 17.630000 57.540000 17.830000 57.740000 ;
        RECT 17.630000 57.950000 17.830000 58.150000 ;
        RECT 17.630000 58.360000 17.830000 58.560000 ;
        RECT 17.630000 58.770000 17.830000 58.970000 ;
        RECT 17.630000 59.180000 17.830000 59.380000 ;
        RECT 17.630000 59.590000 17.830000 59.790000 ;
        RECT 17.630000 60.000000 17.830000 60.200000 ;
        RECT 17.630000 60.410000 17.830000 60.610000 ;
        RECT 18.035000 56.310000 18.235000 56.510000 ;
        RECT 18.035000 56.720000 18.235000 56.920000 ;
        RECT 18.035000 57.130000 18.235000 57.330000 ;
        RECT 18.035000 57.540000 18.235000 57.740000 ;
        RECT 18.035000 57.950000 18.235000 58.150000 ;
        RECT 18.035000 58.360000 18.235000 58.560000 ;
        RECT 18.035000 58.770000 18.235000 58.970000 ;
        RECT 18.035000 59.180000 18.235000 59.380000 ;
        RECT 18.035000 59.590000 18.235000 59.790000 ;
        RECT 18.035000 60.000000 18.235000 60.200000 ;
        RECT 18.035000 60.410000 18.235000 60.610000 ;
        RECT 18.440000 56.310000 18.640000 56.510000 ;
        RECT 18.440000 56.720000 18.640000 56.920000 ;
        RECT 18.440000 57.130000 18.640000 57.330000 ;
        RECT 18.440000 57.540000 18.640000 57.740000 ;
        RECT 18.440000 57.950000 18.640000 58.150000 ;
        RECT 18.440000 58.360000 18.640000 58.560000 ;
        RECT 18.440000 58.770000 18.640000 58.970000 ;
        RECT 18.440000 59.180000 18.640000 59.380000 ;
        RECT 18.440000 59.590000 18.640000 59.790000 ;
        RECT 18.440000 60.000000 18.640000 60.200000 ;
        RECT 18.440000 60.410000 18.640000 60.610000 ;
        RECT 18.845000 56.310000 19.045000 56.510000 ;
        RECT 18.845000 56.720000 19.045000 56.920000 ;
        RECT 18.845000 57.130000 19.045000 57.330000 ;
        RECT 18.845000 57.540000 19.045000 57.740000 ;
        RECT 18.845000 57.950000 19.045000 58.150000 ;
        RECT 18.845000 58.360000 19.045000 58.560000 ;
        RECT 18.845000 58.770000 19.045000 58.970000 ;
        RECT 18.845000 59.180000 19.045000 59.380000 ;
        RECT 18.845000 59.590000 19.045000 59.790000 ;
        RECT 18.845000 60.000000 19.045000 60.200000 ;
        RECT 18.845000 60.410000 19.045000 60.610000 ;
        RECT 19.250000 56.310000 19.450000 56.510000 ;
        RECT 19.250000 56.720000 19.450000 56.920000 ;
        RECT 19.250000 57.130000 19.450000 57.330000 ;
        RECT 19.250000 57.540000 19.450000 57.740000 ;
        RECT 19.250000 57.950000 19.450000 58.150000 ;
        RECT 19.250000 58.360000 19.450000 58.560000 ;
        RECT 19.250000 58.770000 19.450000 58.970000 ;
        RECT 19.250000 59.180000 19.450000 59.380000 ;
        RECT 19.250000 59.590000 19.450000 59.790000 ;
        RECT 19.250000 60.000000 19.450000 60.200000 ;
        RECT 19.250000 60.410000 19.450000 60.610000 ;
        RECT 19.655000 56.310000 19.855000 56.510000 ;
        RECT 19.655000 56.720000 19.855000 56.920000 ;
        RECT 19.655000 57.130000 19.855000 57.330000 ;
        RECT 19.655000 57.540000 19.855000 57.740000 ;
        RECT 19.655000 57.950000 19.855000 58.150000 ;
        RECT 19.655000 58.360000 19.855000 58.560000 ;
        RECT 19.655000 58.770000 19.855000 58.970000 ;
        RECT 19.655000 59.180000 19.855000 59.380000 ;
        RECT 19.655000 59.590000 19.855000 59.790000 ;
        RECT 19.655000 60.000000 19.855000 60.200000 ;
        RECT 19.655000 60.410000 19.855000 60.610000 ;
        RECT 20.060000 56.310000 20.260000 56.510000 ;
        RECT 20.060000 56.720000 20.260000 56.920000 ;
        RECT 20.060000 57.130000 20.260000 57.330000 ;
        RECT 20.060000 57.540000 20.260000 57.740000 ;
        RECT 20.060000 57.950000 20.260000 58.150000 ;
        RECT 20.060000 58.360000 20.260000 58.560000 ;
        RECT 20.060000 58.770000 20.260000 58.970000 ;
        RECT 20.060000 59.180000 20.260000 59.380000 ;
        RECT 20.060000 59.590000 20.260000 59.790000 ;
        RECT 20.060000 60.000000 20.260000 60.200000 ;
        RECT 20.060000 60.410000 20.260000 60.610000 ;
        RECT 20.465000 56.310000 20.665000 56.510000 ;
        RECT 20.465000 56.720000 20.665000 56.920000 ;
        RECT 20.465000 57.130000 20.665000 57.330000 ;
        RECT 20.465000 57.540000 20.665000 57.740000 ;
        RECT 20.465000 57.950000 20.665000 58.150000 ;
        RECT 20.465000 58.360000 20.665000 58.560000 ;
        RECT 20.465000 58.770000 20.665000 58.970000 ;
        RECT 20.465000 59.180000 20.665000 59.380000 ;
        RECT 20.465000 59.590000 20.665000 59.790000 ;
        RECT 20.465000 60.000000 20.665000 60.200000 ;
        RECT 20.465000 60.410000 20.665000 60.610000 ;
        RECT 20.870000 56.310000 21.070000 56.510000 ;
        RECT 20.870000 56.720000 21.070000 56.920000 ;
        RECT 20.870000 57.130000 21.070000 57.330000 ;
        RECT 20.870000 57.540000 21.070000 57.740000 ;
        RECT 20.870000 57.950000 21.070000 58.150000 ;
        RECT 20.870000 58.360000 21.070000 58.560000 ;
        RECT 20.870000 58.770000 21.070000 58.970000 ;
        RECT 20.870000 59.180000 21.070000 59.380000 ;
        RECT 20.870000 59.590000 21.070000 59.790000 ;
        RECT 20.870000 60.000000 21.070000 60.200000 ;
        RECT 20.870000 60.410000 21.070000 60.610000 ;
        RECT 21.275000 56.310000 21.475000 56.510000 ;
        RECT 21.275000 56.720000 21.475000 56.920000 ;
        RECT 21.275000 57.130000 21.475000 57.330000 ;
        RECT 21.275000 57.540000 21.475000 57.740000 ;
        RECT 21.275000 57.950000 21.475000 58.150000 ;
        RECT 21.275000 58.360000 21.475000 58.560000 ;
        RECT 21.275000 58.770000 21.475000 58.970000 ;
        RECT 21.275000 59.180000 21.475000 59.380000 ;
        RECT 21.275000 59.590000 21.475000 59.790000 ;
        RECT 21.275000 60.000000 21.475000 60.200000 ;
        RECT 21.275000 60.410000 21.475000 60.610000 ;
        RECT 21.680000 56.310000 21.880000 56.510000 ;
        RECT 21.680000 56.720000 21.880000 56.920000 ;
        RECT 21.680000 57.130000 21.880000 57.330000 ;
        RECT 21.680000 57.540000 21.880000 57.740000 ;
        RECT 21.680000 57.950000 21.880000 58.150000 ;
        RECT 21.680000 58.360000 21.880000 58.560000 ;
        RECT 21.680000 58.770000 21.880000 58.970000 ;
        RECT 21.680000 59.180000 21.880000 59.380000 ;
        RECT 21.680000 59.590000 21.880000 59.790000 ;
        RECT 21.680000 60.000000 21.880000 60.200000 ;
        RECT 21.680000 60.410000 21.880000 60.610000 ;
        RECT 22.085000 56.310000 22.285000 56.510000 ;
        RECT 22.085000 56.720000 22.285000 56.920000 ;
        RECT 22.085000 57.130000 22.285000 57.330000 ;
        RECT 22.085000 57.540000 22.285000 57.740000 ;
        RECT 22.085000 57.950000 22.285000 58.150000 ;
        RECT 22.085000 58.360000 22.285000 58.560000 ;
        RECT 22.085000 58.770000 22.285000 58.970000 ;
        RECT 22.085000 59.180000 22.285000 59.380000 ;
        RECT 22.085000 59.590000 22.285000 59.790000 ;
        RECT 22.085000 60.000000 22.285000 60.200000 ;
        RECT 22.085000 60.410000 22.285000 60.610000 ;
        RECT 22.490000 56.310000 22.690000 56.510000 ;
        RECT 22.490000 56.720000 22.690000 56.920000 ;
        RECT 22.490000 57.130000 22.690000 57.330000 ;
        RECT 22.490000 57.540000 22.690000 57.740000 ;
        RECT 22.490000 57.950000 22.690000 58.150000 ;
        RECT 22.490000 58.360000 22.690000 58.560000 ;
        RECT 22.490000 58.770000 22.690000 58.970000 ;
        RECT 22.490000 59.180000 22.690000 59.380000 ;
        RECT 22.490000 59.590000 22.690000 59.790000 ;
        RECT 22.490000 60.000000 22.690000 60.200000 ;
        RECT 22.490000 60.410000 22.690000 60.610000 ;
        RECT 22.895000 56.310000 23.095000 56.510000 ;
        RECT 22.895000 56.720000 23.095000 56.920000 ;
        RECT 22.895000 57.130000 23.095000 57.330000 ;
        RECT 22.895000 57.540000 23.095000 57.740000 ;
        RECT 22.895000 57.950000 23.095000 58.150000 ;
        RECT 22.895000 58.360000 23.095000 58.560000 ;
        RECT 22.895000 58.770000 23.095000 58.970000 ;
        RECT 22.895000 59.180000 23.095000 59.380000 ;
        RECT 22.895000 59.590000 23.095000 59.790000 ;
        RECT 22.895000 60.000000 23.095000 60.200000 ;
        RECT 22.895000 60.410000 23.095000 60.610000 ;
        RECT 23.300000 56.310000 23.500000 56.510000 ;
        RECT 23.300000 56.720000 23.500000 56.920000 ;
        RECT 23.300000 57.130000 23.500000 57.330000 ;
        RECT 23.300000 57.540000 23.500000 57.740000 ;
        RECT 23.300000 57.950000 23.500000 58.150000 ;
        RECT 23.300000 58.360000 23.500000 58.560000 ;
        RECT 23.300000 58.770000 23.500000 58.970000 ;
        RECT 23.300000 59.180000 23.500000 59.380000 ;
        RECT 23.300000 59.590000 23.500000 59.790000 ;
        RECT 23.300000 60.000000 23.500000 60.200000 ;
        RECT 23.300000 60.410000 23.500000 60.610000 ;
        RECT 23.705000 56.310000 23.905000 56.510000 ;
        RECT 23.705000 56.720000 23.905000 56.920000 ;
        RECT 23.705000 57.130000 23.905000 57.330000 ;
        RECT 23.705000 57.540000 23.905000 57.740000 ;
        RECT 23.705000 57.950000 23.905000 58.150000 ;
        RECT 23.705000 58.360000 23.905000 58.560000 ;
        RECT 23.705000 58.770000 23.905000 58.970000 ;
        RECT 23.705000 59.180000 23.905000 59.380000 ;
        RECT 23.705000 59.590000 23.905000 59.790000 ;
        RECT 23.705000 60.000000 23.905000 60.200000 ;
        RECT 23.705000 60.410000 23.905000 60.610000 ;
        RECT 24.110000 56.310000 24.310000 56.510000 ;
        RECT 24.110000 56.720000 24.310000 56.920000 ;
        RECT 24.110000 57.130000 24.310000 57.330000 ;
        RECT 24.110000 57.540000 24.310000 57.740000 ;
        RECT 24.110000 57.950000 24.310000 58.150000 ;
        RECT 24.110000 58.360000 24.310000 58.560000 ;
        RECT 24.110000 58.770000 24.310000 58.970000 ;
        RECT 24.110000 59.180000 24.310000 59.380000 ;
        RECT 24.110000 59.590000 24.310000 59.790000 ;
        RECT 24.110000 60.000000 24.310000 60.200000 ;
        RECT 24.110000 60.410000 24.310000 60.610000 ;
        RECT 50.845000 56.310000 51.045000 56.510000 ;
        RECT 50.845000 56.720000 51.045000 56.920000 ;
        RECT 50.845000 57.130000 51.045000 57.330000 ;
        RECT 50.845000 57.540000 51.045000 57.740000 ;
        RECT 50.845000 57.950000 51.045000 58.150000 ;
        RECT 50.845000 58.360000 51.045000 58.560000 ;
        RECT 50.845000 58.770000 51.045000 58.970000 ;
        RECT 50.845000 59.180000 51.045000 59.380000 ;
        RECT 50.845000 59.590000 51.045000 59.790000 ;
        RECT 50.845000 60.000000 51.045000 60.200000 ;
        RECT 50.845000 60.410000 51.045000 60.610000 ;
        RECT 51.255000 56.310000 51.455000 56.510000 ;
        RECT 51.255000 56.720000 51.455000 56.920000 ;
        RECT 51.255000 57.130000 51.455000 57.330000 ;
        RECT 51.255000 57.540000 51.455000 57.740000 ;
        RECT 51.255000 57.950000 51.455000 58.150000 ;
        RECT 51.255000 58.360000 51.455000 58.560000 ;
        RECT 51.255000 58.770000 51.455000 58.970000 ;
        RECT 51.255000 59.180000 51.455000 59.380000 ;
        RECT 51.255000 59.590000 51.455000 59.790000 ;
        RECT 51.255000 60.000000 51.455000 60.200000 ;
        RECT 51.255000 60.410000 51.455000 60.610000 ;
        RECT 51.665000 56.310000 51.865000 56.510000 ;
        RECT 51.665000 56.720000 51.865000 56.920000 ;
        RECT 51.665000 57.130000 51.865000 57.330000 ;
        RECT 51.665000 57.540000 51.865000 57.740000 ;
        RECT 51.665000 57.950000 51.865000 58.150000 ;
        RECT 51.665000 58.360000 51.865000 58.560000 ;
        RECT 51.665000 58.770000 51.865000 58.970000 ;
        RECT 51.665000 59.180000 51.865000 59.380000 ;
        RECT 51.665000 59.590000 51.865000 59.790000 ;
        RECT 51.665000 60.000000 51.865000 60.200000 ;
        RECT 51.665000 60.410000 51.865000 60.610000 ;
        RECT 52.075000 56.310000 52.275000 56.510000 ;
        RECT 52.075000 56.720000 52.275000 56.920000 ;
        RECT 52.075000 57.130000 52.275000 57.330000 ;
        RECT 52.075000 57.540000 52.275000 57.740000 ;
        RECT 52.075000 57.950000 52.275000 58.150000 ;
        RECT 52.075000 58.360000 52.275000 58.560000 ;
        RECT 52.075000 58.770000 52.275000 58.970000 ;
        RECT 52.075000 59.180000 52.275000 59.380000 ;
        RECT 52.075000 59.590000 52.275000 59.790000 ;
        RECT 52.075000 60.000000 52.275000 60.200000 ;
        RECT 52.075000 60.410000 52.275000 60.610000 ;
        RECT 52.485000 56.310000 52.685000 56.510000 ;
        RECT 52.485000 56.720000 52.685000 56.920000 ;
        RECT 52.485000 57.130000 52.685000 57.330000 ;
        RECT 52.485000 57.540000 52.685000 57.740000 ;
        RECT 52.485000 57.950000 52.685000 58.150000 ;
        RECT 52.485000 58.360000 52.685000 58.560000 ;
        RECT 52.485000 58.770000 52.685000 58.970000 ;
        RECT 52.485000 59.180000 52.685000 59.380000 ;
        RECT 52.485000 59.590000 52.685000 59.790000 ;
        RECT 52.485000 60.000000 52.685000 60.200000 ;
        RECT 52.485000 60.410000 52.685000 60.610000 ;
        RECT 52.895000 56.310000 53.095000 56.510000 ;
        RECT 52.895000 56.720000 53.095000 56.920000 ;
        RECT 52.895000 57.130000 53.095000 57.330000 ;
        RECT 52.895000 57.540000 53.095000 57.740000 ;
        RECT 52.895000 57.950000 53.095000 58.150000 ;
        RECT 52.895000 58.360000 53.095000 58.560000 ;
        RECT 52.895000 58.770000 53.095000 58.970000 ;
        RECT 52.895000 59.180000 53.095000 59.380000 ;
        RECT 52.895000 59.590000 53.095000 59.790000 ;
        RECT 52.895000 60.000000 53.095000 60.200000 ;
        RECT 52.895000 60.410000 53.095000 60.610000 ;
        RECT 53.305000 56.310000 53.505000 56.510000 ;
        RECT 53.305000 56.720000 53.505000 56.920000 ;
        RECT 53.305000 57.130000 53.505000 57.330000 ;
        RECT 53.305000 57.540000 53.505000 57.740000 ;
        RECT 53.305000 57.950000 53.505000 58.150000 ;
        RECT 53.305000 58.360000 53.505000 58.560000 ;
        RECT 53.305000 58.770000 53.505000 58.970000 ;
        RECT 53.305000 59.180000 53.505000 59.380000 ;
        RECT 53.305000 59.590000 53.505000 59.790000 ;
        RECT 53.305000 60.000000 53.505000 60.200000 ;
        RECT 53.305000 60.410000 53.505000 60.610000 ;
        RECT 53.715000 56.310000 53.915000 56.510000 ;
        RECT 53.715000 56.720000 53.915000 56.920000 ;
        RECT 53.715000 57.130000 53.915000 57.330000 ;
        RECT 53.715000 57.540000 53.915000 57.740000 ;
        RECT 53.715000 57.950000 53.915000 58.150000 ;
        RECT 53.715000 58.360000 53.915000 58.560000 ;
        RECT 53.715000 58.770000 53.915000 58.970000 ;
        RECT 53.715000 59.180000 53.915000 59.380000 ;
        RECT 53.715000 59.590000 53.915000 59.790000 ;
        RECT 53.715000 60.000000 53.915000 60.200000 ;
        RECT 53.715000 60.410000 53.915000 60.610000 ;
        RECT 54.125000 56.310000 54.325000 56.510000 ;
        RECT 54.125000 56.720000 54.325000 56.920000 ;
        RECT 54.125000 57.130000 54.325000 57.330000 ;
        RECT 54.125000 57.540000 54.325000 57.740000 ;
        RECT 54.125000 57.950000 54.325000 58.150000 ;
        RECT 54.125000 58.360000 54.325000 58.560000 ;
        RECT 54.125000 58.770000 54.325000 58.970000 ;
        RECT 54.125000 59.180000 54.325000 59.380000 ;
        RECT 54.125000 59.590000 54.325000 59.790000 ;
        RECT 54.125000 60.000000 54.325000 60.200000 ;
        RECT 54.125000 60.410000 54.325000 60.610000 ;
        RECT 54.535000 56.310000 54.735000 56.510000 ;
        RECT 54.535000 56.720000 54.735000 56.920000 ;
        RECT 54.535000 57.130000 54.735000 57.330000 ;
        RECT 54.535000 57.540000 54.735000 57.740000 ;
        RECT 54.535000 57.950000 54.735000 58.150000 ;
        RECT 54.535000 58.360000 54.735000 58.560000 ;
        RECT 54.535000 58.770000 54.735000 58.970000 ;
        RECT 54.535000 59.180000 54.735000 59.380000 ;
        RECT 54.535000 59.590000 54.735000 59.790000 ;
        RECT 54.535000 60.000000 54.735000 60.200000 ;
        RECT 54.535000 60.410000 54.735000 60.610000 ;
        RECT 54.945000 56.310000 55.145000 56.510000 ;
        RECT 54.945000 56.720000 55.145000 56.920000 ;
        RECT 54.945000 57.130000 55.145000 57.330000 ;
        RECT 54.945000 57.540000 55.145000 57.740000 ;
        RECT 54.945000 57.950000 55.145000 58.150000 ;
        RECT 54.945000 58.360000 55.145000 58.560000 ;
        RECT 54.945000 58.770000 55.145000 58.970000 ;
        RECT 54.945000 59.180000 55.145000 59.380000 ;
        RECT 54.945000 59.590000 55.145000 59.790000 ;
        RECT 54.945000 60.000000 55.145000 60.200000 ;
        RECT 54.945000 60.410000 55.145000 60.610000 ;
        RECT 55.355000 56.310000 55.555000 56.510000 ;
        RECT 55.355000 56.720000 55.555000 56.920000 ;
        RECT 55.355000 57.130000 55.555000 57.330000 ;
        RECT 55.355000 57.540000 55.555000 57.740000 ;
        RECT 55.355000 57.950000 55.555000 58.150000 ;
        RECT 55.355000 58.360000 55.555000 58.560000 ;
        RECT 55.355000 58.770000 55.555000 58.970000 ;
        RECT 55.355000 59.180000 55.555000 59.380000 ;
        RECT 55.355000 59.590000 55.555000 59.790000 ;
        RECT 55.355000 60.000000 55.555000 60.200000 ;
        RECT 55.355000 60.410000 55.555000 60.610000 ;
        RECT 55.765000 56.310000 55.965000 56.510000 ;
        RECT 55.765000 56.720000 55.965000 56.920000 ;
        RECT 55.765000 57.130000 55.965000 57.330000 ;
        RECT 55.765000 57.540000 55.965000 57.740000 ;
        RECT 55.765000 57.950000 55.965000 58.150000 ;
        RECT 55.765000 58.360000 55.965000 58.560000 ;
        RECT 55.765000 58.770000 55.965000 58.970000 ;
        RECT 55.765000 59.180000 55.965000 59.380000 ;
        RECT 55.765000 59.590000 55.965000 59.790000 ;
        RECT 55.765000 60.000000 55.965000 60.200000 ;
        RECT 55.765000 60.410000 55.965000 60.610000 ;
        RECT 56.175000 56.310000 56.375000 56.510000 ;
        RECT 56.175000 56.720000 56.375000 56.920000 ;
        RECT 56.175000 57.130000 56.375000 57.330000 ;
        RECT 56.175000 57.540000 56.375000 57.740000 ;
        RECT 56.175000 57.950000 56.375000 58.150000 ;
        RECT 56.175000 58.360000 56.375000 58.560000 ;
        RECT 56.175000 58.770000 56.375000 58.970000 ;
        RECT 56.175000 59.180000 56.375000 59.380000 ;
        RECT 56.175000 59.590000 56.375000 59.790000 ;
        RECT 56.175000 60.000000 56.375000 60.200000 ;
        RECT 56.175000 60.410000 56.375000 60.610000 ;
        RECT 56.585000 56.310000 56.785000 56.510000 ;
        RECT 56.585000 56.720000 56.785000 56.920000 ;
        RECT 56.585000 57.130000 56.785000 57.330000 ;
        RECT 56.585000 57.540000 56.785000 57.740000 ;
        RECT 56.585000 57.950000 56.785000 58.150000 ;
        RECT 56.585000 58.360000 56.785000 58.560000 ;
        RECT 56.585000 58.770000 56.785000 58.970000 ;
        RECT 56.585000 59.180000 56.785000 59.380000 ;
        RECT 56.585000 59.590000 56.785000 59.790000 ;
        RECT 56.585000 60.000000 56.785000 60.200000 ;
        RECT 56.585000 60.410000 56.785000 60.610000 ;
        RECT 56.990000 56.310000 57.190000 56.510000 ;
        RECT 56.990000 56.720000 57.190000 56.920000 ;
        RECT 56.990000 57.130000 57.190000 57.330000 ;
        RECT 56.990000 57.540000 57.190000 57.740000 ;
        RECT 56.990000 57.950000 57.190000 58.150000 ;
        RECT 56.990000 58.360000 57.190000 58.560000 ;
        RECT 56.990000 58.770000 57.190000 58.970000 ;
        RECT 56.990000 59.180000 57.190000 59.380000 ;
        RECT 56.990000 59.590000 57.190000 59.790000 ;
        RECT 56.990000 60.000000 57.190000 60.200000 ;
        RECT 56.990000 60.410000 57.190000 60.610000 ;
        RECT 57.395000 56.310000 57.595000 56.510000 ;
        RECT 57.395000 56.720000 57.595000 56.920000 ;
        RECT 57.395000 57.130000 57.595000 57.330000 ;
        RECT 57.395000 57.540000 57.595000 57.740000 ;
        RECT 57.395000 57.950000 57.595000 58.150000 ;
        RECT 57.395000 58.360000 57.595000 58.560000 ;
        RECT 57.395000 58.770000 57.595000 58.970000 ;
        RECT 57.395000 59.180000 57.595000 59.380000 ;
        RECT 57.395000 59.590000 57.595000 59.790000 ;
        RECT 57.395000 60.000000 57.595000 60.200000 ;
        RECT 57.395000 60.410000 57.595000 60.610000 ;
        RECT 57.800000 56.310000 58.000000 56.510000 ;
        RECT 57.800000 56.720000 58.000000 56.920000 ;
        RECT 57.800000 57.130000 58.000000 57.330000 ;
        RECT 57.800000 57.540000 58.000000 57.740000 ;
        RECT 57.800000 57.950000 58.000000 58.150000 ;
        RECT 57.800000 58.360000 58.000000 58.560000 ;
        RECT 57.800000 58.770000 58.000000 58.970000 ;
        RECT 57.800000 59.180000 58.000000 59.380000 ;
        RECT 57.800000 59.590000 58.000000 59.790000 ;
        RECT 57.800000 60.000000 58.000000 60.200000 ;
        RECT 57.800000 60.410000 58.000000 60.610000 ;
        RECT 58.205000 56.310000 58.405000 56.510000 ;
        RECT 58.205000 56.720000 58.405000 56.920000 ;
        RECT 58.205000 57.130000 58.405000 57.330000 ;
        RECT 58.205000 57.540000 58.405000 57.740000 ;
        RECT 58.205000 57.950000 58.405000 58.150000 ;
        RECT 58.205000 58.360000 58.405000 58.560000 ;
        RECT 58.205000 58.770000 58.405000 58.970000 ;
        RECT 58.205000 59.180000 58.405000 59.380000 ;
        RECT 58.205000 59.590000 58.405000 59.790000 ;
        RECT 58.205000 60.000000 58.405000 60.200000 ;
        RECT 58.205000 60.410000 58.405000 60.610000 ;
        RECT 58.610000 56.310000 58.810000 56.510000 ;
        RECT 58.610000 56.720000 58.810000 56.920000 ;
        RECT 58.610000 57.130000 58.810000 57.330000 ;
        RECT 58.610000 57.540000 58.810000 57.740000 ;
        RECT 58.610000 57.950000 58.810000 58.150000 ;
        RECT 58.610000 58.360000 58.810000 58.560000 ;
        RECT 58.610000 58.770000 58.810000 58.970000 ;
        RECT 58.610000 59.180000 58.810000 59.380000 ;
        RECT 58.610000 59.590000 58.810000 59.790000 ;
        RECT 58.610000 60.000000 58.810000 60.200000 ;
        RECT 58.610000 60.410000 58.810000 60.610000 ;
        RECT 59.015000 56.310000 59.215000 56.510000 ;
        RECT 59.015000 56.720000 59.215000 56.920000 ;
        RECT 59.015000 57.130000 59.215000 57.330000 ;
        RECT 59.015000 57.540000 59.215000 57.740000 ;
        RECT 59.015000 57.950000 59.215000 58.150000 ;
        RECT 59.015000 58.360000 59.215000 58.560000 ;
        RECT 59.015000 58.770000 59.215000 58.970000 ;
        RECT 59.015000 59.180000 59.215000 59.380000 ;
        RECT 59.015000 59.590000 59.215000 59.790000 ;
        RECT 59.015000 60.000000 59.215000 60.200000 ;
        RECT 59.015000 60.410000 59.215000 60.610000 ;
        RECT 59.420000 56.310000 59.620000 56.510000 ;
        RECT 59.420000 56.720000 59.620000 56.920000 ;
        RECT 59.420000 57.130000 59.620000 57.330000 ;
        RECT 59.420000 57.540000 59.620000 57.740000 ;
        RECT 59.420000 57.950000 59.620000 58.150000 ;
        RECT 59.420000 58.360000 59.620000 58.560000 ;
        RECT 59.420000 58.770000 59.620000 58.970000 ;
        RECT 59.420000 59.180000 59.620000 59.380000 ;
        RECT 59.420000 59.590000 59.620000 59.790000 ;
        RECT 59.420000 60.000000 59.620000 60.200000 ;
        RECT 59.420000 60.410000 59.620000 60.610000 ;
        RECT 59.825000 56.310000 60.025000 56.510000 ;
        RECT 59.825000 56.720000 60.025000 56.920000 ;
        RECT 59.825000 57.130000 60.025000 57.330000 ;
        RECT 59.825000 57.540000 60.025000 57.740000 ;
        RECT 59.825000 57.950000 60.025000 58.150000 ;
        RECT 59.825000 58.360000 60.025000 58.560000 ;
        RECT 59.825000 58.770000 60.025000 58.970000 ;
        RECT 59.825000 59.180000 60.025000 59.380000 ;
        RECT 59.825000 59.590000 60.025000 59.790000 ;
        RECT 59.825000 60.000000 60.025000 60.200000 ;
        RECT 59.825000 60.410000 60.025000 60.610000 ;
        RECT 60.230000 56.310000 60.430000 56.510000 ;
        RECT 60.230000 56.720000 60.430000 56.920000 ;
        RECT 60.230000 57.130000 60.430000 57.330000 ;
        RECT 60.230000 57.540000 60.430000 57.740000 ;
        RECT 60.230000 57.950000 60.430000 58.150000 ;
        RECT 60.230000 58.360000 60.430000 58.560000 ;
        RECT 60.230000 58.770000 60.430000 58.970000 ;
        RECT 60.230000 59.180000 60.430000 59.380000 ;
        RECT 60.230000 59.590000 60.430000 59.790000 ;
        RECT 60.230000 60.000000 60.430000 60.200000 ;
        RECT 60.230000 60.410000 60.430000 60.610000 ;
        RECT 60.635000 56.310000 60.835000 56.510000 ;
        RECT 60.635000 56.720000 60.835000 56.920000 ;
        RECT 60.635000 57.130000 60.835000 57.330000 ;
        RECT 60.635000 57.540000 60.835000 57.740000 ;
        RECT 60.635000 57.950000 60.835000 58.150000 ;
        RECT 60.635000 58.360000 60.835000 58.560000 ;
        RECT 60.635000 58.770000 60.835000 58.970000 ;
        RECT 60.635000 59.180000 60.835000 59.380000 ;
        RECT 60.635000 59.590000 60.835000 59.790000 ;
        RECT 60.635000 60.000000 60.835000 60.200000 ;
        RECT 60.635000 60.410000 60.835000 60.610000 ;
        RECT 61.040000 56.310000 61.240000 56.510000 ;
        RECT 61.040000 56.720000 61.240000 56.920000 ;
        RECT 61.040000 57.130000 61.240000 57.330000 ;
        RECT 61.040000 57.540000 61.240000 57.740000 ;
        RECT 61.040000 57.950000 61.240000 58.150000 ;
        RECT 61.040000 58.360000 61.240000 58.560000 ;
        RECT 61.040000 58.770000 61.240000 58.970000 ;
        RECT 61.040000 59.180000 61.240000 59.380000 ;
        RECT 61.040000 59.590000 61.240000 59.790000 ;
        RECT 61.040000 60.000000 61.240000 60.200000 ;
        RECT 61.040000 60.410000 61.240000 60.610000 ;
        RECT 61.445000 56.310000 61.645000 56.510000 ;
        RECT 61.445000 56.720000 61.645000 56.920000 ;
        RECT 61.445000 57.130000 61.645000 57.330000 ;
        RECT 61.445000 57.540000 61.645000 57.740000 ;
        RECT 61.445000 57.950000 61.645000 58.150000 ;
        RECT 61.445000 58.360000 61.645000 58.560000 ;
        RECT 61.445000 58.770000 61.645000 58.970000 ;
        RECT 61.445000 59.180000 61.645000 59.380000 ;
        RECT 61.445000 59.590000 61.645000 59.790000 ;
        RECT 61.445000 60.000000 61.645000 60.200000 ;
        RECT 61.445000 60.410000 61.645000 60.610000 ;
        RECT 61.850000 56.310000 62.050000 56.510000 ;
        RECT 61.850000 56.720000 62.050000 56.920000 ;
        RECT 61.850000 57.130000 62.050000 57.330000 ;
        RECT 61.850000 57.540000 62.050000 57.740000 ;
        RECT 61.850000 57.950000 62.050000 58.150000 ;
        RECT 61.850000 58.360000 62.050000 58.560000 ;
        RECT 61.850000 58.770000 62.050000 58.970000 ;
        RECT 61.850000 59.180000 62.050000 59.380000 ;
        RECT 61.850000 59.590000 62.050000 59.790000 ;
        RECT 61.850000 60.000000 62.050000 60.200000 ;
        RECT 61.850000 60.410000 62.050000 60.610000 ;
        RECT 62.255000 56.310000 62.455000 56.510000 ;
        RECT 62.255000 56.720000 62.455000 56.920000 ;
        RECT 62.255000 57.130000 62.455000 57.330000 ;
        RECT 62.255000 57.540000 62.455000 57.740000 ;
        RECT 62.255000 57.950000 62.455000 58.150000 ;
        RECT 62.255000 58.360000 62.455000 58.560000 ;
        RECT 62.255000 58.770000 62.455000 58.970000 ;
        RECT 62.255000 59.180000 62.455000 59.380000 ;
        RECT 62.255000 59.590000 62.455000 59.790000 ;
        RECT 62.255000 60.000000 62.455000 60.200000 ;
        RECT 62.255000 60.410000 62.455000 60.610000 ;
        RECT 62.660000 56.310000 62.860000 56.510000 ;
        RECT 62.660000 56.720000 62.860000 56.920000 ;
        RECT 62.660000 57.130000 62.860000 57.330000 ;
        RECT 62.660000 57.540000 62.860000 57.740000 ;
        RECT 62.660000 57.950000 62.860000 58.150000 ;
        RECT 62.660000 58.360000 62.860000 58.560000 ;
        RECT 62.660000 58.770000 62.860000 58.970000 ;
        RECT 62.660000 59.180000 62.860000 59.380000 ;
        RECT 62.660000 59.590000 62.860000 59.790000 ;
        RECT 62.660000 60.000000 62.860000 60.200000 ;
        RECT 62.660000 60.410000 62.860000 60.610000 ;
        RECT 63.065000 56.310000 63.265000 56.510000 ;
        RECT 63.065000 56.720000 63.265000 56.920000 ;
        RECT 63.065000 57.130000 63.265000 57.330000 ;
        RECT 63.065000 57.540000 63.265000 57.740000 ;
        RECT 63.065000 57.950000 63.265000 58.150000 ;
        RECT 63.065000 58.360000 63.265000 58.560000 ;
        RECT 63.065000 58.770000 63.265000 58.970000 ;
        RECT 63.065000 59.180000 63.265000 59.380000 ;
        RECT 63.065000 59.590000 63.265000 59.790000 ;
        RECT 63.065000 60.000000 63.265000 60.200000 ;
        RECT 63.065000 60.410000 63.265000 60.610000 ;
        RECT 63.470000 56.310000 63.670000 56.510000 ;
        RECT 63.470000 56.720000 63.670000 56.920000 ;
        RECT 63.470000 57.130000 63.670000 57.330000 ;
        RECT 63.470000 57.540000 63.670000 57.740000 ;
        RECT 63.470000 57.950000 63.670000 58.150000 ;
        RECT 63.470000 58.360000 63.670000 58.560000 ;
        RECT 63.470000 58.770000 63.670000 58.970000 ;
        RECT 63.470000 59.180000 63.670000 59.380000 ;
        RECT 63.470000 59.590000 63.670000 59.790000 ;
        RECT 63.470000 60.000000 63.670000 60.200000 ;
        RECT 63.470000 60.410000 63.670000 60.610000 ;
        RECT 63.875000 56.310000 64.075000 56.510000 ;
        RECT 63.875000 56.720000 64.075000 56.920000 ;
        RECT 63.875000 57.130000 64.075000 57.330000 ;
        RECT 63.875000 57.540000 64.075000 57.740000 ;
        RECT 63.875000 57.950000 64.075000 58.150000 ;
        RECT 63.875000 58.360000 64.075000 58.560000 ;
        RECT 63.875000 58.770000 64.075000 58.970000 ;
        RECT 63.875000 59.180000 64.075000 59.380000 ;
        RECT 63.875000 59.590000 64.075000 59.790000 ;
        RECT 63.875000 60.000000 64.075000 60.200000 ;
        RECT 63.875000 60.410000 64.075000 60.610000 ;
        RECT 64.280000 56.310000 64.480000 56.510000 ;
        RECT 64.280000 56.720000 64.480000 56.920000 ;
        RECT 64.280000 57.130000 64.480000 57.330000 ;
        RECT 64.280000 57.540000 64.480000 57.740000 ;
        RECT 64.280000 57.950000 64.480000 58.150000 ;
        RECT 64.280000 58.360000 64.480000 58.560000 ;
        RECT 64.280000 58.770000 64.480000 58.970000 ;
        RECT 64.280000 59.180000 64.480000 59.380000 ;
        RECT 64.280000 59.590000 64.480000 59.790000 ;
        RECT 64.280000 60.000000 64.480000 60.200000 ;
        RECT 64.280000 60.410000 64.480000 60.610000 ;
        RECT 64.685000 56.310000 64.885000 56.510000 ;
        RECT 64.685000 56.720000 64.885000 56.920000 ;
        RECT 64.685000 57.130000 64.885000 57.330000 ;
        RECT 64.685000 57.540000 64.885000 57.740000 ;
        RECT 64.685000 57.950000 64.885000 58.150000 ;
        RECT 64.685000 58.360000 64.885000 58.560000 ;
        RECT 64.685000 58.770000 64.885000 58.970000 ;
        RECT 64.685000 59.180000 64.885000 59.380000 ;
        RECT 64.685000 59.590000 64.885000 59.790000 ;
        RECT 64.685000 60.000000 64.885000 60.200000 ;
        RECT 64.685000 60.410000 64.885000 60.610000 ;
        RECT 65.090000 56.310000 65.290000 56.510000 ;
        RECT 65.090000 56.720000 65.290000 56.920000 ;
        RECT 65.090000 57.130000 65.290000 57.330000 ;
        RECT 65.090000 57.540000 65.290000 57.740000 ;
        RECT 65.090000 57.950000 65.290000 58.150000 ;
        RECT 65.090000 58.360000 65.290000 58.560000 ;
        RECT 65.090000 58.770000 65.290000 58.970000 ;
        RECT 65.090000 59.180000 65.290000 59.380000 ;
        RECT 65.090000 59.590000 65.290000 59.790000 ;
        RECT 65.090000 60.000000 65.290000 60.200000 ;
        RECT 65.090000 60.410000 65.290000 60.610000 ;
        RECT 65.495000 56.310000 65.695000 56.510000 ;
        RECT 65.495000 56.720000 65.695000 56.920000 ;
        RECT 65.495000 57.130000 65.695000 57.330000 ;
        RECT 65.495000 57.540000 65.695000 57.740000 ;
        RECT 65.495000 57.950000 65.695000 58.150000 ;
        RECT 65.495000 58.360000 65.695000 58.560000 ;
        RECT 65.495000 58.770000 65.695000 58.970000 ;
        RECT 65.495000 59.180000 65.695000 59.380000 ;
        RECT 65.495000 59.590000 65.695000 59.790000 ;
        RECT 65.495000 60.000000 65.695000 60.200000 ;
        RECT 65.495000 60.410000 65.695000 60.610000 ;
        RECT 65.900000 56.310000 66.100000 56.510000 ;
        RECT 65.900000 56.720000 66.100000 56.920000 ;
        RECT 65.900000 57.130000 66.100000 57.330000 ;
        RECT 65.900000 57.540000 66.100000 57.740000 ;
        RECT 65.900000 57.950000 66.100000 58.150000 ;
        RECT 65.900000 58.360000 66.100000 58.560000 ;
        RECT 65.900000 58.770000 66.100000 58.970000 ;
        RECT 65.900000 59.180000 66.100000 59.380000 ;
        RECT 65.900000 59.590000 66.100000 59.790000 ;
        RECT 65.900000 60.000000 66.100000 60.200000 ;
        RECT 65.900000 60.410000 66.100000 60.610000 ;
        RECT 66.305000 56.310000 66.505000 56.510000 ;
        RECT 66.305000 56.720000 66.505000 56.920000 ;
        RECT 66.305000 57.130000 66.505000 57.330000 ;
        RECT 66.305000 57.540000 66.505000 57.740000 ;
        RECT 66.305000 57.950000 66.505000 58.150000 ;
        RECT 66.305000 58.360000 66.505000 58.560000 ;
        RECT 66.305000 58.770000 66.505000 58.970000 ;
        RECT 66.305000 59.180000 66.505000 59.380000 ;
        RECT 66.305000 59.590000 66.505000 59.790000 ;
        RECT 66.305000 60.000000 66.505000 60.200000 ;
        RECT 66.305000 60.410000 66.505000 60.610000 ;
        RECT 66.710000 56.310000 66.910000 56.510000 ;
        RECT 66.710000 56.720000 66.910000 56.920000 ;
        RECT 66.710000 57.130000 66.910000 57.330000 ;
        RECT 66.710000 57.540000 66.910000 57.740000 ;
        RECT 66.710000 57.950000 66.910000 58.150000 ;
        RECT 66.710000 58.360000 66.910000 58.560000 ;
        RECT 66.710000 58.770000 66.910000 58.970000 ;
        RECT 66.710000 59.180000 66.910000 59.380000 ;
        RECT 66.710000 59.590000 66.910000 59.790000 ;
        RECT 66.710000 60.000000 66.910000 60.200000 ;
        RECT 66.710000 60.410000 66.910000 60.610000 ;
        RECT 67.115000 56.310000 67.315000 56.510000 ;
        RECT 67.115000 56.720000 67.315000 56.920000 ;
        RECT 67.115000 57.130000 67.315000 57.330000 ;
        RECT 67.115000 57.540000 67.315000 57.740000 ;
        RECT 67.115000 57.950000 67.315000 58.150000 ;
        RECT 67.115000 58.360000 67.315000 58.560000 ;
        RECT 67.115000 58.770000 67.315000 58.970000 ;
        RECT 67.115000 59.180000 67.315000 59.380000 ;
        RECT 67.115000 59.590000 67.315000 59.790000 ;
        RECT 67.115000 60.000000 67.315000 60.200000 ;
        RECT 67.115000 60.410000 67.315000 60.610000 ;
        RECT 67.520000 56.310000 67.720000 56.510000 ;
        RECT 67.520000 56.720000 67.720000 56.920000 ;
        RECT 67.520000 57.130000 67.720000 57.330000 ;
        RECT 67.520000 57.540000 67.720000 57.740000 ;
        RECT 67.520000 57.950000 67.720000 58.150000 ;
        RECT 67.520000 58.360000 67.720000 58.560000 ;
        RECT 67.520000 58.770000 67.720000 58.970000 ;
        RECT 67.520000 59.180000 67.720000 59.380000 ;
        RECT 67.520000 59.590000 67.720000 59.790000 ;
        RECT 67.520000 60.000000 67.720000 60.200000 ;
        RECT 67.520000 60.410000 67.720000 60.610000 ;
        RECT 67.925000 56.310000 68.125000 56.510000 ;
        RECT 67.925000 56.720000 68.125000 56.920000 ;
        RECT 67.925000 57.130000 68.125000 57.330000 ;
        RECT 67.925000 57.540000 68.125000 57.740000 ;
        RECT 67.925000 57.950000 68.125000 58.150000 ;
        RECT 67.925000 58.360000 68.125000 58.560000 ;
        RECT 67.925000 58.770000 68.125000 58.970000 ;
        RECT 67.925000 59.180000 68.125000 59.380000 ;
        RECT 67.925000 59.590000 68.125000 59.790000 ;
        RECT 67.925000 60.000000 68.125000 60.200000 ;
        RECT 67.925000 60.410000 68.125000 60.610000 ;
        RECT 68.330000 56.310000 68.530000 56.510000 ;
        RECT 68.330000 56.720000 68.530000 56.920000 ;
        RECT 68.330000 57.130000 68.530000 57.330000 ;
        RECT 68.330000 57.540000 68.530000 57.740000 ;
        RECT 68.330000 57.950000 68.530000 58.150000 ;
        RECT 68.330000 58.360000 68.530000 58.560000 ;
        RECT 68.330000 58.770000 68.530000 58.970000 ;
        RECT 68.330000 59.180000 68.530000 59.380000 ;
        RECT 68.330000 59.590000 68.530000 59.790000 ;
        RECT 68.330000 60.000000 68.530000 60.200000 ;
        RECT 68.330000 60.410000 68.530000 60.610000 ;
        RECT 68.735000 56.310000 68.935000 56.510000 ;
        RECT 68.735000 56.720000 68.935000 56.920000 ;
        RECT 68.735000 57.130000 68.935000 57.330000 ;
        RECT 68.735000 57.540000 68.935000 57.740000 ;
        RECT 68.735000 57.950000 68.935000 58.150000 ;
        RECT 68.735000 58.360000 68.935000 58.560000 ;
        RECT 68.735000 58.770000 68.935000 58.970000 ;
        RECT 68.735000 59.180000 68.935000 59.380000 ;
        RECT 68.735000 59.590000 68.935000 59.790000 ;
        RECT 68.735000 60.000000 68.935000 60.200000 ;
        RECT 68.735000 60.410000 68.935000 60.610000 ;
        RECT 69.140000 56.310000 69.340000 56.510000 ;
        RECT 69.140000 56.720000 69.340000 56.920000 ;
        RECT 69.140000 57.130000 69.340000 57.330000 ;
        RECT 69.140000 57.540000 69.340000 57.740000 ;
        RECT 69.140000 57.950000 69.340000 58.150000 ;
        RECT 69.140000 58.360000 69.340000 58.560000 ;
        RECT 69.140000 58.770000 69.340000 58.970000 ;
        RECT 69.140000 59.180000 69.340000 59.380000 ;
        RECT 69.140000 59.590000 69.340000 59.790000 ;
        RECT 69.140000 60.000000 69.340000 60.200000 ;
        RECT 69.140000 60.410000 69.340000 60.610000 ;
        RECT 69.545000 56.310000 69.745000 56.510000 ;
        RECT 69.545000 56.720000 69.745000 56.920000 ;
        RECT 69.545000 57.130000 69.745000 57.330000 ;
        RECT 69.545000 57.540000 69.745000 57.740000 ;
        RECT 69.545000 57.950000 69.745000 58.150000 ;
        RECT 69.545000 58.360000 69.745000 58.560000 ;
        RECT 69.545000 58.770000 69.745000 58.970000 ;
        RECT 69.545000 59.180000 69.745000 59.380000 ;
        RECT 69.545000 59.590000 69.745000 59.790000 ;
        RECT 69.545000 60.000000 69.745000 60.200000 ;
        RECT 69.545000 60.410000 69.745000 60.610000 ;
        RECT 69.950000 56.310000 70.150000 56.510000 ;
        RECT 69.950000 56.720000 70.150000 56.920000 ;
        RECT 69.950000 57.130000 70.150000 57.330000 ;
        RECT 69.950000 57.540000 70.150000 57.740000 ;
        RECT 69.950000 57.950000 70.150000 58.150000 ;
        RECT 69.950000 58.360000 70.150000 58.560000 ;
        RECT 69.950000 58.770000 70.150000 58.970000 ;
        RECT 69.950000 59.180000 70.150000 59.380000 ;
        RECT 69.950000 59.590000 70.150000 59.790000 ;
        RECT 69.950000 60.000000 70.150000 60.200000 ;
        RECT 69.950000 60.410000 70.150000 60.610000 ;
        RECT 70.355000 56.310000 70.555000 56.510000 ;
        RECT 70.355000 56.720000 70.555000 56.920000 ;
        RECT 70.355000 57.130000 70.555000 57.330000 ;
        RECT 70.355000 57.540000 70.555000 57.740000 ;
        RECT 70.355000 57.950000 70.555000 58.150000 ;
        RECT 70.355000 58.360000 70.555000 58.560000 ;
        RECT 70.355000 58.770000 70.555000 58.970000 ;
        RECT 70.355000 59.180000 70.555000 59.380000 ;
        RECT 70.355000 59.590000 70.555000 59.790000 ;
        RECT 70.355000 60.000000 70.555000 60.200000 ;
        RECT 70.355000 60.410000 70.555000 60.610000 ;
        RECT 70.760000 56.310000 70.960000 56.510000 ;
        RECT 70.760000 56.720000 70.960000 56.920000 ;
        RECT 70.760000 57.130000 70.960000 57.330000 ;
        RECT 70.760000 57.540000 70.960000 57.740000 ;
        RECT 70.760000 57.950000 70.960000 58.150000 ;
        RECT 70.760000 58.360000 70.960000 58.560000 ;
        RECT 70.760000 58.770000 70.960000 58.970000 ;
        RECT 70.760000 59.180000 70.960000 59.380000 ;
        RECT 70.760000 59.590000 70.960000 59.790000 ;
        RECT 70.760000 60.000000 70.960000 60.200000 ;
        RECT 70.760000 60.410000 70.960000 60.610000 ;
        RECT 71.165000 56.310000 71.365000 56.510000 ;
        RECT 71.165000 56.720000 71.365000 56.920000 ;
        RECT 71.165000 57.130000 71.365000 57.330000 ;
        RECT 71.165000 57.540000 71.365000 57.740000 ;
        RECT 71.165000 57.950000 71.365000 58.150000 ;
        RECT 71.165000 58.360000 71.365000 58.560000 ;
        RECT 71.165000 58.770000 71.365000 58.970000 ;
        RECT 71.165000 59.180000 71.365000 59.380000 ;
        RECT 71.165000 59.590000 71.365000 59.790000 ;
        RECT 71.165000 60.000000 71.365000 60.200000 ;
        RECT 71.165000 60.410000 71.365000 60.610000 ;
        RECT 71.570000 56.310000 71.770000 56.510000 ;
        RECT 71.570000 56.720000 71.770000 56.920000 ;
        RECT 71.570000 57.130000 71.770000 57.330000 ;
        RECT 71.570000 57.540000 71.770000 57.740000 ;
        RECT 71.570000 57.950000 71.770000 58.150000 ;
        RECT 71.570000 58.360000 71.770000 58.560000 ;
        RECT 71.570000 58.770000 71.770000 58.970000 ;
        RECT 71.570000 59.180000 71.770000 59.380000 ;
        RECT 71.570000 59.590000 71.770000 59.790000 ;
        RECT 71.570000 60.000000 71.770000 60.200000 ;
        RECT 71.570000 60.410000 71.770000 60.610000 ;
        RECT 71.975000 56.310000 72.175000 56.510000 ;
        RECT 71.975000 56.720000 72.175000 56.920000 ;
        RECT 71.975000 57.130000 72.175000 57.330000 ;
        RECT 71.975000 57.540000 72.175000 57.740000 ;
        RECT 71.975000 57.950000 72.175000 58.150000 ;
        RECT 71.975000 58.360000 72.175000 58.560000 ;
        RECT 71.975000 58.770000 72.175000 58.970000 ;
        RECT 71.975000 59.180000 72.175000 59.380000 ;
        RECT 71.975000 59.590000 72.175000 59.790000 ;
        RECT 71.975000 60.000000 72.175000 60.200000 ;
        RECT 71.975000 60.410000 72.175000 60.610000 ;
        RECT 72.380000 56.310000 72.580000 56.510000 ;
        RECT 72.380000 56.720000 72.580000 56.920000 ;
        RECT 72.380000 57.130000 72.580000 57.330000 ;
        RECT 72.380000 57.540000 72.580000 57.740000 ;
        RECT 72.380000 57.950000 72.580000 58.150000 ;
        RECT 72.380000 58.360000 72.580000 58.560000 ;
        RECT 72.380000 58.770000 72.580000 58.970000 ;
        RECT 72.380000 59.180000 72.580000 59.380000 ;
        RECT 72.380000 59.590000 72.580000 59.790000 ;
        RECT 72.380000 60.000000 72.580000 60.200000 ;
        RECT 72.380000 60.410000 72.580000 60.610000 ;
        RECT 72.785000 56.310000 72.985000 56.510000 ;
        RECT 72.785000 56.720000 72.985000 56.920000 ;
        RECT 72.785000 57.130000 72.985000 57.330000 ;
        RECT 72.785000 57.540000 72.985000 57.740000 ;
        RECT 72.785000 57.950000 72.985000 58.150000 ;
        RECT 72.785000 58.360000 72.985000 58.560000 ;
        RECT 72.785000 58.770000 72.985000 58.970000 ;
        RECT 72.785000 59.180000 72.985000 59.380000 ;
        RECT 72.785000 59.590000 72.985000 59.790000 ;
        RECT 72.785000 60.000000 72.985000 60.200000 ;
        RECT 72.785000 60.410000 72.985000 60.610000 ;
        RECT 73.190000 56.310000 73.390000 56.510000 ;
        RECT 73.190000 56.720000 73.390000 56.920000 ;
        RECT 73.190000 57.130000 73.390000 57.330000 ;
        RECT 73.190000 57.540000 73.390000 57.740000 ;
        RECT 73.190000 57.950000 73.390000 58.150000 ;
        RECT 73.190000 58.360000 73.390000 58.560000 ;
        RECT 73.190000 58.770000 73.390000 58.970000 ;
        RECT 73.190000 59.180000 73.390000 59.380000 ;
        RECT 73.190000 59.590000 73.390000 59.790000 ;
        RECT 73.190000 60.000000 73.390000 60.200000 ;
        RECT 73.190000 60.410000 73.390000 60.610000 ;
        RECT 73.595000 56.310000 73.795000 56.510000 ;
        RECT 73.595000 56.720000 73.795000 56.920000 ;
        RECT 73.595000 57.130000 73.795000 57.330000 ;
        RECT 73.595000 57.540000 73.795000 57.740000 ;
        RECT 73.595000 57.950000 73.795000 58.150000 ;
        RECT 73.595000 58.360000 73.795000 58.560000 ;
        RECT 73.595000 58.770000 73.795000 58.970000 ;
        RECT 73.595000 59.180000 73.795000 59.380000 ;
        RECT 73.595000 59.590000 73.795000 59.790000 ;
        RECT 73.595000 60.000000 73.795000 60.200000 ;
        RECT 73.595000 60.410000 73.795000 60.610000 ;
        RECT 74.000000 56.310000 74.200000 56.510000 ;
        RECT 74.000000 56.720000 74.200000 56.920000 ;
        RECT 74.000000 57.130000 74.200000 57.330000 ;
        RECT 74.000000 57.540000 74.200000 57.740000 ;
        RECT 74.000000 57.950000 74.200000 58.150000 ;
        RECT 74.000000 58.360000 74.200000 58.560000 ;
        RECT 74.000000 58.770000 74.200000 58.970000 ;
        RECT 74.000000 59.180000 74.200000 59.380000 ;
        RECT 74.000000 59.590000 74.200000 59.790000 ;
        RECT 74.000000 60.000000 74.200000 60.200000 ;
        RECT 74.000000 60.410000 74.200000 60.610000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 29.885000 1.270000 33.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 29.885000 75.000000 33.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 29.985000 1.270000 33.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 29.985000 75.000000 33.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met1 ;
      RECT 0.000000 0.000000 75.000000 198.000000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 75.000000 198.000000 ;
    LAYER met3 ;
      RECT  0.000000   0.000000 75.000000  23.440000 ;
      RECT  0.000000  28.880000 75.000000  55.840000 ;
      RECT  0.000000  61.080000 75.000000 170.795000 ;
      RECT 13.300000 170.795000 61.645000 198.000000 ;
      RECT 24.800000  23.440000 50.355000  28.880000 ;
      RECT 24.800000  55.840000 50.355000  61.080000 ;
      RECT 74.690000  23.440000 75.000000  28.880000 ;
      RECT 74.690000  55.840000 75.000000  61.080000 ;
    LAYER met4 ;
      RECT  0.000000   5.885000  1.670000   6.485000 ;
      RECT  0.000000  11.935000  1.365000  12.535000 ;
      RECT  0.000000  16.785000  1.365000  17.385000 ;
      RECT  0.000000  22.835000  1.670000  23.435000 ;
      RECT  0.000000  28.885000  1.670000  29.485000 ;
      RECT  0.000000  33.735000  1.670000  34.335000 ;
      RECT  0.000000  38.585000  1.670000  39.185000 ;
      RECT  0.000000  44.635000  1.670000  45.335000 ;
      RECT  0.000000  55.135000  1.670000  55.835000 ;
      RECT  0.000000  61.085000  1.670000  61.685000 ;
      RECT  0.000000  66.935000  1.670000  67.635000 ;
      RECT  0.000000  93.400000 75.000000 173.385000 ;
      RECT  1.365000  11.935000 73.635000  17.385000 ;
      RECT  1.365000  11.935000 73.635000  17.385000 ;
      RECT  1.670000   0.000000 73.330000  11.935000 ;
      RECT  1.670000   0.000000 73.330000  23.435000 ;
      RECT  1.670000   0.000000 73.330000  23.435000 ;
      RECT  1.670000   0.000000 73.330000  23.435000 ;
      RECT  1.670000  17.385000 73.330000  23.435000 ;
      RECT  1.670000  28.885000 73.330000  55.835000 ;
      RECT  1.670000  28.885000 73.330000  55.835000 ;
      RECT  1.670000  28.885000 73.330000  55.835000 ;
      RECT  1.670000  28.885000 73.330000  55.835000 ;
      RECT  1.670000  28.885000 73.330000  55.835000 ;
      RECT  1.670000  61.085000 73.330000  93.400000 ;
      RECT  1.670000  61.085000 73.330000 173.435000 ;
      RECT  1.670000  61.085000 73.330000 173.435000 ;
      RECT  1.670000  61.085000 73.330000 173.435000 ;
      RECT  1.670000 173.385000 73.330000 173.435000 ;
      RECT 13.300000  61.085000 61.675000 198.000000 ;
      RECT 13.300000 173.435000 61.675000 198.000000 ;
      RECT 24.775000   0.000000 50.380000  61.085000 ;
      RECT 24.775000   0.000000 50.380000 198.000000 ;
      RECT 24.775000  23.435000 50.380000  28.885000 ;
      RECT 24.775000  55.835000 50.380000  61.085000 ;
      RECT 73.330000   5.885000 75.000000   6.485000 ;
      RECT 73.330000  22.835000 75.000000  23.435000 ;
      RECT 73.330000  28.885000 75.000000  29.485000 ;
      RECT 73.330000  33.735000 75.000000  34.335000 ;
      RECT 73.330000  38.585000 75.000000  39.185000 ;
      RECT 73.330000  44.635000 75.000000  45.335000 ;
      RECT 73.330000  55.135000 75.000000  55.835000 ;
      RECT 73.330000  61.085000 75.000000  61.685000 ;
      RECT 73.330000  66.935000 75.000000  67.635000 ;
      RECT 73.635000  11.935000 75.000000  12.535000 ;
      RECT 73.635000  16.785000 75.000000  17.385000 ;
    LAYER met5 ;
      RECT 0.000000  93.785000 75.000000 172.985000 ;
      RECT 1.765000  12.235000 73.235000  17.085000 ;
      RECT 2.070000   0.000000 72.930000  12.235000 ;
      RECT 2.070000  17.085000 72.930000  93.785000 ;
      RECT 2.070000 172.985000 72.930000 198.000000 ;
  END
END sky130_fd_io__overlay_vssio_lvc
END LIBRARY
