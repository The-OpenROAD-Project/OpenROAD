module ram_8x7 (R0_addr,
    R0_en,
    R0_clk,
    R0_data,
    W0_addr,
    W0_en,
    W0_clk,
    W0_data);
 input [2:0] R0_addr;
 input R0_en;
 input R0_clk;
 output [6:0] R0_data;
 input [2:0] W0_addr;
 input W0_en;
 input W0_clk;
 input [6:0] W0_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;

 DFFHQNx1_ASAP7_75t_R \Memory[0][0]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_056_),
    .QN(_055_));
 DFFHQNx1_ASAP7_75t_R \Memory[0][1]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_057_),
    .QN(_054_));
 DFFHQNx1_ASAP7_75t_R \Memory[0][2]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_058_),
    .QN(_053_));
 DFFHQNx1_ASAP7_75t_R \Memory[0][3]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_059_),
    .QN(_052_));
 DFFHQNx1_ASAP7_75t_R \Memory[0][4]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_060_),
    .QN(_051_));
 DFFHQNx1_ASAP7_75t_R \Memory[0][5]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_061_),
    .QN(_050_));
 DFFHQNx1_ASAP7_75t_R \Memory[0][6]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_062_),
    .QN(_049_));
 DFFHQNx1_ASAP7_75t_R \Memory[1][0]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_063_),
    .QN(_048_));
 DFFHQNx1_ASAP7_75t_R \Memory[1][1]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_064_),
    .QN(_047_));
 DFFHQNx1_ASAP7_75t_R \Memory[1][2]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_065_),
    .QN(_046_));
 DFFHQNx1_ASAP7_75t_R \Memory[1][3]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_066_),
    .QN(_045_));
 DFFHQNx1_ASAP7_75t_R \Memory[1][4]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_067_),
    .QN(_044_));
 DFFHQNx1_ASAP7_75t_R \Memory[1][5]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_068_),
    .QN(_043_));
 DFFHQNx1_ASAP7_75t_R \Memory[1][6]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_069_),
    .QN(_042_));
 DFFHQNx1_ASAP7_75t_R \Memory[2][0]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_070_),
    .QN(_041_));
 DFFHQNx1_ASAP7_75t_R \Memory[2][1]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_071_),
    .QN(_040_));
 DFFHQNx1_ASAP7_75t_R \Memory[2][2]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_072_),
    .QN(_039_));
 DFFHQNx1_ASAP7_75t_R \Memory[2][3]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_073_),
    .QN(_038_));
 DFFHQNx1_ASAP7_75t_R \Memory[2][4]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_074_),
    .QN(_037_));
 DFFHQNx1_ASAP7_75t_R \Memory[2][5]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_075_),
    .QN(_036_));
 DFFHQNx1_ASAP7_75t_R \Memory[2][6]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_076_),
    .QN(_035_));
 DFFHQNx1_ASAP7_75t_R \Memory[3][0]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_077_),
    .QN(_034_));
 DFFHQNx1_ASAP7_75t_R \Memory[3][1]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_078_),
    .QN(_033_));
 DFFHQNx1_ASAP7_75t_R \Memory[3][2]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_079_),
    .QN(_032_));
 DFFHQNx1_ASAP7_75t_R \Memory[3][3]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_080_),
    .QN(_031_));
 DFFHQNx1_ASAP7_75t_R \Memory[3][4]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_081_),
    .QN(_030_));
 DFFHQNx1_ASAP7_75t_R \Memory[3][5]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_082_),
    .QN(_029_));
 DFFHQNx1_ASAP7_75t_R \Memory[3][6]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_083_),
    .QN(_028_));
 DFFHQNx1_ASAP7_75t_R \Memory[4][0]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_084_),
    .QN(_027_));
 DFFHQNx1_ASAP7_75t_R \Memory[4][1]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_085_),
    .QN(_026_));
 DFFHQNx1_ASAP7_75t_R \Memory[4][2]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_086_),
    .QN(_025_));
 DFFHQNx1_ASAP7_75t_R \Memory[4][3]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_087_),
    .QN(_024_));
 DFFHQNx1_ASAP7_75t_R \Memory[4][4]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_088_),
    .QN(_023_));
 DFFHQNx1_ASAP7_75t_R \Memory[4][5]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_089_),
    .QN(_022_));
 DFFHQNx1_ASAP7_75t_R \Memory[4][6]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_090_),
    .QN(_021_));
 DFFHQNx1_ASAP7_75t_R \Memory[5][0]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_091_),
    .QN(_020_));
 DFFHQNx1_ASAP7_75t_R \Memory[5][1]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_092_),
    .QN(_019_));
 DFFHQNx1_ASAP7_75t_R \Memory[5][2]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_093_),
    .QN(_018_));
 DFFHQNx1_ASAP7_75t_R \Memory[5][3]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_094_),
    .QN(_017_));
 DFFHQNx1_ASAP7_75t_R \Memory[5][4]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_095_),
    .QN(_016_));
 DFFHQNx1_ASAP7_75t_R \Memory[5][5]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_096_),
    .QN(_015_));
 DFFHQNx1_ASAP7_75t_R \Memory[5][6]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_097_),
    .QN(_014_));
 DFFHQNx1_ASAP7_75t_R \Memory[6][0]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_098_),
    .QN(_013_));
 DFFHQNx1_ASAP7_75t_R \Memory[6][1]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_099_),
    .QN(_012_));
 DFFHQNx1_ASAP7_75t_R \Memory[6][2]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_100_),
    .QN(_011_));
 DFFHQNx1_ASAP7_75t_R \Memory[6][3]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_101_),
    .QN(_010_));
 DFFHQNx1_ASAP7_75t_R \Memory[6][4]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_102_),
    .QN(_009_));
 DFFHQNx1_ASAP7_75t_R \Memory[6][5]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_103_),
    .QN(_008_));
 DFFHQNx1_ASAP7_75t_R \Memory[6][6]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_104_),
    .QN(_007_));
 DFFHQNx1_ASAP7_75t_R \Memory[7][0]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_105_),
    .QN(_006_));
 DFFHQNx1_ASAP7_75t_R \Memory[7][1]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_106_),
    .QN(_005_));
 DFFHQNx1_ASAP7_75t_R \Memory[7][2]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_107_),
    .QN(_004_));
 DFFHQNx1_ASAP7_75t_R \Memory[7][3]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_108_),
    .QN(_003_));
 DFFHQNx1_ASAP7_75t_R \Memory[7][4]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_109_),
    .QN(_002_));
 DFFHQNx1_ASAP7_75t_R \Memory[7][5]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_110_),
    .QN(_001_));
 DFFHQNx1_ASAP7_75t_R \Memory[7][6]$_DFFE_PP_  (.CLK(W0_clk),
    .D(_111_),
    .QN(_000_));
 INVx1_ASAP7_75t_R _284_ (.A(W0_addr[0]),
    .Y(_112_));
 NOR2x1_ASAP7_75t_R _285_ (.A(W0_addr[2]),
    .B(W0_addr[1]),
    .Y(_113_));
 AND3x2_ASAP7_75t_R _286_ (.A(_112_),
    .B(W0_en),
    .C(_113_),
    .Y(_114_));
 BUFx3_ASAP7_75t_R _287_ (.A(_114_),
    .Y(_115_));
 NOR2x1_ASAP7_75t_R _288_ (.A(_055_),
    .B(_115_),
    .Y(_116_));
 AO21x1_ASAP7_75t_R _289_ (.A1(W0_data[0]),
    .A2(_115_),
    .B(_116_),
    .Y(_056_));
 NOR2x1_ASAP7_75t_R _290_ (.A(_054_),
    .B(_115_),
    .Y(_117_));
 AO21x1_ASAP7_75t_R _291_ (.A1(W0_data[1]),
    .A2(_115_),
    .B(_117_),
    .Y(_057_));
 NOR2x1_ASAP7_75t_R _292_ (.A(_053_),
    .B(_115_),
    .Y(_118_));
 AO21x1_ASAP7_75t_R _293_ (.A1(W0_data[2]),
    .A2(_115_),
    .B(_118_),
    .Y(_058_));
 NOR2x1_ASAP7_75t_R _294_ (.A(_052_),
    .B(_114_),
    .Y(_119_));
 AO21x1_ASAP7_75t_R _295_ (.A1(W0_data[3]),
    .A2(_115_),
    .B(_119_),
    .Y(_059_));
 NOR2x1_ASAP7_75t_R _296_ (.A(_051_),
    .B(_114_),
    .Y(_120_));
 AO21x1_ASAP7_75t_R _297_ (.A1(W0_data[4]),
    .A2(_115_),
    .B(_120_),
    .Y(_060_));
 NOR2x1_ASAP7_75t_R _298_ (.A(_050_),
    .B(_114_),
    .Y(_121_));
 AO21x1_ASAP7_75t_R _299_ (.A1(W0_data[5]),
    .A2(_115_),
    .B(_121_),
    .Y(_061_));
 NOR2x1_ASAP7_75t_R _300_ (.A(_049_),
    .B(_114_),
    .Y(_122_));
 AO21x1_ASAP7_75t_R _301_ (.A1(W0_data[6]),
    .A2(_115_),
    .B(_122_),
    .Y(_062_));
 AND3x2_ASAP7_75t_R _302_ (.A(W0_addr[0]),
    .B(W0_en),
    .C(_113_),
    .Y(_123_));
 BUFx3_ASAP7_75t_R _303_ (.A(_123_),
    .Y(_124_));
 NOR2x1_ASAP7_75t_R _304_ (.A(_048_),
    .B(_124_),
    .Y(_125_));
 AO21x1_ASAP7_75t_R _305_ (.A1(W0_data[0]),
    .A2(_124_),
    .B(_125_),
    .Y(_063_));
 NOR2x1_ASAP7_75t_R _306_ (.A(_047_),
    .B(_124_),
    .Y(_126_));
 AO21x1_ASAP7_75t_R _307_ (.A1(W0_data[1]),
    .A2(_124_),
    .B(_126_),
    .Y(_064_));
 NOR2x1_ASAP7_75t_R _308_ (.A(_046_),
    .B(_124_),
    .Y(_127_));
 AO21x1_ASAP7_75t_R _309_ (.A1(W0_data[2]),
    .A2(_124_),
    .B(_127_),
    .Y(_065_));
 NOR2x1_ASAP7_75t_R _310_ (.A(_045_),
    .B(_123_),
    .Y(_128_));
 AO21x1_ASAP7_75t_R _311_ (.A1(W0_data[3]),
    .A2(_124_),
    .B(_128_),
    .Y(_066_));
 NOR2x1_ASAP7_75t_R _312_ (.A(_044_),
    .B(_123_),
    .Y(_129_));
 AO21x1_ASAP7_75t_R _313_ (.A1(W0_data[4]),
    .A2(_124_),
    .B(_129_),
    .Y(_067_));
 NOR2x1_ASAP7_75t_R _314_ (.A(_043_),
    .B(_123_),
    .Y(_130_));
 AO21x1_ASAP7_75t_R _315_ (.A1(W0_data[5]),
    .A2(_124_),
    .B(_130_),
    .Y(_068_));
 NOR2x1_ASAP7_75t_R _316_ (.A(_042_),
    .B(_123_),
    .Y(_131_));
 AO21x1_ASAP7_75t_R _317_ (.A1(W0_data[6]),
    .A2(_124_),
    .B(_131_),
    .Y(_069_));
 INVx2_ASAP7_75t_R _318_ (.A(W0_addr[1]),
    .Y(_132_));
 INVx2_ASAP7_75t_R _319_ (.A(W0_en),
    .Y(_133_));
 OR4x2_ASAP7_75t_R _320_ (.A(W0_addr[2]),
    .B(_132_),
    .C(W0_addr[0]),
    .D(_133_),
    .Y(_134_));
 BUFx6f_ASAP7_75t_R _321_ (.A(_134_),
    .Y(_135_));
 NAND2x1_ASAP7_75t_R _322_ (.A(_041_),
    .B(_135_),
    .Y(_136_));
 OA21x2_ASAP7_75t_R _323_ (.A1(W0_data[0]),
    .A2(_135_),
    .B(_136_),
    .Y(_070_));
 NAND2x1_ASAP7_75t_R _324_ (.A(_040_),
    .B(_135_),
    .Y(_137_));
 OA21x2_ASAP7_75t_R _325_ (.A1(W0_data[1]),
    .A2(_135_),
    .B(_137_),
    .Y(_071_));
 NAND2x1_ASAP7_75t_R _326_ (.A(_039_),
    .B(_135_),
    .Y(_138_));
 OA21x2_ASAP7_75t_R _327_ (.A1(W0_data[2]),
    .A2(_135_),
    .B(_138_),
    .Y(_072_));
 NAND2x1_ASAP7_75t_R _328_ (.A(_038_),
    .B(_134_),
    .Y(_139_));
 OA21x2_ASAP7_75t_R _329_ (.A1(W0_data[3]),
    .A2(_135_),
    .B(_139_),
    .Y(_073_));
 NAND2x1_ASAP7_75t_R _330_ (.A(_037_),
    .B(_134_),
    .Y(_140_));
 OA21x2_ASAP7_75t_R _331_ (.A1(W0_data[4]),
    .A2(_135_),
    .B(_140_),
    .Y(_074_));
 NAND2x1_ASAP7_75t_R _332_ (.A(_036_),
    .B(_134_),
    .Y(_141_));
 OA21x2_ASAP7_75t_R _333_ (.A1(W0_data[5]),
    .A2(_135_),
    .B(_141_),
    .Y(_075_));
 NAND2x1_ASAP7_75t_R _334_ (.A(_035_),
    .B(_134_),
    .Y(_142_));
 OA21x2_ASAP7_75t_R _335_ (.A1(W0_data[6]),
    .A2(_135_),
    .B(_142_),
    .Y(_076_));
 INVx1_ASAP7_75t_R _336_ (.A(W0_addr[2]),
    .Y(_143_));
 AND4x2_ASAP7_75t_R _337_ (.A(_143_),
    .B(W0_addr[1]),
    .C(W0_addr[0]),
    .D(W0_en),
    .Y(_144_));
 BUFx3_ASAP7_75t_R _338_ (.A(_144_),
    .Y(_145_));
 NOR2x1_ASAP7_75t_R _339_ (.A(_034_),
    .B(_145_),
    .Y(_146_));
 AO21x1_ASAP7_75t_R _340_ (.A1(W0_data[0]),
    .A2(_145_),
    .B(_146_),
    .Y(_077_));
 NOR2x1_ASAP7_75t_R _341_ (.A(_033_),
    .B(_145_),
    .Y(_147_));
 AO21x1_ASAP7_75t_R _342_ (.A1(W0_data[1]),
    .A2(_145_),
    .B(_147_),
    .Y(_078_));
 NOR2x1_ASAP7_75t_R _343_ (.A(_032_),
    .B(_145_),
    .Y(_148_));
 AO21x1_ASAP7_75t_R _344_ (.A1(W0_data[2]),
    .A2(_145_),
    .B(_148_),
    .Y(_079_));
 NOR2x1_ASAP7_75t_R _345_ (.A(_031_),
    .B(_144_),
    .Y(_149_));
 AO21x1_ASAP7_75t_R _346_ (.A1(W0_data[3]),
    .A2(_145_),
    .B(_149_),
    .Y(_080_));
 NOR2x1_ASAP7_75t_R _347_ (.A(_030_),
    .B(_144_),
    .Y(_150_));
 AO21x1_ASAP7_75t_R _348_ (.A1(W0_data[4]),
    .A2(_145_),
    .B(_150_),
    .Y(_081_));
 NOR2x1_ASAP7_75t_R _349_ (.A(_029_),
    .B(_144_),
    .Y(_151_));
 AO21x1_ASAP7_75t_R _350_ (.A1(W0_data[5]),
    .A2(_145_),
    .B(_151_),
    .Y(_082_));
 NOR2x1_ASAP7_75t_R _351_ (.A(_028_),
    .B(_144_),
    .Y(_152_));
 AO21x1_ASAP7_75t_R _352_ (.A1(W0_data[6]),
    .A2(_145_),
    .B(_152_),
    .Y(_083_));
 OR4x2_ASAP7_75t_R _353_ (.A(_143_),
    .B(W0_addr[1]),
    .C(W0_addr[0]),
    .D(_133_),
    .Y(_153_));
 BUFx6f_ASAP7_75t_R _354_ (.A(_153_),
    .Y(_154_));
 NAND2x1_ASAP7_75t_R _355_ (.A(_027_),
    .B(_154_),
    .Y(_155_));
 OA21x2_ASAP7_75t_R _356_ (.A1(W0_data[0]),
    .A2(_154_),
    .B(_155_),
    .Y(_084_));
 NAND2x1_ASAP7_75t_R _357_ (.A(_026_),
    .B(_154_),
    .Y(_156_));
 OA21x2_ASAP7_75t_R _358_ (.A1(W0_data[1]),
    .A2(_154_),
    .B(_156_),
    .Y(_085_));
 NAND2x1_ASAP7_75t_R _359_ (.A(_025_),
    .B(_154_),
    .Y(_157_));
 OA21x2_ASAP7_75t_R _360_ (.A1(W0_data[2]),
    .A2(_154_),
    .B(_157_),
    .Y(_086_));
 NAND2x1_ASAP7_75t_R _361_ (.A(_024_),
    .B(_153_),
    .Y(_158_));
 OA21x2_ASAP7_75t_R _362_ (.A1(W0_data[3]),
    .A2(_154_),
    .B(_158_),
    .Y(_087_));
 NAND2x1_ASAP7_75t_R _363_ (.A(_023_),
    .B(_153_),
    .Y(_159_));
 OA21x2_ASAP7_75t_R _364_ (.A1(W0_data[4]),
    .A2(_154_),
    .B(_159_),
    .Y(_088_));
 NAND2x1_ASAP7_75t_R _365_ (.A(_022_),
    .B(_153_),
    .Y(_160_));
 OA21x2_ASAP7_75t_R _366_ (.A1(W0_data[5]),
    .A2(_154_),
    .B(_160_),
    .Y(_089_));
 NAND2x1_ASAP7_75t_R _367_ (.A(_021_),
    .B(_153_),
    .Y(_161_));
 OA21x2_ASAP7_75t_R _368_ (.A1(W0_data[6]),
    .A2(_154_),
    .B(_161_),
    .Y(_090_));
 AND4x2_ASAP7_75t_R _369_ (.A(W0_addr[2]),
    .B(_132_),
    .C(W0_addr[0]),
    .D(W0_en),
    .Y(_162_));
 BUFx3_ASAP7_75t_R _370_ (.A(_162_),
    .Y(_163_));
 NOR2x1_ASAP7_75t_R _371_ (.A(_020_),
    .B(_163_),
    .Y(_164_));
 AO21x1_ASAP7_75t_R _372_ (.A1(W0_data[0]),
    .A2(_163_),
    .B(_164_),
    .Y(_091_));
 NOR2x1_ASAP7_75t_R _373_ (.A(_019_),
    .B(_163_),
    .Y(_165_));
 AO21x1_ASAP7_75t_R _374_ (.A1(W0_data[1]),
    .A2(_163_),
    .B(_165_),
    .Y(_092_));
 NOR2x1_ASAP7_75t_R _375_ (.A(_018_),
    .B(_163_),
    .Y(_166_));
 AO21x1_ASAP7_75t_R _376_ (.A1(W0_data[2]),
    .A2(_163_),
    .B(_166_),
    .Y(_093_));
 NOR2x1_ASAP7_75t_R _377_ (.A(_017_),
    .B(_162_),
    .Y(_167_));
 AO21x1_ASAP7_75t_R _378_ (.A1(W0_data[3]),
    .A2(_163_),
    .B(_167_),
    .Y(_094_));
 NOR2x1_ASAP7_75t_R _379_ (.A(_016_),
    .B(_162_),
    .Y(_168_));
 AO21x1_ASAP7_75t_R _380_ (.A1(W0_data[4]),
    .A2(_163_),
    .B(_168_),
    .Y(_095_));
 NOR2x1_ASAP7_75t_R _381_ (.A(_015_),
    .B(_162_),
    .Y(_169_));
 AO21x1_ASAP7_75t_R _382_ (.A1(W0_data[5]),
    .A2(_163_),
    .B(_169_),
    .Y(_096_));
 NOR2x1_ASAP7_75t_R _383_ (.A(_014_),
    .B(_162_),
    .Y(_170_));
 AO21x1_ASAP7_75t_R _384_ (.A1(W0_data[6]),
    .A2(_163_),
    .B(_170_),
    .Y(_097_));
 OR4x2_ASAP7_75t_R _385_ (.A(_143_),
    .B(_132_),
    .C(W0_addr[0]),
    .D(_133_),
    .Y(_171_));
 BUFx6f_ASAP7_75t_R _386_ (.A(_171_),
    .Y(_172_));
 NAND2x1_ASAP7_75t_R _387_ (.A(_013_),
    .B(_172_),
    .Y(_173_));
 OA21x2_ASAP7_75t_R _388_ (.A1(W0_data[0]),
    .A2(_172_),
    .B(_173_),
    .Y(_098_));
 NAND2x1_ASAP7_75t_R _389_ (.A(_012_),
    .B(_172_),
    .Y(_174_));
 OA21x2_ASAP7_75t_R _390_ (.A1(W0_data[1]),
    .A2(_172_),
    .B(_174_),
    .Y(_099_));
 NAND2x1_ASAP7_75t_R _391_ (.A(_011_),
    .B(_172_),
    .Y(_175_));
 OA21x2_ASAP7_75t_R _392_ (.A1(W0_data[2]),
    .A2(_172_),
    .B(_175_),
    .Y(_100_));
 NAND2x1_ASAP7_75t_R _393_ (.A(_010_),
    .B(_171_),
    .Y(_176_));
 OA21x2_ASAP7_75t_R _394_ (.A1(W0_data[3]),
    .A2(_172_),
    .B(_176_),
    .Y(_101_));
 NAND2x1_ASAP7_75t_R _395_ (.A(_009_),
    .B(_171_),
    .Y(_177_));
 OA21x2_ASAP7_75t_R _396_ (.A1(W0_data[4]),
    .A2(_172_),
    .B(_177_),
    .Y(_102_));
 NAND2x1_ASAP7_75t_R _397_ (.A(_008_),
    .B(_171_),
    .Y(_178_));
 OA21x2_ASAP7_75t_R _398_ (.A1(W0_data[5]),
    .A2(_172_),
    .B(_178_),
    .Y(_103_));
 NAND2x1_ASAP7_75t_R _399_ (.A(_007_),
    .B(_171_),
    .Y(_179_));
 OA21x2_ASAP7_75t_R _400_ (.A1(W0_data[6]),
    .A2(_172_),
    .B(_179_),
    .Y(_104_));
 AND4x1_ASAP7_75t_R _401_ (.A(W0_addr[2]),
    .B(W0_addr[1]),
    .C(W0_addr[0]),
    .D(W0_en),
    .Y(_180_));
 BUFx3_ASAP7_75t_R _402_ (.A(_180_),
    .Y(_181_));
 NOR2x1_ASAP7_75t_R _403_ (.A(_006_),
    .B(_181_),
    .Y(_182_));
 AO21x1_ASAP7_75t_R _404_ (.A1(W0_data[0]),
    .A2(_181_),
    .B(_182_),
    .Y(_105_));
 NOR2x1_ASAP7_75t_R _405_ (.A(_005_),
    .B(_181_),
    .Y(_183_));
 AO21x1_ASAP7_75t_R _406_ (.A1(W0_data[1]),
    .A2(_181_),
    .B(_183_),
    .Y(_106_));
 NOR2x1_ASAP7_75t_R _407_ (.A(_004_),
    .B(_181_),
    .Y(_184_));
 AO21x1_ASAP7_75t_R _408_ (.A1(W0_data[2]),
    .A2(_181_),
    .B(_184_),
    .Y(_107_));
 NOR2x1_ASAP7_75t_R _409_ (.A(_003_),
    .B(_180_),
    .Y(_185_));
 AO21x1_ASAP7_75t_R _410_ (.A1(W0_data[3]),
    .A2(_181_),
    .B(_185_),
    .Y(_108_));
 NOR2x1_ASAP7_75t_R _411_ (.A(_002_),
    .B(_180_),
    .Y(_186_));
 AO21x1_ASAP7_75t_R _412_ (.A1(W0_data[4]),
    .A2(_181_),
    .B(_186_),
    .Y(_109_));
 NOR2x1_ASAP7_75t_R _413_ (.A(_001_),
    .B(_180_),
    .Y(_187_));
 AO21x1_ASAP7_75t_R _414_ (.A1(W0_data[5]),
    .A2(_181_),
    .B(_187_),
    .Y(_110_));
 NOR2x1_ASAP7_75t_R _415_ (.A(_000_),
    .B(_180_),
    .Y(_188_));
 AO21x1_ASAP7_75t_R _416_ (.A1(W0_data[6]),
    .A2(_181_),
    .B(_188_),
    .Y(_111_));
 BUFx6f_ASAP7_75t_R _417_ (.A(R0_addr[0]),
    .Y(_189_));
 BUFx2_ASAP7_75t_R _418_ (.A(_189_),
    .Y(_190_));
 INVx1_ASAP7_75t_R _419_ (.A(_013_),
    .Y(_191_));
 BUFx2_ASAP7_75t_R _420_ (.A(R0_addr[0]),
    .Y(_192_));
 NAND2x1_ASAP7_75t_R _421_ (.A(_192_),
    .B(_006_),
    .Y(_193_));
 AND2x2_ASAP7_75t_R _422_ (.A(R0_addr[1]),
    .B(R0_addr[2]),
    .Y(_194_));
 OA211x2_ASAP7_75t_R _423_ (.A1(_190_),
    .A2(_191_),
    .B(_193_),
    .C(_194_),
    .Y(_195_));
 INVx1_ASAP7_75t_R _424_ (.A(_027_),
    .Y(_196_));
 BUFx12f_ASAP7_75t_R _425_ (.A(_189_),
    .Y(_197_));
 NAND2x1_ASAP7_75t_R _426_ (.A(_197_),
    .B(_020_),
    .Y(_198_));
 INVx1_ASAP7_75t_R _427_ (.A(R0_addr[1]),
    .Y(_199_));
 AND2x2_ASAP7_75t_R _428_ (.A(_199_),
    .B(R0_addr[2]),
    .Y(_200_));
 OA211x2_ASAP7_75t_R _429_ (.A1(_190_),
    .A2(_196_),
    .B(_198_),
    .C(_200_),
    .Y(_201_));
 BUFx2_ASAP7_75t_R _430_ (.A(_189_),
    .Y(_202_));
 INVx1_ASAP7_75t_R _431_ (.A(_041_),
    .Y(_203_));
 BUFx12f_ASAP7_75t_R _432_ (.A(_189_),
    .Y(_204_));
 NAND2x1_ASAP7_75t_R _433_ (.A(_204_),
    .B(_034_),
    .Y(_205_));
 NOR2x1_ASAP7_75t_R _434_ (.A(_199_),
    .B(R0_addr[2]),
    .Y(_206_));
 OA211x2_ASAP7_75t_R _435_ (.A1(_202_),
    .A2(_203_),
    .B(_205_),
    .C(_206_),
    .Y(_207_));
 INVx1_ASAP7_75t_R _436_ (.A(_055_),
    .Y(_208_));
 NAND2x1_ASAP7_75t_R _437_ (.A(_204_),
    .B(_048_),
    .Y(_209_));
 NOR2x1_ASAP7_75t_R _438_ (.A(R0_addr[1]),
    .B(R0_addr[2]),
    .Y(_210_));
 OA211x2_ASAP7_75t_R _439_ (.A1(_192_),
    .A2(_208_),
    .B(_209_),
    .C(_210_),
    .Y(_211_));
 OR4x1_ASAP7_75t_R _440_ (.A(_195_),
    .B(_201_),
    .C(_207_),
    .D(_211_),
    .Y(R0_data[0]));
 INVx1_ASAP7_75t_R _441_ (.A(_012_),
    .Y(_212_));
 NAND2x1_ASAP7_75t_R _442_ (.A(_192_),
    .B(_005_),
    .Y(_213_));
 OA211x2_ASAP7_75t_R _443_ (.A1(_190_),
    .A2(_212_),
    .B(_194_),
    .C(_213_),
    .Y(_214_));
 INVx1_ASAP7_75t_R _444_ (.A(_026_),
    .Y(_215_));
 NAND2x1_ASAP7_75t_R _445_ (.A(_197_),
    .B(_019_),
    .Y(_216_));
 OA211x2_ASAP7_75t_R _446_ (.A1(_190_),
    .A2(_215_),
    .B(_200_),
    .C(_216_),
    .Y(_217_));
 INVx1_ASAP7_75t_R _447_ (.A(_040_),
    .Y(_218_));
 NAND2x1_ASAP7_75t_R _448_ (.A(_204_),
    .B(_033_),
    .Y(_219_));
 OA211x2_ASAP7_75t_R _449_ (.A1(_202_),
    .A2(_218_),
    .B(_206_),
    .C(_219_),
    .Y(_220_));
 INVx1_ASAP7_75t_R _450_ (.A(_054_),
    .Y(_221_));
 NAND2x1_ASAP7_75t_R _451_ (.A(_189_),
    .B(_047_),
    .Y(_222_));
 OA211x2_ASAP7_75t_R _452_ (.A1(_192_),
    .A2(_221_),
    .B(_210_),
    .C(_222_),
    .Y(_223_));
 OR4x1_ASAP7_75t_R _453_ (.A(_214_),
    .B(_217_),
    .C(_220_),
    .D(_223_),
    .Y(R0_data[1]));
 INVx1_ASAP7_75t_R _454_ (.A(_011_),
    .Y(_224_));
 NAND2x1_ASAP7_75t_R _455_ (.A(_197_),
    .B(_004_),
    .Y(_225_));
 OA211x2_ASAP7_75t_R _456_ (.A1(_190_),
    .A2(_224_),
    .B(_194_),
    .C(_225_),
    .Y(_226_));
 INVx1_ASAP7_75t_R _457_ (.A(_025_),
    .Y(_227_));
 NAND2x1_ASAP7_75t_R _458_ (.A(_197_),
    .B(_018_),
    .Y(_228_));
 OA211x2_ASAP7_75t_R _459_ (.A1(_190_),
    .A2(_227_),
    .B(_200_),
    .C(_228_),
    .Y(_229_));
 INVx1_ASAP7_75t_R _460_ (.A(_039_),
    .Y(_230_));
 NAND2x1_ASAP7_75t_R _461_ (.A(_204_),
    .B(_032_),
    .Y(_231_));
 OA211x2_ASAP7_75t_R _462_ (.A1(_202_),
    .A2(_230_),
    .B(_206_),
    .C(_231_),
    .Y(_232_));
 INVx1_ASAP7_75t_R _463_ (.A(_053_),
    .Y(_233_));
 NAND2x1_ASAP7_75t_R _464_ (.A(_189_),
    .B(_046_),
    .Y(_234_));
 OA211x2_ASAP7_75t_R _465_ (.A1(_192_),
    .A2(_233_),
    .B(_210_),
    .C(_234_),
    .Y(_235_));
 OR4x1_ASAP7_75t_R _466_ (.A(_226_),
    .B(_229_),
    .C(_232_),
    .D(_235_),
    .Y(R0_data[2]));
 INVx1_ASAP7_75t_R _467_ (.A(_010_),
    .Y(_236_));
 NAND2x1_ASAP7_75t_R _468_ (.A(_197_),
    .B(_003_),
    .Y(_237_));
 OA211x2_ASAP7_75t_R _469_ (.A1(_190_),
    .A2(_236_),
    .B(_194_),
    .C(_237_),
    .Y(_238_));
 INVx1_ASAP7_75t_R _470_ (.A(_024_),
    .Y(_239_));
 NAND2x1_ASAP7_75t_R _471_ (.A(_197_),
    .B(_017_),
    .Y(_240_));
 OA211x2_ASAP7_75t_R _472_ (.A1(_202_),
    .A2(_239_),
    .B(_200_),
    .C(_240_),
    .Y(_241_));
 INVx1_ASAP7_75t_R _473_ (.A(_038_),
    .Y(_242_));
 NAND2x1_ASAP7_75t_R _474_ (.A(_204_),
    .B(_031_),
    .Y(_243_));
 OA211x2_ASAP7_75t_R _475_ (.A1(_202_),
    .A2(_242_),
    .B(_206_),
    .C(_243_),
    .Y(_244_));
 INVx1_ASAP7_75t_R _476_ (.A(_052_),
    .Y(_245_));
 NAND2x1_ASAP7_75t_R _477_ (.A(_189_),
    .B(_045_),
    .Y(_246_));
 OA211x2_ASAP7_75t_R _478_ (.A1(_192_),
    .A2(_245_),
    .B(_210_),
    .C(_246_),
    .Y(_247_));
 OR4x1_ASAP7_75t_R _479_ (.A(_238_),
    .B(_241_),
    .C(_244_),
    .D(_247_),
    .Y(R0_data[3]));
 INVx1_ASAP7_75t_R _480_ (.A(_009_),
    .Y(_248_));
 NAND2x1_ASAP7_75t_R _481_ (.A(_197_),
    .B(_002_),
    .Y(_249_));
 OA211x2_ASAP7_75t_R _482_ (.A1(_190_),
    .A2(_248_),
    .B(_194_),
    .C(_249_),
    .Y(_250_));
 INVx1_ASAP7_75t_R _483_ (.A(_023_),
    .Y(_251_));
 NAND2x1_ASAP7_75t_R _484_ (.A(_197_),
    .B(_016_),
    .Y(_252_));
 OA211x2_ASAP7_75t_R _485_ (.A1(_202_),
    .A2(_251_),
    .B(_200_),
    .C(_252_),
    .Y(_253_));
 INVx1_ASAP7_75t_R _486_ (.A(_037_),
    .Y(_254_));
 NAND2x1_ASAP7_75t_R _487_ (.A(_204_),
    .B(_030_),
    .Y(_255_));
 OA211x2_ASAP7_75t_R _488_ (.A1(_202_),
    .A2(_254_),
    .B(_206_),
    .C(_255_),
    .Y(_256_));
 INVx1_ASAP7_75t_R _489_ (.A(_051_),
    .Y(_257_));
 NAND2x1_ASAP7_75t_R _490_ (.A(_189_),
    .B(_044_),
    .Y(_258_));
 OA211x2_ASAP7_75t_R _491_ (.A1(_192_),
    .A2(_257_),
    .B(_210_),
    .C(_258_),
    .Y(_259_));
 OR4x1_ASAP7_75t_R _492_ (.A(_250_),
    .B(_253_),
    .C(_256_),
    .D(_259_),
    .Y(R0_data[4]));
 INVx1_ASAP7_75t_R _493_ (.A(_008_),
    .Y(_260_));
 NAND2x1_ASAP7_75t_R _494_ (.A(_197_),
    .B(_001_),
    .Y(_261_));
 OA211x2_ASAP7_75t_R _495_ (.A1(_190_),
    .A2(_260_),
    .B(_194_),
    .C(_261_),
    .Y(_262_));
 INVx1_ASAP7_75t_R _496_ (.A(_022_),
    .Y(_263_));
 NAND2x1_ASAP7_75t_R _497_ (.A(_204_),
    .B(_015_),
    .Y(_264_));
 OA211x2_ASAP7_75t_R _498_ (.A1(_202_),
    .A2(_263_),
    .B(_200_),
    .C(_264_),
    .Y(_265_));
 INVx1_ASAP7_75t_R _499_ (.A(_036_),
    .Y(_266_));
 NAND2x1_ASAP7_75t_R _500_ (.A(_204_),
    .B(_029_),
    .Y(_267_));
 OA211x2_ASAP7_75t_R _501_ (.A1(_202_),
    .A2(_266_),
    .B(_206_),
    .C(_267_),
    .Y(_268_));
 INVx1_ASAP7_75t_R _502_ (.A(_050_),
    .Y(_269_));
 NAND2x1_ASAP7_75t_R _503_ (.A(_189_),
    .B(_043_),
    .Y(_270_));
 OA211x2_ASAP7_75t_R _504_ (.A1(_192_),
    .A2(_269_),
    .B(_210_),
    .C(_270_),
    .Y(_271_));
 OR4x1_ASAP7_75t_R _505_ (.A(_262_),
    .B(_265_),
    .C(_268_),
    .D(_271_),
    .Y(R0_data[5]));
 INVx1_ASAP7_75t_R _506_ (.A(_007_),
    .Y(_272_));
 NAND2x1_ASAP7_75t_R _507_ (.A(_197_),
    .B(_000_),
    .Y(_273_));
 OA211x2_ASAP7_75t_R _508_ (.A1(_190_),
    .A2(_272_),
    .B(_194_),
    .C(_273_),
    .Y(_274_));
 INVx1_ASAP7_75t_R _509_ (.A(_021_),
    .Y(_275_));
 NAND2x1_ASAP7_75t_R _510_ (.A(_204_),
    .B(_014_),
    .Y(_276_));
 OA211x2_ASAP7_75t_R _511_ (.A1(_202_),
    .A2(_275_),
    .B(_200_),
    .C(_276_),
    .Y(_277_));
 INVx1_ASAP7_75t_R _512_ (.A(_035_),
    .Y(_278_));
 NAND2x1_ASAP7_75t_R _513_ (.A(_204_),
    .B(_028_),
    .Y(_279_));
 OA211x2_ASAP7_75t_R _514_ (.A1(_192_),
    .A2(_278_),
    .B(_206_),
    .C(_279_),
    .Y(_280_));
 INVx1_ASAP7_75t_R _515_ (.A(_049_),
    .Y(_281_));
 NAND2x1_ASAP7_75t_R _516_ (.A(_189_),
    .B(_042_),
    .Y(_282_));
 OA211x2_ASAP7_75t_R _517_ (.A1(_192_),
    .A2(_281_),
    .B(_210_),
    .C(_282_),
    .Y(_283_));
 OR4x1_ASAP7_75t_R _518_ (.A(_274_),
    .B(_277_),
    .C(_280_),
    .D(_283_),
    .Y(R0_data[6]));
endmodule
