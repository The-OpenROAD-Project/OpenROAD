module gcd (clk,
    req_rdy,
    req_val,
    reset,
    resp_rdy,
    resp_val,
    req_msg,
    resp_msg);
 input clk;
 output req_rdy;
 input req_val;
 input reset;
 input resp_rdy;
 output resp_val;
 input [31:0] req_msg;
 output [15:0] resp_msg;

 INV_X1 _440_ (.A(_109_),
    .ZN(_142_));
 AND3_X1 _441_ (.A1(_142_),
    .A2(_108_),
    .A3(_059_),
    .ZN(_423_));
 XOR2_X1 _442_ (.A(_110_),
    .B(_126_),
    .Z(_406_));
 NOR4_X1 _443_ (.A1(_139_),
    .A2(_138_),
    .A3(_137_),
    .A4(_136_),
    .ZN(_143_));
 INV_X1 _444_ (.A(_135_),
    .ZN(_144_));
 INV_X1 _445_ (.A(_134_),
    .ZN(_145_));
 NOR2_X1 _446_ (.A1(_133_),
    .A2(_126_),
    .ZN(_146_));
 NAND4_X1 _447_ (.A1(_143_),
    .A2(_144_),
    .A3(_145_),
    .A4(_146_),
    .ZN(_147_));
 NOR4_X1 _448_ (.A1(_128_),
    .A2(_127_),
    .A3(_141_),
    .A4(_140_),
    .ZN(_148_));
 NOR4_X1 _449_ (.A1(_132_),
    .A2(_131_),
    .A3(_130_),
    .A4(_129_),
    .ZN(_149_));
 NAND2_X1 _450_ (.A1(_148_),
    .A2(_149_),
    .ZN(_150_));
 NOR2_X1 _451_ (.A1(_147_),
    .A2(_150_),
    .ZN(_151_));
 INV_X1 _452_ (.A(_405_),
    .ZN(_152_));
 INV_X1 _453_ (.A(_058_),
    .ZN(_153_));
 NAND3_X1 _454_ (.A1(_151_),
    .A2(_152_),
    .A3(_153_),
    .ZN(_154_));
 AND2_X1 _455_ (.A1(_423_),
    .A2(_422_),
    .ZN(_155_));
 OR3_X1 _456_ (.A1(_155_),
    .A2(_405_),
    .A3(_057_),
    .ZN(_156_));
 NAND2_X1 _457_ (.A1(_154_),
    .A2(_156_),
    .ZN(_055_));
 OAI211_X2 _458_ (.A(_152_),
    .B(_153_),
    .C1(_147_),
    .C2(_150_),
    .ZN(_157_));
 INV_X2 _459_ (.A(_059_),
    .ZN(_158_));
 BUF_X4 _460_ (.A(_158_),
    .Z(_159_));
 BUF_X4 _461_ (.A(_403_),
    .Z(_160_));
 NAND4_X1 _462_ (.A1(_152_),
    .A2(_159_),
    .A3(_160_),
    .A4(_404_),
    .ZN(_161_));
 NAND2_X1 _463_ (.A1(_157_),
    .A2(_161_),
    .ZN(_056_));
 NAND3_X1 _464_ (.A1(_423_),
    .A2(_152_),
    .A3(_422_),
    .ZN(_162_));
 NOR2_X1 _465_ (.A1(_162_),
    .A2(_057_),
    .ZN(_163_));
 AOI211_X4 _466_ (.A(_405_),
    .B(_059_),
    .C1(_403_),
    .C2(_404_),
    .ZN(_164_));
 OR3_X1 _467_ (.A1(_163_),
    .A2(_405_),
    .A3(_164_),
    .ZN(_054_));
 BUF_X4 _468_ (.A(_142_),
    .Z(_165_));
 OAI21_X1 _469_ (.A(_378_),
    .B1(_165_),
    .B2(_159_),
    .ZN(_166_));
 INV_X1 _470_ (.A(_116_),
    .ZN(_167_));
 NAND2_X1 _471_ (.A1(_167_),
    .A2(_132_),
    .ZN(_168_));
 XNOR2_X2 _472_ (.A(_123_),
    .B(_139_),
    .ZN(_169_));
 XNOR2_X2 _473_ (.A(_122_),
    .B(_138_),
    .ZN(_170_));
 AND2_X4 _474_ (.A1(_169_),
    .A2(_170_),
    .ZN(_171_));
 XNOR2_X2 _475_ (.A(_119_),
    .B(_135_),
    .ZN(_172_));
 XNOR2_X2 _476_ (.A(_118_),
    .B(_134_),
    .ZN(_173_));
 AND2_X2 _477_ (.A1(_172_),
    .A2(_173_),
    .ZN(_174_));
 XNOR2_X2 _478_ (.A(_121_),
    .B(_137_),
    .ZN(_175_));
 XNOR2_X2 _479_ (.A(_120_),
    .B(_136_),
    .ZN(_176_));
 AND2_X4 _480_ (.A1(_175_),
    .A2(_176_),
    .ZN(_177_));
 NAND3_X2 _481_ (.A1(_171_),
    .A2(_174_),
    .A3(_177_),
    .ZN(_178_));
 INV_X4 _482_ (.A(_133_),
    .ZN(_179_));
 AND2_X1 _483_ (.A1(_179_),
    .A2(_117_),
    .ZN(_180_));
 NOR2_X1 _484_ (.A1(_179_),
    .A2(_117_),
    .ZN(_181_));
 INV_X1 _485_ (.A(_110_),
    .ZN(_182_));
 NOR3_X1 _486_ (.A1(_181_),
    .A2(_182_),
    .A3(_126_),
    .ZN(_183_));
 OR3_X4 _487_ (.A1(_178_),
    .A2(_180_),
    .A3(_183_),
    .ZN(_184_));
 INV_X1 _488_ (.A(_120_),
    .ZN(_185_));
 AND3_X1 _489_ (.A1(_175_),
    .A2(_185_),
    .A3(_136_),
    .ZN(_186_));
 INV_X1 _490_ (.A(_121_),
    .ZN(_187_));
 AND2_X1 _491_ (.A1(_187_),
    .A2(_137_),
    .ZN(_188_));
 OAI21_X1 _492_ (.A(_171_),
    .B1(_186_),
    .B2(_188_),
    .ZN(_189_));
 INV_X1 _493_ (.A(_139_),
    .ZN(_190_));
 NOR2_X1 _494_ (.A1(_190_),
    .A2(_123_),
    .ZN(_191_));
 INV_X1 _495_ (.A(_191_),
    .ZN(_192_));
 INV_X1 _496_ (.A(_122_),
    .ZN(_193_));
 NAND3_X1 _497_ (.A1(_169_),
    .A2(_193_),
    .A3(_138_),
    .ZN(_194_));
 AND3_X1 _498_ (.A1(_189_),
    .A2(_192_),
    .A3(_194_),
    .ZN(_195_));
 NOR2_X1 _499_ (.A1(_144_),
    .A2(_119_),
    .ZN(_196_));
 AOI211_X4 _500_ (.A(_118_),
    .B(_145_),
    .C1(_119_),
    .C2(_144_),
    .ZN(_197_));
 OAI211_X2 _501_ (.A(_171_),
    .B(_177_),
    .C1(_196_),
    .C2(_197_),
    .ZN(_198_));
 NAND3_X1 _502_ (.A1(_184_),
    .A2(_195_),
    .A3(_198_),
    .ZN(_199_));
 XNOR2_X2 _503_ (.A(_111_),
    .B(_127_),
    .ZN(_200_));
 XNOR2_X2 _504_ (.A(_112_),
    .B(_128_),
    .ZN(_201_));
 AND2_X1 _505_ (.A1(_200_),
    .A2(_201_),
    .ZN(_202_));
 XNOR2_X1 _506_ (.A(_125_),
    .B(_141_),
    .ZN(_203_));
 XNOR2_X1 _507_ (.A(_124_),
    .B(_140_),
    .ZN(_204_));
 AND3_X1 _508_ (.A1(_202_),
    .A2(_203_),
    .A3(_204_),
    .ZN(_205_));
 XNOR2_X1 _509_ (.A(_115_),
    .B(_131_),
    .ZN(_206_));
 XNOR2_X1 _510_ (.A(_116_),
    .B(_132_),
    .ZN(_207_));
 NAND2_X1 _511_ (.A1(_206_),
    .A2(_207_),
    .ZN(_208_));
 XNOR2_X1 _512_ (.A(_114_),
    .B(_130_),
    .ZN(_209_));
 INV_X1 _513_ (.A(_209_),
    .ZN(_210_));
 XNOR2_X2 _514_ (.A(_113_),
    .B(_129_),
    .ZN(_211_));
 INV_X1 _515_ (.A(_211_),
    .ZN(_212_));
 NOR3_X2 _516_ (.A1(_208_),
    .A2(_210_),
    .A3(_212_),
    .ZN(_213_));
 AND2_X4 _517_ (.A1(_205_),
    .A2(_213_),
    .ZN(_214_));
 NAND2_X1 _518_ (.A1(_199_),
    .A2(_214_),
    .ZN(_215_));
 INV_X1 _519_ (.A(_124_),
    .ZN(_216_));
 AND3_X1 _520_ (.A1(_203_),
    .A2(_216_),
    .A3(_140_),
    .ZN(_217_));
 INV_X1 _521_ (.A(_125_),
    .ZN(_218_));
 AND2_X1 _522_ (.A1(_218_),
    .A2(_141_),
    .ZN(_219_));
 OAI21_X1 _523_ (.A(_202_),
    .B1(_217_),
    .B2(_219_),
    .ZN(_220_));
 INV_X1 _524_ (.A(_112_),
    .ZN(_221_));
 NOR2_X1 _525_ (.A1(_221_),
    .A2(_128_),
    .ZN(_222_));
 INV_X1 _526_ (.A(_111_),
    .ZN(_223_));
 AOI22_X1 _527_ (.A1(_221_),
    .A2(_128_),
    .B1(_223_),
    .B2(_127_),
    .ZN(_224_));
 OAI21_X1 _528_ (.A(_220_),
    .B1(_222_),
    .B2(_224_),
    .ZN(_225_));
 NAND2_X1 _529_ (.A1(_225_),
    .A2(_213_),
    .ZN(_226_));
 INV_X1 _530_ (.A(_115_),
    .ZN(_227_));
 NAND3_X1 _531_ (.A1(_207_),
    .A2(_227_),
    .A3(_131_),
    .ZN(_228_));
 AND4_X4 _532_ (.A1(_168_),
    .A2(_215_),
    .A3(_226_),
    .A4(_228_),
    .ZN(_229_));
 AND2_X1 _533_ (.A1(_109_),
    .A2(_059_),
    .ZN(_230_));
 INV_X1 _534_ (.A(_114_),
    .ZN(_231_));
 NOR2_X1 _535_ (.A1(_231_),
    .A2(_130_),
    .ZN(_232_));
 INV_X1 _536_ (.A(_113_),
    .ZN(_233_));
 AOI22_X1 _537_ (.A1(_231_),
    .A2(_130_),
    .B1(_233_),
    .B2(_129_),
    .ZN(_234_));
 OR3_X1 _538_ (.A1(_208_),
    .A2(_232_),
    .A3(_234_),
    .ZN(_235_));
 NAND4_X1 _539_ (.A1(_229_),
    .A2(_406_),
    .A3(_230_),
    .A4(_235_),
    .ZN(_236_));
 AND2_X1 _540_ (.A1(_171_),
    .A2(_177_),
    .ZN(_237_));
 NAND4_X1 _541_ (.A1(_205_),
    .A2(_237_),
    .A3(_213_),
    .A4(_174_),
    .ZN(_238_));
 XNOR2_X1 _542_ (.A(_117_),
    .B(_133_),
    .ZN(_239_));
 INV_X1 _543_ (.A(_239_),
    .ZN(_240_));
 NOR3_X2 _544_ (.A1(_238_),
    .A2(_406_),
    .A3(_240_),
    .ZN(_241_));
 AOI21_X4 _545_ (.A(_241_),
    .B1(_229_),
    .B2(_235_),
    .ZN(_242_));
 NAND2_X4 _546_ (.A1(_242_),
    .A2(_109_),
    .ZN(_243_));
 OR2_X4 _547_ (.A1(_243_),
    .A2(_158_),
    .ZN(_244_));
 BUF_X16 _548_ (.A(_244_),
    .Z(_245_));
 BUF_X32 _549_ (.A(_245_),
    .Z(_246_));
 OAI211_X2 _550_ (.A(_166_),
    .B(_236_),
    .C1(_246_),
    .C2(_060_),
    .ZN(_247_));
 OR2_X1 _551_ (.A1(_109_),
    .A2(_403_),
    .ZN(_248_));
 BUF_X4 _552_ (.A(_248_),
    .Z(_249_));
 BUF_X4 _553_ (.A(_249_),
    .Z(_250_));
 MUX2_X1 _554_ (.A(_110_),
    .B(_247_),
    .S(_250_),
    .Z(_076_));
 OAI21_X1 _555_ (.A(_379_),
    .B1(_165_),
    .B2(_159_),
    .ZN(_251_));
 INV_X1 _556_ (.A(_230_),
    .ZN(_252_));
 NOR2_X4 _557_ (.A1(_242_),
    .A2(_252_),
    .ZN(_253_));
 BUF_X2 _558_ (.A(_253_),
    .Z(_254_));
 NAND2_X1 _559_ (.A1(_182_),
    .A2(_126_),
    .ZN(_255_));
 XOR2_X1 _560_ (.A(_239_),
    .B(_255_),
    .Z(_413_));
 NAND2_X1 _561_ (.A1(_254_),
    .A2(_413_),
    .ZN(_256_));
 OAI211_X2 _562_ (.A(_251_),
    .B(_256_),
    .C1(_246_),
    .C2(_061_),
    .ZN(_257_));
 MUX2_X1 _563_ (.A(_117_),
    .B(_257_),
    .S(_250_),
    .Z(_083_));
 OAI21_X1 _564_ (.A(_380_),
    .B1(_165_),
    .B2(_159_),
    .ZN(_258_));
 AOI21_X1 _565_ (.A(_180_),
    .B1(_239_),
    .B2(_255_),
    .ZN(_259_));
 XNOR2_X1 _566_ (.A(_259_),
    .B(_173_),
    .ZN(_414_));
 NAND2_X1 _567_ (.A1(_254_),
    .A2(_414_),
    .ZN(_260_));
 OAI211_X2 _568_ (.A(_258_),
    .B(_260_),
    .C1(_246_),
    .C2(_062_),
    .ZN(_261_));
 MUX2_X1 _569_ (.A(_118_),
    .B(_261_),
    .S(_250_),
    .Z(_084_));
 OAI21_X1 _570_ (.A(_381_),
    .B1(_165_),
    .B2(_159_),
    .ZN(_262_));
 INV_X1 _571_ (.A(_259_),
    .ZN(_263_));
 AND2_X1 _572_ (.A1(_263_),
    .A2(_173_),
    .ZN(_264_));
 AND2_X1 _573_ (.A1(_145_),
    .A2(_118_),
    .ZN(_265_));
 NOR2_X1 _574_ (.A1(_264_),
    .A2(_265_),
    .ZN(_266_));
 XNOR2_X1 _575_ (.A(_266_),
    .B(_172_),
    .ZN(_415_));
 NAND2_X1 _576_ (.A1(_254_),
    .A2(_415_),
    .ZN(_267_));
 OAI211_X2 _577_ (.A(_262_),
    .B(_267_),
    .C1(_246_),
    .C2(_063_),
    .ZN(_268_));
 MUX2_X1 _578_ (.A(_119_),
    .B(_268_),
    .S(_250_),
    .Z(_085_));
 OAI21_X1 _579_ (.A(_383_),
    .B1(_165_),
    .B2(_159_),
    .ZN(_269_));
 AND2_X1 _580_ (.A1(_172_),
    .A2(_265_),
    .ZN(_270_));
 AOI21_X4 _581_ (.A(_270_),
    .B1(_119_),
    .B2(_144_),
    .ZN(_271_));
 NAND2_X1 _582_ (.A1(_263_),
    .A2(_174_),
    .ZN(_272_));
 NAND2_X2 _583_ (.A1(_271_),
    .A2(_272_),
    .ZN(_273_));
 XOR2_X1 _584_ (.A(_273_),
    .B(_176_),
    .Z(_416_));
 NAND2_X1 _585_ (.A1(_254_),
    .A2(_416_),
    .ZN(_274_));
 OAI211_X2 _586_ (.A(_269_),
    .B(_274_),
    .C1(_246_),
    .C2(_064_),
    .ZN(_275_));
 MUX2_X1 _587_ (.A(_120_),
    .B(_275_),
    .S(_250_),
    .Z(_086_));
 OAI21_X1 _588_ (.A(_384_),
    .B1(_165_),
    .B2(_159_),
    .ZN(_276_));
 AND2_X1 _589_ (.A1(_273_),
    .A2(_176_),
    .ZN(_277_));
 NOR2_X1 _590_ (.A1(_185_),
    .A2(_136_),
    .ZN(_278_));
 NOR3_X1 _591_ (.A1(_277_),
    .A2(_175_),
    .A3(_278_),
    .ZN(_279_));
 AOI221_X4 _592_ (.A(_279_),
    .B1(_175_),
    .B2(_278_),
    .C1(_177_),
    .C2(_273_),
    .ZN(_417_));
 NAND2_X1 _593_ (.A1(_254_),
    .A2(_417_),
    .ZN(_280_));
 OAI211_X2 _594_ (.A(_276_),
    .B(_280_),
    .C1(_246_),
    .C2(_065_),
    .ZN(_281_));
 MUX2_X1 _595_ (.A(_121_),
    .B(_281_),
    .S(_250_),
    .Z(_087_));
 OAI21_X1 _596_ (.A(_385_),
    .B1(_165_),
    .B2(_159_),
    .ZN(_282_));
 NAND2_X1 _597_ (.A1(_175_),
    .A2(_278_),
    .ZN(_283_));
 OAI21_X1 _598_ (.A(_283_),
    .B1(_187_),
    .B2(_137_),
    .ZN(_284_));
 AOI21_X1 _599_ (.A(_284_),
    .B1(_273_),
    .B2(_177_),
    .ZN(_285_));
 XNOR2_X1 _600_ (.A(_285_),
    .B(_170_),
    .ZN(_418_));
 NAND2_X1 _601_ (.A1(_254_),
    .A2(_418_),
    .ZN(_286_));
 OAI211_X2 _602_ (.A(_282_),
    .B(_286_),
    .C1(_246_),
    .C2(_066_),
    .ZN(_287_));
 MUX2_X1 _603_ (.A(_122_),
    .B(_287_),
    .S(_249_),
    .Z(_088_));
 OAI21_X1 _604_ (.A(_386_),
    .B1(_165_),
    .B2(_158_),
    .ZN(_288_));
 AND2_X1 _605_ (.A1(_193_),
    .A2(_138_),
    .ZN(_289_));
 NOR2_X1 _606_ (.A1(_193_),
    .A2(_138_),
    .ZN(_290_));
 NOR3_X1 _607_ (.A1(_285_),
    .A2(_289_),
    .A3(_290_),
    .ZN(_291_));
 NOR2_X1 _608_ (.A1(_291_),
    .A2(_290_),
    .ZN(_292_));
 XNOR2_X1 _609_ (.A(_292_),
    .B(_169_),
    .ZN(_419_));
 NAND2_X1 _610_ (.A1(_254_),
    .A2(_419_),
    .ZN(_293_));
 OAI211_X2 _611_ (.A(_288_),
    .B(_293_),
    .C1(_246_),
    .C2(_067_),
    .ZN(_294_));
 MUX2_X1 _612_ (.A(_123_),
    .B(_294_),
    .S(_249_),
    .Z(_089_));
 OAI21_X1 _613_ (.A(_387_),
    .B1(_142_),
    .B2(_158_),
    .ZN(_295_));
 NAND2_X2 _614_ (.A1(_273_),
    .A2(_237_),
    .ZN(_296_));
 AND2_X1 _615_ (.A1(_169_),
    .A2(_290_),
    .ZN(_297_));
 AOI221_X2 _616_ (.A(_297_),
    .B1(_123_),
    .B2(_190_),
    .C1(_284_),
    .C2(_171_),
    .ZN(_298_));
 NAND2_X2 _617_ (.A1(_296_),
    .A2(_298_),
    .ZN(_299_));
 XOR2_X1 _618_ (.A(_299_),
    .B(_204_),
    .Z(_420_));
 NAND2_X1 _619_ (.A1(_254_),
    .A2(_420_),
    .ZN(_300_));
 OAI211_X2 _620_ (.A(_295_),
    .B(_300_),
    .C1(_246_),
    .C2(_068_),
    .ZN(_301_));
 MUX2_X1 _621_ (.A(_124_),
    .B(_301_),
    .S(_249_),
    .Z(_090_));
 AND3_X1 _622_ (.A1(_299_),
    .A2(_203_),
    .A3(_204_),
    .ZN(_302_));
 AND2_X1 _623_ (.A1(_299_),
    .A2(_204_),
    .ZN(_303_));
 NOR2_X1 _624_ (.A1(_216_),
    .A2(_140_),
    .ZN(_304_));
 NOR3_X1 _625_ (.A1(_303_),
    .A2(_203_),
    .A3(_304_),
    .ZN(_305_));
 AOI211_X4 _626_ (.A(_302_),
    .B(_305_),
    .C1(_203_),
    .C2(_304_),
    .ZN(_421_));
 NAND2_X1 _627_ (.A1(_421_),
    .A2(_253_),
    .ZN(_306_));
 OAI21_X1 _628_ (.A(_388_),
    .B1(_142_),
    .B2(_158_),
    .ZN(_307_));
 OAI211_X2 _629_ (.A(_306_),
    .B(_307_),
    .C1(_245_),
    .C2(_069_),
    .ZN(_308_));
 MUX2_X1 _630_ (.A(_125_),
    .B(_308_),
    .S(_249_),
    .Z(_091_));
 OAI21_X1 _631_ (.A(_389_),
    .B1(_142_),
    .B2(_158_),
    .ZN(_309_));
 NOR2_X1 _632_ (.A1(_218_),
    .A2(_141_),
    .ZN(_310_));
 AOI21_X1 _633_ (.A(_310_),
    .B1(_203_),
    .B2(_304_),
    .ZN(_311_));
 INV_X1 _634_ (.A(_311_),
    .ZN(_312_));
 NOR2_X1 _635_ (.A1(_302_),
    .A2(_312_),
    .ZN(_313_));
 XNOR2_X1 _636_ (.A(_313_),
    .B(_200_),
    .ZN(_407_));
 NAND2_X1 _637_ (.A1(_253_),
    .A2(_407_),
    .ZN(_314_));
 OAI211_X2 _638_ (.A(_309_),
    .B(_314_),
    .C1(_245_),
    .C2(_070_),
    .ZN(_315_));
 MUX2_X1 _639_ (.A(_111_),
    .B(_315_),
    .S(_249_),
    .Z(_077_));
 OAI21_X1 _640_ (.A(_390_),
    .B1(_165_),
    .B2(_159_),
    .ZN(_316_));
 OAI21_X4 _641_ (.A(_316_),
    .B1(_246_),
    .B2(_071_),
    .ZN(_317_));
 OAI21_X1 _642_ (.A(_200_),
    .B1(_302_),
    .B2(_312_),
    .ZN(_318_));
 NOR2_X1 _643_ (.A1(_223_),
    .A2(_127_),
    .ZN(_319_));
 INV_X1 _644_ (.A(_319_),
    .ZN(_320_));
 NAND2_X1 _645_ (.A1(_318_),
    .A2(_320_),
    .ZN(_321_));
 INV_X1 _646_ (.A(_201_),
    .ZN(_322_));
 XNOR2_X1 _647_ (.A(_321_),
    .B(_322_),
    .ZN(_408_));
 AND2_X1 _648_ (.A1(_408_),
    .A2(_254_),
    .ZN(_323_));
 OAI21_X2 _649_ (.A(_250_),
    .B1(_317_),
    .B2(_323_),
    .ZN(_324_));
 OAI21_X1 _650_ (.A(_324_),
    .B1(_221_),
    .B2(_250_),
    .ZN(_078_));
 OAI21_X1 _651_ (.A(_391_),
    .B1(_142_),
    .B2(_158_),
    .ZN(_325_));
 AND2_X2 _652_ (.A1(_299_),
    .A2(_205_),
    .ZN(_326_));
 AND3_X1 _653_ (.A1(_312_),
    .A2(_200_),
    .A3(_201_),
    .ZN(_327_));
 NAND2_X1 _654_ (.A1(_201_),
    .A2(_319_),
    .ZN(_328_));
 OAI21_X1 _655_ (.A(_328_),
    .B1(_221_),
    .B2(_128_),
    .ZN(_329_));
 NOR3_X4 _656_ (.A1(_326_),
    .A2(_327_),
    .A3(_329_),
    .ZN(_330_));
 XNOR2_X1 _657_ (.A(_330_),
    .B(_211_),
    .ZN(_409_));
 NAND2_X1 _658_ (.A1(_253_),
    .A2(_409_),
    .ZN(_331_));
 OAI211_X2 _659_ (.A(_325_),
    .B(_331_),
    .C1(_245_),
    .C2(_072_),
    .ZN(_332_));
 MUX2_X1 _660_ (.A(_113_),
    .B(_332_),
    .S(_249_),
    .Z(_079_));
 NOR2_X1 _661_ (.A1(_330_),
    .A2(_212_),
    .ZN(_333_));
 NOR2_X1 _662_ (.A1(_233_),
    .A2(_129_),
    .ZN(_334_));
 NOR2_X2 _663_ (.A1(_333_),
    .A2(_334_),
    .ZN(_335_));
 XNOR2_X1 _664_ (.A(_335_),
    .B(_209_),
    .ZN(_410_));
 NAND2_X1 _665_ (.A1(_410_),
    .A2(_253_),
    .ZN(_336_));
 OAI21_X1 _666_ (.A(_392_),
    .B1(_142_),
    .B2(_158_),
    .ZN(_337_));
 OAI211_X2 _667_ (.A(_336_),
    .B(_337_),
    .C1(_073_),
    .C2(_245_),
    .ZN(_338_));
 MUX2_X1 _668_ (.A(_114_),
    .B(_338_),
    .S(_249_),
    .Z(_080_));
 OR3_X4 _669_ (.A1(_330_),
    .A2(_210_),
    .A3(_212_),
    .ZN(_339_));
 INV_X1 _670_ (.A(_206_),
    .ZN(_340_));
 AOI22_X1 _671_ (.A1(_209_),
    .A2(_334_),
    .B1(_114_),
    .B2(_073_),
    .ZN(_341_));
 AND3_X4 _672_ (.A1(_339_),
    .A2(_340_),
    .A3(_341_),
    .ZN(_342_));
 AOI21_X4 _673_ (.A(_340_),
    .B1(_339_),
    .B2(_341_),
    .ZN(_343_));
 NOR2_X1 _674_ (.A1(_342_),
    .A2(_343_),
    .ZN(_411_));
 NAND2_X1 _675_ (.A1(_411_),
    .A2(_253_),
    .ZN(_344_));
 OAI21_X1 _676_ (.A(_394_),
    .B1(_142_),
    .B2(_158_),
    .ZN(_345_));
 OAI211_X2 _677_ (.A(_344_),
    .B(_345_),
    .C1(_074_),
    .C2(_245_),
    .ZN(_346_));
 MUX2_X1 _678_ (.A(_115_),
    .B(_346_),
    .S(_249_),
    .Z(_081_));
 NOR2_X1 _679_ (.A1(_227_),
    .A2(_131_),
    .ZN(_347_));
 NOR2_X4 _680_ (.A1(_343_),
    .A2(_347_),
    .ZN(_348_));
 XNOR2_X1 _681_ (.A(_348_),
    .B(_207_),
    .ZN(_412_));
 AND2_X2 _682_ (.A1(_412_),
    .A2(_254_),
    .ZN(_349_));
 OAI21_X1 _683_ (.A(_395_),
    .B1(_165_),
    .B2(_159_),
    .ZN(_350_));
 OAI21_X1 _684_ (.A(_350_),
    .B1(_245_),
    .B2(_075_),
    .ZN(_351_));
 OAI21_X1 _685_ (.A(_250_),
    .B1(_349_),
    .B2(_351_),
    .ZN(_352_));
 OAI21_X1 _686_ (.A(_352_),
    .B1(_167_),
    .B2(_250_),
    .ZN(_082_));
 MUX2_X1 _687_ (.A(_110_),
    .B(_371_),
    .S(_160_),
    .Z(_353_));
 NAND2_X2 _688_ (.A1(_243_),
    .A2(_059_),
    .ZN(_354_));
 BUF_X4 _689_ (.A(_354_),
    .Z(_355_));
 MUX2_X1 _690_ (.A(_126_),
    .B(_353_),
    .S(_355_),
    .Z(_092_));
 MUX2_X1 _691_ (.A(_117_),
    .B(_382_),
    .S(_160_),
    .Z(_356_));
 MUX2_X1 _692_ (.A(_133_),
    .B(_356_),
    .S(_355_),
    .Z(_099_));
 MUX2_X1 _693_ (.A(_118_),
    .B(_393_),
    .S(_160_),
    .Z(_357_));
 MUX2_X1 _694_ (.A(_134_),
    .B(_357_),
    .S(_355_),
    .Z(_100_));
 MUX2_X1 _695_ (.A(_119_),
    .B(_396_),
    .S(_160_),
    .Z(_358_));
 MUX2_X1 _696_ (.A(_135_),
    .B(_358_),
    .S(_355_),
    .Z(_101_));
 MUX2_X1 _697_ (.A(_120_),
    .B(_397_),
    .S(_160_),
    .Z(_359_));
 MUX2_X1 _698_ (.A(_136_),
    .B(_359_),
    .S(_355_),
    .Z(_102_));
 MUX2_X1 _699_ (.A(_121_),
    .B(_398_),
    .S(_160_),
    .Z(_360_));
 MUX2_X1 _700_ (.A(_137_),
    .B(_360_),
    .S(_355_),
    .Z(_103_));
 MUX2_X1 _701_ (.A(_122_),
    .B(_399_),
    .S(_160_),
    .Z(_361_));
 MUX2_X1 _702_ (.A(_138_),
    .B(_361_),
    .S(_355_),
    .Z(_104_));
 MUX2_X1 _703_ (.A(_123_),
    .B(_400_),
    .S(_160_),
    .Z(_362_));
 MUX2_X1 _704_ (.A(_139_),
    .B(_362_),
    .S(_355_),
    .Z(_105_));
 MUX2_X1 _705_ (.A(_124_),
    .B(_401_),
    .S(_160_),
    .Z(_363_));
 MUX2_X1 _706_ (.A(_140_),
    .B(_363_),
    .S(_355_),
    .Z(_106_));
 MUX2_X1 _707_ (.A(_125_),
    .B(_402_),
    .S(_403_),
    .Z(_364_));
 MUX2_X1 _708_ (.A(_141_),
    .B(_364_),
    .S(_355_),
    .Z(_107_));
 MUX2_X1 _709_ (.A(_111_),
    .B(_372_),
    .S(_403_),
    .Z(_365_));
 MUX2_X1 _710_ (.A(_127_),
    .B(_365_),
    .S(_354_),
    .Z(_093_));
 MUX2_X1 _711_ (.A(_112_),
    .B(_373_),
    .S(_403_),
    .Z(_366_));
 MUX2_X1 _712_ (.A(_128_),
    .B(_366_),
    .S(_354_),
    .Z(_094_));
 MUX2_X1 _713_ (.A(_113_),
    .B(_374_),
    .S(_403_),
    .Z(_367_));
 MUX2_X1 _714_ (.A(_129_),
    .B(_367_),
    .S(_354_),
    .Z(_095_));
 MUX2_X1 _715_ (.A(_114_),
    .B(_375_),
    .S(_403_),
    .Z(_368_));
 MUX2_X1 _716_ (.A(_130_),
    .B(_368_),
    .S(_354_),
    .Z(_096_));
 MUX2_X1 _717_ (.A(_115_),
    .B(_376_),
    .S(_403_),
    .Z(_369_));
 MUX2_X1 _718_ (.A(_131_),
    .B(_369_),
    .S(_354_),
    .Z(_097_));
 MUX2_X1 _719_ (.A(_116_),
    .B(_377_),
    .S(_403_),
    .Z(_370_));
 MUX2_X1 _720_ (.A(_132_),
    .B(_370_),
    .S(_354_),
    .Z(_098_));
 BUF_X1 _721_ (.A(reset),
    .Z(_405_));
 BUF_X1 _722_ (.A(\ctrl.state.out[2] ),
    .Z(_109_));
 BUF_X1 _723_ (.A(\ctrl.state.out[1] ),
    .Z(_108_));
 BUF_X1 _724_ (.A(_005_),
    .Z(_059_));
 BUF_X1 _725_ (.A(_423_),
    .Z(resp_val));
 BUF_X1 _726_ (.A(resp_rdy),
    .Z(_422_));
 BUF_X1 _727_ (.A(\dpath.a_lt_b$in0[15] ),
    .Z(_116_));
 BUF_X1 _728_ (.A(\dpath.a_lt_b$in1[15] ),
    .Z(_132_));
 BUF_X1 _729_ (.A(\dpath.a_lt_b$in0[14] ),
    .Z(_115_));
 BUF_X1 _730_ (.A(\dpath.a_lt_b$in1[14] ),
    .Z(_131_));
 BUF_X1 _731_ (.A(\dpath.a_lt_b$in0[13] ),
    .Z(_114_));
 BUF_X1 _732_ (.A(\dpath.a_lt_b$in1[13] ),
    .Z(_130_));
 BUF_X1 _733_ (.A(\dpath.a_lt_b$in0[12] ),
    .Z(_113_));
 BUF_X1 _734_ (.A(\dpath.a_lt_b$in1[12] ),
    .Z(_129_));
 BUF_X1 _735_ (.A(\dpath.a_lt_b$in0[11] ),
    .Z(_112_));
 BUF_X1 _736_ (.A(\dpath.a_lt_b$in1[11] ),
    .Z(_128_));
 BUF_X1 _737_ (.A(\dpath.a_lt_b$in0[10] ),
    .Z(_111_));
 BUF_X1 _738_ (.A(\dpath.a_lt_b$in1[10] ),
    .Z(_127_));
 BUF_X1 _739_ (.A(\dpath.a_lt_b$in0[9] ),
    .Z(_125_));
 BUF_X1 _740_ (.A(\dpath.a_lt_b$in1[9] ),
    .Z(_141_));
 BUF_X1 _741_ (.A(\dpath.a_lt_b$in0[8] ),
    .Z(_124_));
 BUF_X1 _742_ (.A(\dpath.a_lt_b$in1[8] ),
    .Z(_140_));
 BUF_X1 _743_ (.A(\dpath.a_lt_b$in0[7] ),
    .Z(_123_));
 BUF_X1 _744_ (.A(\dpath.a_lt_b$in1[7] ),
    .Z(_139_));
 BUF_X1 _745_ (.A(\dpath.a_lt_b$in0[6] ),
    .Z(_122_));
 BUF_X1 _746_ (.A(\dpath.a_lt_b$in1[6] ),
    .Z(_138_));
 BUF_X1 _747_ (.A(\dpath.a_lt_b$in0[5] ),
    .Z(_121_));
 BUF_X1 _748_ (.A(\dpath.a_lt_b$in1[5] ),
    .Z(_137_));
 BUF_X1 _749_ (.A(\dpath.a_lt_b$in0[4] ),
    .Z(_120_));
 BUF_X1 _750_ (.A(\dpath.a_lt_b$in1[4] ),
    .Z(_136_));
 BUF_X1 _751_ (.A(\dpath.a_lt_b$in0[3] ),
    .Z(_119_));
 BUF_X1 _752_ (.A(\dpath.a_lt_b$in1[3] ),
    .Z(_135_));
 BUF_X1 _753_ (.A(\dpath.a_lt_b$in0[2] ),
    .Z(_118_));
 BUF_X1 _754_ (.A(\dpath.a_lt_b$in1[2] ),
    .Z(_134_));
 BUF_X1 _755_ (.A(\dpath.a_lt_b$in0[1] ),
    .Z(_117_));
 BUF_X1 _756_ (.A(\dpath.a_lt_b$in1[1] ),
    .Z(_133_));
 BUF_X1 _757_ (.A(\dpath.a_lt_b$in0[0] ),
    .Z(_110_));
 BUF_X1 _758_ (.A(\dpath.a_lt_b$in1[0] ),
    .Z(_126_));
 BUF_X1 _759_ (.A(_406_),
    .Z(resp_msg[0]));
 BUF_X1 _760_ (.A(_004_),
    .Z(_058_));
 BUF_X1 _761_ (.A(_003_),
    .Z(_057_));
 BUF_X1 _762_ (.A(_055_),
    .Z(_001_));
 BUF_X1 _763_ (.A(req_rdy),
    .Z(_403_));
 BUF_X1 _764_ (.A(req_val),
    .Z(_404_));
 BUF_X1 _765_ (.A(_056_),
    .Z(_002_));
 BUF_X1 _766_ (.A(_054_),
    .Z(_000_));
 BUF_X1 _767_ (.A(_006_),
    .Z(_060_));
 BUF_X1 _768_ (.A(req_msg[16]),
    .Z(_378_));
 BUF_X1 _769_ (.A(_076_),
    .Z(_022_));
 BUF_X1 _770_ (.A(_007_),
    .Z(_061_));
 BUF_X1 _771_ (.A(req_msg[17]),
    .Z(_379_));
 BUF_X1 _772_ (.A(_083_),
    .Z(_029_));
 BUF_X1 _773_ (.A(_008_),
    .Z(_062_));
 BUF_X1 _774_ (.A(req_msg[18]),
    .Z(_380_));
 BUF_X1 _775_ (.A(_084_),
    .Z(_030_));
 BUF_X1 _776_ (.A(_009_),
    .Z(_063_));
 BUF_X1 _777_ (.A(req_msg[19]),
    .Z(_381_));
 BUF_X1 _778_ (.A(_085_),
    .Z(_031_));
 BUF_X1 _779_ (.A(_010_),
    .Z(_064_));
 BUF_X1 _780_ (.A(req_msg[20]),
    .Z(_383_));
 BUF_X1 _781_ (.A(_086_),
    .Z(_032_));
 BUF_X1 _782_ (.A(_011_),
    .Z(_065_));
 BUF_X1 _783_ (.A(req_msg[21]),
    .Z(_384_));
 BUF_X1 _784_ (.A(_087_),
    .Z(_033_));
 BUF_X1 _785_ (.A(_012_),
    .Z(_066_));
 BUF_X1 _786_ (.A(req_msg[22]),
    .Z(_385_));
 BUF_X1 _787_ (.A(_088_),
    .Z(_034_));
 BUF_X1 _788_ (.A(_013_),
    .Z(_067_));
 BUF_X1 _789_ (.A(req_msg[23]),
    .Z(_386_));
 BUF_X1 _790_ (.A(_089_),
    .Z(_035_));
 BUF_X1 _791_ (.A(_014_),
    .Z(_068_));
 BUF_X1 _792_ (.A(req_msg[24]),
    .Z(_387_));
 BUF_X1 _793_ (.A(_090_),
    .Z(_036_));
 BUF_X1 _794_ (.A(_015_),
    .Z(_069_));
 BUF_X1 _795_ (.A(req_msg[25]),
    .Z(_388_));
 BUF_X1 _796_ (.A(_091_),
    .Z(_037_));
 BUF_X1 _797_ (.A(_016_),
    .Z(_070_));
 BUF_X1 _798_ (.A(req_msg[26]),
    .Z(_389_));
 BUF_X1 _799_ (.A(_077_),
    .Z(_023_));
 BUF_X1 _800_ (.A(_017_),
    .Z(_071_));
 BUF_X1 _801_ (.A(req_msg[27]),
    .Z(_390_));
 BUF_X1 _802_ (.A(_078_),
    .Z(_024_));
 BUF_X1 _803_ (.A(_018_),
    .Z(_072_));
 BUF_X1 _804_ (.A(req_msg[28]),
    .Z(_391_));
 BUF_X1 _805_ (.A(_079_),
    .Z(_025_));
 BUF_X1 _806_ (.A(_019_),
    .Z(_073_));
 BUF_X1 _807_ (.A(req_msg[29]),
    .Z(_392_));
 BUF_X1 _808_ (.A(_080_),
    .Z(_026_));
 BUF_X1 _809_ (.A(_020_),
    .Z(_074_));
 BUF_X1 _810_ (.A(req_msg[30]),
    .Z(_394_));
 BUF_X1 _811_ (.A(_081_),
    .Z(_027_));
 BUF_X1 _812_ (.A(_021_),
    .Z(_075_));
 BUF_X1 _813_ (.A(req_msg[31]),
    .Z(_395_));
 BUF_X1 _814_ (.A(_082_),
    .Z(_028_));
 BUF_X1 _815_ (.A(req_msg[0]),
    .Z(_371_));
 BUF_X1 _816_ (.A(_092_),
    .Z(_038_));
 BUF_X1 _817_ (.A(req_msg[1]),
    .Z(_382_));
 BUF_X1 _818_ (.A(_099_),
    .Z(_045_));
 BUF_X1 _819_ (.A(req_msg[2]),
    .Z(_393_));
 BUF_X1 _820_ (.A(_100_),
    .Z(_046_));
 BUF_X1 _821_ (.A(req_msg[3]),
    .Z(_396_));
 BUF_X1 _822_ (.A(_101_),
    .Z(_047_));
 BUF_X1 _823_ (.A(req_msg[4]),
    .Z(_397_));
 BUF_X1 _824_ (.A(_102_),
    .Z(_048_));
 BUF_X1 _825_ (.A(req_msg[5]),
    .Z(_398_));
 BUF_X1 _826_ (.A(_103_),
    .Z(_049_));
 BUF_X1 _827_ (.A(req_msg[6]),
    .Z(_399_));
 BUF_X1 _828_ (.A(_104_),
    .Z(_050_));
 BUF_X1 _829_ (.A(req_msg[7]),
    .Z(_400_));
 BUF_X1 _830_ (.A(_105_),
    .Z(_051_));
 BUF_X1 _831_ (.A(req_msg[8]),
    .Z(_401_));
 BUF_X1 _832_ (.A(_106_),
    .Z(_052_));
 BUF_X1 _833_ (.A(req_msg[9]),
    .Z(_402_));
 BUF_X1 _834_ (.A(_107_),
    .Z(_053_));
 BUF_X1 _835_ (.A(req_msg[10]),
    .Z(_372_));
 BUF_X1 _836_ (.A(_093_),
    .Z(_039_));
 BUF_X1 _837_ (.A(req_msg[11]),
    .Z(_373_));
 BUF_X1 _838_ (.A(_094_),
    .Z(_040_));
 BUF_X1 _839_ (.A(req_msg[12]),
    .Z(_374_));
 BUF_X1 _840_ (.A(_095_),
    .Z(_041_));
 BUF_X1 _841_ (.A(req_msg[13]),
    .Z(_375_));
 BUF_X1 _842_ (.A(_096_),
    .Z(_042_));
 BUF_X1 _843_ (.A(req_msg[14]),
    .Z(_376_));
 BUF_X1 _844_ (.A(_097_),
    .Z(_043_));
 BUF_X1 _845_ (.A(req_msg[15]),
    .Z(_377_));
 BUF_X1 _846_ (.A(_098_),
    .Z(_044_));
 BUF_X1 _847_ (.A(_413_),
    .Z(resp_msg[1]));
 BUF_X1 _848_ (.A(_414_),
    .Z(resp_msg[2]));
 BUF_X1 _849_ (.A(_415_),
    .Z(resp_msg[3]));
 BUF_X1 _850_ (.A(_416_),
    .Z(resp_msg[4]));
 BUF_X1 _851_ (.A(_417_),
    .Z(resp_msg[5]));
 BUF_X1 _852_ (.A(_418_),
    .Z(resp_msg[6]));
 BUF_X1 _853_ (.A(_419_),
    .Z(resp_msg[7]));
 BUF_X1 _854_ (.A(_420_),
    .Z(resp_msg[8]));
 BUF_X1 _855_ (.A(_421_),
    .Z(resp_msg[9]));
 BUF_X1 _856_ (.A(_407_),
    .Z(resp_msg[10]));
 BUF_X1 _857_ (.A(_408_),
    .Z(resp_msg[11]));
 BUF_X1 _858_ (.A(_409_),
    .Z(resp_msg[12]));
 BUF_X1 _859_ (.A(_410_),
    .Z(resp_msg[13]));
 BUF_X1 _860_ (.A(_411_),
    .Z(resp_msg[14]));
 BUF_X1 _861_ (.A(_412_),
    .Z(resp_msg[15]));
 DFF_X1 _862_ (.D(_000_),
    .CK(clk),
    .Q(req_rdy),
    .QN(_005_));
 DFF_X1 _863_ (.D(_001_),
    .CK(clk),
    .Q(\ctrl.state.out[1] ),
    .QN(_003_));
 DFF_X1 _864_ (.D(_002_),
    .CK(clk),
    .Q(\ctrl.state.out[2] ),
    .QN(_004_));
 DFF_X1 _865_ (.D(_022_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in0[0] ),
    .QN(_424_));
 DFF_X1 _866_ (.D(_029_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in0[1] ),
    .QN(_425_));
 DFF_X1 _867_ (.D(_030_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in0[2] ),
    .QN(_426_));
 DFF_X1 _868_ (.D(_031_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in0[3] ),
    .QN(_427_));
 DFF_X1 _869_ (.D(_032_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in0[4] ),
    .QN(_428_));
 DFF_X1 _870_ (.D(_033_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in0[5] ),
    .QN(_429_));
 DFF_X1 _871_ (.D(_034_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in0[6] ),
    .QN(_430_));
 DFF_X1 _872_ (.D(_035_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in0[7] ),
    .QN(_431_));
 DFF_X1 _873_ (.D(_036_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in0[8] ),
    .QN(_432_));
 DFF_X1 _874_ (.D(_037_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in0[9] ),
    .QN(_433_));
 DFF_X1 _875_ (.D(_023_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in0[10] ),
    .QN(_434_));
 DFF_X1 _876_ (.D(_024_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in0[11] ),
    .QN(_435_));
 DFF_X1 _877_ (.D(_025_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in0[12] ),
    .QN(_436_));
 DFF_X1 _878_ (.D(_026_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in0[13] ),
    .QN(_437_));
 DFF_X1 _879_ (.D(_027_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in0[14] ),
    .QN(_438_));
 DFF_X1 _880_ (.D(_028_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in0[15] ),
    .QN(_439_));
 DFF_X1 _881_ (.D(_038_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in1[0] ),
    .QN(_006_));
 DFF_X1 _882_ (.D(_045_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in1[1] ),
    .QN(_007_));
 DFF_X1 _883_ (.D(_046_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in1[2] ),
    .QN(_008_));
 DFF_X1 _884_ (.D(_047_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in1[3] ),
    .QN(_009_));
 DFF_X1 _885_ (.D(_048_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in1[4] ),
    .QN(_010_));
 DFF_X1 _886_ (.D(_049_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in1[5] ),
    .QN(_011_));
 DFF_X1 _887_ (.D(_050_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in1[6] ),
    .QN(_012_));
 DFF_X1 _888_ (.D(_051_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in1[7] ),
    .QN(_013_));
 DFF_X1 _889_ (.D(_052_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in1[8] ),
    .QN(_014_));
 DFF_X1 _890_ (.D(_053_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in1[9] ),
    .QN(_015_));
 DFF_X1 _891_ (.D(_039_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in1[10] ),
    .QN(_016_));
 DFF_X1 _892_ (.D(_040_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in1[11] ),
    .QN(_017_));
 DFF_X1 _893_ (.D(_041_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in1[12] ),
    .QN(_018_));
 DFF_X1 _894_ (.D(_042_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in1[13] ),
    .QN(_019_));
 DFF_X1 _895_ (.D(_043_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in1[14] ),
    .QN(_020_));
 DFF_X1 _896_ (.D(_044_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in1[15] ),
    .QN(_021_));
endmodule
