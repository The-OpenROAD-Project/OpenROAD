VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram45_256x16
  FOREIGN fakeram45_256x16 0 0 ;
  SYMMETRY X Y ;
  SIZE 57.570 BY 133.000 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.165 0.070 4.235 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.265 0.070 6.335 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.465 0.070 10.535 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.565 0.070 12.635 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.665 0.070 14.735 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.765 0.070 16.835 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.865 0.070 18.935 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.065 0.070 23.135 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.165 0.070 25.235 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.265 0.070 27.335 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.365 0.070 29.435 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.465 0.070 31.535 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.565 0.070 33.635 ;
    END
  END w_mask_in[15]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.615 0.070 34.685 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.715 0.070 36.785 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.815 0.070 38.885 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.915 0.070 40.985 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.015 0.070 43.085 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.115 0.070 45.185 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.215 0.070 47.285 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.315 0.070 49.385 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.415 0.070 51.485 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.515 0.070 53.585 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.615 0.070 55.685 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.715 0.070 57.785 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.815 0.070 59.885 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.915 0.070 61.985 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.015 0.070 64.085 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.115 0.070 66.185 ;
    END
  END rd_out[15]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.165 0.070 67.235 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.265 0.070 69.335 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.365 0.070 71.435 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.465 0.070 73.535 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.565 0.070 75.635 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.665 0.070 77.735 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.765 0.070 79.835 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.865 0.070 81.935 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.965 0.070 84.035 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.065 0.070 86.135 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.165 0.070 88.235 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.265 0.070 90.335 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.365 0.070 92.435 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.465 0.070 94.535 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.565 0.070 96.635 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.665 0.070 98.735 ;
    END
  END wd_in[15]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.715 0.070 99.785 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.815 0.070 101.885 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.915 0.070 103.985 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.015 0.070 106.085 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.115 0.070 108.185 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.215 0.070 110.285 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.315 0.070 112.385 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.415 0.070 114.485 ;
    END
  END addr_in[7]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.465 0.070 115.535 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.565 0.070 117.635 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.665 0.070 119.735 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.960 2.100 2.240 130.900 ;
      RECT 5.320 2.100 5.600 130.900 ;
      RECT 8.680 2.100 8.960 130.900 ;
      RECT 12.040 2.100 12.320 130.900 ;
      RECT 15.400 2.100 15.680 130.900 ;
      RECT 18.760 2.100 19.040 130.900 ;
      RECT 22.120 2.100 22.400 130.900 ;
      RECT 25.480 2.100 25.760 130.900 ;
      RECT 28.840 2.100 29.120 130.900 ;
      RECT 32.200 2.100 32.480 130.900 ;
      RECT 35.560 2.100 35.840 130.900 ;
      RECT 38.920 2.100 39.200 130.900 ;
      RECT 42.280 2.100 42.560 130.900 ;
      RECT 45.640 2.100 45.920 130.900 ;
      RECT 49.000 2.100 49.280 130.900 ;
      RECT 52.360 2.100 52.640 130.900 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 3.640 2.100 3.920 130.900 ;
      RECT 7.000 2.100 7.280 130.900 ;
      RECT 10.360 2.100 10.640 130.900 ;
      RECT 13.720 2.100 14.000 130.900 ;
      RECT 17.080 2.100 17.360 130.900 ;
      RECT 20.440 2.100 20.720 130.900 ;
      RECT 23.800 2.100 24.080 130.900 ;
      RECT 27.160 2.100 27.440 130.900 ;
      RECT 30.520 2.100 30.800 130.900 ;
      RECT 33.880 2.100 34.160 130.900 ;
      RECT 37.240 2.100 37.520 130.900 ;
      RECT 40.600 2.100 40.880 130.900 ;
      RECT 43.960 2.100 44.240 130.900 ;
      RECT 47.320 2.100 47.600 130.900 ;
      RECT 50.680 2.100 50.960 130.900 ;
      RECT 54.040 2.100 54.320 130.900 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 57.570 133.000 ;
    LAYER metal2 ;
    RECT 0 0 57.570 133.000 ;
    LAYER metal3 ;
    RECT 0.070 0 57.570 133.000 ;
    RECT 0 0.000 0.070 2.065 ;
    RECT 0 2.135 0.070 4.165 ;
    RECT 0 4.235 0.070 6.265 ;
    RECT 0 6.335 0.070 8.365 ;
    RECT 0 8.435 0.070 10.465 ;
    RECT 0 10.535 0.070 12.565 ;
    RECT 0 12.635 0.070 14.665 ;
    RECT 0 14.735 0.070 16.765 ;
    RECT 0 16.835 0.070 18.865 ;
    RECT 0 18.935 0.070 20.965 ;
    RECT 0 21.035 0.070 23.065 ;
    RECT 0 23.135 0.070 25.165 ;
    RECT 0 25.235 0.070 27.265 ;
    RECT 0 27.335 0.070 29.365 ;
    RECT 0 29.435 0.070 31.465 ;
    RECT 0 31.535 0.070 33.565 ;
    RECT 0 33.635 0.070 34.615 ;
    RECT 0 34.685 0.070 36.715 ;
    RECT 0 36.785 0.070 38.815 ;
    RECT 0 38.885 0.070 40.915 ;
    RECT 0 40.985 0.070 43.015 ;
    RECT 0 43.085 0.070 45.115 ;
    RECT 0 45.185 0.070 47.215 ;
    RECT 0 47.285 0.070 49.315 ;
    RECT 0 49.385 0.070 51.415 ;
    RECT 0 51.485 0.070 53.515 ;
    RECT 0 53.585 0.070 55.615 ;
    RECT 0 55.685 0.070 57.715 ;
    RECT 0 57.785 0.070 59.815 ;
    RECT 0 59.885 0.070 61.915 ;
    RECT 0 61.985 0.070 64.015 ;
    RECT 0 64.085 0.070 66.115 ;
    RECT 0 66.185 0.070 67.165 ;
    RECT 0 67.235 0.070 69.265 ;
    RECT 0 69.335 0.070 71.365 ;
    RECT 0 71.435 0.070 73.465 ;
    RECT 0 73.535 0.070 75.565 ;
    RECT 0 75.635 0.070 77.665 ;
    RECT 0 77.735 0.070 79.765 ;
    RECT 0 79.835 0.070 81.865 ;
    RECT 0 81.935 0.070 83.965 ;
    RECT 0 84.035 0.070 86.065 ;
    RECT 0 86.135 0.070 88.165 ;
    RECT 0 88.235 0.070 90.265 ;
    RECT 0 90.335 0.070 92.365 ;
    RECT 0 92.435 0.070 94.465 ;
    RECT 0 94.535 0.070 96.565 ;
    RECT 0 96.635 0.070 98.665 ;
    RECT 0 98.735 0.070 99.715 ;
    RECT 0 99.785 0.070 101.815 ;
    RECT 0 101.885 0.070 103.915 ;
    RECT 0 103.985 0.070 106.015 ;
    RECT 0 106.085 0.070 108.115 ;
    RECT 0 108.185 0.070 110.215 ;
    RECT 0 110.285 0.070 112.315 ;
    RECT 0 112.385 0.070 114.415 ;
    RECT 0 114.485 0.070 115.465 ;
    RECT 0 115.535 0.070 117.565 ;
    RECT 0 117.635 0.070 119.665 ;
    RECT 0 119.735 0.070 133.000 ;
    LAYER metal4 ;
    RECT 0 0 57.570 2.100 ;
    RECT 0 130.900 57.570 133.000 ;
    RECT 0.000 2.100 1.960 130.900 ;
    RECT 2.240 2.100 3.640 130.900 ;
    RECT 3.920 2.100 5.320 130.900 ;
    RECT 5.600 2.100 7.000 130.900 ;
    RECT 7.280 2.100 8.680 130.900 ;
    RECT 8.960 2.100 10.360 130.900 ;
    RECT 10.640 2.100 12.040 130.900 ;
    RECT 12.320 2.100 13.720 130.900 ;
    RECT 14.000 2.100 15.400 130.900 ;
    RECT 15.680 2.100 17.080 130.900 ;
    RECT 17.360 2.100 18.760 130.900 ;
    RECT 19.040 2.100 20.440 130.900 ;
    RECT 20.720 2.100 22.120 130.900 ;
    RECT 22.400 2.100 23.800 130.900 ;
    RECT 24.080 2.100 25.480 130.900 ;
    RECT 25.760 2.100 27.160 130.900 ;
    RECT 27.440 2.100 28.840 130.900 ;
    RECT 29.120 2.100 30.520 130.900 ;
    RECT 30.800 2.100 32.200 130.900 ;
    RECT 32.480 2.100 33.880 130.900 ;
    RECT 34.160 2.100 35.560 130.900 ;
    RECT 35.840 2.100 37.240 130.900 ;
    RECT 37.520 2.100 38.920 130.900 ;
    RECT 39.200 2.100 40.600 130.900 ;
    RECT 40.880 2.100 42.280 130.900 ;
    RECT 42.560 2.100 43.960 130.900 ;
    RECT 44.240 2.100 45.640 130.900 ;
    RECT 45.920 2.100 47.320 130.900 ;
    RECT 47.600 2.100 49.000 130.900 ;
    RECT 49.280 2.100 50.680 130.900 ;
    RECT 50.960 2.100 52.360 130.900 ;
    RECT 52.640 2.100 54.040 130.900 ;
    RECT 54.320 2.100 57.570 130.900 ;
    LAYER OVERLAP ;
    RECT 0 0 57.570 133.000 ;
  END
END fakeram45_256x16

END LIBRARY
