# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_io__overlay_vssd_lvc
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 198 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 51.125000 1.270000 54.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.125000 75.000000 54.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 46.365000 1.270000 49.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 46.365000 75.000000 49.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 6.885000 1.270000 11.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 6.885000 75.000000 11.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 6.985000 1.270000 11.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 6.985000 75.000000 11.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 0.035000 1.270000 5.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 0.035000 75.000000 5.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 0.135000 1.270000 5.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 0.135000 75.000000 5.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 12.935000 0.965000 16.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035000 12.935000 75.000000 16.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 13.035000 0.965000 16.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 13.035000 75.000000 16.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 17.785000 1.270000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 68.035000 1.270000 93.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 17.785000 75.000000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 68.035000 75.000000 93.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 17.885000 1.270000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 68.035000 1.270000 92.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 17.885000 75.000000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 68.035000 75.000000 92.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 62.085000 1.270000 66.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 62.085000 75.000000 66.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 62.185000 1.270000 66.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 62.185000 75.000000 66.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 34.735000 1.270000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 45.735000 1.270000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 49.645000 1.270000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 54.405000 1.270000 54.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 34.735000 75.000000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 45.735000 75.000000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 49.645000 75.000000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 54.405000 75.000000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 34.840000 1.270000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 45.735000 1.270000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 34.840000 75.000000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 45.735000 75.000000 54.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.500000 39.590000 24.500000 44.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755000 39.590000 74.700000 44.230000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 39.585000 24.475000 44.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.780000 39.585000 75.000000 44.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 39.685000 1.270000 44.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 39.685000 75.000000 44.135000 ;
    END
    PORT
      LAYER via3 ;
        RECT  0.590000 39.660000  0.790000 39.860000 ;
        RECT  0.590000 40.090000  0.790000 40.290000 ;
        RECT  0.590000 40.520000  0.790000 40.720000 ;
        RECT  0.590000 40.950000  0.790000 41.150000 ;
        RECT  0.590000 41.380000  0.790000 41.580000 ;
        RECT  0.590000 41.810000  0.790000 42.010000 ;
        RECT  0.590000 42.240000  0.790000 42.440000 ;
        RECT  0.590000 42.670000  0.790000 42.870000 ;
        RECT  0.590000 43.100000  0.790000 43.300000 ;
        RECT  0.590000 43.530000  0.790000 43.730000 ;
        RECT  0.590000 43.960000  0.790000 44.160000 ;
        RECT  0.995000 39.660000  1.195000 39.860000 ;
        RECT  0.995000 40.090000  1.195000 40.290000 ;
        RECT  0.995000 40.520000  1.195000 40.720000 ;
        RECT  0.995000 40.950000  1.195000 41.150000 ;
        RECT  0.995000 41.380000  1.195000 41.580000 ;
        RECT  0.995000 41.810000  1.195000 42.010000 ;
        RECT  0.995000 42.240000  1.195000 42.440000 ;
        RECT  0.995000 42.670000  1.195000 42.870000 ;
        RECT  0.995000 43.100000  1.195000 43.300000 ;
        RECT  0.995000 43.530000  1.195000 43.730000 ;
        RECT  0.995000 43.960000  1.195000 44.160000 ;
        RECT  1.400000 39.660000  1.600000 39.860000 ;
        RECT  1.400000 40.090000  1.600000 40.290000 ;
        RECT  1.400000 40.520000  1.600000 40.720000 ;
        RECT  1.400000 40.950000  1.600000 41.150000 ;
        RECT  1.400000 41.380000  1.600000 41.580000 ;
        RECT  1.400000 41.810000  1.600000 42.010000 ;
        RECT  1.400000 42.240000  1.600000 42.440000 ;
        RECT  1.400000 42.670000  1.600000 42.870000 ;
        RECT  1.400000 43.100000  1.600000 43.300000 ;
        RECT  1.400000 43.530000  1.600000 43.730000 ;
        RECT  1.400000 43.960000  1.600000 44.160000 ;
        RECT  1.805000 39.660000  2.005000 39.860000 ;
        RECT  1.805000 40.090000  2.005000 40.290000 ;
        RECT  1.805000 40.520000  2.005000 40.720000 ;
        RECT  1.805000 40.950000  2.005000 41.150000 ;
        RECT  1.805000 41.380000  2.005000 41.580000 ;
        RECT  1.805000 41.810000  2.005000 42.010000 ;
        RECT  1.805000 42.240000  2.005000 42.440000 ;
        RECT  1.805000 42.670000  2.005000 42.870000 ;
        RECT  1.805000 43.100000  2.005000 43.300000 ;
        RECT  1.805000 43.530000  2.005000 43.730000 ;
        RECT  1.805000 43.960000  2.005000 44.160000 ;
        RECT  2.210000 39.660000  2.410000 39.860000 ;
        RECT  2.210000 40.090000  2.410000 40.290000 ;
        RECT  2.210000 40.520000  2.410000 40.720000 ;
        RECT  2.210000 40.950000  2.410000 41.150000 ;
        RECT  2.210000 41.380000  2.410000 41.580000 ;
        RECT  2.210000 41.810000  2.410000 42.010000 ;
        RECT  2.210000 42.240000  2.410000 42.440000 ;
        RECT  2.210000 42.670000  2.410000 42.870000 ;
        RECT  2.210000 43.100000  2.410000 43.300000 ;
        RECT  2.210000 43.530000  2.410000 43.730000 ;
        RECT  2.210000 43.960000  2.410000 44.160000 ;
        RECT  2.610000 39.660000  2.810000 39.860000 ;
        RECT  2.610000 40.090000  2.810000 40.290000 ;
        RECT  2.610000 40.520000  2.810000 40.720000 ;
        RECT  2.610000 40.950000  2.810000 41.150000 ;
        RECT  2.610000 41.380000  2.810000 41.580000 ;
        RECT  2.610000 41.810000  2.810000 42.010000 ;
        RECT  2.610000 42.240000  2.810000 42.440000 ;
        RECT  2.610000 42.670000  2.810000 42.870000 ;
        RECT  2.610000 43.100000  2.810000 43.300000 ;
        RECT  2.610000 43.530000  2.810000 43.730000 ;
        RECT  2.610000 43.960000  2.810000 44.160000 ;
        RECT  3.010000 39.660000  3.210000 39.860000 ;
        RECT  3.010000 40.090000  3.210000 40.290000 ;
        RECT  3.010000 40.520000  3.210000 40.720000 ;
        RECT  3.010000 40.950000  3.210000 41.150000 ;
        RECT  3.010000 41.380000  3.210000 41.580000 ;
        RECT  3.010000 41.810000  3.210000 42.010000 ;
        RECT  3.010000 42.240000  3.210000 42.440000 ;
        RECT  3.010000 42.670000  3.210000 42.870000 ;
        RECT  3.010000 43.100000  3.210000 43.300000 ;
        RECT  3.010000 43.530000  3.210000 43.730000 ;
        RECT  3.010000 43.960000  3.210000 44.160000 ;
        RECT  3.410000 39.660000  3.610000 39.860000 ;
        RECT  3.410000 40.090000  3.610000 40.290000 ;
        RECT  3.410000 40.520000  3.610000 40.720000 ;
        RECT  3.410000 40.950000  3.610000 41.150000 ;
        RECT  3.410000 41.380000  3.610000 41.580000 ;
        RECT  3.410000 41.810000  3.610000 42.010000 ;
        RECT  3.410000 42.240000  3.610000 42.440000 ;
        RECT  3.410000 42.670000  3.610000 42.870000 ;
        RECT  3.410000 43.100000  3.610000 43.300000 ;
        RECT  3.410000 43.530000  3.610000 43.730000 ;
        RECT  3.410000 43.960000  3.610000 44.160000 ;
        RECT  3.810000 39.660000  4.010000 39.860000 ;
        RECT  3.810000 40.090000  4.010000 40.290000 ;
        RECT  3.810000 40.520000  4.010000 40.720000 ;
        RECT  3.810000 40.950000  4.010000 41.150000 ;
        RECT  3.810000 41.380000  4.010000 41.580000 ;
        RECT  3.810000 41.810000  4.010000 42.010000 ;
        RECT  3.810000 42.240000  4.010000 42.440000 ;
        RECT  3.810000 42.670000  4.010000 42.870000 ;
        RECT  3.810000 43.100000  4.010000 43.300000 ;
        RECT  3.810000 43.530000  4.010000 43.730000 ;
        RECT  3.810000 43.960000  4.010000 44.160000 ;
        RECT  4.210000 39.660000  4.410000 39.860000 ;
        RECT  4.210000 40.090000  4.410000 40.290000 ;
        RECT  4.210000 40.520000  4.410000 40.720000 ;
        RECT  4.210000 40.950000  4.410000 41.150000 ;
        RECT  4.210000 41.380000  4.410000 41.580000 ;
        RECT  4.210000 41.810000  4.410000 42.010000 ;
        RECT  4.210000 42.240000  4.410000 42.440000 ;
        RECT  4.210000 42.670000  4.410000 42.870000 ;
        RECT  4.210000 43.100000  4.410000 43.300000 ;
        RECT  4.210000 43.530000  4.410000 43.730000 ;
        RECT  4.210000 43.960000  4.410000 44.160000 ;
        RECT  4.610000 39.660000  4.810000 39.860000 ;
        RECT  4.610000 40.090000  4.810000 40.290000 ;
        RECT  4.610000 40.520000  4.810000 40.720000 ;
        RECT  4.610000 40.950000  4.810000 41.150000 ;
        RECT  4.610000 41.380000  4.810000 41.580000 ;
        RECT  4.610000 41.810000  4.810000 42.010000 ;
        RECT  4.610000 42.240000  4.810000 42.440000 ;
        RECT  4.610000 42.670000  4.810000 42.870000 ;
        RECT  4.610000 43.100000  4.810000 43.300000 ;
        RECT  4.610000 43.530000  4.810000 43.730000 ;
        RECT  4.610000 43.960000  4.810000 44.160000 ;
        RECT  5.010000 39.660000  5.210000 39.860000 ;
        RECT  5.010000 40.090000  5.210000 40.290000 ;
        RECT  5.010000 40.520000  5.210000 40.720000 ;
        RECT  5.010000 40.950000  5.210000 41.150000 ;
        RECT  5.010000 41.380000  5.210000 41.580000 ;
        RECT  5.010000 41.810000  5.210000 42.010000 ;
        RECT  5.010000 42.240000  5.210000 42.440000 ;
        RECT  5.010000 42.670000  5.210000 42.870000 ;
        RECT  5.010000 43.100000  5.210000 43.300000 ;
        RECT  5.010000 43.530000  5.210000 43.730000 ;
        RECT  5.010000 43.960000  5.210000 44.160000 ;
        RECT  5.410000 39.660000  5.610000 39.860000 ;
        RECT  5.410000 40.090000  5.610000 40.290000 ;
        RECT  5.410000 40.520000  5.610000 40.720000 ;
        RECT  5.410000 40.950000  5.610000 41.150000 ;
        RECT  5.410000 41.380000  5.610000 41.580000 ;
        RECT  5.410000 41.810000  5.610000 42.010000 ;
        RECT  5.410000 42.240000  5.610000 42.440000 ;
        RECT  5.410000 42.670000  5.610000 42.870000 ;
        RECT  5.410000 43.100000  5.610000 43.300000 ;
        RECT  5.410000 43.530000  5.610000 43.730000 ;
        RECT  5.410000 43.960000  5.610000 44.160000 ;
        RECT  5.810000 39.660000  6.010000 39.860000 ;
        RECT  5.810000 40.090000  6.010000 40.290000 ;
        RECT  5.810000 40.520000  6.010000 40.720000 ;
        RECT  5.810000 40.950000  6.010000 41.150000 ;
        RECT  5.810000 41.380000  6.010000 41.580000 ;
        RECT  5.810000 41.810000  6.010000 42.010000 ;
        RECT  5.810000 42.240000  6.010000 42.440000 ;
        RECT  5.810000 42.670000  6.010000 42.870000 ;
        RECT  5.810000 43.100000  6.010000 43.300000 ;
        RECT  5.810000 43.530000  6.010000 43.730000 ;
        RECT  5.810000 43.960000  6.010000 44.160000 ;
        RECT  6.210000 39.660000  6.410000 39.860000 ;
        RECT  6.210000 40.090000  6.410000 40.290000 ;
        RECT  6.210000 40.520000  6.410000 40.720000 ;
        RECT  6.210000 40.950000  6.410000 41.150000 ;
        RECT  6.210000 41.380000  6.410000 41.580000 ;
        RECT  6.210000 41.810000  6.410000 42.010000 ;
        RECT  6.210000 42.240000  6.410000 42.440000 ;
        RECT  6.210000 42.670000  6.410000 42.870000 ;
        RECT  6.210000 43.100000  6.410000 43.300000 ;
        RECT  6.210000 43.530000  6.410000 43.730000 ;
        RECT  6.210000 43.960000  6.410000 44.160000 ;
        RECT  6.610000 39.660000  6.810000 39.860000 ;
        RECT  6.610000 40.090000  6.810000 40.290000 ;
        RECT  6.610000 40.520000  6.810000 40.720000 ;
        RECT  6.610000 40.950000  6.810000 41.150000 ;
        RECT  6.610000 41.380000  6.810000 41.580000 ;
        RECT  6.610000 41.810000  6.810000 42.010000 ;
        RECT  6.610000 42.240000  6.810000 42.440000 ;
        RECT  6.610000 42.670000  6.810000 42.870000 ;
        RECT  6.610000 43.100000  6.810000 43.300000 ;
        RECT  6.610000 43.530000  6.810000 43.730000 ;
        RECT  6.610000 43.960000  6.810000 44.160000 ;
        RECT  7.010000 39.660000  7.210000 39.860000 ;
        RECT  7.010000 40.090000  7.210000 40.290000 ;
        RECT  7.010000 40.520000  7.210000 40.720000 ;
        RECT  7.010000 40.950000  7.210000 41.150000 ;
        RECT  7.010000 41.380000  7.210000 41.580000 ;
        RECT  7.010000 41.810000  7.210000 42.010000 ;
        RECT  7.010000 42.240000  7.210000 42.440000 ;
        RECT  7.010000 42.670000  7.210000 42.870000 ;
        RECT  7.010000 43.100000  7.210000 43.300000 ;
        RECT  7.010000 43.530000  7.210000 43.730000 ;
        RECT  7.010000 43.960000  7.210000 44.160000 ;
        RECT  7.410000 39.660000  7.610000 39.860000 ;
        RECT  7.410000 40.090000  7.610000 40.290000 ;
        RECT  7.410000 40.520000  7.610000 40.720000 ;
        RECT  7.410000 40.950000  7.610000 41.150000 ;
        RECT  7.410000 41.380000  7.610000 41.580000 ;
        RECT  7.410000 41.810000  7.610000 42.010000 ;
        RECT  7.410000 42.240000  7.610000 42.440000 ;
        RECT  7.410000 42.670000  7.610000 42.870000 ;
        RECT  7.410000 43.100000  7.610000 43.300000 ;
        RECT  7.410000 43.530000  7.610000 43.730000 ;
        RECT  7.410000 43.960000  7.610000 44.160000 ;
        RECT  7.810000 39.660000  8.010000 39.860000 ;
        RECT  7.810000 40.090000  8.010000 40.290000 ;
        RECT  7.810000 40.520000  8.010000 40.720000 ;
        RECT  7.810000 40.950000  8.010000 41.150000 ;
        RECT  7.810000 41.380000  8.010000 41.580000 ;
        RECT  7.810000 41.810000  8.010000 42.010000 ;
        RECT  7.810000 42.240000  8.010000 42.440000 ;
        RECT  7.810000 42.670000  8.010000 42.870000 ;
        RECT  7.810000 43.100000  8.010000 43.300000 ;
        RECT  7.810000 43.530000  8.010000 43.730000 ;
        RECT  7.810000 43.960000  8.010000 44.160000 ;
        RECT  8.210000 39.660000  8.410000 39.860000 ;
        RECT  8.210000 40.090000  8.410000 40.290000 ;
        RECT  8.210000 40.520000  8.410000 40.720000 ;
        RECT  8.210000 40.950000  8.410000 41.150000 ;
        RECT  8.210000 41.380000  8.410000 41.580000 ;
        RECT  8.210000 41.810000  8.410000 42.010000 ;
        RECT  8.210000 42.240000  8.410000 42.440000 ;
        RECT  8.210000 42.670000  8.410000 42.870000 ;
        RECT  8.210000 43.100000  8.410000 43.300000 ;
        RECT  8.210000 43.530000  8.410000 43.730000 ;
        RECT  8.210000 43.960000  8.410000 44.160000 ;
        RECT  8.610000 39.660000  8.810000 39.860000 ;
        RECT  8.610000 40.090000  8.810000 40.290000 ;
        RECT  8.610000 40.520000  8.810000 40.720000 ;
        RECT  8.610000 40.950000  8.810000 41.150000 ;
        RECT  8.610000 41.380000  8.810000 41.580000 ;
        RECT  8.610000 41.810000  8.810000 42.010000 ;
        RECT  8.610000 42.240000  8.810000 42.440000 ;
        RECT  8.610000 42.670000  8.810000 42.870000 ;
        RECT  8.610000 43.100000  8.810000 43.300000 ;
        RECT  8.610000 43.530000  8.810000 43.730000 ;
        RECT  8.610000 43.960000  8.810000 44.160000 ;
        RECT  9.010000 39.660000  9.210000 39.860000 ;
        RECT  9.010000 40.090000  9.210000 40.290000 ;
        RECT  9.010000 40.520000  9.210000 40.720000 ;
        RECT  9.010000 40.950000  9.210000 41.150000 ;
        RECT  9.010000 41.380000  9.210000 41.580000 ;
        RECT  9.010000 41.810000  9.210000 42.010000 ;
        RECT  9.010000 42.240000  9.210000 42.440000 ;
        RECT  9.010000 42.670000  9.210000 42.870000 ;
        RECT  9.010000 43.100000  9.210000 43.300000 ;
        RECT  9.010000 43.530000  9.210000 43.730000 ;
        RECT  9.010000 43.960000  9.210000 44.160000 ;
        RECT  9.410000 39.660000  9.610000 39.860000 ;
        RECT  9.410000 40.090000  9.610000 40.290000 ;
        RECT  9.410000 40.520000  9.610000 40.720000 ;
        RECT  9.410000 40.950000  9.610000 41.150000 ;
        RECT  9.410000 41.380000  9.610000 41.580000 ;
        RECT  9.410000 41.810000  9.610000 42.010000 ;
        RECT  9.410000 42.240000  9.610000 42.440000 ;
        RECT  9.410000 42.670000  9.610000 42.870000 ;
        RECT  9.410000 43.100000  9.610000 43.300000 ;
        RECT  9.410000 43.530000  9.610000 43.730000 ;
        RECT  9.410000 43.960000  9.610000 44.160000 ;
        RECT  9.810000 39.660000 10.010000 39.860000 ;
        RECT  9.810000 40.090000 10.010000 40.290000 ;
        RECT  9.810000 40.520000 10.010000 40.720000 ;
        RECT  9.810000 40.950000 10.010000 41.150000 ;
        RECT  9.810000 41.380000 10.010000 41.580000 ;
        RECT  9.810000 41.810000 10.010000 42.010000 ;
        RECT  9.810000 42.240000 10.010000 42.440000 ;
        RECT  9.810000 42.670000 10.010000 42.870000 ;
        RECT  9.810000 43.100000 10.010000 43.300000 ;
        RECT  9.810000 43.530000 10.010000 43.730000 ;
        RECT  9.810000 43.960000 10.010000 44.160000 ;
        RECT 10.210000 39.660000 10.410000 39.860000 ;
        RECT 10.210000 40.090000 10.410000 40.290000 ;
        RECT 10.210000 40.520000 10.410000 40.720000 ;
        RECT 10.210000 40.950000 10.410000 41.150000 ;
        RECT 10.210000 41.380000 10.410000 41.580000 ;
        RECT 10.210000 41.810000 10.410000 42.010000 ;
        RECT 10.210000 42.240000 10.410000 42.440000 ;
        RECT 10.210000 42.670000 10.410000 42.870000 ;
        RECT 10.210000 43.100000 10.410000 43.300000 ;
        RECT 10.210000 43.530000 10.410000 43.730000 ;
        RECT 10.210000 43.960000 10.410000 44.160000 ;
        RECT 10.610000 39.660000 10.810000 39.860000 ;
        RECT 10.610000 40.090000 10.810000 40.290000 ;
        RECT 10.610000 40.520000 10.810000 40.720000 ;
        RECT 10.610000 40.950000 10.810000 41.150000 ;
        RECT 10.610000 41.380000 10.810000 41.580000 ;
        RECT 10.610000 41.810000 10.810000 42.010000 ;
        RECT 10.610000 42.240000 10.810000 42.440000 ;
        RECT 10.610000 42.670000 10.810000 42.870000 ;
        RECT 10.610000 43.100000 10.810000 43.300000 ;
        RECT 10.610000 43.530000 10.810000 43.730000 ;
        RECT 10.610000 43.960000 10.810000 44.160000 ;
        RECT 11.010000 39.660000 11.210000 39.860000 ;
        RECT 11.010000 40.090000 11.210000 40.290000 ;
        RECT 11.010000 40.520000 11.210000 40.720000 ;
        RECT 11.010000 40.950000 11.210000 41.150000 ;
        RECT 11.010000 41.380000 11.210000 41.580000 ;
        RECT 11.010000 41.810000 11.210000 42.010000 ;
        RECT 11.010000 42.240000 11.210000 42.440000 ;
        RECT 11.010000 42.670000 11.210000 42.870000 ;
        RECT 11.010000 43.100000 11.210000 43.300000 ;
        RECT 11.010000 43.530000 11.210000 43.730000 ;
        RECT 11.010000 43.960000 11.210000 44.160000 ;
        RECT 11.410000 39.660000 11.610000 39.860000 ;
        RECT 11.410000 40.090000 11.610000 40.290000 ;
        RECT 11.410000 40.520000 11.610000 40.720000 ;
        RECT 11.410000 40.950000 11.610000 41.150000 ;
        RECT 11.410000 41.380000 11.610000 41.580000 ;
        RECT 11.410000 41.810000 11.610000 42.010000 ;
        RECT 11.410000 42.240000 11.610000 42.440000 ;
        RECT 11.410000 42.670000 11.610000 42.870000 ;
        RECT 11.410000 43.100000 11.610000 43.300000 ;
        RECT 11.410000 43.530000 11.610000 43.730000 ;
        RECT 11.410000 43.960000 11.610000 44.160000 ;
        RECT 11.810000 39.660000 12.010000 39.860000 ;
        RECT 11.810000 40.090000 12.010000 40.290000 ;
        RECT 11.810000 40.520000 12.010000 40.720000 ;
        RECT 11.810000 40.950000 12.010000 41.150000 ;
        RECT 11.810000 41.380000 12.010000 41.580000 ;
        RECT 11.810000 41.810000 12.010000 42.010000 ;
        RECT 11.810000 42.240000 12.010000 42.440000 ;
        RECT 11.810000 42.670000 12.010000 42.870000 ;
        RECT 11.810000 43.100000 12.010000 43.300000 ;
        RECT 11.810000 43.530000 12.010000 43.730000 ;
        RECT 11.810000 43.960000 12.010000 44.160000 ;
        RECT 12.210000 39.660000 12.410000 39.860000 ;
        RECT 12.210000 40.090000 12.410000 40.290000 ;
        RECT 12.210000 40.520000 12.410000 40.720000 ;
        RECT 12.210000 40.950000 12.410000 41.150000 ;
        RECT 12.210000 41.380000 12.410000 41.580000 ;
        RECT 12.210000 41.810000 12.410000 42.010000 ;
        RECT 12.210000 42.240000 12.410000 42.440000 ;
        RECT 12.210000 42.670000 12.410000 42.870000 ;
        RECT 12.210000 43.100000 12.410000 43.300000 ;
        RECT 12.210000 43.530000 12.410000 43.730000 ;
        RECT 12.210000 43.960000 12.410000 44.160000 ;
        RECT 12.610000 39.660000 12.810000 39.860000 ;
        RECT 12.610000 40.090000 12.810000 40.290000 ;
        RECT 12.610000 40.520000 12.810000 40.720000 ;
        RECT 12.610000 40.950000 12.810000 41.150000 ;
        RECT 12.610000 41.380000 12.810000 41.580000 ;
        RECT 12.610000 41.810000 12.810000 42.010000 ;
        RECT 12.610000 42.240000 12.810000 42.440000 ;
        RECT 12.610000 42.670000 12.810000 42.870000 ;
        RECT 12.610000 43.100000 12.810000 43.300000 ;
        RECT 12.610000 43.530000 12.810000 43.730000 ;
        RECT 12.610000 43.960000 12.810000 44.160000 ;
        RECT 13.010000 39.660000 13.210000 39.860000 ;
        RECT 13.010000 40.090000 13.210000 40.290000 ;
        RECT 13.010000 40.520000 13.210000 40.720000 ;
        RECT 13.010000 40.950000 13.210000 41.150000 ;
        RECT 13.010000 41.380000 13.210000 41.580000 ;
        RECT 13.010000 41.810000 13.210000 42.010000 ;
        RECT 13.010000 42.240000 13.210000 42.440000 ;
        RECT 13.010000 42.670000 13.210000 42.870000 ;
        RECT 13.010000 43.100000 13.210000 43.300000 ;
        RECT 13.010000 43.530000 13.210000 43.730000 ;
        RECT 13.010000 43.960000 13.210000 44.160000 ;
        RECT 13.410000 39.660000 13.610000 39.860000 ;
        RECT 13.410000 40.090000 13.610000 40.290000 ;
        RECT 13.410000 40.520000 13.610000 40.720000 ;
        RECT 13.410000 40.950000 13.610000 41.150000 ;
        RECT 13.410000 41.380000 13.610000 41.580000 ;
        RECT 13.410000 41.810000 13.610000 42.010000 ;
        RECT 13.410000 42.240000 13.610000 42.440000 ;
        RECT 13.410000 42.670000 13.610000 42.870000 ;
        RECT 13.410000 43.100000 13.610000 43.300000 ;
        RECT 13.410000 43.530000 13.610000 43.730000 ;
        RECT 13.410000 43.960000 13.610000 44.160000 ;
        RECT 13.810000 39.660000 14.010000 39.860000 ;
        RECT 13.810000 40.090000 14.010000 40.290000 ;
        RECT 13.810000 40.520000 14.010000 40.720000 ;
        RECT 13.810000 40.950000 14.010000 41.150000 ;
        RECT 13.810000 41.380000 14.010000 41.580000 ;
        RECT 13.810000 41.810000 14.010000 42.010000 ;
        RECT 13.810000 42.240000 14.010000 42.440000 ;
        RECT 13.810000 42.670000 14.010000 42.870000 ;
        RECT 13.810000 43.100000 14.010000 43.300000 ;
        RECT 13.810000 43.530000 14.010000 43.730000 ;
        RECT 13.810000 43.960000 14.010000 44.160000 ;
        RECT 14.210000 39.660000 14.410000 39.860000 ;
        RECT 14.210000 40.090000 14.410000 40.290000 ;
        RECT 14.210000 40.520000 14.410000 40.720000 ;
        RECT 14.210000 40.950000 14.410000 41.150000 ;
        RECT 14.210000 41.380000 14.410000 41.580000 ;
        RECT 14.210000 41.810000 14.410000 42.010000 ;
        RECT 14.210000 42.240000 14.410000 42.440000 ;
        RECT 14.210000 42.670000 14.410000 42.870000 ;
        RECT 14.210000 43.100000 14.410000 43.300000 ;
        RECT 14.210000 43.530000 14.410000 43.730000 ;
        RECT 14.210000 43.960000 14.410000 44.160000 ;
        RECT 14.610000 39.660000 14.810000 39.860000 ;
        RECT 14.610000 40.090000 14.810000 40.290000 ;
        RECT 14.610000 40.520000 14.810000 40.720000 ;
        RECT 14.610000 40.950000 14.810000 41.150000 ;
        RECT 14.610000 41.380000 14.810000 41.580000 ;
        RECT 14.610000 41.810000 14.810000 42.010000 ;
        RECT 14.610000 42.240000 14.810000 42.440000 ;
        RECT 14.610000 42.670000 14.810000 42.870000 ;
        RECT 14.610000 43.100000 14.810000 43.300000 ;
        RECT 14.610000 43.530000 14.810000 43.730000 ;
        RECT 14.610000 43.960000 14.810000 44.160000 ;
        RECT 15.010000 39.660000 15.210000 39.860000 ;
        RECT 15.010000 40.090000 15.210000 40.290000 ;
        RECT 15.010000 40.520000 15.210000 40.720000 ;
        RECT 15.010000 40.950000 15.210000 41.150000 ;
        RECT 15.010000 41.380000 15.210000 41.580000 ;
        RECT 15.010000 41.810000 15.210000 42.010000 ;
        RECT 15.010000 42.240000 15.210000 42.440000 ;
        RECT 15.010000 42.670000 15.210000 42.870000 ;
        RECT 15.010000 43.100000 15.210000 43.300000 ;
        RECT 15.010000 43.530000 15.210000 43.730000 ;
        RECT 15.010000 43.960000 15.210000 44.160000 ;
        RECT 15.410000 39.660000 15.610000 39.860000 ;
        RECT 15.410000 40.090000 15.610000 40.290000 ;
        RECT 15.410000 40.520000 15.610000 40.720000 ;
        RECT 15.410000 40.950000 15.610000 41.150000 ;
        RECT 15.410000 41.380000 15.610000 41.580000 ;
        RECT 15.410000 41.810000 15.610000 42.010000 ;
        RECT 15.410000 42.240000 15.610000 42.440000 ;
        RECT 15.410000 42.670000 15.610000 42.870000 ;
        RECT 15.410000 43.100000 15.610000 43.300000 ;
        RECT 15.410000 43.530000 15.610000 43.730000 ;
        RECT 15.410000 43.960000 15.610000 44.160000 ;
        RECT 15.810000 39.660000 16.010000 39.860000 ;
        RECT 15.810000 40.090000 16.010000 40.290000 ;
        RECT 15.810000 40.520000 16.010000 40.720000 ;
        RECT 15.810000 40.950000 16.010000 41.150000 ;
        RECT 15.810000 41.380000 16.010000 41.580000 ;
        RECT 15.810000 41.810000 16.010000 42.010000 ;
        RECT 15.810000 42.240000 16.010000 42.440000 ;
        RECT 15.810000 42.670000 16.010000 42.870000 ;
        RECT 15.810000 43.100000 16.010000 43.300000 ;
        RECT 15.810000 43.530000 16.010000 43.730000 ;
        RECT 15.810000 43.960000 16.010000 44.160000 ;
        RECT 16.210000 39.660000 16.410000 39.860000 ;
        RECT 16.210000 40.090000 16.410000 40.290000 ;
        RECT 16.210000 40.520000 16.410000 40.720000 ;
        RECT 16.210000 40.950000 16.410000 41.150000 ;
        RECT 16.210000 41.380000 16.410000 41.580000 ;
        RECT 16.210000 41.810000 16.410000 42.010000 ;
        RECT 16.210000 42.240000 16.410000 42.440000 ;
        RECT 16.210000 42.670000 16.410000 42.870000 ;
        RECT 16.210000 43.100000 16.410000 43.300000 ;
        RECT 16.210000 43.530000 16.410000 43.730000 ;
        RECT 16.210000 43.960000 16.410000 44.160000 ;
        RECT 16.610000 39.660000 16.810000 39.860000 ;
        RECT 16.610000 40.090000 16.810000 40.290000 ;
        RECT 16.610000 40.520000 16.810000 40.720000 ;
        RECT 16.610000 40.950000 16.810000 41.150000 ;
        RECT 16.610000 41.380000 16.810000 41.580000 ;
        RECT 16.610000 41.810000 16.810000 42.010000 ;
        RECT 16.610000 42.240000 16.810000 42.440000 ;
        RECT 16.610000 42.670000 16.810000 42.870000 ;
        RECT 16.610000 43.100000 16.810000 43.300000 ;
        RECT 16.610000 43.530000 16.810000 43.730000 ;
        RECT 16.610000 43.960000 16.810000 44.160000 ;
        RECT 17.010000 39.660000 17.210000 39.860000 ;
        RECT 17.010000 40.090000 17.210000 40.290000 ;
        RECT 17.010000 40.520000 17.210000 40.720000 ;
        RECT 17.010000 40.950000 17.210000 41.150000 ;
        RECT 17.010000 41.380000 17.210000 41.580000 ;
        RECT 17.010000 41.810000 17.210000 42.010000 ;
        RECT 17.010000 42.240000 17.210000 42.440000 ;
        RECT 17.010000 42.670000 17.210000 42.870000 ;
        RECT 17.010000 43.100000 17.210000 43.300000 ;
        RECT 17.010000 43.530000 17.210000 43.730000 ;
        RECT 17.010000 43.960000 17.210000 44.160000 ;
        RECT 17.410000 39.660000 17.610000 39.860000 ;
        RECT 17.410000 40.090000 17.610000 40.290000 ;
        RECT 17.410000 40.520000 17.610000 40.720000 ;
        RECT 17.410000 40.950000 17.610000 41.150000 ;
        RECT 17.410000 41.380000 17.610000 41.580000 ;
        RECT 17.410000 41.810000 17.610000 42.010000 ;
        RECT 17.410000 42.240000 17.610000 42.440000 ;
        RECT 17.410000 42.670000 17.610000 42.870000 ;
        RECT 17.410000 43.100000 17.610000 43.300000 ;
        RECT 17.410000 43.530000 17.610000 43.730000 ;
        RECT 17.410000 43.960000 17.610000 44.160000 ;
        RECT 17.810000 39.660000 18.010000 39.860000 ;
        RECT 17.810000 40.090000 18.010000 40.290000 ;
        RECT 17.810000 40.520000 18.010000 40.720000 ;
        RECT 17.810000 40.950000 18.010000 41.150000 ;
        RECT 17.810000 41.380000 18.010000 41.580000 ;
        RECT 17.810000 41.810000 18.010000 42.010000 ;
        RECT 17.810000 42.240000 18.010000 42.440000 ;
        RECT 17.810000 42.670000 18.010000 42.870000 ;
        RECT 17.810000 43.100000 18.010000 43.300000 ;
        RECT 17.810000 43.530000 18.010000 43.730000 ;
        RECT 17.810000 43.960000 18.010000 44.160000 ;
        RECT 18.210000 39.660000 18.410000 39.860000 ;
        RECT 18.210000 40.090000 18.410000 40.290000 ;
        RECT 18.210000 40.520000 18.410000 40.720000 ;
        RECT 18.210000 40.950000 18.410000 41.150000 ;
        RECT 18.210000 41.380000 18.410000 41.580000 ;
        RECT 18.210000 41.810000 18.410000 42.010000 ;
        RECT 18.210000 42.240000 18.410000 42.440000 ;
        RECT 18.210000 42.670000 18.410000 42.870000 ;
        RECT 18.210000 43.100000 18.410000 43.300000 ;
        RECT 18.210000 43.530000 18.410000 43.730000 ;
        RECT 18.210000 43.960000 18.410000 44.160000 ;
        RECT 18.610000 39.660000 18.810000 39.860000 ;
        RECT 18.610000 40.090000 18.810000 40.290000 ;
        RECT 18.610000 40.520000 18.810000 40.720000 ;
        RECT 18.610000 40.950000 18.810000 41.150000 ;
        RECT 18.610000 41.380000 18.810000 41.580000 ;
        RECT 18.610000 41.810000 18.810000 42.010000 ;
        RECT 18.610000 42.240000 18.810000 42.440000 ;
        RECT 18.610000 42.670000 18.810000 42.870000 ;
        RECT 18.610000 43.100000 18.810000 43.300000 ;
        RECT 18.610000 43.530000 18.810000 43.730000 ;
        RECT 18.610000 43.960000 18.810000 44.160000 ;
        RECT 19.010000 39.660000 19.210000 39.860000 ;
        RECT 19.010000 40.090000 19.210000 40.290000 ;
        RECT 19.010000 40.520000 19.210000 40.720000 ;
        RECT 19.010000 40.950000 19.210000 41.150000 ;
        RECT 19.010000 41.380000 19.210000 41.580000 ;
        RECT 19.010000 41.810000 19.210000 42.010000 ;
        RECT 19.010000 42.240000 19.210000 42.440000 ;
        RECT 19.010000 42.670000 19.210000 42.870000 ;
        RECT 19.010000 43.100000 19.210000 43.300000 ;
        RECT 19.010000 43.530000 19.210000 43.730000 ;
        RECT 19.010000 43.960000 19.210000 44.160000 ;
        RECT 19.410000 39.660000 19.610000 39.860000 ;
        RECT 19.410000 40.090000 19.610000 40.290000 ;
        RECT 19.410000 40.520000 19.610000 40.720000 ;
        RECT 19.410000 40.950000 19.610000 41.150000 ;
        RECT 19.410000 41.380000 19.610000 41.580000 ;
        RECT 19.410000 41.810000 19.610000 42.010000 ;
        RECT 19.410000 42.240000 19.610000 42.440000 ;
        RECT 19.410000 42.670000 19.610000 42.870000 ;
        RECT 19.410000 43.100000 19.610000 43.300000 ;
        RECT 19.410000 43.530000 19.610000 43.730000 ;
        RECT 19.410000 43.960000 19.610000 44.160000 ;
        RECT 19.810000 39.660000 20.010000 39.860000 ;
        RECT 19.810000 40.090000 20.010000 40.290000 ;
        RECT 19.810000 40.520000 20.010000 40.720000 ;
        RECT 19.810000 40.950000 20.010000 41.150000 ;
        RECT 19.810000 41.380000 20.010000 41.580000 ;
        RECT 19.810000 41.810000 20.010000 42.010000 ;
        RECT 19.810000 42.240000 20.010000 42.440000 ;
        RECT 19.810000 42.670000 20.010000 42.870000 ;
        RECT 19.810000 43.100000 20.010000 43.300000 ;
        RECT 19.810000 43.530000 20.010000 43.730000 ;
        RECT 19.810000 43.960000 20.010000 44.160000 ;
        RECT 20.210000 39.660000 20.410000 39.860000 ;
        RECT 20.210000 40.090000 20.410000 40.290000 ;
        RECT 20.210000 40.520000 20.410000 40.720000 ;
        RECT 20.210000 40.950000 20.410000 41.150000 ;
        RECT 20.210000 41.380000 20.410000 41.580000 ;
        RECT 20.210000 41.810000 20.410000 42.010000 ;
        RECT 20.210000 42.240000 20.410000 42.440000 ;
        RECT 20.210000 42.670000 20.410000 42.870000 ;
        RECT 20.210000 43.100000 20.410000 43.300000 ;
        RECT 20.210000 43.530000 20.410000 43.730000 ;
        RECT 20.210000 43.960000 20.410000 44.160000 ;
        RECT 20.610000 39.660000 20.810000 39.860000 ;
        RECT 20.610000 40.090000 20.810000 40.290000 ;
        RECT 20.610000 40.520000 20.810000 40.720000 ;
        RECT 20.610000 40.950000 20.810000 41.150000 ;
        RECT 20.610000 41.380000 20.810000 41.580000 ;
        RECT 20.610000 41.810000 20.810000 42.010000 ;
        RECT 20.610000 42.240000 20.810000 42.440000 ;
        RECT 20.610000 42.670000 20.810000 42.870000 ;
        RECT 20.610000 43.100000 20.810000 43.300000 ;
        RECT 20.610000 43.530000 20.810000 43.730000 ;
        RECT 20.610000 43.960000 20.810000 44.160000 ;
        RECT 21.010000 39.660000 21.210000 39.860000 ;
        RECT 21.010000 40.090000 21.210000 40.290000 ;
        RECT 21.010000 40.520000 21.210000 40.720000 ;
        RECT 21.010000 40.950000 21.210000 41.150000 ;
        RECT 21.010000 41.380000 21.210000 41.580000 ;
        RECT 21.010000 41.810000 21.210000 42.010000 ;
        RECT 21.010000 42.240000 21.210000 42.440000 ;
        RECT 21.010000 42.670000 21.210000 42.870000 ;
        RECT 21.010000 43.100000 21.210000 43.300000 ;
        RECT 21.010000 43.530000 21.210000 43.730000 ;
        RECT 21.010000 43.960000 21.210000 44.160000 ;
        RECT 21.410000 39.660000 21.610000 39.860000 ;
        RECT 21.410000 40.090000 21.610000 40.290000 ;
        RECT 21.410000 40.520000 21.610000 40.720000 ;
        RECT 21.410000 40.950000 21.610000 41.150000 ;
        RECT 21.410000 41.380000 21.610000 41.580000 ;
        RECT 21.410000 41.810000 21.610000 42.010000 ;
        RECT 21.410000 42.240000 21.610000 42.440000 ;
        RECT 21.410000 42.670000 21.610000 42.870000 ;
        RECT 21.410000 43.100000 21.610000 43.300000 ;
        RECT 21.410000 43.530000 21.610000 43.730000 ;
        RECT 21.410000 43.960000 21.610000 44.160000 ;
        RECT 21.810000 39.660000 22.010000 39.860000 ;
        RECT 21.810000 40.090000 22.010000 40.290000 ;
        RECT 21.810000 40.520000 22.010000 40.720000 ;
        RECT 21.810000 40.950000 22.010000 41.150000 ;
        RECT 21.810000 41.380000 22.010000 41.580000 ;
        RECT 21.810000 41.810000 22.010000 42.010000 ;
        RECT 21.810000 42.240000 22.010000 42.440000 ;
        RECT 21.810000 42.670000 22.010000 42.870000 ;
        RECT 21.810000 43.100000 22.010000 43.300000 ;
        RECT 21.810000 43.530000 22.010000 43.730000 ;
        RECT 21.810000 43.960000 22.010000 44.160000 ;
        RECT 22.210000 39.660000 22.410000 39.860000 ;
        RECT 22.210000 40.090000 22.410000 40.290000 ;
        RECT 22.210000 40.520000 22.410000 40.720000 ;
        RECT 22.210000 40.950000 22.410000 41.150000 ;
        RECT 22.210000 41.380000 22.410000 41.580000 ;
        RECT 22.210000 41.810000 22.410000 42.010000 ;
        RECT 22.210000 42.240000 22.410000 42.440000 ;
        RECT 22.210000 42.670000 22.410000 42.870000 ;
        RECT 22.210000 43.100000 22.410000 43.300000 ;
        RECT 22.210000 43.530000 22.410000 43.730000 ;
        RECT 22.210000 43.960000 22.410000 44.160000 ;
        RECT 22.610000 39.660000 22.810000 39.860000 ;
        RECT 22.610000 40.090000 22.810000 40.290000 ;
        RECT 22.610000 40.520000 22.810000 40.720000 ;
        RECT 22.610000 40.950000 22.810000 41.150000 ;
        RECT 22.610000 41.380000 22.810000 41.580000 ;
        RECT 22.610000 41.810000 22.810000 42.010000 ;
        RECT 22.610000 42.240000 22.810000 42.440000 ;
        RECT 22.610000 42.670000 22.810000 42.870000 ;
        RECT 22.610000 43.100000 22.810000 43.300000 ;
        RECT 22.610000 43.530000 22.810000 43.730000 ;
        RECT 22.610000 43.960000 22.810000 44.160000 ;
        RECT 23.010000 39.660000 23.210000 39.860000 ;
        RECT 23.010000 40.090000 23.210000 40.290000 ;
        RECT 23.010000 40.520000 23.210000 40.720000 ;
        RECT 23.010000 40.950000 23.210000 41.150000 ;
        RECT 23.010000 41.380000 23.210000 41.580000 ;
        RECT 23.010000 41.810000 23.210000 42.010000 ;
        RECT 23.010000 42.240000 23.210000 42.440000 ;
        RECT 23.010000 42.670000 23.210000 42.870000 ;
        RECT 23.010000 43.100000 23.210000 43.300000 ;
        RECT 23.010000 43.530000 23.210000 43.730000 ;
        RECT 23.010000 43.960000 23.210000 44.160000 ;
        RECT 23.410000 39.660000 23.610000 39.860000 ;
        RECT 23.410000 40.090000 23.610000 40.290000 ;
        RECT 23.410000 40.520000 23.610000 40.720000 ;
        RECT 23.410000 40.950000 23.610000 41.150000 ;
        RECT 23.410000 41.380000 23.610000 41.580000 ;
        RECT 23.410000 41.810000 23.610000 42.010000 ;
        RECT 23.410000 42.240000 23.610000 42.440000 ;
        RECT 23.410000 42.670000 23.610000 42.870000 ;
        RECT 23.410000 43.100000 23.610000 43.300000 ;
        RECT 23.410000 43.530000 23.610000 43.730000 ;
        RECT 23.410000 43.960000 23.610000 44.160000 ;
        RECT 23.810000 39.660000 24.010000 39.860000 ;
        RECT 23.810000 40.090000 24.010000 40.290000 ;
        RECT 23.810000 40.520000 24.010000 40.720000 ;
        RECT 23.810000 40.950000 24.010000 41.150000 ;
        RECT 23.810000 41.380000 24.010000 41.580000 ;
        RECT 23.810000 41.810000 24.010000 42.010000 ;
        RECT 23.810000 42.240000 24.010000 42.440000 ;
        RECT 23.810000 42.670000 24.010000 42.870000 ;
        RECT 23.810000 43.100000 24.010000 43.300000 ;
        RECT 23.810000 43.530000 24.010000 43.730000 ;
        RECT 23.810000 43.960000 24.010000 44.160000 ;
        RECT 24.210000 39.660000 24.410000 39.860000 ;
        RECT 24.210000 40.090000 24.410000 40.290000 ;
        RECT 24.210000 40.520000 24.410000 40.720000 ;
        RECT 24.210000 40.950000 24.410000 41.150000 ;
        RECT 24.210000 41.380000 24.410000 41.580000 ;
        RECT 24.210000 41.810000 24.410000 42.010000 ;
        RECT 24.210000 42.240000 24.410000 42.440000 ;
        RECT 24.210000 42.670000 24.410000 42.870000 ;
        RECT 24.210000 43.100000 24.410000 43.300000 ;
        RECT 24.210000 43.530000 24.410000 43.730000 ;
        RECT 24.210000 43.960000 24.410000 44.160000 ;
        RECT 50.845000 39.660000 51.045000 39.860000 ;
        RECT 50.845000 40.090000 51.045000 40.290000 ;
        RECT 50.845000 40.520000 51.045000 40.720000 ;
        RECT 50.845000 40.950000 51.045000 41.150000 ;
        RECT 50.845000 41.380000 51.045000 41.580000 ;
        RECT 50.845000 41.810000 51.045000 42.010000 ;
        RECT 50.845000 42.240000 51.045000 42.440000 ;
        RECT 50.845000 42.670000 51.045000 42.870000 ;
        RECT 50.845000 43.100000 51.045000 43.300000 ;
        RECT 50.845000 43.530000 51.045000 43.730000 ;
        RECT 50.845000 43.960000 51.045000 44.160000 ;
        RECT 51.255000 39.660000 51.455000 39.860000 ;
        RECT 51.255000 40.090000 51.455000 40.290000 ;
        RECT 51.255000 40.520000 51.455000 40.720000 ;
        RECT 51.255000 40.950000 51.455000 41.150000 ;
        RECT 51.255000 41.380000 51.455000 41.580000 ;
        RECT 51.255000 41.810000 51.455000 42.010000 ;
        RECT 51.255000 42.240000 51.455000 42.440000 ;
        RECT 51.255000 42.670000 51.455000 42.870000 ;
        RECT 51.255000 43.100000 51.455000 43.300000 ;
        RECT 51.255000 43.530000 51.455000 43.730000 ;
        RECT 51.255000 43.960000 51.455000 44.160000 ;
        RECT 51.665000 39.660000 51.865000 39.860000 ;
        RECT 51.665000 40.090000 51.865000 40.290000 ;
        RECT 51.665000 40.520000 51.865000 40.720000 ;
        RECT 51.665000 40.950000 51.865000 41.150000 ;
        RECT 51.665000 41.380000 51.865000 41.580000 ;
        RECT 51.665000 41.810000 51.865000 42.010000 ;
        RECT 51.665000 42.240000 51.865000 42.440000 ;
        RECT 51.665000 42.670000 51.865000 42.870000 ;
        RECT 51.665000 43.100000 51.865000 43.300000 ;
        RECT 51.665000 43.530000 51.865000 43.730000 ;
        RECT 51.665000 43.960000 51.865000 44.160000 ;
        RECT 52.075000 39.660000 52.275000 39.860000 ;
        RECT 52.075000 40.090000 52.275000 40.290000 ;
        RECT 52.075000 40.520000 52.275000 40.720000 ;
        RECT 52.075000 40.950000 52.275000 41.150000 ;
        RECT 52.075000 41.380000 52.275000 41.580000 ;
        RECT 52.075000 41.810000 52.275000 42.010000 ;
        RECT 52.075000 42.240000 52.275000 42.440000 ;
        RECT 52.075000 42.670000 52.275000 42.870000 ;
        RECT 52.075000 43.100000 52.275000 43.300000 ;
        RECT 52.075000 43.530000 52.275000 43.730000 ;
        RECT 52.075000 43.960000 52.275000 44.160000 ;
        RECT 52.485000 39.660000 52.685000 39.860000 ;
        RECT 52.485000 40.090000 52.685000 40.290000 ;
        RECT 52.485000 40.520000 52.685000 40.720000 ;
        RECT 52.485000 40.950000 52.685000 41.150000 ;
        RECT 52.485000 41.380000 52.685000 41.580000 ;
        RECT 52.485000 41.810000 52.685000 42.010000 ;
        RECT 52.485000 42.240000 52.685000 42.440000 ;
        RECT 52.485000 42.670000 52.685000 42.870000 ;
        RECT 52.485000 43.100000 52.685000 43.300000 ;
        RECT 52.485000 43.530000 52.685000 43.730000 ;
        RECT 52.485000 43.960000 52.685000 44.160000 ;
        RECT 52.895000 39.660000 53.095000 39.860000 ;
        RECT 52.895000 40.090000 53.095000 40.290000 ;
        RECT 52.895000 40.520000 53.095000 40.720000 ;
        RECT 52.895000 40.950000 53.095000 41.150000 ;
        RECT 52.895000 41.380000 53.095000 41.580000 ;
        RECT 52.895000 41.810000 53.095000 42.010000 ;
        RECT 52.895000 42.240000 53.095000 42.440000 ;
        RECT 52.895000 42.670000 53.095000 42.870000 ;
        RECT 52.895000 43.100000 53.095000 43.300000 ;
        RECT 52.895000 43.530000 53.095000 43.730000 ;
        RECT 52.895000 43.960000 53.095000 44.160000 ;
        RECT 53.305000 39.660000 53.505000 39.860000 ;
        RECT 53.305000 40.090000 53.505000 40.290000 ;
        RECT 53.305000 40.520000 53.505000 40.720000 ;
        RECT 53.305000 40.950000 53.505000 41.150000 ;
        RECT 53.305000 41.380000 53.505000 41.580000 ;
        RECT 53.305000 41.810000 53.505000 42.010000 ;
        RECT 53.305000 42.240000 53.505000 42.440000 ;
        RECT 53.305000 42.670000 53.505000 42.870000 ;
        RECT 53.305000 43.100000 53.505000 43.300000 ;
        RECT 53.305000 43.530000 53.505000 43.730000 ;
        RECT 53.305000 43.960000 53.505000 44.160000 ;
        RECT 53.715000 39.660000 53.915000 39.860000 ;
        RECT 53.715000 40.090000 53.915000 40.290000 ;
        RECT 53.715000 40.520000 53.915000 40.720000 ;
        RECT 53.715000 40.950000 53.915000 41.150000 ;
        RECT 53.715000 41.380000 53.915000 41.580000 ;
        RECT 53.715000 41.810000 53.915000 42.010000 ;
        RECT 53.715000 42.240000 53.915000 42.440000 ;
        RECT 53.715000 42.670000 53.915000 42.870000 ;
        RECT 53.715000 43.100000 53.915000 43.300000 ;
        RECT 53.715000 43.530000 53.915000 43.730000 ;
        RECT 53.715000 43.960000 53.915000 44.160000 ;
        RECT 54.125000 39.660000 54.325000 39.860000 ;
        RECT 54.125000 40.090000 54.325000 40.290000 ;
        RECT 54.125000 40.520000 54.325000 40.720000 ;
        RECT 54.125000 40.950000 54.325000 41.150000 ;
        RECT 54.125000 41.380000 54.325000 41.580000 ;
        RECT 54.125000 41.810000 54.325000 42.010000 ;
        RECT 54.125000 42.240000 54.325000 42.440000 ;
        RECT 54.125000 42.670000 54.325000 42.870000 ;
        RECT 54.125000 43.100000 54.325000 43.300000 ;
        RECT 54.125000 43.530000 54.325000 43.730000 ;
        RECT 54.125000 43.960000 54.325000 44.160000 ;
        RECT 54.535000 39.660000 54.735000 39.860000 ;
        RECT 54.535000 40.090000 54.735000 40.290000 ;
        RECT 54.535000 40.520000 54.735000 40.720000 ;
        RECT 54.535000 40.950000 54.735000 41.150000 ;
        RECT 54.535000 41.380000 54.735000 41.580000 ;
        RECT 54.535000 41.810000 54.735000 42.010000 ;
        RECT 54.535000 42.240000 54.735000 42.440000 ;
        RECT 54.535000 42.670000 54.735000 42.870000 ;
        RECT 54.535000 43.100000 54.735000 43.300000 ;
        RECT 54.535000 43.530000 54.735000 43.730000 ;
        RECT 54.535000 43.960000 54.735000 44.160000 ;
        RECT 54.945000 39.660000 55.145000 39.860000 ;
        RECT 54.945000 40.090000 55.145000 40.290000 ;
        RECT 54.945000 40.520000 55.145000 40.720000 ;
        RECT 54.945000 40.950000 55.145000 41.150000 ;
        RECT 54.945000 41.380000 55.145000 41.580000 ;
        RECT 54.945000 41.810000 55.145000 42.010000 ;
        RECT 54.945000 42.240000 55.145000 42.440000 ;
        RECT 54.945000 42.670000 55.145000 42.870000 ;
        RECT 54.945000 43.100000 55.145000 43.300000 ;
        RECT 54.945000 43.530000 55.145000 43.730000 ;
        RECT 54.945000 43.960000 55.145000 44.160000 ;
        RECT 55.355000 39.660000 55.555000 39.860000 ;
        RECT 55.355000 40.090000 55.555000 40.290000 ;
        RECT 55.355000 40.520000 55.555000 40.720000 ;
        RECT 55.355000 40.950000 55.555000 41.150000 ;
        RECT 55.355000 41.380000 55.555000 41.580000 ;
        RECT 55.355000 41.810000 55.555000 42.010000 ;
        RECT 55.355000 42.240000 55.555000 42.440000 ;
        RECT 55.355000 42.670000 55.555000 42.870000 ;
        RECT 55.355000 43.100000 55.555000 43.300000 ;
        RECT 55.355000 43.530000 55.555000 43.730000 ;
        RECT 55.355000 43.960000 55.555000 44.160000 ;
        RECT 55.765000 39.660000 55.965000 39.860000 ;
        RECT 55.765000 40.090000 55.965000 40.290000 ;
        RECT 55.765000 40.520000 55.965000 40.720000 ;
        RECT 55.765000 40.950000 55.965000 41.150000 ;
        RECT 55.765000 41.380000 55.965000 41.580000 ;
        RECT 55.765000 41.810000 55.965000 42.010000 ;
        RECT 55.765000 42.240000 55.965000 42.440000 ;
        RECT 55.765000 42.670000 55.965000 42.870000 ;
        RECT 55.765000 43.100000 55.965000 43.300000 ;
        RECT 55.765000 43.530000 55.965000 43.730000 ;
        RECT 55.765000 43.960000 55.965000 44.160000 ;
        RECT 56.175000 39.660000 56.375000 39.860000 ;
        RECT 56.175000 40.090000 56.375000 40.290000 ;
        RECT 56.175000 40.520000 56.375000 40.720000 ;
        RECT 56.175000 40.950000 56.375000 41.150000 ;
        RECT 56.175000 41.380000 56.375000 41.580000 ;
        RECT 56.175000 41.810000 56.375000 42.010000 ;
        RECT 56.175000 42.240000 56.375000 42.440000 ;
        RECT 56.175000 42.670000 56.375000 42.870000 ;
        RECT 56.175000 43.100000 56.375000 43.300000 ;
        RECT 56.175000 43.530000 56.375000 43.730000 ;
        RECT 56.175000 43.960000 56.375000 44.160000 ;
        RECT 56.585000 39.660000 56.785000 39.860000 ;
        RECT 56.585000 40.090000 56.785000 40.290000 ;
        RECT 56.585000 40.520000 56.785000 40.720000 ;
        RECT 56.585000 40.950000 56.785000 41.150000 ;
        RECT 56.585000 41.380000 56.785000 41.580000 ;
        RECT 56.585000 41.810000 56.785000 42.010000 ;
        RECT 56.585000 42.240000 56.785000 42.440000 ;
        RECT 56.585000 42.670000 56.785000 42.870000 ;
        RECT 56.585000 43.100000 56.785000 43.300000 ;
        RECT 56.585000 43.530000 56.785000 43.730000 ;
        RECT 56.585000 43.960000 56.785000 44.160000 ;
        RECT 56.995000 39.660000 57.195000 39.860000 ;
        RECT 56.995000 40.090000 57.195000 40.290000 ;
        RECT 56.995000 40.520000 57.195000 40.720000 ;
        RECT 56.995000 40.950000 57.195000 41.150000 ;
        RECT 56.995000 41.380000 57.195000 41.580000 ;
        RECT 56.995000 41.810000 57.195000 42.010000 ;
        RECT 56.995000 42.240000 57.195000 42.440000 ;
        RECT 56.995000 42.670000 57.195000 42.870000 ;
        RECT 56.995000 43.100000 57.195000 43.300000 ;
        RECT 56.995000 43.530000 57.195000 43.730000 ;
        RECT 56.995000 43.960000 57.195000 44.160000 ;
        RECT 57.400000 39.660000 57.600000 39.860000 ;
        RECT 57.400000 40.090000 57.600000 40.290000 ;
        RECT 57.400000 40.520000 57.600000 40.720000 ;
        RECT 57.400000 40.950000 57.600000 41.150000 ;
        RECT 57.400000 41.380000 57.600000 41.580000 ;
        RECT 57.400000 41.810000 57.600000 42.010000 ;
        RECT 57.400000 42.240000 57.600000 42.440000 ;
        RECT 57.400000 42.670000 57.600000 42.870000 ;
        RECT 57.400000 43.100000 57.600000 43.300000 ;
        RECT 57.400000 43.530000 57.600000 43.730000 ;
        RECT 57.400000 43.960000 57.600000 44.160000 ;
        RECT 57.805000 39.660000 58.005000 39.860000 ;
        RECT 57.805000 40.090000 58.005000 40.290000 ;
        RECT 57.805000 40.520000 58.005000 40.720000 ;
        RECT 57.805000 40.950000 58.005000 41.150000 ;
        RECT 57.805000 41.380000 58.005000 41.580000 ;
        RECT 57.805000 41.810000 58.005000 42.010000 ;
        RECT 57.805000 42.240000 58.005000 42.440000 ;
        RECT 57.805000 42.670000 58.005000 42.870000 ;
        RECT 57.805000 43.100000 58.005000 43.300000 ;
        RECT 57.805000 43.530000 58.005000 43.730000 ;
        RECT 57.805000 43.960000 58.005000 44.160000 ;
        RECT 58.210000 39.660000 58.410000 39.860000 ;
        RECT 58.210000 40.090000 58.410000 40.290000 ;
        RECT 58.210000 40.520000 58.410000 40.720000 ;
        RECT 58.210000 40.950000 58.410000 41.150000 ;
        RECT 58.210000 41.380000 58.410000 41.580000 ;
        RECT 58.210000 41.810000 58.410000 42.010000 ;
        RECT 58.210000 42.240000 58.410000 42.440000 ;
        RECT 58.210000 42.670000 58.410000 42.870000 ;
        RECT 58.210000 43.100000 58.410000 43.300000 ;
        RECT 58.210000 43.530000 58.410000 43.730000 ;
        RECT 58.210000 43.960000 58.410000 44.160000 ;
        RECT 58.615000 39.660000 58.815000 39.860000 ;
        RECT 58.615000 40.090000 58.815000 40.290000 ;
        RECT 58.615000 40.520000 58.815000 40.720000 ;
        RECT 58.615000 40.950000 58.815000 41.150000 ;
        RECT 58.615000 41.380000 58.815000 41.580000 ;
        RECT 58.615000 41.810000 58.815000 42.010000 ;
        RECT 58.615000 42.240000 58.815000 42.440000 ;
        RECT 58.615000 42.670000 58.815000 42.870000 ;
        RECT 58.615000 43.100000 58.815000 43.300000 ;
        RECT 58.615000 43.530000 58.815000 43.730000 ;
        RECT 58.615000 43.960000 58.815000 44.160000 ;
        RECT 59.020000 39.660000 59.220000 39.860000 ;
        RECT 59.020000 40.090000 59.220000 40.290000 ;
        RECT 59.020000 40.520000 59.220000 40.720000 ;
        RECT 59.020000 40.950000 59.220000 41.150000 ;
        RECT 59.020000 41.380000 59.220000 41.580000 ;
        RECT 59.020000 41.810000 59.220000 42.010000 ;
        RECT 59.020000 42.240000 59.220000 42.440000 ;
        RECT 59.020000 42.670000 59.220000 42.870000 ;
        RECT 59.020000 43.100000 59.220000 43.300000 ;
        RECT 59.020000 43.530000 59.220000 43.730000 ;
        RECT 59.020000 43.960000 59.220000 44.160000 ;
        RECT 59.425000 39.660000 59.625000 39.860000 ;
        RECT 59.425000 40.090000 59.625000 40.290000 ;
        RECT 59.425000 40.520000 59.625000 40.720000 ;
        RECT 59.425000 40.950000 59.625000 41.150000 ;
        RECT 59.425000 41.380000 59.625000 41.580000 ;
        RECT 59.425000 41.810000 59.625000 42.010000 ;
        RECT 59.425000 42.240000 59.625000 42.440000 ;
        RECT 59.425000 42.670000 59.625000 42.870000 ;
        RECT 59.425000 43.100000 59.625000 43.300000 ;
        RECT 59.425000 43.530000 59.625000 43.730000 ;
        RECT 59.425000 43.960000 59.625000 44.160000 ;
        RECT 59.830000 39.660000 60.030000 39.860000 ;
        RECT 59.830000 40.090000 60.030000 40.290000 ;
        RECT 59.830000 40.520000 60.030000 40.720000 ;
        RECT 59.830000 40.950000 60.030000 41.150000 ;
        RECT 59.830000 41.380000 60.030000 41.580000 ;
        RECT 59.830000 41.810000 60.030000 42.010000 ;
        RECT 59.830000 42.240000 60.030000 42.440000 ;
        RECT 59.830000 42.670000 60.030000 42.870000 ;
        RECT 59.830000 43.100000 60.030000 43.300000 ;
        RECT 59.830000 43.530000 60.030000 43.730000 ;
        RECT 59.830000 43.960000 60.030000 44.160000 ;
        RECT 60.235000 39.660000 60.435000 39.860000 ;
        RECT 60.235000 40.090000 60.435000 40.290000 ;
        RECT 60.235000 40.520000 60.435000 40.720000 ;
        RECT 60.235000 40.950000 60.435000 41.150000 ;
        RECT 60.235000 41.380000 60.435000 41.580000 ;
        RECT 60.235000 41.810000 60.435000 42.010000 ;
        RECT 60.235000 42.240000 60.435000 42.440000 ;
        RECT 60.235000 42.670000 60.435000 42.870000 ;
        RECT 60.235000 43.100000 60.435000 43.300000 ;
        RECT 60.235000 43.530000 60.435000 43.730000 ;
        RECT 60.235000 43.960000 60.435000 44.160000 ;
        RECT 60.640000 39.660000 60.840000 39.860000 ;
        RECT 60.640000 40.090000 60.840000 40.290000 ;
        RECT 60.640000 40.520000 60.840000 40.720000 ;
        RECT 60.640000 40.950000 60.840000 41.150000 ;
        RECT 60.640000 41.380000 60.840000 41.580000 ;
        RECT 60.640000 41.810000 60.840000 42.010000 ;
        RECT 60.640000 42.240000 60.840000 42.440000 ;
        RECT 60.640000 42.670000 60.840000 42.870000 ;
        RECT 60.640000 43.100000 60.840000 43.300000 ;
        RECT 60.640000 43.530000 60.840000 43.730000 ;
        RECT 60.640000 43.960000 60.840000 44.160000 ;
        RECT 61.045000 39.660000 61.245000 39.860000 ;
        RECT 61.045000 40.090000 61.245000 40.290000 ;
        RECT 61.045000 40.520000 61.245000 40.720000 ;
        RECT 61.045000 40.950000 61.245000 41.150000 ;
        RECT 61.045000 41.380000 61.245000 41.580000 ;
        RECT 61.045000 41.810000 61.245000 42.010000 ;
        RECT 61.045000 42.240000 61.245000 42.440000 ;
        RECT 61.045000 42.670000 61.245000 42.870000 ;
        RECT 61.045000 43.100000 61.245000 43.300000 ;
        RECT 61.045000 43.530000 61.245000 43.730000 ;
        RECT 61.045000 43.960000 61.245000 44.160000 ;
        RECT 61.450000 39.660000 61.650000 39.860000 ;
        RECT 61.450000 40.090000 61.650000 40.290000 ;
        RECT 61.450000 40.520000 61.650000 40.720000 ;
        RECT 61.450000 40.950000 61.650000 41.150000 ;
        RECT 61.450000 41.380000 61.650000 41.580000 ;
        RECT 61.450000 41.810000 61.650000 42.010000 ;
        RECT 61.450000 42.240000 61.650000 42.440000 ;
        RECT 61.450000 42.670000 61.650000 42.870000 ;
        RECT 61.450000 43.100000 61.650000 43.300000 ;
        RECT 61.450000 43.530000 61.650000 43.730000 ;
        RECT 61.450000 43.960000 61.650000 44.160000 ;
        RECT 61.855000 39.660000 62.055000 39.860000 ;
        RECT 61.855000 40.090000 62.055000 40.290000 ;
        RECT 61.855000 40.520000 62.055000 40.720000 ;
        RECT 61.855000 40.950000 62.055000 41.150000 ;
        RECT 61.855000 41.380000 62.055000 41.580000 ;
        RECT 61.855000 41.810000 62.055000 42.010000 ;
        RECT 61.855000 42.240000 62.055000 42.440000 ;
        RECT 61.855000 42.670000 62.055000 42.870000 ;
        RECT 61.855000 43.100000 62.055000 43.300000 ;
        RECT 61.855000 43.530000 62.055000 43.730000 ;
        RECT 61.855000 43.960000 62.055000 44.160000 ;
        RECT 62.260000 39.660000 62.460000 39.860000 ;
        RECT 62.260000 40.090000 62.460000 40.290000 ;
        RECT 62.260000 40.520000 62.460000 40.720000 ;
        RECT 62.260000 40.950000 62.460000 41.150000 ;
        RECT 62.260000 41.380000 62.460000 41.580000 ;
        RECT 62.260000 41.810000 62.460000 42.010000 ;
        RECT 62.260000 42.240000 62.460000 42.440000 ;
        RECT 62.260000 42.670000 62.460000 42.870000 ;
        RECT 62.260000 43.100000 62.460000 43.300000 ;
        RECT 62.260000 43.530000 62.460000 43.730000 ;
        RECT 62.260000 43.960000 62.460000 44.160000 ;
        RECT 62.665000 39.660000 62.865000 39.860000 ;
        RECT 62.665000 40.090000 62.865000 40.290000 ;
        RECT 62.665000 40.520000 62.865000 40.720000 ;
        RECT 62.665000 40.950000 62.865000 41.150000 ;
        RECT 62.665000 41.380000 62.865000 41.580000 ;
        RECT 62.665000 41.810000 62.865000 42.010000 ;
        RECT 62.665000 42.240000 62.865000 42.440000 ;
        RECT 62.665000 42.670000 62.865000 42.870000 ;
        RECT 62.665000 43.100000 62.865000 43.300000 ;
        RECT 62.665000 43.530000 62.865000 43.730000 ;
        RECT 62.665000 43.960000 62.865000 44.160000 ;
        RECT 63.070000 39.660000 63.270000 39.860000 ;
        RECT 63.070000 40.090000 63.270000 40.290000 ;
        RECT 63.070000 40.520000 63.270000 40.720000 ;
        RECT 63.070000 40.950000 63.270000 41.150000 ;
        RECT 63.070000 41.380000 63.270000 41.580000 ;
        RECT 63.070000 41.810000 63.270000 42.010000 ;
        RECT 63.070000 42.240000 63.270000 42.440000 ;
        RECT 63.070000 42.670000 63.270000 42.870000 ;
        RECT 63.070000 43.100000 63.270000 43.300000 ;
        RECT 63.070000 43.530000 63.270000 43.730000 ;
        RECT 63.070000 43.960000 63.270000 44.160000 ;
        RECT 63.475000 39.660000 63.675000 39.860000 ;
        RECT 63.475000 40.090000 63.675000 40.290000 ;
        RECT 63.475000 40.520000 63.675000 40.720000 ;
        RECT 63.475000 40.950000 63.675000 41.150000 ;
        RECT 63.475000 41.380000 63.675000 41.580000 ;
        RECT 63.475000 41.810000 63.675000 42.010000 ;
        RECT 63.475000 42.240000 63.675000 42.440000 ;
        RECT 63.475000 42.670000 63.675000 42.870000 ;
        RECT 63.475000 43.100000 63.675000 43.300000 ;
        RECT 63.475000 43.530000 63.675000 43.730000 ;
        RECT 63.475000 43.960000 63.675000 44.160000 ;
        RECT 63.880000 39.660000 64.080000 39.860000 ;
        RECT 63.880000 40.090000 64.080000 40.290000 ;
        RECT 63.880000 40.520000 64.080000 40.720000 ;
        RECT 63.880000 40.950000 64.080000 41.150000 ;
        RECT 63.880000 41.380000 64.080000 41.580000 ;
        RECT 63.880000 41.810000 64.080000 42.010000 ;
        RECT 63.880000 42.240000 64.080000 42.440000 ;
        RECT 63.880000 42.670000 64.080000 42.870000 ;
        RECT 63.880000 43.100000 64.080000 43.300000 ;
        RECT 63.880000 43.530000 64.080000 43.730000 ;
        RECT 63.880000 43.960000 64.080000 44.160000 ;
        RECT 64.285000 39.660000 64.485000 39.860000 ;
        RECT 64.285000 40.090000 64.485000 40.290000 ;
        RECT 64.285000 40.520000 64.485000 40.720000 ;
        RECT 64.285000 40.950000 64.485000 41.150000 ;
        RECT 64.285000 41.380000 64.485000 41.580000 ;
        RECT 64.285000 41.810000 64.485000 42.010000 ;
        RECT 64.285000 42.240000 64.485000 42.440000 ;
        RECT 64.285000 42.670000 64.485000 42.870000 ;
        RECT 64.285000 43.100000 64.485000 43.300000 ;
        RECT 64.285000 43.530000 64.485000 43.730000 ;
        RECT 64.285000 43.960000 64.485000 44.160000 ;
        RECT 64.690000 39.660000 64.890000 39.860000 ;
        RECT 64.690000 40.090000 64.890000 40.290000 ;
        RECT 64.690000 40.520000 64.890000 40.720000 ;
        RECT 64.690000 40.950000 64.890000 41.150000 ;
        RECT 64.690000 41.380000 64.890000 41.580000 ;
        RECT 64.690000 41.810000 64.890000 42.010000 ;
        RECT 64.690000 42.240000 64.890000 42.440000 ;
        RECT 64.690000 42.670000 64.890000 42.870000 ;
        RECT 64.690000 43.100000 64.890000 43.300000 ;
        RECT 64.690000 43.530000 64.890000 43.730000 ;
        RECT 64.690000 43.960000 64.890000 44.160000 ;
        RECT 65.095000 39.660000 65.295000 39.860000 ;
        RECT 65.095000 40.090000 65.295000 40.290000 ;
        RECT 65.095000 40.520000 65.295000 40.720000 ;
        RECT 65.095000 40.950000 65.295000 41.150000 ;
        RECT 65.095000 41.380000 65.295000 41.580000 ;
        RECT 65.095000 41.810000 65.295000 42.010000 ;
        RECT 65.095000 42.240000 65.295000 42.440000 ;
        RECT 65.095000 42.670000 65.295000 42.870000 ;
        RECT 65.095000 43.100000 65.295000 43.300000 ;
        RECT 65.095000 43.530000 65.295000 43.730000 ;
        RECT 65.095000 43.960000 65.295000 44.160000 ;
        RECT 65.500000 39.660000 65.700000 39.860000 ;
        RECT 65.500000 40.090000 65.700000 40.290000 ;
        RECT 65.500000 40.520000 65.700000 40.720000 ;
        RECT 65.500000 40.950000 65.700000 41.150000 ;
        RECT 65.500000 41.380000 65.700000 41.580000 ;
        RECT 65.500000 41.810000 65.700000 42.010000 ;
        RECT 65.500000 42.240000 65.700000 42.440000 ;
        RECT 65.500000 42.670000 65.700000 42.870000 ;
        RECT 65.500000 43.100000 65.700000 43.300000 ;
        RECT 65.500000 43.530000 65.700000 43.730000 ;
        RECT 65.500000 43.960000 65.700000 44.160000 ;
        RECT 65.905000 39.660000 66.105000 39.860000 ;
        RECT 65.905000 40.090000 66.105000 40.290000 ;
        RECT 65.905000 40.520000 66.105000 40.720000 ;
        RECT 65.905000 40.950000 66.105000 41.150000 ;
        RECT 65.905000 41.380000 66.105000 41.580000 ;
        RECT 65.905000 41.810000 66.105000 42.010000 ;
        RECT 65.905000 42.240000 66.105000 42.440000 ;
        RECT 65.905000 42.670000 66.105000 42.870000 ;
        RECT 65.905000 43.100000 66.105000 43.300000 ;
        RECT 65.905000 43.530000 66.105000 43.730000 ;
        RECT 65.905000 43.960000 66.105000 44.160000 ;
        RECT 66.310000 39.660000 66.510000 39.860000 ;
        RECT 66.310000 40.090000 66.510000 40.290000 ;
        RECT 66.310000 40.520000 66.510000 40.720000 ;
        RECT 66.310000 40.950000 66.510000 41.150000 ;
        RECT 66.310000 41.380000 66.510000 41.580000 ;
        RECT 66.310000 41.810000 66.510000 42.010000 ;
        RECT 66.310000 42.240000 66.510000 42.440000 ;
        RECT 66.310000 42.670000 66.510000 42.870000 ;
        RECT 66.310000 43.100000 66.510000 43.300000 ;
        RECT 66.310000 43.530000 66.510000 43.730000 ;
        RECT 66.310000 43.960000 66.510000 44.160000 ;
        RECT 66.715000 39.660000 66.915000 39.860000 ;
        RECT 66.715000 40.090000 66.915000 40.290000 ;
        RECT 66.715000 40.520000 66.915000 40.720000 ;
        RECT 66.715000 40.950000 66.915000 41.150000 ;
        RECT 66.715000 41.380000 66.915000 41.580000 ;
        RECT 66.715000 41.810000 66.915000 42.010000 ;
        RECT 66.715000 42.240000 66.915000 42.440000 ;
        RECT 66.715000 42.670000 66.915000 42.870000 ;
        RECT 66.715000 43.100000 66.915000 43.300000 ;
        RECT 66.715000 43.530000 66.915000 43.730000 ;
        RECT 66.715000 43.960000 66.915000 44.160000 ;
        RECT 67.120000 39.660000 67.320000 39.860000 ;
        RECT 67.120000 40.090000 67.320000 40.290000 ;
        RECT 67.120000 40.520000 67.320000 40.720000 ;
        RECT 67.120000 40.950000 67.320000 41.150000 ;
        RECT 67.120000 41.380000 67.320000 41.580000 ;
        RECT 67.120000 41.810000 67.320000 42.010000 ;
        RECT 67.120000 42.240000 67.320000 42.440000 ;
        RECT 67.120000 42.670000 67.320000 42.870000 ;
        RECT 67.120000 43.100000 67.320000 43.300000 ;
        RECT 67.120000 43.530000 67.320000 43.730000 ;
        RECT 67.120000 43.960000 67.320000 44.160000 ;
        RECT 67.525000 39.660000 67.725000 39.860000 ;
        RECT 67.525000 40.090000 67.725000 40.290000 ;
        RECT 67.525000 40.520000 67.725000 40.720000 ;
        RECT 67.525000 40.950000 67.725000 41.150000 ;
        RECT 67.525000 41.380000 67.725000 41.580000 ;
        RECT 67.525000 41.810000 67.725000 42.010000 ;
        RECT 67.525000 42.240000 67.725000 42.440000 ;
        RECT 67.525000 42.670000 67.725000 42.870000 ;
        RECT 67.525000 43.100000 67.725000 43.300000 ;
        RECT 67.525000 43.530000 67.725000 43.730000 ;
        RECT 67.525000 43.960000 67.725000 44.160000 ;
        RECT 67.930000 39.660000 68.130000 39.860000 ;
        RECT 67.930000 40.090000 68.130000 40.290000 ;
        RECT 67.930000 40.520000 68.130000 40.720000 ;
        RECT 67.930000 40.950000 68.130000 41.150000 ;
        RECT 67.930000 41.380000 68.130000 41.580000 ;
        RECT 67.930000 41.810000 68.130000 42.010000 ;
        RECT 67.930000 42.240000 68.130000 42.440000 ;
        RECT 67.930000 42.670000 68.130000 42.870000 ;
        RECT 67.930000 43.100000 68.130000 43.300000 ;
        RECT 67.930000 43.530000 68.130000 43.730000 ;
        RECT 67.930000 43.960000 68.130000 44.160000 ;
        RECT 68.335000 39.660000 68.535000 39.860000 ;
        RECT 68.335000 40.090000 68.535000 40.290000 ;
        RECT 68.335000 40.520000 68.535000 40.720000 ;
        RECT 68.335000 40.950000 68.535000 41.150000 ;
        RECT 68.335000 41.380000 68.535000 41.580000 ;
        RECT 68.335000 41.810000 68.535000 42.010000 ;
        RECT 68.335000 42.240000 68.535000 42.440000 ;
        RECT 68.335000 42.670000 68.535000 42.870000 ;
        RECT 68.335000 43.100000 68.535000 43.300000 ;
        RECT 68.335000 43.530000 68.535000 43.730000 ;
        RECT 68.335000 43.960000 68.535000 44.160000 ;
        RECT 68.740000 39.660000 68.940000 39.860000 ;
        RECT 68.740000 40.090000 68.940000 40.290000 ;
        RECT 68.740000 40.520000 68.940000 40.720000 ;
        RECT 68.740000 40.950000 68.940000 41.150000 ;
        RECT 68.740000 41.380000 68.940000 41.580000 ;
        RECT 68.740000 41.810000 68.940000 42.010000 ;
        RECT 68.740000 42.240000 68.940000 42.440000 ;
        RECT 68.740000 42.670000 68.940000 42.870000 ;
        RECT 68.740000 43.100000 68.940000 43.300000 ;
        RECT 68.740000 43.530000 68.940000 43.730000 ;
        RECT 68.740000 43.960000 68.940000 44.160000 ;
        RECT 69.145000 39.660000 69.345000 39.860000 ;
        RECT 69.145000 40.090000 69.345000 40.290000 ;
        RECT 69.145000 40.520000 69.345000 40.720000 ;
        RECT 69.145000 40.950000 69.345000 41.150000 ;
        RECT 69.145000 41.380000 69.345000 41.580000 ;
        RECT 69.145000 41.810000 69.345000 42.010000 ;
        RECT 69.145000 42.240000 69.345000 42.440000 ;
        RECT 69.145000 42.670000 69.345000 42.870000 ;
        RECT 69.145000 43.100000 69.345000 43.300000 ;
        RECT 69.145000 43.530000 69.345000 43.730000 ;
        RECT 69.145000 43.960000 69.345000 44.160000 ;
        RECT 69.550000 39.660000 69.750000 39.860000 ;
        RECT 69.550000 40.090000 69.750000 40.290000 ;
        RECT 69.550000 40.520000 69.750000 40.720000 ;
        RECT 69.550000 40.950000 69.750000 41.150000 ;
        RECT 69.550000 41.380000 69.750000 41.580000 ;
        RECT 69.550000 41.810000 69.750000 42.010000 ;
        RECT 69.550000 42.240000 69.750000 42.440000 ;
        RECT 69.550000 42.670000 69.750000 42.870000 ;
        RECT 69.550000 43.100000 69.750000 43.300000 ;
        RECT 69.550000 43.530000 69.750000 43.730000 ;
        RECT 69.550000 43.960000 69.750000 44.160000 ;
        RECT 69.955000 39.660000 70.155000 39.860000 ;
        RECT 69.955000 40.090000 70.155000 40.290000 ;
        RECT 69.955000 40.520000 70.155000 40.720000 ;
        RECT 69.955000 40.950000 70.155000 41.150000 ;
        RECT 69.955000 41.380000 70.155000 41.580000 ;
        RECT 69.955000 41.810000 70.155000 42.010000 ;
        RECT 69.955000 42.240000 70.155000 42.440000 ;
        RECT 69.955000 42.670000 70.155000 42.870000 ;
        RECT 69.955000 43.100000 70.155000 43.300000 ;
        RECT 69.955000 43.530000 70.155000 43.730000 ;
        RECT 69.955000 43.960000 70.155000 44.160000 ;
        RECT 70.360000 39.660000 70.560000 39.860000 ;
        RECT 70.360000 40.090000 70.560000 40.290000 ;
        RECT 70.360000 40.520000 70.560000 40.720000 ;
        RECT 70.360000 40.950000 70.560000 41.150000 ;
        RECT 70.360000 41.380000 70.560000 41.580000 ;
        RECT 70.360000 41.810000 70.560000 42.010000 ;
        RECT 70.360000 42.240000 70.560000 42.440000 ;
        RECT 70.360000 42.670000 70.560000 42.870000 ;
        RECT 70.360000 43.100000 70.560000 43.300000 ;
        RECT 70.360000 43.530000 70.560000 43.730000 ;
        RECT 70.360000 43.960000 70.560000 44.160000 ;
        RECT 70.765000 39.660000 70.965000 39.860000 ;
        RECT 70.765000 40.090000 70.965000 40.290000 ;
        RECT 70.765000 40.520000 70.965000 40.720000 ;
        RECT 70.765000 40.950000 70.965000 41.150000 ;
        RECT 70.765000 41.380000 70.965000 41.580000 ;
        RECT 70.765000 41.810000 70.965000 42.010000 ;
        RECT 70.765000 42.240000 70.965000 42.440000 ;
        RECT 70.765000 42.670000 70.965000 42.870000 ;
        RECT 70.765000 43.100000 70.965000 43.300000 ;
        RECT 70.765000 43.530000 70.965000 43.730000 ;
        RECT 70.765000 43.960000 70.965000 44.160000 ;
        RECT 71.170000 39.660000 71.370000 39.860000 ;
        RECT 71.170000 40.090000 71.370000 40.290000 ;
        RECT 71.170000 40.520000 71.370000 40.720000 ;
        RECT 71.170000 40.950000 71.370000 41.150000 ;
        RECT 71.170000 41.380000 71.370000 41.580000 ;
        RECT 71.170000 41.810000 71.370000 42.010000 ;
        RECT 71.170000 42.240000 71.370000 42.440000 ;
        RECT 71.170000 42.670000 71.370000 42.870000 ;
        RECT 71.170000 43.100000 71.370000 43.300000 ;
        RECT 71.170000 43.530000 71.370000 43.730000 ;
        RECT 71.170000 43.960000 71.370000 44.160000 ;
        RECT 71.575000 39.660000 71.775000 39.860000 ;
        RECT 71.575000 40.090000 71.775000 40.290000 ;
        RECT 71.575000 40.520000 71.775000 40.720000 ;
        RECT 71.575000 40.950000 71.775000 41.150000 ;
        RECT 71.575000 41.380000 71.775000 41.580000 ;
        RECT 71.575000 41.810000 71.775000 42.010000 ;
        RECT 71.575000 42.240000 71.775000 42.440000 ;
        RECT 71.575000 42.670000 71.775000 42.870000 ;
        RECT 71.575000 43.100000 71.775000 43.300000 ;
        RECT 71.575000 43.530000 71.775000 43.730000 ;
        RECT 71.575000 43.960000 71.775000 44.160000 ;
        RECT 71.980000 39.660000 72.180000 39.860000 ;
        RECT 71.980000 40.090000 72.180000 40.290000 ;
        RECT 71.980000 40.520000 72.180000 40.720000 ;
        RECT 71.980000 40.950000 72.180000 41.150000 ;
        RECT 71.980000 41.380000 72.180000 41.580000 ;
        RECT 71.980000 41.810000 72.180000 42.010000 ;
        RECT 71.980000 42.240000 72.180000 42.440000 ;
        RECT 71.980000 42.670000 72.180000 42.870000 ;
        RECT 71.980000 43.100000 72.180000 43.300000 ;
        RECT 71.980000 43.530000 72.180000 43.730000 ;
        RECT 71.980000 43.960000 72.180000 44.160000 ;
        RECT 72.385000 39.660000 72.585000 39.860000 ;
        RECT 72.385000 40.090000 72.585000 40.290000 ;
        RECT 72.385000 40.520000 72.585000 40.720000 ;
        RECT 72.385000 40.950000 72.585000 41.150000 ;
        RECT 72.385000 41.380000 72.585000 41.580000 ;
        RECT 72.385000 41.810000 72.585000 42.010000 ;
        RECT 72.385000 42.240000 72.585000 42.440000 ;
        RECT 72.385000 42.670000 72.585000 42.870000 ;
        RECT 72.385000 43.100000 72.585000 43.300000 ;
        RECT 72.385000 43.530000 72.585000 43.730000 ;
        RECT 72.385000 43.960000 72.585000 44.160000 ;
        RECT 72.790000 39.660000 72.990000 39.860000 ;
        RECT 72.790000 40.090000 72.990000 40.290000 ;
        RECT 72.790000 40.520000 72.990000 40.720000 ;
        RECT 72.790000 40.950000 72.990000 41.150000 ;
        RECT 72.790000 41.380000 72.990000 41.580000 ;
        RECT 72.790000 41.810000 72.990000 42.010000 ;
        RECT 72.790000 42.240000 72.990000 42.440000 ;
        RECT 72.790000 42.670000 72.990000 42.870000 ;
        RECT 72.790000 43.100000 72.990000 43.300000 ;
        RECT 72.790000 43.530000 72.990000 43.730000 ;
        RECT 72.790000 43.960000 72.990000 44.160000 ;
        RECT 73.195000 39.660000 73.395000 39.860000 ;
        RECT 73.195000 40.090000 73.395000 40.290000 ;
        RECT 73.195000 40.520000 73.395000 40.720000 ;
        RECT 73.195000 40.950000 73.395000 41.150000 ;
        RECT 73.195000 41.380000 73.395000 41.580000 ;
        RECT 73.195000 41.810000 73.395000 42.010000 ;
        RECT 73.195000 42.240000 73.395000 42.440000 ;
        RECT 73.195000 42.670000 73.395000 42.870000 ;
        RECT 73.195000 43.100000 73.395000 43.300000 ;
        RECT 73.195000 43.530000 73.395000 43.730000 ;
        RECT 73.195000 43.960000 73.395000 44.160000 ;
        RECT 73.600000 39.660000 73.800000 39.860000 ;
        RECT 73.600000 40.090000 73.800000 40.290000 ;
        RECT 73.600000 40.520000 73.800000 40.720000 ;
        RECT 73.600000 40.950000 73.800000 41.150000 ;
        RECT 73.600000 41.380000 73.800000 41.580000 ;
        RECT 73.600000 41.810000 73.800000 42.010000 ;
        RECT 73.600000 42.240000 73.800000 42.440000 ;
        RECT 73.600000 42.670000 73.800000 42.870000 ;
        RECT 73.600000 43.100000 73.800000 43.300000 ;
        RECT 73.600000 43.530000 73.800000 43.730000 ;
        RECT 73.600000 43.960000 73.800000 44.160000 ;
        RECT 74.005000 39.660000 74.205000 39.860000 ;
        RECT 74.005000 40.090000 74.205000 40.290000 ;
        RECT 74.005000 40.520000 74.205000 40.720000 ;
        RECT 74.005000 40.950000 74.205000 41.150000 ;
        RECT 74.005000 41.380000 74.205000 41.580000 ;
        RECT 74.005000 41.810000 74.205000 42.010000 ;
        RECT 74.005000 42.240000 74.205000 42.440000 ;
        RECT 74.005000 42.670000 74.205000 42.870000 ;
        RECT 74.005000 43.100000 74.205000 43.300000 ;
        RECT 74.005000 43.530000 74.205000 43.730000 ;
        RECT 74.005000 43.960000 74.205000 44.160000 ;
        RECT 74.410000 39.660000 74.610000 39.860000 ;
        RECT 74.410000 40.090000 74.610000 40.290000 ;
        RECT 74.410000 40.520000 74.610000 40.720000 ;
        RECT 74.410000 40.950000 74.610000 41.150000 ;
        RECT 74.410000 41.380000 74.610000 41.580000 ;
        RECT 74.410000 41.810000 74.610000 42.010000 ;
        RECT 74.410000 42.240000 74.610000 42.440000 ;
        RECT 74.410000 42.670000 74.610000 42.870000 ;
        RECT 74.410000 43.100000 74.610000 43.300000 ;
        RECT 74.410000 43.530000 74.610000 43.730000 ;
        RECT 74.410000 43.960000 74.610000 44.160000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 23.835000 1.270000 28.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 23.835000 75.000000 28.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 23.935000 1.270000 28.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 23.935000 75.000000 28.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 56.235000 1.270000 60.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 56.235000 75.000000 60.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 56.335000 1.270000 60.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 56.335000 75.000000 60.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 29.885000 1.270000 33.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 29.885000 75.000000 33.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 29.985000 1.270000 33.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 29.985000 75.000000 33.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met1 ;
      RECT 0.000000 0.000000 75.000000 198.000000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 75.000000 198.000000 ;
    LAYER met3 ;
      RECT  0.000000  0.000000 75.000000  39.190000 ;
      RECT  0.000000 44.630000 75.000000 198.000000 ;
      RECT 24.900000 39.190000 50.355000  44.630000 ;
    LAYER met4 ;
      RECT  0.000000   5.885000  1.670000   6.485000 ;
      RECT  0.000000  11.935000  1.365000  12.535000 ;
      RECT  0.000000  16.785000  1.365000  17.385000 ;
      RECT  0.000000  22.835000  1.670000  23.435000 ;
      RECT  0.000000  28.885000  1.670000  29.485000 ;
      RECT  0.000000  33.735000  1.670000  34.335000 ;
      RECT  0.000000  38.585000  1.670000  39.185000 ;
      RECT  0.000000  44.635000  1.670000  45.335000 ;
      RECT  0.000000  55.135000  1.670000  55.835000 ;
      RECT  0.000000  61.085000  1.670000  61.685000 ;
      RECT  0.000000  66.935000  1.670000  67.635000 ;
      RECT  0.000000  93.400000 75.000000 173.385000 ;
      RECT  1.365000  11.935000 73.635000  17.385000 ;
      RECT  1.670000   0.000000 73.330000  11.935000 ;
      RECT  1.670000  17.385000 73.330000  39.185000 ;
      RECT  1.670000  44.635000 73.330000  93.400000 ;
      RECT  1.670000 173.385000 73.330000 198.000000 ;
      RECT 24.875000  39.185000 50.380000  44.635000 ;
      RECT 73.330000   5.885000 75.000000   6.485000 ;
      RECT 73.330000  22.835000 75.000000  23.435000 ;
      RECT 73.330000  28.885000 75.000000  29.485000 ;
      RECT 73.330000  33.735000 75.000000  34.335000 ;
      RECT 73.330000  38.585000 75.000000  39.185000 ;
      RECT 73.330000  44.635000 75.000000  45.335000 ;
      RECT 73.330000  55.135000 75.000000  55.835000 ;
      RECT 73.330000  61.085000 75.000000  61.685000 ;
      RECT 73.330000  66.935000 75.000000  67.635000 ;
      RECT 73.635000  11.935000 75.000000  12.535000 ;
      RECT 73.635000  16.785000 75.000000  17.385000 ;
    LAYER met5 ;
      RECT 0.000000  93.785000 75.000000 172.985000 ;
      RECT 1.765000  12.235000 73.235000  17.085000 ;
      RECT 2.070000   0.000000 72.930000  12.235000 ;
      RECT 2.070000  17.085000 72.930000  93.785000 ;
      RECT 2.070000 172.985000 72.930000 198.000000 ;
  END
END sky130_fd_io__overlay_vssd_lvc
END LIBRARY
