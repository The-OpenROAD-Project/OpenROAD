VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  LIBRARY LEF58_CELLEDGESPACINGTABLE STRING
    "CELLEDGESPACINGTABLE
      EDGETYPE VERTICAL_EDGE_1 VERTICAL_EDGE_1 0.1
      EDGETYPE VERTICAL_EDGE_2 VERTICAL_EDGE_2 0.5 ; " ;

END PROPERTYDEFINITIONS