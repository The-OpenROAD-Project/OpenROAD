VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO array_tile
  FOREIGN array_tile 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 300 BY 300 ;
  CLASS BLOCK ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
      RECT 0.000 299.86 0.14 300.00 ;
    END
  END clk
  PIN e_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
      RECT 299.93 100.00 300.00 100.07 ;
    END
  END e_in
  PIN e_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
      RECT 299.93 100.14 300.00 100.21 ;
    END
  END e_out
  PIN w_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.14 0.070 100.21 ;
    END
  END w_in
  PIN w_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.00 0.070 100.07 ;
    END
  END w_out
  OBS
    LAYER metal1 ;
    RECT 0 0 300 300 ;
    LAYER metal2 ;
    RECT 0 0 300 300 ;
    LAYER metal3 ;
    RECT 0 0 300 300 ;
    LAYER metal4 ;
    RECT 0 0 300 300 ;
    LAYER metal5 ;
    RECT 0 0 300 300 ;
  END
END array_tile

END LIBRARY
