VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO cus_tg_mux41_buf
  CLASS CORE ;
  FOREIGN cus_tg_mux41_buf ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN S0
    ANTENNAGATEAREA 0.216000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.980 1.310 2.300 1.570 ;
        RECT 2.035 0.800 2.245 1.310 ;
        RECT 1.995 0.480 2.255 0.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.145 1.550 0.375 1.700 ;
        RECT 1.980 1.550 2.300 1.570 ;
        RECT 0.145 1.410 2.300 1.550 ;
        RECT 1.980 1.310 2.300 1.410 ;
      LAYER via ;
        RECT 2.010 1.310 2.270 1.570 ;
    END
  END S0
  PIN S1N
    ANTENNAGATEAREA 0.108000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 4.720 1.875 5.070 1.925 ;
        RECT 3.925 1.735 5.070 1.875 ;
        RECT 3.925 1.360 4.095 1.735 ;
        RECT 4.720 1.675 5.070 1.735 ;
        RECT 3.865 1.130 4.155 1.360 ;
    END
  END S1N
  PIN S1
    ANTENNAGATEAREA 0.108000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 4.720 1.195 5.075 1.465 ;
    END
  END S1
  PIN S0N
    ANTENNAGATEAREA 0.216000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 3.155 1.480 3.445 1.570 ;
        RECT 2.905 1.340 3.445 1.480 ;
        RECT 0.145 1.170 0.375 1.200 ;
        RECT 2.905 1.170 3.045 1.340 ;
        RECT 0.145 1.030 3.045 1.170 ;
        RECT 0.145 0.910 0.375 1.030 ;
        RECT 1.635 0.940 1.925 1.030 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.695 0.890 1.865 1.220 ;
      LAYER mcon ;
        RECT 1.695 0.970 1.865 1.140 ;
    END
  END S0N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.635 2.910 ;
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.420 -0.085 0.590 0.085 ;
    END
  END VNB
  PIN A2
    ANTENNADIFFAREA 0.187200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.035 0.255 2.205 2.465 ;
    END
  END A2
  PIN A1
    ANTENNADIFFAREA 0.190800 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355 0.255 1.525 2.465 ;
    END
  END A1
  PIN X
    ANTENNADIFFAREA 0.383600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.060 1.765 6.265 2.465 ;
        RECT 6.075 0.255 6.265 1.765 ;
    END
  END X
  PIN A3
    ANTENNADIFFAREA 0.190800 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.875 0.255 3.045 2.465 ;
    END
  END A3
  PIN A0
    ANTENNADIFFAREA 0.187200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.255 0.685 2.465 ;
    END
  END A0
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.175 1.390 0.345 1.720 ;
        RECT 0.175 0.890 0.345 1.220 ;
        RECT 0.935 0.255 1.105 2.465 ;
        RECT 2.455 0.255 2.625 2.465 ;
        RECT 3.215 1.290 3.385 1.620 ;
        RECT 3.215 0.790 3.385 1.120 ;
        RECT 3.585 0.255 3.755 2.465 ;
        RECT 4.005 2.110 4.175 2.465 ;
        RECT 3.925 1.030 4.095 1.360 ;
        RECT 3.995 0.690 4.175 0.860 ;
        RECT 4.005 0.255 4.175 0.690 ;
        RECT 4.425 0.255 4.595 2.465 ;
        RECT 5.165 2.135 5.435 2.465 ;
        RECT 4.765 1.725 5.095 1.895 ;
        RECT 4.765 1.245 5.095 1.415 ;
        RECT 5.265 1.410 5.435 2.135 ;
        RECT 5.635 1.775 5.860 2.635 ;
        RECT 5.735 1.410 5.905 1.490 ;
        RECT 5.265 1.240 5.905 1.410 ;
        RECT 4.825 0.685 4.995 1.015 ;
        RECT 5.265 0.605 5.435 1.240 ;
        RECT 5.735 1.160 5.905 1.240 ;
        RECT 5.165 0.255 5.435 0.605 ;
        RECT 5.655 0.085 5.905 0.945 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 0.935 1.720 1.105 1.890 ;
        RECT 0.175 1.470 0.345 1.640 ;
        RECT 0.175 0.970 0.345 1.140 ;
        RECT 3.585 1.770 3.755 1.940 ;
        RECT 3.215 1.370 3.385 1.540 ;
        RECT 3.215 0.870 3.385 1.040 ;
        RECT 2.455 0.410 2.625 0.580 ;
        RECT 3.925 1.160 4.095 1.330 ;
        RECT 4.825 1.725 4.995 1.895 ;
        RECT 4.825 1.245 4.995 1.415 ;
        RECT 4.825 0.765 4.995 0.935 ;
        RECT 4.425 0.410 4.595 0.580 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
      LAYER met1 ;
        RECT 3.940 2.020 4.260 2.340 ;
        RECT 0.875 1.850 1.165 1.920 ;
        RECT 3.555 1.850 3.785 2.000 ;
        RECT 0.875 1.710 3.785 1.850 ;
        RECT 0.875 1.690 1.165 1.710 ;
        RECT 3.185 0.890 3.415 1.100 ;
        RECT 2.065 0.810 3.415 0.890 ;
        RECT 3.910 0.960 4.230 0.990 ;
        RECT 4.765 0.960 5.030 0.995 ;
        RECT 2.065 0.800 3.385 0.810 ;
        RECT 1.995 0.750 3.385 0.800 ;
        RECT 3.910 0.790 5.030 0.960 ;
        RECT 1.995 0.480 2.255 0.750 ;
        RECT 3.910 0.660 4.230 0.790 ;
        RECT 4.795 0.705 5.030 0.790 ;
        RECT 2.395 0.520 2.685 0.610 ;
        RECT 4.365 0.520 4.655 0.610 ;
        RECT 2.395 0.380 4.655 0.520 ;
      LAYER via ;
        RECT 3.970 2.055 4.230 2.315 ;
        RECT 1.995 0.510 2.255 0.770 ;
        RECT 3.940 0.725 4.200 0.985 ;
      LAYER met2 ;
        RECT 3.920 2.050 4.260 2.340 ;
        RECT 4.005 0.990 4.155 2.050 ;
        RECT 3.910 0.720 4.230 0.990 ;
  END
END cus_tg_mux41_buf
MACRO BlockRAM_1KB
  CLASS BLOCK ;
  SIZE 530.3800 BY 470.9000 ;
  FOREIGN BlockRAM_1KB 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.5654 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 238.92 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.406 LAYER met4  ;
    ANTENNAMAXAREACAR 74.7629 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 377.112 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 9.4700 0.0000 9.8500 0.7200 ;
    END
  END clk
  PIN rd_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.731 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.547 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 11.0753 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 55.2055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 128.692 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 686.824 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.8952 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 31.592 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 97.5600 0.7200 97.9400 ;
    END
  END rd_addr[7]
  PIN rd_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1654 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.719 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 11.2965 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.3115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 130.024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 693.928 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.949 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.016 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 94.1600 0.7200 94.5400 ;
    END
  END rd_addr[6]
  PIN rd_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2498 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.141 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 10.2745 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.2015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 133.081 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 710.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.501 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.96 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 90.7600 0.7200 91.1400 ;
    END
  END rd_addr[5]
  PIN rd_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7968 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.876 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.8521 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.0895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 37.426 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 200.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.193 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.984 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 87.7000 0.7200 88.0800 ;
    END
  END rd_addr[4]
  PIN rd_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8472 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.128 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.8469 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.0635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 45.368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 242.584 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 84.3000 0.7200 84.6800 ;
    END
  END rd_addr[3]
  PIN rd_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.5966 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 87.801 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6145 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.7568 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 85.128 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 81.2400 0.7200 81.6200 ;
    END
  END rd_addr[2]
  PIN rd_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3142 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.463 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2645 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.196 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.4538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 104.224 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 77.8400 0.7200 78.2200 ;
    END
  END rd_addr[1]
  PIN rd_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1854 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.819 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 28.9435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 144.546 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.217 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 49.466 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 264.44 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 74.7800 0.7200 75.1600 ;
    END
  END rd_addr[0]
  PIN rd_data[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.243 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.107 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.4288 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 237.424 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 291.0200 0.7200 291.4000 ;
    END
  END rd_data[31]
  PIN rd_data[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.998 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.0988 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.258 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 287.6200 0.7200 288.0000 ;
    END
  END rd_data[30]
  PIN rd_data[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.298 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 261.345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0736 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.25 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 284.2200 0.7200 284.6000 ;
    END
  END rd_data[29]
  PIN rd_data[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6508 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.146 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.0924 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.226 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 280.8200 0.7200 281.2000 ;
    END
  END rd_data[28]
  PIN rd_data[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.277 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.277 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.8684 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 134.106 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 277.4200 0.7200 277.8000 ;
    END
  END rd_data[27]
  PIN rd_data[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0638 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.211 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.8852 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 134.19 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 274.0200 0.7200 274.4000 ;
    END
  END rd_data[26]
  PIN rd_data[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.121 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.497 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 28.7108 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 143.318 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 270.6200 0.7200 271.0000 ;
    END
  END rd_data[25]
  PIN rd_data[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 43.6166 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 217.938 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1684 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.724 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 267.2200 0.7200 267.6000 ;
    END
  END rd_data[24]
  PIN rd_data[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8132 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.958 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 29.4864 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 147.196 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 263.8200 0.7200 264.2000 ;
    END
  END rd_data[23]
  PIN rd_data[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 43.8112 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 218.911 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4876 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.32 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 260.4200 0.7200 260.8000 ;
    END
  END rd_data[22]
  PIN rd_data[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3142 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.463 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.3612 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.57 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 257.0200 0.7200 257.4000 ;
    END
  END rd_data[21]
  PIN rd_data[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.705 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4475 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.6704 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.116 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 253.6200 0.7200 254.0000 ;
    END
  END rd_data[20]
  PIN rd_data[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 38.7222 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 193.466 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5496 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.63 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 250.2200 0.7200 250.6000 ;
    END
  END rd_data[19]
  PIN rd_data[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 37.5154 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 187.432 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1684 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.724 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 246.8200 0.7200 247.2000 ;
    END
  END rd_data[18]
  PIN rd_data[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.434 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 67.025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6924 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.344 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 243.4200 0.7200 243.8000 ;
    END
  END rd_data[17]
  PIN rd_data[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.1314 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 50.512 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4072 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.918 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 240.0200 0.7200 240.4000 ;
    END
  END rd_data[16]
  PIN rd_data[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 35.6901 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 178.28 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.539 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.6108 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 67.728 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 58.4600 0.7200 58.8400 ;
    END
  END rd_data[15]
  PIN rd_data[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1854 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.819 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6645 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.5908 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.088 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 108.503 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 579.152 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 55.0600 0.7200 55.4400 ;
    END
  END rd_data[14]
  PIN rd_data[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 58.9858 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 294.784 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.392 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 52.0000 0.7200 52.3800 ;
    END
  END rd_data[13]
  PIN rd_data[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8136 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.96 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 19.0679 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 95.1685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.1418 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.36 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.6968 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 233.52 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 48.6000 0.7200 48.9800 ;
    END
  END rd_data[12]
  PIN rd_data[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.354 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.7364 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.446 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 45.5400 0.7200 45.9200 ;
    END
  END rd_data[11]
  PIN rd_data[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4502 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.143 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 41.6961 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 208.31 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.194 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.5228 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 200.592 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 42.1400 0.7200 42.5200 ;
    END
  END rd_data[10]
  PIN rd_data[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.5318 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 52.514 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.3596 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.68 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 39.0800 0.7200 39.4600 ;
    END
  END rd_data[9]
  PIN rd_data[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.143 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.57 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.6228 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.878 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 35.6800 0.7200 36.0600 ;
    END
  END rd_data[8]
  PIN rd_data[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4006 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.858 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 12.5159 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 62.4085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.2448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 65.776 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 32.2800 0.7200 32.6600 ;
    END
  END rd_data[7]
  PIN rd_data[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4398 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.091 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 22.2613 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 111.136 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.974 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 78.9756 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 422.144 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 29.2200 0.7200 29.6000 ;
    END
  END rd_data[6]
  PIN rd_data[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2071 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 124.559 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 664.784 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 25.8200 0.7200 26.2000 ;
    END
  END rd_data[5]
  PIN rd_data[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6242 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.976 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 28.1119 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 140.388 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 23.3028 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 124.752 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 22.7600 0.7200 23.1400 ;
    END
  END rd_data[4]
  PIN rd_data[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.375 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.767 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1595 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 126.533 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 675.312 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 19.3600 0.7200 19.7400 ;
    END
  END rd_data[3]
  PIN rd_data[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.053 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.157 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0957 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.3075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.6998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 105.536 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 16.3000 0.7200 16.6800 ;
    END
  END rd_data[2]
  PIN rd_data[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8452 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.081 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.9544 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.654 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 12.9000 0.7200 13.2800 ;
    END
  END rd_data[1]
  PIN rd_data[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8514 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.112 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 33.2328 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 165.928 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 9.8400 0.7200 10.2200 ;
    END
  END rd_data[0]
  PIN wr_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.535 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.567 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 16.5437 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 82.5475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.3792 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.84 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 325.0200 0.7200 325.4000 ;
    END
  END wr_addr[7]
  PIN wr_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9424 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.604 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 16.4555 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 82.1065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.6922 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.176 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 321.6200 0.7200 322.0000 ;
    END
  END wr_addr[6]
  PIN wr_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5896 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.84 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 17.4957 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 87.3075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.6472 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.936 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 318.2200 0.7200 318.6000 ;
    END
  END wr_addr[5]
  PIN wr_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0194 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.989 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 17.9045 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 89.3515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.8042 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.44 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 314.8200 0.7200 315.2000 ;
    END
  END wr_addr[4]
  PIN wr_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7618 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.701 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 18.4813 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 92.2355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.0652 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.832 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 311.4200 0.7200 311.8000 ;
    END
  END wr_addr[3]
  PIN wr_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5686 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.735 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 18.5485 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 92.5715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.9412 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.504 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 308.0200 0.7200 308.4000 ;
    END
  END wr_addr[2]
  PIN wr_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1514 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.649 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 19.5395 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 97.4085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.4682 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.648 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 304.6200 0.7200 305.0000 ;
    END
  END wr_addr[1]
  PIN wr_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7958 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.871 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 41.5701 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 207.68 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.38 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 157.16 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.7932 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.048 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 301.2200 0.7200 301.6000 ;
    END
  END wr_addr[0]
  PIN wr_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1854 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.819 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 22.4443 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 111.815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 32.5174 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 175.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 19.8381 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 94.9206 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 379.4200 0.7200 379.8000 ;
    END
  END wr_data[31]
  PIN wr_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7958 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.871 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.8581 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.8835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 61.6966 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 332.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 20.9651 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 101.456 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 376.0200 0.7200 376.4000 ;
    END
  END wr_data[30]
  PIN wr_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5378 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.581 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 36.4379 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 181.311 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.7896 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.152 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 16.5413 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 73.6627 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 372.6200 0.7200 373.0000 ;
    END
  END wr_data[29]
  PIN wr_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2466 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.6277 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.9675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.8212 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.928 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 64.7762 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 326.206 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 369.2200 0.7200 369.6000 ;
    END
  END wr_data[28]
  PIN wr_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3754 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.769 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.3131 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.3945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.2712 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.328 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 97.7 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 500.488 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 365.8200 0.7200 366.2000 ;
    END
  END wr_data[27]
  PIN wr_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7006 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.395 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 32.6755 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 162.97 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.3268 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.88 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 98.4048 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 479.968 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 362.4200 0.7200 362.8000 ;
    END
  END wr_data[26]
  PIN wr_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9242 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.513 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 11.3283 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.2345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.5892 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 65.1425 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 322.181 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 359.0200 0.7200 359.4000 ;
    END
  END wr_data[25]
  PIN wr_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7282 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.533 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 24.6657 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 122.686 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 51.3658 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 274.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 21.3313 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 105.395 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 355.6200 0.7200 356.0000 ;
    END
  END wr_data[24]
  PIN wr_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3382 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.583 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 16.7571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 83.1425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.7948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 22.3032 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 103.187 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 352.2200 0.7200 352.6000 ;
    END
  END wr_data[23]
  PIN wr_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1482 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.633 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 9.6079 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.7505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 67.8556 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 365.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 29.819 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 146.286 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 348.8200 0.7200 349.2000 ;
    END
  END wr_data[22]
  PIN wr_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7184 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.484 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.7991 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.8245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 56.6158 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 302.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 18.1746 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 86.869 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 345.4200 0.7200 345.8000 ;
    END
  END wr_data[21]
  PIN wr_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0478 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.094 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 21.0596 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 104.944 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met2  ;
    ANTENNAMAXAREACAR 68.6338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 324.821 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 342.0200 0.7200 342.4000 ;
    END
  END wr_data[20]
  PIN wr_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3418 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.601 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.2447 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.9345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 52.426 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 280.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 23.9254 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 117.171 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 338.6200 0.7200 339.0000 ;
    END
  END wr_data[19]
  PIN wr_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0226 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 38.1569 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 190.614 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.3326 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 78.754 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 390.413 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 335.2200 0.7200 335.6000 ;
    END
  END wr_data[18]
  PIN wr_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 22.303 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 111.37 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met1  ;
    ANTENNAMAXAREACAR 45.2432 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 225.253 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7552 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.442 LAYER met2  ;
    ANTENNAGATEAREA 1.737 LAYER met2  ;
    ANTENNAMAXAREACAR 46.2537 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 230.113 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.318651 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 331.8200 0.7200 332.2000 ;
    END
  END wr_data[17]
  PIN wr_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1854 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.819 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.2996 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.83 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.494 LAYER met2  ;
    ANTENNAMAXAREACAR 17.9576 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 71.563 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 328.4200 0.7200 328.8000 ;
    END
  END wr_data[16]
  PIN wr_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.1594 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 155.652 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2337 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 14.271 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 55.0417 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.566667 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 149.2400 0.7200 149.6200 ;
    END
  END wr_data[15]
  PIN wr_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7282 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.533 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 19.232 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 95.816 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 81.4706 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 388.746 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 146.1800 0.7200 146.5600 ;
    END
  END wr_data[14]
  PIN wr_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 28.869 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 144.2 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.7304 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.426 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 15.9881 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 61.8016 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 142.7800 0.7200 143.1600 ;
    END
  END wr_data[13]
  PIN wr_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3142 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.463 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.252 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.916 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 24.7722 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 104.718 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 139.7200 0.7200 140.1000 ;
    END
  END wr_data[12]
  PIN wr_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.8114 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 128.912 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.7256 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.284 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 19.9373 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 81.0794 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 136.3200 0.7200 136.7000 ;
    END
  END wr_data[11]
  PIN wr_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3624 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.704 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 17.118 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 85.246 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 74.2944 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 352.329 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 133.2600 0.7200 133.6400 ;
    END
  END wr_data[10]
  PIN wr_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9826 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 15.4282 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 76.797 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 67.5889 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 318.802 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 129.8600 0.7200 130.2400 ;
    END
  END wr_data[9]
  PIN wr_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3554 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.669 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 14.6848 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.08 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 64.1278 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 301.496 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 126.8000 0.7200 127.1800 ;
    END
  END wr_data[8]
  PIN wr_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2806 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.295 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 12.7421 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 63.4305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.539 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.0776 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 48.56 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 102.545 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 534.679 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.636111 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 123.4000 0.7200 123.7800 ;
    END
  END wr_data[7]
  PIN wr_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 23.192 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 115.815 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1621 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.4446 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.184 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 90.7286 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 465.871 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 120.0000 0.7200 120.3800 ;
    END
  END wr_data[6]
  PIN wr_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1514 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.649 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.6035 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.8465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 53.7344 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 287.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.7496 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.56 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 73.9726 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 375.226 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.85635 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 116.9400 0.7200 117.3200 ;
    END
  END wr_data[5]
  PIN wr_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3142 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.463 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 11.8129 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 58.7755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 39.682 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 212.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.0014 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.04 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 52.8111 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 265.355 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 113.5400 0.7200 113.9200 ;
    END
  END wr_data[4]
  PIN wr_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6434 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.109 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.8655 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.0385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.5424 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.688 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 55.8738 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 274.573 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.7802 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.312 LAYER met4  ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 58.9698 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 291.685 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 110.4800 0.7200 110.8600 ;
    END
  END wr_data[3]
  PIN wr_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.746 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.622 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 10.1821 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.7395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 37.912 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 202.664 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.19902 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.2 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 101.091 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 519.442 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 107.0800 0.7200 107.4600 ;
    END
  END wr_data[2]
  PIN wr_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9728 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.756 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.0815 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.2365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.9464 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 69.664 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 109.004 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 565.885 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 104.0200 0.7200 104.4000 ;
    END
  END wr_data[1]
  PIN wr_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0834 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.309 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 9.0523 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.0905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 32.989 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 176.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.3666 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.768 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 66.8746 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 340.891 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 100.6200 0.7200 101.0000 ;
    END
  END wr_data[0]
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9994 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.889 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.72 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.912 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.611 LAYER met2  ;
    ANTENNAMAXAREACAR 7.06741 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 33.3716 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 61.5200 0.7200 61.9000 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4362 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.073 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.3692 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.384 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.242 LAYER met2  ;
    ANTENNAMAXAREACAR 41.3357 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 200.564 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 64.9200 0.7200 65.3000 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0708 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.246 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 54.8256 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 273.784 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met2  ;
    ANTENNAMAXAREACAR 56.0919 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 278.048 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 68.3200 0.7200 68.7000 ;
    END
  END C2
  PIN C3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2378 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.044 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 50.7788 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 253.54 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met2  ;
    ANTENNAMAXAREACAR 71.967 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 348.799 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 71.3800 0.7200 71.7600 ;
    END
  END C3
  PIN C4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.135 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 40.53 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5234 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.499 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 1.69495 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 6.99697 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 294.4200 0.7200 294.8000 ;
    END
  END C4
  PIN C5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.4924 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 62.1145 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.756 LAYER met1  ;
    ANTENNAMAXAREACAR 19.8176 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 86.0985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAMAXCUTCAR 0.144444 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.2451 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.5925 LAYER met2  ;
    ANTENNAGATEAREA 2.52 LAYER met2  ;
    ANTENNAMAXAREACAR 21.1053 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 92.286 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.219841 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.7188 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 148.304 LAYER met3  ;
    ANTENNAGATEAREA 8.064 LAYER met3  ;
    ANTENNAMAXAREACAR 24.5427 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 110.677 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.300469 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 297.8200 0.7200 298.2000 ;
    END
  END C5
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 528.7800 462.6800 530.3800 464.2800 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.0000 462.6800 1.6000 464.2800 ;
    END
    PORT
      LAYER met3 ;
        RECT 528.7800 5.4300 530.3800 7.0300 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.0000 5.4300 1.6000 7.0300 ;
    END
    PORT
      LAYER met4 ;
        RECT 523.2200 469.3000 524.8200 470.9000 ;
    END
    PORT
      LAYER met4 ;
        RECT 523.2200 0.0000 524.8200 1.6000 ;
    END
    PORT
      LAYER met4 ;
        RECT 5.5600 469.3000 7.1600 470.9000 ;
    END
    PORT
      LAYER met4 ;
        RECT 5.5600 0.0000 7.1600 1.6000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.0000 5.4300 530.3800 7.0300 ;
        RECT 0.0000 462.6800 530.3800 464.2800 ;
        RECT 5.5600 9.6200 7.1600 10.1000 ;
        RECT 5.5600 15.0600 7.1600 15.5400 ;
        RECT 5.5600 20.5000 7.1600 20.9800 ;
        RECT 5.5600 25.9400 7.1600 26.4200 ;
        RECT 5.5600 31.3800 7.1600 31.8600 ;
        RECT 5.5600 69.4600 7.1600 69.9400 ;
        RECT 5.5600 36.8200 7.1600 37.3000 ;
        RECT 5.5600 42.2600 7.1600 42.7400 ;
        RECT 5.5600 47.7000 7.1600 48.1800 ;
        RECT 5.5600 53.1400 7.1600 53.6200 ;
        RECT 5.5600 58.5800 7.1600 59.0600 ;
        RECT 5.5600 64.0200 7.1600 64.5000 ;
        RECT 5.5600 74.9000 7.1600 75.3800 ;
        RECT 5.5600 80.3400 7.1600 80.8200 ;
        RECT 5.5600 85.7800 7.1600 86.2600 ;
        RECT 5.5600 91.2200 7.1600 91.7000 ;
        RECT 5.5600 96.6600 7.1600 97.1400 ;
        RECT 5.5600 102.1000 7.1600 102.5800 ;
        RECT 5.5600 107.5400 7.1600 108.0200 ;
        RECT 5.5600 112.9800 7.1600 113.4600 ;
        RECT 5.5600 118.4200 7.1600 118.9000 ;
        RECT 5.5600 123.8600 7.1600 124.3400 ;
        RECT 5.5600 129.3000 7.1600 129.7800 ;
        RECT 5.5600 134.7400 7.1600 135.2200 ;
        RECT 5.5600 140.1800 7.1600 140.6600 ;
        RECT 5.5600 145.6200 7.1600 146.1000 ;
        RECT 5.5600 151.0600 7.1600 151.5400 ;
        RECT 5.5600 156.5000 7.1600 156.9800 ;
        RECT 5.5600 161.9400 7.1600 162.4200 ;
        RECT 5.5600 167.3800 7.1600 167.8600 ;
        RECT 5.5600 172.8200 7.1600 173.3000 ;
        RECT 5.5600 178.2600 7.1600 178.7400 ;
        RECT 5.5600 183.7000 7.1600 184.1800 ;
        RECT 5.5600 189.1400 7.1600 189.6200 ;
        RECT 5.5600 194.5800 7.1600 195.0600 ;
        RECT 5.5600 200.0200 7.1600 200.5000 ;
        RECT 5.5600 205.4600 7.1600 205.9400 ;
        RECT 5.5600 210.9000 7.1600 211.3800 ;
        RECT 5.5600 216.3400 7.1600 216.8200 ;
        RECT 5.5600 221.7800 7.1600 222.2600 ;
        RECT 5.5600 227.2200 7.1600 227.7000 ;
        RECT 5.5600 232.6600 7.1600 233.1400 ;
        RECT 523.2200 9.6200 524.8200 10.1000 ;
        RECT 523.2200 15.0600 524.8200 15.5400 ;
        RECT 523.2200 20.5000 524.8200 20.9800 ;
        RECT 523.2200 25.9400 524.8200 26.4200 ;
        RECT 523.2200 31.3800 524.8200 31.8600 ;
        RECT 523.2200 69.4600 524.8200 69.9400 ;
        RECT 523.2200 36.8200 524.8200 37.3000 ;
        RECT 523.2200 42.2600 524.8200 42.7400 ;
        RECT 523.2200 47.7000 524.8200 48.1800 ;
        RECT 523.2200 53.1400 524.8200 53.6200 ;
        RECT 523.2200 58.5800 524.8200 59.0600 ;
        RECT 523.2200 64.0200 524.8200 64.5000 ;
        RECT 523.2200 74.9000 524.8200 75.3800 ;
        RECT 523.2200 80.3400 524.8200 80.8200 ;
        RECT 523.2200 85.7800 524.8200 86.2600 ;
        RECT 523.2200 91.2200 524.8200 91.7000 ;
        RECT 523.2200 96.6600 524.8200 97.1400 ;
        RECT 523.2200 102.1000 524.8200 102.5800 ;
        RECT 523.2200 107.5400 524.8200 108.0200 ;
        RECT 523.2200 112.9800 524.8200 113.4600 ;
        RECT 523.2200 118.4200 524.8200 118.9000 ;
        RECT 523.2200 123.8600 524.8200 124.3400 ;
        RECT 523.2200 129.3000 524.8200 129.7800 ;
        RECT 523.2200 134.7400 524.8200 135.2200 ;
        RECT 523.2200 140.1800 524.8200 140.6600 ;
        RECT 523.2200 145.6200 524.8200 146.1000 ;
        RECT 523.2200 151.0600 524.8200 151.5400 ;
        RECT 523.2200 156.5000 524.8200 156.9800 ;
        RECT 523.2200 161.9400 524.8200 162.4200 ;
        RECT 523.2200 167.3800 524.8200 167.8600 ;
        RECT 523.2200 172.8200 524.8200 173.3000 ;
        RECT 523.2200 178.2600 524.8200 178.7400 ;
        RECT 523.2200 183.7000 524.8200 184.1800 ;
        RECT 523.2200 189.1400 524.8200 189.6200 ;
        RECT 523.2200 194.5800 524.8200 195.0600 ;
        RECT 523.2200 200.0200 524.8200 200.5000 ;
        RECT 523.2200 205.4600 524.8200 205.9400 ;
        RECT 523.2200 210.9000 524.8200 211.3800 ;
        RECT 523.2200 216.3400 524.8200 216.8200 ;
        RECT 523.2200 221.7800 524.8200 222.2600 ;
        RECT 523.2200 227.2200 524.8200 227.7000 ;
        RECT 523.2200 232.6600 524.8200 233.1400 ;
        RECT 5.5600 238.1000 7.1600 238.5800 ;
        RECT 5.5600 243.5400 7.1600 244.0200 ;
        RECT 5.5600 248.9800 7.1600 249.4600 ;
        RECT 5.5600 259.8600 7.1600 260.3400 ;
        RECT 5.5600 254.4200 7.1600 254.9000 ;
        RECT 5.5600 265.3000 7.1600 265.7800 ;
        RECT 5.5600 270.7400 7.1600 271.2200 ;
        RECT 5.5600 276.1800 7.1600 276.6600 ;
        RECT 5.5600 281.6200 7.1600 282.1000 ;
        RECT 5.5600 287.0600 7.1600 287.5400 ;
        RECT 5.5600 292.5000 7.1600 292.9800 ;
        RECT 5.5600 297.9400 7.1600 298.4200 ;
        RECT 5.5600 303.3800 7.1600 303.8600 ;
        RECT 5.5600 308.8200 7.1600 309.3000 ;
        RECT 5.5600 314.2600 7.1600 314.7400 ;
        RECT 5.5600 319.7000 7.1600 320.1800 ;
        RECT 5.5600 325.1400 7.1600 325.6200 ;
        RECT 5.5600 330.5800 7.1600 331.0600 ;
        RECT 5.5600 336.0200 7.1600 336.5000 ;
        RECT 5.5600 341.4600 7.1600 341.9400 ;
        RECT 5.5600 346.9000 7.1600 347.3800 ;
        RECT 5.5600 352.3400 7.1600 352.8200 ;
        RECT 5.5600 357.7800 7.1600 358.2600 ;
        RECT 5.5600 363.2200 7.1600 363.7000 ;
        RECT 5.5600 433.9400 7.1600 434.4200 ;
        RECT 5.5600 368.6600 7.1600 369.1400 ;
        RECT 5.5600 374.1000 7.1600 374.5800 ;
        RECT 5.5600 379.5400 7.1600 380.0200 ;
        RECT 5.5600 384.9800 7.1600 385.4600 ;
        RECT 5.5600 390.4200 7.1600 390.9000 ;
        RECT 5.5600 395.8600 7.1600 396.3400 ;
        RECT 5.5600 417.6200 7.1600 418.1000 ;
        RECT 5.5600 401.3000 7.1600 401.7800 ;
        RECT 5.5600 406.7400 7.1600 407.2200 ;
        RECT 5.5600 412.1800 7.1600 412.6600 ;
        RECT 5.5600 423.0600 7.1600 423.5400 ;
        RECT 5.5600 428.5000 7.1600 428.9800 ;
        RECT 30.2500 429.6100 31.6200 431.2100 ;
        RECT 5.5600 439.3800 7.1600 439.8600 ;
        RECT 5.5600 444.8200 7.1600 445.3000 ;
        RECT 5.5600 450.2600 7.1600 450.7400 ;
        RECT 5.5600 455.7000 7.1600 456.1800 ;
        RECT 523.2200 238.1000 524.8200 238.5800 ;
        RECT 523.2200 243.5400 524.8200 244.0200 ;
        RECT 523.2200 248.9800 524.8200 249.4600 ;
        RECT 523.2200 259.8600 524.8200 260.3400 ;
        RECT 523.2200 254.4200 524.8200 254.9000 ;
        RECT 523.2200 265.3000 524.8200 265.7800 ;
        RECT 523.2200 270.7400 524.8200 271.2200 ;
        RECT 523.2200 276.1800 524.8200 276.6600 ;
        RECT 523.2200 281.6200 524.8200 282.1000 ;
        RECT 523.2200 287.0600 524.8200 287.5400 ;
        RECT 523.2200 292.5000 524.8200 292.9800 ;
        RECT 523.2200 297.9400 524.8200 298.4200 ;
        RECT 523.2200 303.3800 524.8200 303.8600 ;
        RECT 523.2200 308.8200 524.8200 309.3000 ;
        RECT 523.2200 314.2600 524.8200 314.7400 ;
        RECT 523.2200 319.7000 524.8200 320.1800 ;
        RECT 523.2200 325.1400 524.8200 325.6200 ;
        RECT 523.2200 330.5800 524.8200 331.0600 ;
        RECT 523.2200 336.0200 524.8200 336.5000 ;
        RECT 523.2200 341.4600 524.8200 341.9400 ;
        RECT 523.2200 346.9000 524.8200 347.3800 ;
        RECT 523.2200 352.3400 524.8200 352.8200 ;
        RECT 523.2200 357.7800 524.8200 358.2600 ;
        RECT 523.2200 363.2200 524.8200 363.7000 ;
        RECT 523.2200 433.9400 524.8200 434.4200 ;
        RECT 523.2200 368.6600 524.8200 369.1400 ;
        RECT 523.2200 374.1000 524.8200 374.5800 ;
        RECT 523.2200 379.5400 524.8200 380.0200 ;
        RECT 523.2200 384.9800 524.8200 385.4600 ;
        RECT 523.2200 390.4200 524.8200 390.9000 ;
        RECT 523.2200 395.8600 524.8200 396.3400 ;
        RECT 523.2200 417.6200 524.8200 418.1000 ;
        RECT 523.2200 401.3000 524.8200 401.7800 ;
        RECT 523.2200 406.7400 524.8200 407.2200 ;
        RECT 523.2200 412.1800 524.8200 412.6600 ;
        RECT 523.2200 423.0600 524.8200 423.5400 ;
        RECT 523.2200 428.5000 524.8200 428.9800 ;
        RECT 523.2200 439.3800 524.8200 439.8600 ;
        RECT 523.2200 444.8200 524.8200 445.3000 ;
        RECT 523.2200 450.2600 524.8200 450.7400 ;
        RECT 523.2200 455.7000 524.8200 456.1800 ;
      LAYER met4 ;
        RECT 5.5600 0.0000 7.1600 470.9000 ;
        RECT 523.2200 0.0000 524.8200 470.9000 ;
        RECT 30.2250 429.6100 31.6450 431.2100 ;
    END
# end of P/G power stripe data as pin


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met3 ;
        RECT 29.8800 429.5400 500.1400 431.2800 ;
      LAYER met3 ;
        RECT 29.8800 43.3000 500.1400 45.0400 ;
      LAYER met4 ;
        RECT 29.8800 43.3000 31.6200 431.2800 ;
      LAYER met4 ;
        RECT 498.4000 43.3000 500.1400 431.2800 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 528.7800 465.2800 530.3800 466.8800 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.0000 465.2800 1.6000 466.8800 ;
    END
    PORT
      LAYER met3 ;
        RECT 528.7800 2.8300 530.3800 4.4300 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.0000 2.8300 1.6000 4.4300 ;
    END
    PORT
      LAYER met4 ;
        RECT 525.8200 469.3000 527.4200 470.9000 ;
    END
    PORT
      LAYER met4 ;
        RECT 525.8200 0.0000 527.4200 1.6000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.9600 469.3000 4.5600 470.9000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.9600 0.0000 4.5600 1.6000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.0000 2.8300 530.3800 4.4300 ;
        RECT 0.0000 465.2800 530.3800 466.8800 ;
        RECT 2.9600 235.3800 4.5600 235.8600 ;
        RECT 525.8200 235.3800 527.4200 235.8600 ;
        RECT 2.9600 12.3400 4.5600 12.8200 ;
        RECT 2.9600 17.7800 4.5600 18.2600 ;
        RECT 2.9600 23.2200 4.5600 23.7000 ;
        RECT 2.9600 28.6600 4.5600 29.1400 ;
        RECT 2.9600 34.1000 4.5600 34.5800 ;
        RECT 2.9600 39.5400 4.5600 40.0200 ;
        RECT 2.9600 44.9800 4.5600 45.4600 ;
        RECT 2.9600 50.4200 4.5600 50.9000 ;
        RECT 2.9600 61.3000 4.5600 61.7800 ;
        RECT 2.9600 55.8600 4.5600 56.3400 ;
        RECT 2.9600 66.7400 4.5600 67.2200 ;
        RECT 2.9600 77.6200 4.5600 78.1000 ;
        RECT 2.9600 72.1800 4.5600 72.6600 ;
        RECT 2.9600 83.0600 4.5600 83.5400 ;
        RECT 2.9600 93.9400 4.5600 94.4200 ;
        RECT 2.9600 88.5000 4.5600 88.9800 ;
        RECT 2.9600 99.3800 4.5600 99.8600 ;
        RECT 2.9600 110.2600 4.5600 110.7400 ;
        RECT 2.9600 104.8200 4.5600 105.3000 ;
        RECT 2.9600 115.7000 4.5600 116.1800 ;
        RECT 2.9600 126.5800 4.5600 127.0600 ;
        RECT 2.9600 121.1400 4.5600 121.6200 ;
        RECT 2.9600 132.0200 4.5600 132.5000 ;
        RECT 2.9600 142.9000 4.5600 143.3800 ;
        RECT 2.9600 137.4600 4.5600 137.9400 ;
        RECT 2.9600 148.3400 4.5600 148.8200 ;
        RECT 2.9600 159.2200 4.5600 159.7000 ;
        RECT 2.9600 153.7800 4.5600 154.2600 ;
        RECT 2.9600 164.6600 4.5600 165.1400 ;
        RECT 2.9600 175.5400 4.5600 176.0200 ;
        RECT 2.9600 170.1000 4.5600 170.5800 ;
        RECT 2.9600 180.9800 4.5600 181.4600 ;
        RECT 2.9600 191.8600 4.5600 192.3400 ;
        RECT 2.9600 186.4200 4.5600 186.9000 ;
        RECT 2.9600 197.3000 4.5600 197.7800 ;
        RECT 2.9600 208.1800 4.5600 208.6600 ;
        RECT 2.9600 202.7400 4.5600 203.2200 ;
        RECT 2.9600 213.6200 4.5600 214.1000 ;
        RECT 2.9600 224.5000 4.5600 224.9800 ;
        RECT 2.9600 219.0600 4.5600 219.5400 ;
        RECT 2.9600 229.9400 4.5600 230.4200 ;
        RECT 525.8200 12.3400 527.4200 12.8200 ;
        RECT 525.8200 17.7800 527.4200 18.2600 ;
        RECT 525.8200 23.2200 527.4200 23.7000 ;
        RECT 525.8200 28.6600 527.4200 29.1400 ;
        RECT 525.8200 34.1000 527.4200 34.5800 ;
        RECT 525.8200 39.5400 527.4200 40.0200 ;
        RECT 525.8200 44.9800 527.4200 45.4600 ;
        RECT 525.8200 50.4200 527.4200 50.9000 ;
        RECT 525.8200 61.3000 527.4200 61.7800 ;
        RECT 525.8200 55.8600 527.4200 56.3400 ;
        RECT 525.8200 66.7400 527.4200 67.2200 ;
        RECT 525.8200 77.6200 527.4200 78.1000 ;
        RECT 525.8200 72.1800 527.4200 72.6600 ;
        RECT 525.8200 83.0600 527.4200 83.5400 ;
        RECT 525.8200 93.9400 527.4200 94.4200 ;
        RECT 525.8200 88.5000 527.4200 88.9800 ;
        RECT 525.8200 99.3800 527.4200 99.8600 ;
        RECT 525.8200 110.2600 527.4200 110.7400 ;
        RECT 525.8200 104.8200 527.4200 105.3000 ;
        RECT 525.8200 115.7000 527.4200 116.1800 ;
        RECT 525.8200 126.5800 527.4200 127.0600 ;
        RECT 525.8200 121.1400 527.4200 121.6200 ;
        RECT 525.8200 132.0200 527.4200 132.5000 ;
        RECT 525.8200 142.9000 527.4200 143.3800 ;
        RECT 525.8200 137.4600 527.4200 137.9400 ;
        RECT 525.8200 148.3400 527.4200 148.8200 ;
        RECT 525.8200 159.2200 527.4200 159.7000 ;
        RECT 525.8200 153.7800 527.4200 154.2600 ;
        RECT 525.8200 164.6600 527.4200 165.1400 ;
        RECT 525.8200 175.5400 527.4200 176.0200 ;
        RECT 525.8200 170.1000 527.4200 170.5800 ;
        RECT 525.8200 180.9800 527.4200 181.4600 ;
        RECT 525.8200 191.8600 527.4200 192.3400 ;
        RECT 525.8200 186.4200 527.4200 186.9000 ;
        RECT 525.8200 197.3000 527.4200 197.7800 ;
        RECT 525.8200 208.1800 527.4200 208.6600 ;
        RECT 525.8200 202.7400 527.4200 203.2200 ;
        RECT 525.8200 213.6200 527.4200 214.1000 ;
        RECT 525.8200 224.5000 527.4200 224.9800 ;
        RECT 525.8200 219.0600 527.4200 219.5400 ;
        RECT 525.8200 229.9400 527.4200 230.4200 ;
        RECT 2.9600 251.7000 4.5600 252.1800 ;
        RECT 2.9600 246.2600 4.5600 246.7400 ;
        RECT 2.9600 240.8200 4.5600 241.3000 ;
        RECT 2.9600 257.1400 4.5600 257.6200 ;
        RECT 2.9600 262.5800 4.5600 263.0600 ;
        RECT 2.9600 268.0200 4.5600 268.5000 ;
        RECT 2.9600 273.4600 4.5600 273.9400 ;
        RECT 2.9600 278.9000 4.5600 279.3800 ;
        RECT 2.9600 284.3400 4.5600 284.8200 ;
        RECT 2.9600 289.7800 4.5600 290.2600 ;
        RECT 2.9600 295.2200 4.5600 295.7000 ;
        RECT 2.9600 300.6600 4.5600 301.1400 ;
        RECT 2.9600 306.1000 4.5600 306.5800 ;
        RECT 2.9600 311.5400 4.5600 312.0200 ;
        RECT 2.9600 316.9800 4.5600 317.4600 ;
        RECT 2.9600 322.4200 4.5600 322.9000 ;
        RECT 2.9600 327.8600 4.5600 328.3400 ;
        RECT 2.9600 333.3000 4.5600 333.7800 ;
        RECT 2.9600 338.7400 4.5600 339.2200 ;
        RECT 2.9600 344.1800 4.5600 344.6600 ;
        RECT 2.9600 349.6200 4.5600 350.1000 ;
        RECT 2.9600 355.0600 4.5600 355.5400 ;
        RECT 2.9600 360.5000 4.5600 360.9800 ;
        RECT 2.9600 365.9400 4.5600 366.4200 ;
        RECT 26.8500 433.0100 28.2200 434.6100 ;
        RECT 2.9600 371.3800 4.5600 371.8600 ;
        RECT 2.9600 376.8200 4.5600 377.3000 ;
        RECT 2.9600 382.2600 4.5600 382.7400 ;
        RECT 2.9600 387.7000 4.5600 388.1800 ;
        RECT 2.9600 393.1400 4.5600 393.6200 ;
        RECT 2.9600 398.5800 4.5600 399.0600 ;
        RECT 2.9600 409.4600 4.5600 409.9400 ;
        RECT 2.9600 404.0200 4.5600 404.5000 ;
        RECT 2.9600 414.9000 4.5600 415.3800 ;
        RECT 2.9600 425.7800 4.5600 426.2600 ;
        RECT 2.9600 420.3400 4.5600 420.8200 ;
        RECT 2.9600 431.2200 4.5600 431.7000 ;
        RECT 2.9600 436.6600 4.5600 437.1400 ;
        RECT 2.9600 442.1000 4.5600 442.5800 ;
        RECT 2.9600 447.5400 4.5600 448.0200 ;
        RECT 2.9600 452.9800 4.5600 453.4600 ;
        RECT 2.9600 458.4200 4.5600 458.9000 ;
        RECT 525.8200 251.7000 527.4200 252.1800 ;
        RECT 525.8200 246.2600 527.4200 246.7400 ;
        RECT 525.8200 240.8200 527.4200 241.3000 ;
        RECT 525.8200 257.1400 527.4200 257.6200 ;
        RECT 525.8200 262.5800 527.4200 263.0600 ;
        RECT 525.8200 268.0200 527.4200 268.5000 ;
        RECT 525.8200 273.4600 527.4200 273.9400 ;
        RECT 525.8200 278.9000 527.4200 279.3800 ;
        RECT 525.8200 284.3400 527.4200 284.8200 ;
        RECT 525.8200 289.7800 527.4200 290.2600 ;
        RECT 525.8200 295.2200 527.4200 295.7000 ;
        RECT 525.8200 300.6600 527.4200 301.1400 ;
        RECT 525.8200 306.1000 527.4200 306.5800 ;
        RECT 525.8200 311.5400 527.4200 312.0200 ;
        RECT 525.8200 316.9800 527.4200 317.4600 ;
        RECT 525.8200 322.4200 527.4200 322.9000 ;
        RECT 525.8200 327.8600 527.4200 328.3400 ;
        RECT 525.8200 333.3000 527.4200 333.7800 ;
        RECT 525.8200 338.7400 527.4200 339.2200 ;
        RECT 525.8200 344.1800 527.4200 344.6600 ;
        RECT 525.8200 349.6200 527.4200 350.1000 ;
        RECT 525.8200 355.0600 527.4200 355.5400 ;
        RECT 525.8200 360.5000 527.4200 360.9800 ;
        RECT 525.8200 365.9400 527.4200 366.4200 ;
        RECT 525.8200 371.3800 527.4200 371.8600 ;
        RECT 525.8200 376.8200 527.4200 377.3000 ;
        RECT 525.8200 382.2600 527.4200 382.7400 ;
        RECT 525.8200 387.7000 527.4200 388.1800 ;
        RECT 525.8200 393.1400 527.4200 393.6200 ;
        RECT 525.8200 398.5800 527.4200 399.0600 ;
        RECT 525.8200 409.4600 527.4200 409.9400 ;
        RECT 525.8200 404.0200 527.4200 404.5000 ;
        RECT 525.8200 414.9000 527.4200 415.3800 ;
        RECT 525.8200 425.7800 527.4200 426.2600 ;
        RECT 525.8200 420.3400 527.4200 420.8200 ;
        RECT 525.8200 431.2200 527.4200 431.7000 ;
        RECT 525.8200 436.6600 527.4200 437.1400 ;
        RECT 525.8200 442.1000 527.4200 442.5800 ;
        RECT 525.8200 447.5400 527.4200 448.0200 ;
        RECT 525.8200 452.9800 527.4200 453.4600 ;
        RECT 525.8200 458.4200 527.4200 458.9000 ;
      LAYER met4 ;
        RECT 2.9600 0.0000 4.5600 470.9000 ;
        RECT 525.8200 0.0000 527.4200 470.9000 ;
        RECT 26.8250 433.0100 28.2450 434.6100 ;
    END
# end of P/G power stripe data as pin


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 501.8000 39.9000 503.5400 434.6800 ;
      LAYER met3 ;
        RECT 26.4800 39.9000 503.5400 41.6400 ;
      LAYER met3 ;
        RECT 26.4800 432.9400 503.5400 434.6800 ;
      LAYER met4 ;
        RECT 26.4800 39.9000 28.2200 434.6800 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vssd1
  OBS
    LAYER li1 ;
      RECT 0.0000 0.0000 530.3800 470.9000 ;
    LAYER met1 ;
      RECT 0.0000 379.9400 530.3800 470.9000 ;
      RECT 0.8600 379.2800 530.3800 379.9400 ;
      RECT 0.0000 376.5400 530.3800 379.2800 ;
      RECT 0.8600 375.8800 530.3800 376.5400 ;
      RECT 0.0000 373.1400 530.3800 375.8800 ;
      RECT 0.8600 372.4800 530.3800 373.1400 ;
      RECT 0.0000 369.7400 530.3800 372.4800 ;
      RECT 0.8600 369.0800 530.3800 369.7400 ;
      RECT 0.0000 366.3400 530.3800 369.0800 ;
      RECT 0.8600 365.6800 530.3800 366.3400 ;
      RECT 0.0000 362.9400 530.3800 365.6800 ;
      RECT 0.8600 362.2800 530.3800 362.9400 ;
      RECT 0.0000 359.5400 530.3800 362.2800 ;
      RECT 0.8600 358.8800 530.3800 359.5400 ;
      RECT 0.0000 356.1400 530.3800 358.8800 ;
      RECT 0.8600 355.4800 530.3800 356.1400 ;
      RECT 0.0000 352.7400 530.3800 355.4800 ;
      RECT 0.8600 352.0800 530.3800 352.7400 ;
      RECT 0.0000 349.3400 530.3800 352.0800 ;
      RECT 0.8600 348.6800 530.3800 349.3400 ;
      RECT 0.0000 345.9400 530.3800 348.6800 ;
      RECT 0.8600 345.2800 530.3800 345.9400 ;
      RECT 0.0000 342.5400 530.3800 345.2800 ;
      RECT 0.8600 341.8800 530.3800 342.5400 ;
      RECT 0.0000 339.1400 530.3800 341.8800 ;
      RECT 0.8600 338.4800 530.3800 339.1400 ;
      RECT 0.0000 335.7400 530.3800 338.4800 ;
      RECT 0.8600 335.0800 530.3800 335.7400 ;
      RECT 0.0000 332.3400 530.3800 335.0800 ;
      RECT 0.8600 331.6800 530.3800 332.3400 ;
      RECT 0.0000 328.9400 530.3800 331.6800 ;
      RECT 0.8600 328.2800 530.3800 328.9400 ;
      RECT 0.0000 325.5400 530.3800 328.2800 ;
      RECT 0.8600 324.8800 530.3800 325.5400 ;
      RECT 0.0000 322.1400 530.3800 324.8800 ;
      RECT 0.8600 321.4800 530.3800 322.1400 ;
      RECT 0.0000 318.7400 530.3800 321.4800 ;
      RECT 0.8600 318.0800 530.3800 318.7400 ;
      RECT 0.0000 315.3400 530.3800 318.0800 ;
      RECT 0.8600 314.6800 530.3800 315.3400 ;
      RECT 0.0000 311.9400 530.3800 314.6800 ;
      RECT 0.8600 311.2800 530.3800 311.9400 ;
      RECT 0.0000 308.5400 530.3800 311.2800 ;
      RECT 0.8600 307.8800 530.3800 308.5400 ;
      RECT 0.0000 305.1400 530.3800 307.8800 ;
      RECT 0.8600 304.4800 530.3800 305.1400 ;
      RECT 0.0000 301.7400 530.3800 304.4800 ;
      RECT 0.8600 301.0800 530.3800 301.7400 ;
      RECT 0.0000 298.3400 530.3800 301.0800 ;
      RECT 0.8600 297.6800 530.3800 298.3400 ;
      RECT 0.0000 294.9400 530.3800 297.6800 ;
      RECT 0.8600 294.2800 530.3800 294.9400 ;
      RECT 0.0000 291.5400 530.3800 294.2800 ;
      RECT 0.8600 290.8800 530.3800 291.5400 ;
      RECT 0.0000 288.1400 530.3800 290.8800 ;
      RECT 0.8600 287.4800 530.3800 288.1400 ;
      RECT 0.0000 284.7400 530.3800 287.4800 ;
      RECT 0.8600 284.0800 530.3800 284.7400 ;
      RECT 0.0000 281.3400 530.3800 284.0800 ;
      RECT 0.8600 280.6800 530.3800 281.3400 ;
      RECT 0.0000 277.9400 530.3800 280.6800 ;
      RECT 0.8600 277.2800 530.3800 277.9400 ;
      RECT 0.0000 274.5400 530.3800 277.2800 ;
      RECT 0.8600 273.8800 530.3800 274.5400 ;
      RECT 0.0000 271.1400 530.3800 273.8800 ;
      RECT 0.8600 270.4800 530.3800 271.1400 ;
      RECT 0.0000 267.7400 530.3800 270.4800 ;
      RECT 0.8600 267.0800 530.3800 267.7400 ;
      RECT 0.0000 264.3400 530.3800 267.0800 ;
      RECT 0.8600 263.6800 530.3800 264.3400 ;
      RECT 0.0000 260.9400 530.3800 263.6800 ;
      RECT 0.8600 260.2800 530.3800 260.9400 ;
      RECT 0.0000 257.5400 530.3800 260.2800 ;
      RECT 0.8600 256.8800 530.3800 257.5400 ;
      RECT 0.0000 254.1400 530.3800 256.8800 ;
      RECT 0.8600 253.4800 530.3800 254.1400 ;
      RECT 0.0000 250.7400 530.3800 253.4800 ;
      RECT 0.8600 250.0800 530.3800 250.7400 ;
      RECT 0.0000 247.3400 530.3800 250.0800 ;
      RECT 0.8600 246.6800 530.3800 247.3400 ;
      RECT 0.0000 243.9400 530.3800 246.6800 ;
      RECT 0.8600 243.2800 530.3800 243.9400 ;
      RECT 0.0000 240.5400 530.3800 243.2800 ;
      RECT 0.8600 239.8800 530.3800 240.5400 ;
      RECT 0.0000 149.7600 530.3800 239.8800 ;
      RECT 0.8600 149.1000 530.3800 149.7600 ;
      RECT 0.0000 146.7000 530.3800 149.1000 ;
      RECT 0.8600 146.0400 530.3800 146.7000 ;
      RECT 0.0000 143.3000 530.3800 146.0400 ;
      RECT 0.8600 142.6400 530.3800 143.3000 ;
      RECT 0.0000 140.2400 530.3800 142.6400 ;
      RECT 0.8600 139.5800 530.3800 140.2400 ;
      RECT 0.0000 136.8400 530.3800 139.5800 ;
      RECT 0.8600 136.1800 530.3800 136.8400 ;
      RECT 0.0000 133.7800 530.3800 136.1800 ;
      RECT 0.8600 133.1200 530.3800 133.7800 ;
      RECT 0.0000 130.3800 530.3800 133.1200 ;
      RECT 0.8600 129.7200 530.3800 130.3800 ;
      RECT 0.0000 127.3200 530.3800 129.7200 ;
      RECT 0.8600 126.6600 530.3800 127.3200 ;
      RECT 0.0000 123.9200 530.3800 126.6600 ;
      RECT 0.8600 123.2600 530.3800 123.9200 ;
      RECT 0.0000 120.5200 530.3800 123.2600 ;
      RECT 0.8600 119.8600 530.3800 120.5200 ;
      RECT 0.0000 117.4600 530.3800 119.8600 ;
      RECT 0.8600 116.8000 530.3800 117.4600 ;
      RECT 0.0000 114.0600 530.3800 116.8000 ;
      RECT 0.8600 113.4000 530.3800 114.0600 ;
      RECT 0.0000 111.0000 530.3800 113.4000 ;
      RECT 0.8600 110.3400 530.3800 111.0000 ;
      RECT 0.0000 107.6000 530.3800 110.3400 ;
      RECT 0.8600 106.9400 530.3800 107.6000 ;
      RECT 0.0000 104.5400 530.3800 106.9400 ;
      RECT 0.8600 103.8800 530.3800 104.5400 ;
      RECT 0.0000 101.1400 530.3800 103.8800 ;
      RECT 0.8600 100.4800 530.3800 101.1400 ;
      RECT 0.0000 98.0800 530.3800 100.4800 ;
      RECT 0.8600 97.4200 530.3800 98.0800 ;
      RECT 0.0000 94.6800 530.3800 97.4200 ;
      RECT 0.8600 94.0200 530.3800 94.6800 ;
      RECT 0.0000 91.2800 530.3800 94.0200 ;
      RECT 0.8600 90.6200 530.3800 91.2800 ;
      RECT 0.0000 88.2200 530.3800 90.6200 ;
      RECT 0.8600 87.5600 530.3800 88.2200 ;
      RECT 0.0000 84.8200 530.3800 87.5600 ;
      RECT 0.8600 84.1600 530.3800 84.8200 ;
      RECT 0.0000 81.7600 530.3800 84.1600 ;
      RECT 0.8600 81.1000 530.3800 81.7600 ;
      RECT 0.0000 78.3600 530.3800 81.1000 ;
      RECT 0.8600 77.7000 530.3800 78.3600 ;
      RECT 0.0000 75.3000 530.3800 77.7000 ;
      RECT 0.8600 74.6400 530.3800 75.3000 ;
      RECT 0.0000 71.9000 530.3800 74.6400 ;
      RECT 0.8600 71.2400 530.3800 71.9000 ;
      RECT 0.0000 68.8400 530.3800 71.2400 ;
      RECT 0.8600 68.1800 530.3800 68.8400 ;
      RECT 0.0000 65.4400 530.3800 68.1800 ;
      RECT 0.8600 64.7800 530.3800 65.4400 ;
      RECT 0.0000 62.0400 530.3800 64.7800 ;
      RECT 0.8600 61.3800 530.3800 62.0400 ;
      RECT 0.0000 58.9800 530.3800 61.3800 ;
      RECT 0.8600 58.3200 530.3800 58.9800 ;
      RECT 0.0000 55.5800 530.3800 58.3200 ;
      RECT 0.8600 54.9200 530.3800 55.5800 ;
      RECT 0.0000 52.5200 530.3800 54.9200 ;
      RECT 0.8600 51.8600 530.3800 52.5200 ;
      RECT 0.0000 49.1200 530.3800 51.8600 ;
      RECT 0.8600 48.4600 530.3800 49.1200 ;
      RECT 0.0000 46.0600 530.3800 48.4600 ;
      RECT 0.8600 45.4000 530.3800 46.0600 ;
      RECT 0.0000 42.6600 530.3800 45.4000 ;
      RECT 0.8600 42.0000 530.3800 42.6600 ;
      RECT 0.0000 39.6000 530.3800 42.0000 ;
      RECT 0.8600 38.9400 530.3800 39.6000 ;
      RECT 0.0000 36.2000 530.3800 38.9400 ;
      RECT 0.8600 35.5400 530.3800 36.2000 ;
      RECT 0.0000 32.8000 530.3800 35.5400 ;
      RECT 0.8600 32.1400 530.3800 32.8000 ;
      RECT 0.0000 29.7400 530.3800 32.1400 ;
      RECT 0.8600 29.0800 530.3800 29.7400 ;
      RECT 0.0000 26.3400 530.3800 29.0800 ;
      RECT 0.8600 25.6800 530.3800 26.3400 ;
      RECT 0.0000 23.2800 530.3800 25.6800 ;
      RECT 0.8600 22.6200 530.3800 23.2800 ;
      RECT 0.0000 19.8800 530.3800 22.6200 ;
      RECT 0.8600 19.2200 530.3800 19.8800 ;
      RECT 0.0000 16.8200 530.3800 19.2200 ;
      RECT 0.8600 16.1600 530.3800 16.8200 ;
      RECT 0.0000 13.4200 530.3800 16.1600 ;
      RECT 0.8600 12.7600 530.3800 13.4200 ;
      RECT 0.0000 10.3600 530.3800 12.7600 ;
      RECT 0.8600 9.7000 530.3800 10.3600 ;
      RECT 0.0000 0.0000 530.3800 9.7000 ;
    LAYER met2 ;
      RECT 0.0000 0.0000 530.3800 470.9000 ;
    LAYER met3 ;
      RECT 0.0000 467.1800 530.3800 470.9000 ;
      RECT 0.0000 464.5800 530.3800 464.9800 ;
      RECT 0.0000 459.2000 530.3800 462.3800 ;
      RECT 527.7200 458.1200 530.3800 459.2000 ;
      RECT 4.8600 458.1200 525.5200 459.2000 ;
      RECT 0.0000 458.1200 2.6600 459.2000 ;
      RECT 0.0000 456.4800 530.3800 458.1200 ;
      RECT 525.1200 455.4000 530.3800 456.4800 ;
      RECT 7.4600 455.4000 522.9200 456.4800 ;
      RECT 0.0000 455.4000 5.2600 456.4800 ;
      RECT 0.0000 453.7600 530.3800 455.4000 ;
      RECT 527.7200 452.6800 530.3800 453.7600 ;
      RECT 4.8600 452.6800 525.5200 453.7600 ;
      RECT 0.0000 452.6800 2.6600 453.7600 ;
      RECT 0.0000 451.0400 530.3800 452.6800 ;
      RECT 525.1200 449.9600 530.3800 451.0400 ;
      RECT 7.4600 449.9600 522.9200 451.0400 ;
      RECT 0.0000 449.9600 5.2600 451.0400 ;
      RECT 0.0000 448.3200 530.3800 449.9600 ;
      RECT 527.7200 447.2400 530.3800 448.3200 ;
      RECT 4.8600 447.2400 525.5200 448.3200 ;
      RECT 0.0000 447.2400 2.6600 448.3200 ;
      RECT 0.0000 445.6000 530.3800 447.2400 ;
      RECT 525.1200 444.5200 530.3800 445.6000 ;
      RECT 7.4600 444.5200 522.9200 445.6000 ;
      RECT 0.0000 444.5200 5.2600 445.6000 ;
      RECT 0.0000 442.8800 530.3800 444.5200 ;
      RECT 527.7200 441.8000 530.3800 442.8800 ;
      RECT 4.8600 441.8000 525.5200 442.8800 ;
      RECT 0.0000 441.8000 2.6600 442.8800 ;
      RECT 0.0000 440.1600 530.3800 441.8000 ;
      RECT 525.1200 439.0800 530.3800 440.1600 ;
      RECT 7.4600 439.0800 522.9200 440.1600 ;
      RECT 0.0000 439.0800 5.2600 440.1600 ;
      RECT 0.0000 437.4400 530.3800 439.0800 ;
      RECT 527.7200 436.3600 530.3800 437.4400 ;
      RECT 4.8600 436.3600 525.5200 437.4400 ;
      RECT 0.0000 436.3600 2.6600 437.4400 ;
      RECT 0.0000 434.9100 530.3800 436.3600 ;
      RECT 28.5200 434.7200 530.3800 434.9100 ;
      RECT 0.0000 434.7200 26.5500 434.9100 ;
      RECT 525.1200 433.6400 530.3800 434.7200 ;
      RECT 28.5200 433.6400 522.9200 434.7200 ;
      RECT 7.4600 433.6400 26.5500 434.7200 ;
      RECT 0.0000 433.6400 5.2600 434.7200 ;
      RECT 28.5200 432.7100 530.3800 433.6400 ;
      RECT 0.0000 432.7100 26.5500 433.6400 ;
      RECT 0.0000 432.0000 530.3800 432.7100 ;
      RECT 4.8600 431.5100 525.5200 432.0000 ;
      RECT 527.7200 430.9200 530.3800 432.0000 ;
      RECT 31.9200 430.9200 525.5200 431.5100 ;
      RECT 4.8600 430.9200 29.9500 431.5100 ;
      RECT 0.0000 430.9200 2.6600 432.0000 ;
      RECT 31.9200 429.3100 530.3800 430.9200 ;
      RECT 0.0000 429.3100 29.9500 430.9200 ;
      RECT 0.0000 429.2800 530.3800 429.3100 ;
      RECT 525.1200 428.2000 530.3800 429.2800 ;
      RECT 7.4600 428.2000 522.9200 429.2800 ;
      RECT 0.0000 428.2000 5.2600 429.2800 ;
      RECT 0.0000 426.5600 530.3800 428.2000 ;
      RECT 527.7200 425.4800 530.3800 426.5600 ;
      RECT 4.8600 425.4800 525.5200 426.5600 ;
      RECT 0.0000 425.4800 2.6600 426.5600 ;
      RECT 0.0000 423.8400 530.3800 425.4800 ;
      RECT 525.1200 422.7600 530.3800 423.8400 ;
      RECT 7.4600 422.7600 522.9200 423.8400 ;
      RECT 0.0000 422.7600 5.2600 423.8400 ;
      RECT 0.0000 421.1200 530.3800 422.7600 ;
      RECT 527.7200 420.0400 530.3800 421.1200 ;
      RECT 4.8600 420.0400 525.5200 421.1200 ;
      RECT 0.0000 420.0400 2.6600 421.1200 ;
      RECT 0.0000 418.4000 530.3800 420.0400 ;
      RECT 525.1200 417.3200 530.3800 418.4000 ;
      RECT 7.4600 417.3200 522.9200 418.4000 ;
      RECT 0.0000 417.3200 5.2600 418.4000 ;
      RECT 0.0000 415.6800 530.3800 417.3200 ;
      RECT 527.7200 414.6000 530.3800 415.6800 ;
      RECT 4.8600 414.6000 525.5200 415.6800 ;
      RECT 0.0000 414.6000 2.6600 415.6800 ;
      RECT 0.0000 412.9600 530.3800 414.6000 ;
      RECT 525.1200 411.8800 530.3800 412.9600 ;
      RECT 7.4600 411.8800 522.9200 412.9600 ;
      RECT 0.0000 411.8800 5.2600 412.9600 ;
      RECT 0.0000 410.2400 530.3800 411.8800 ;
      RECT 527.7200 409.1600 530.3800 410.2400 ;
      RECT 4.8600 409.1600 525.5200 410.2400 ;
      RECT 0.0000 409.1600 2.6600 410.2400 ;
      RECT 0.0000 407.5200 530.3800 409.1600 ;
      RECT 525.1200 406.4400 530.3800 407.5200 ;
      RECT 7.4600 406.4400 522.9200 407.5200 ;
      RECT 0.0000 406.4400 5.2600 407.5200 ;
      RECT 0.0000 404.8000 530.3800 406.4400 ;
      RECT 527.7200 403.7200 530.3800 404.8000 ;
      RECT 4.8600 403.7200 525.5200 404.8000 ;
      RECT 0.0000 403.7200 2.6600 404.8000 ;
      RECT 0.0000 402.0800 530.3800 403.7200 ;
      RECT 525.1200 401.0000 530.3800 402.0800 ;
      RECT 7.4600 401.0000 522.9200 402.0800 ;
      RECT 0.0000 401.0000 5.2600 402.0800 ;
      RECT 0.0000 399.3600 530.3800 401.0000 ;
      RECT 527.7200 398.2800 530.3800 399.3600 ;
      RECT 4.8600 398.2800 525.5200 399.3600 ;
      RECT 0.0000 398.2800 2.6600 399.3600 ;
      RECT 0.0000 396.6400 530.3800 398.2800 ;
      RECT 525.1200 395.5600 530.3800 396.6400 ;
      RECT 7.4600 395.5600 522.9200 396.6400 ;
      RECT 0.0000 395.5600 5.2600 396.6400 ;
      RECT 0.0000 393.9200 530.3800 395.5600 ;
      RECT 527.7200 392.8400 530.3800 393.9200 ;
      RECT 4.8600 392.8400 525.5200 393.9200 ;
      RECT 0.0000 392.8400 2.6600 393.9200 ;
      RECT 0.0000 391.2000 530.3800 392.8400 ;
      RECT 525.1200 390.1200 530.3800 391.2000 ;
      RECT 7.4600 390.1200 522.9200 391.2000 ;
      RECT 0.0000 390.1200 5.2600 391.2000 ;
      RECT 0.0000 388.4800 530.3800 390.1200 ;
      RECT 527.7200 387.4000 530.3800 388.4800 ;
      RECT 4.8600 387.4000 525.5200 388.4800 ;
      RECT 0.0000 387.4000 2.6600 388.4800 ;
      RECT 0.0000 385.7600 530.3800 387.4000 ;
      RECT 525.1200 384.6800 530.3800 385.7600 ;
      RECT 7.4600 384.6800 522.9200 385.7600 ;
      RECT 0.0000 384.6800 5.2600 385.7600 ;
      RECT 0.0000 383.0400 530.3800 384.6800 ;
      RECT 527.7200 381.9600 530.3800 383.0400 ;
      RECT 4.8600 381.9600 525.5200 383.0400 ;
      RECT 0.0000 381.9600 2.6600 383.0400 ;
      RECT 0.0000 380.3200 530.3800 381.9600 ;
      RECT 525.1200 379.2400 530.3800 380.3200 ;
      RECT 7.4600 379.2400 522.9200 380.3200 ;
      RECT 0.0000 379.2400 5.2600 380.3200 ;
      RECT 0.0000 377.6000 530.3800 379.2400 ;
      RECT 527.7200 376.5200 530.3800 377.6000 ;
      RECT 4.8600 376.5200 525.5200 377.6000 ;
      RECT 0.0000 376.5200 2.6600 377.6000 ;
      RECT 0.0000 374.8800 530.3800 376.5200 ;
      RECT 525.1200 373.8000 530.3800 374.8800 ;
      RECT 7.4600 373.8000 522.9200 374.8800 ;
      RECT 0.0000 373.8000 5.2600 374.8800 ;
      RECT 0.0000 372.1600 530.3800 373.8000 ;
      RECT 527.7200 371.0800 530.3800 372.1600 ;
      RECT 4.8600 371.0800 525.5200 372.1600 ;
      RECT 0.0000 371.0800 2.6600 372.1600 ;
      RECT 0.0000 369.4400 530.3800 371.0800 ;
      RECT 525.1200 368.3600 530.3800 369.4400 ;
      RECT 7.4600 368.3600 522.9200 369.4400 ;
      RECT 0.0000 368.3600 5.2600 369.4400 ;
      RECT 0.0000 366.7200 530.3800 368.3600 ;
      RECT 527.7200 365.6400 530.3800 366.7200 ;
      RECT 4.8600 365.6400 525.5200 366.7200 ;
      RECT 0.0000 365.6400 2.6600 366.7200 ;
      RECT 0.0000 364.0000 530.3800 365.6400 ;
      RECT 525.1200 362.9200 530.3800 364.0000 ;
      RECT 7.4600 362.9200 522.9200 364.0000 ;
      RECT 0.0000 362.9200 5.2600 364.0000 ;
      RECT 0.0000 361.2800 530.3800 362.9200 ;
      RECT 527.7200 360.2000 530.3800 361.2800 ;
      RECT 4.8600 360.2000 525.5200 361.2800 ;
      RECT 0.0000 360.2000 2.6600 361.2800 ;
      RECT 0.0000 358.5600 530.3800 360.2000 ;
      RECT 525.1200 357.4800 530.3800 358.5600 ;
      RECT 7.4600 357.4800 522.9200 358.5600 ;
      RECT 0.0000 357.4800 5.2600 358.5600 ;
      RECT 0.0000 355.8400 530.3800 357.4800 ;
      RECT 527.7200 354.7600 530.3800 355.8400 ;
      RECT 4.8600 354.7600 525.5200 355.8400 ;
      RECT 0.0000 354.7600 2.6600 355.8400 ;
      RECT 0.0000 353.1200 530.3800 354.7600 ;
      RECT 525.1200 352.0400 530.3800 353.1200 ;
      RECT 7.4600 352.0400 522.9200 353.1200 ;
      RECT 0.0000 352.0400 5.2600 353.1200 ;
      RECT 0.0000 350.4000 530.3800 352.0400 ;
      RECT 527.7200 349.3200 530.3800 350.4000 ;
      RECT 4.8600 349.3200 525.5200 350.4000 ;
      RECT 0.0000 349.3200 2.6600 350.4000 ;
      RECT 0.0000 347.6800 530.3800 349.3200 ;
      RECT 525.1200 346.6000 530.3800 347.6800 ;
      RECT 7.4600 346.6000 522.9200 347.6800 ;
      RECT 0.0000 346.6000 5.2600 347.6800 ;
      RECT 0.0000 344.9600 530.3800 346.6000 ;
      RECT 527.7200 343.8800 530.3800 344.9600 ;
      RECT 4.8600 343.8800 525.5200 344.9600 ;
      RECT 0.0000 343.8800 2.6600 344.9600 ;
      RECT 0.0000 342.2400 530.3800 343.8800 ;
      RECT 525.1200 341.1600 530.3800 342.2400 ;
      RECT 7.4600 341.1600 522.9200 342.2400 ;
      RECT 0.0000 341.1600 5.2600 342.2400 ;
      RECT 0.0000 339.5200 530.3800 341.1600 ;
      RECT 527.7200 338.4400 530.3800 339.5200 ;
      RECT 4.8600 338.4400 525.5200 339.5200 ;
      RECT 0.0000 338.4400 2.6600 339.5200 ;
      RECT 0.0000 336.8000 530.3800 338.4400 ;
      RECT 525.1200 335.7200 530.3800 336.8000 ;
      RECT 7.4600 335.7200 522.9200 336.8000 ;
      RECT 0.0000 335.7200 5.2600 336.8000 ;
      RECT 0.0000 334.0800 530.3800 335.7200 ;
      RECT 527.7200 333.0000 530.3800 334.0800 ;
      RECT 4.8600 333.0000 525.5200 334.0800 ;
      RECT 0.0000 333.0000 2.6600 334.0800 ;
      RECT 0.0000 331.3600 530.3800 333.0000 ;
      RECT 525.1200 330.2800 530.3800 331.3600 ;
      RECT 7.4600 330.2800 522.9200 331.3600 ;
      RECT 0.0000 330.2800 5.2600 331.3600 ;
      RECT 0.0000 328.6400 530.3800 330.2800 ;
      RECT 527.7200 327.5600 530.3800 328.6400 ;
      RECT 4.8600 327.5600 525.5200 328.6400 ;
      RECT 0.0000 327.5600 2.6600 328.6400 ;
      RECT 0.0000 325.9200 530.3800 327.5600 ;
      RECT 525.1200 324.8400 530.3800 325.9200 ;
      RECT 7.4600 324.8400 522.9200 325.9200 ;
      RECT 0.0000 324.8400 5.2600 325.9200 ;
      RECT 0.0000 323.2000 530.3800 324.8400 ;
      RECT 527.7200 322.1200 530.3800 323.2000 ;
      RECT 4.8600 322.1200 525.5200 323.2000 ;
      RECT 0.0000 322.1200 2.6600 323.2000 ;
      RECT 0.0000 320.4800 530.3800 322.1200 ;
      RECT 525.1200 319.4000 530.3800 320.4800 ;
      RECT 7.4600 319.4000 522.9200 320.4800 ;
      RECT 0.0000 319.4000 5.2600 320.4800 ;
      RECT 0.0000 317.7600 530.3800 319.4000 ;
      RECT 527.7200 316.6800 530.3800 317.7600 ;
      RECT 4.8600 316.6800 525.5200 317.7600 ;
      RECT 0.0000 316.6800 2.6600 317.7600 ;
      RECT 0.0000 315.0400 530.3800 316.6800 ;
      RECT 525.1200 313.9600 530.3800 315.0400 ;
      RECT 7.4600 313.9600 522.9200 315.0400 ;
      RECT 0.0000 313.9600 5.2600 315.0400 ;
      RECT 0.0000 312.3200 530.3800 313.9600 ;
      RECT 527.7200 311.2400 530.3800 312.3200 ;
      RECT 4.8600 311.2400 525.5200 312.3200 ;
      RECT 0.0000 311.2400 2.6600 312.3200 ;
      RECT 0.0000 309.6000 530.3800 311.2400 ;
      RECT 525.1200 308.5200 530.3800 309.6000 ;
      RECT 7.4600 308.5200 522.9200 309.6000 ;
      RECT 0.0000 308.5200 5.2600 309.6000 ;
      RECT 0.0000 306.8800 530.3800 308.5200 ;
      RECT 527.7200 305.8000 530.3800 306.8800 ;
      RECT 4.8600 305.8000 525.5200 306.8800 ;
      RECT 0.0000 305.8000 2.6600 306.8800 ;
      RECT 0.0000 304.1600 530.3800 305.8000 ;
      RECT 525.1200 303.0800 530.3800 304.1600 ;
      RECT 7.4600 303.0800 522.9200 304.1600 ;
      RECT 0.0000 303.0800 5.2600 304.1600 ;
      RECT 0.0000 301.4400 530.3800 303.0800 ;
      RECT 527.7200 300.3600 530.3800 301.4400 ;
      RECT 4.8600 300.3600 525.5200 301.4400 ;
      RECT 0.0000 300.3600 2.6600 301.4400 ;
      RECT 0.0000 298.7200 530.3800 300.3600 ;
      RECT 525.1200 297.6400 530.3800 298.7200 ;
      RECT 7.4600 297.6400 522.9200 298.7200 ;
      RECT 0.0000 297.6400 5.2600 298.7200 ;
      RECT 0.0000 296.0000 530.3800 297.6400 ;
      RECT 527.7200 294.9200 530.3800 296.0000 ;
      RECT 4.8600 294.9200 525.5200 296.0000 ;
      RECT 0.0000 294.9200 2.6600 296.0000 ;
      RECT 0.0000 293.2800 530.3800 294.9200 ;
      RECT 525.1200 292.2000 530.3800 293.2800 ;
      RECT 7.4600 292.2000 522.9200 293.2800 ;
      RECT 0.0000 292.2000 5.2600 293.2800 ;
      RECT 0.0000 290.5600 530.3800 292.2000 ;
      RECT 527.7200 289.4800 530.3800 290.5600 ;
      RECT 4.8600 289.4800 525.5200 290.5600 ;
      RECT 0.0000 289.4800 2.6600 290.5600 ;
      RECT 0.0000 287.8400 530.3800 289.4800 ;
      RECT 525.1200 286.7600 530.3800 287.8400 ;
      RECT 7.4600 286.7600 522.9200 287.8400 ;
      RECT 0.0000 286.7600 5.2600 287.8400 ;
      RECT 0.0000 285.1200 530.3800 286.7600 ;
      RECT 527.7200 284.0400 530.3800 285.1200 ;
      RECT 4.8600 284.0400 525.5200 285.1200 ;
      RECT 0.0000 284.0400 2.6600 285.1200 ;
      RECT 0.0000 282.4000 530.3800 284.0400 ;
      RECT 525.1200 281.3200 530.3800 282.4000 ;
      RECT 7.4600 281.3200 522.9200 282.4000 ;
      RECT 0.0000 281.3200 5.2600 282.4000 ;
      RECT 0.0000 279.6800 530.3800 281.3200 ;
      RECT 527.7200 278.6000 530.3800 279.6800 ;
      RECT 4.8600 278.6000 525.5200 279.6800 ;
      RECT 0.0000 278.6000 2.6600 279.6800 ;
      RECT 0.0000 276.9600 530.3800 278.6000 ;
      RECT 525.1200 275.8800 530.3800 276.9600 ;
      RECT 7.4600 275.8800 522.9200 276.9600 ;
      RECT 0.0000 275.8800 5.2600 276.9600 ;
      RECT 0.0000 274.2400 530.3800 275.8800 ;
      RECT 527.7200 273.1600 530.3800 274.2400 ;
      RECT 4.8600 273.1600 525.5200 274.2400 ;
      RECT 0.0000 273.1600 2.6600 274.2400 ;
      RECT 0.0000 271.5200 530.3800 273.1600 ;
      RECT 525.1200 270.4400 530.3800 271.5200 ;
      RECT 7.4600 270.4400 522.9200 271.5200 ;
      RECT 0.0000 270.4400 5.2600 271.5200 ;
      RECT 0.0000 268.8000 530.3800 270.4400 ;
      RECT 527.7200 267.7200 530.3800 268.8000 ;
      RECT 4.8600 267.7200 525.5200 268.8000 ;
      RECT 0.0000 267.7200 2.6600 268.8000 ;
      RECT 0.0000 266.0800 530.3800 267.7200 ;
      RECT 525.1200 265.0000 530.3800 266.0800 ;
      RECT 7.4600 265.0000 522.9200 266.0800 ;
      RECT 0.0000 265.0000 5.2600 266.0800 ;
      RECT 0.0000 263.3600 530.3800 265.0000 ;
      RECT 527.7200 262.2800 530.3800 263.3600 ;
      RECT 4.8600 262.2800 525.5200 263.3600 ;
      RECT 0.0000 262.2800 2.6600 263.3600 ;
      RECT 0.0000 260.6400 530.3800 262.2800 ;
      RECT 525.1200 259.5600 530.3800 260.6400 ;
      RECT 7.4600 259.5600 522.9200 260.6400 ;
      RECT 0.0000 259.5600 5.2600 260.6400 ;
      RECT 0.0000 257.9200 530.3800 259.5600 ;
      RECT 527.7200 256.8400 530.3800 257.9200 ;
      RECT 4.8600 256.8400 525.5200 257.9200 ;
      RECT 0.0000 256.8400 2.6600 257.9200 ;
      RECT 0.0000 255.2000 530.3800 256.8400 ;
      RECT 525.1200 254.1200 530.3800 255.2000 ;
      RECT 7.4600 254.1200 522.9200 255.2000 ;
      RECT 0.0000 254.1200 5.2600 255.2000 ;
      RECT 0.0000 252.4800 530.3800 254.1200 ;
      RECT 527.7200 251.4000 530.3800 252.4800 ;
      RECT 4.8600 251.4000 525.5200 252.4800 ;
      RECT 0.0000 251.4000 2.6600 252.4800 ;
      RECT 0.0000 249.7600 530.3800 251.4000 ;
      RECT 525.1200 248.6800 530.3800 249.7600 ;
      RECT 7.4600 248.6800 522.9200 249.7600 ;
      RECT 0.0000 248.6800 5.2600 249.7600 ;
      RECT 0.0000 247.0400 530.3800 248.6800 ;
      RECT 527.7200 245.9600 530.3800 247.0400 ;
      RECT 4.8600 245.9600 525.5200 247.0400 ;
      RECT 0.0000 245.9600 2.6600 247.0400 ;
      RECT 0.0000 244.3200 530.3800 245.9600 ;
      RECT 525.1200 243.2400 530.3800 244.3200 ;
      RECT 7.4600 243.2400 522.9200 244.3200 ;
      RECT 0.0000 243.2400 5.2600 244.3200 ;
      RECT 0.0000 241.6000 530.3800 243.2400 ;
      RECT 527.7200 240.5200 530.3800 241.6000 ;
      RECT 4.8600 240.5200 525.5200 241.6000 ;
      RECT 0.0000 240.5200 2.6600 241.6000 ;
      RECT 0.0000 238.8800 530.3800 240.5200 ;
      RECT 525.1200 237.8000 530.3800 238.8800 ;
      RECT 7.4600 237.8000 522.9200 238.8800 ;
      RECT 0.0000 237.8000 5.2600 238.8800 ;
      RECT 0.0000 236.1600 530.3800 237.8000 ;
      RECT 527.7200 235.0800 530.3800 236.1600 ;
      RECT 4.8600 235.0800 525.5200 236.1600 ;
      RECT 0.0000 235.0800 2.6600 236.1600 ;
      RECT 0.0000 233.4400 530.3800 235.0800 ;
      RECT 525.1200 232.3600 530.3800 233.4400 ;
      RECT 7.4600 232.3600 522.9200 233.4400 ;
      RECT 0.0000 232.3600 5.2600 233.4400 ;
      RECT 0.0000 230.7200 530.3800 232.3600 ;
      RECT 527.7200 229.6400 530.3800 230.7200 ;
      RECT 4.8600 229.6400 525.5200 230.7200 ;
      RECT 0.0000 229.6400 2.6600 230.7200 ;
      RECT 0.0000 228.0000 530.3800 229.6400 ;
      RECT 525.1200 226.9200 530.3800 228.0000 ;
      RECT 7.4600 226.9200 522.9200 228.0000 ;
      RECT 0.0000 226.9200 5.2600 228.0000 ;
      RECT 0.0000 225.2800 530.3800 226.9200 ;
      RECT 527.7200 224.2000 530.3800 225.2800 ;
      RECT 4.8600 224.2000 525.5200 225.2800 ;
      RECT 0.0000 224.2000 2.6600 225.2800 ;
      RECT 0.0000 222.5600 530.3800 224.2000 ;
      RECT 525.1200 221.4800 530.3800 222.5600 ;
      RECT 7.4600 221.4800 522.9200 222.5600 ;
      RECT 0.0000 221.4800 5.2600 222.5600 ;
      RECT 0.0000 219.8400 530.3800 221.4800 ;
      RECT 527.7200 218.7600 530.3800 219.8400 ;
      RECT 4.8600 218.7600 525.5200 219.8400 ;
      RECT 0.0000 218.7600 2.6600 219.8400 ;
      RECT 0.0000 217.1200 530.3800 218.7600 ;
      RECT 525.1200 216.0400 530.3800 217.1200 ;
      RECT 7.4600 216.0400 522.9200 217.1200 ;
      RECT 0.0000 216.0400 5.2600 217.1200 ;
      RECT 0.0000 214.4000 530.3800 216.0400 ;
      RECT 527.7200 213.3200 530.3800 214.4000 ;
      RECT 4.8600 213.3200 525.5200 214.4000 ;
      RECT 0.0000 213.3200 2.6600 214.4000 ;
      RECT 0.0000 211.6800 530.3800 213.3200 ;
      RECT 525.1200 210.6000 530.3800 211.6800 ;
      RECT 7.4600 210.6000 522.9200 211.6800 ;
      RECT 0.0000 210.6000 5.2600 211.6800 ;
      RECT 0.0000 208.9600 530.3800 210.6000 ;
      RECT 527.7200 207.8800 530.3800 208.9600 ;
      RECT 4.8600 207.8800 525.5200 208.9600 ;
      RECT 0.0000 207.8800 2.6600 208.9600 ;
      RECT 0.0000 206.2400 530.3800 207.8800 ;
      RECT 525.1200 205.1600 530.3800 206.2400 ;
      RECT 7.4600 205.1600 522.9200 206.2400 ;
      RECT 0.0000 205.1600 5.2600 206.2400 ;
      RECT 0.0000 203.5200 530.3800 205.1600 ;
      RECT 527.7200 202.4400 530.3800 203.5200 ;
      RECT 4.8600 202.4400 525.5200 203.5200 ;
      RECT 0.0000 202.4400 2.6600 203.5200 ;
      RECT 0.0000 200.8000 530.3800 202.4400 ;
      RECT 525.1200 199.7200 530.3800 200.8000 ;
      RECT 7.4600 199.7200 522.9200 200.8000 ;
      RECT 0.0000 199.7200 5.2600 200.8000 ;
      RECT 0.0000 198.0800 530.3800 199.7200 ;
      RECT 527.7200 197.0000 530.3800 198.0800 ;
      RECT 4.8600 197.0000 525.5200 198.0800 ;
      RECT 0.0000 197.0000 2.6600 198.0800 ;
      RECT 0.0000 195.3600 530.3800 197.0000 ;
      RECT 525.1200 194.2800 530.3800 195.3600 ;
      RECT 7.4600 194.2800 522.9200 195.3600 ;
      RECT 0.0000 194.2800 5.2600 195.3600 ;
      RECT 0.0000 192.6400 530.3800 194.2800 ;
      RECT 527.7200 191.5600 530.3800 192.6400 ;
      RECT 4.8600 191.5600 525.5200 192.6400 ;
      RECT 0.0000 191.5600 2.6600 192.6400 ;
      RECT 0.0000 189.9200 530.3800 191.5600 ;
      RECT 525.1200 188.8400 530.3800 189.9200 ;
      RECT 7.4600 188.8400 522.9200 189.9200 ;
      RECT 0.0000 188.8400 5.2600 189.9200 ;
      RECT 0.0000 187.2000 530.3800 188.8400 ;
      RECT 527.7200 186.1200 530.3800 187.2000 ;
      RECT 4.8600 186.1200 525.5200 187.2000 ;
      RECT 0.0000 186.1200 2.6600 187.2000 ;
      RECT 0.0000 184.4800 530.3800 186.1200 ;
      RECT 525.1200 183.4000 530.3800 184.4800 ;
      RECT 7.4600 183.4000 522.9200 184.4800 ;
      RECT 0.0000 183.4000 5.2600 184.4800 ;
      RECT 0.0000 181.7600 530.3800 183.4000 ;
      RECT 527.7200 180.6800 530.3800 181.7600 ;
      RECT 4.8600 180.6800 525.5200 181.7600 ;
      RECT 0.0000 180.6800 2.6600 181.7600 ;
      RECT 0.0000 179.0400 530.3800 180.6800 ;
      RECT 525.1200 177.9600 530.3800 179.0400 ;
      RECT 7.4600 177.9600 522.9200 179.0400 ;
      RECT 0.0000 177.9600 5.2600 179.0400 ;
      RECT 0.0000 176.3200 530.3800 177.9600 ;
      RECT 527.7200 175.2400 530.3800 176.3200 ;
      RECT 4.8600 175.2400 525.5200 176.3200 ;
      RECT 0.0000 175.2400 2.6600 176.3200 ;
      RECT 0.0000 173.6000 530.3800 175.2400 ;
      RECT 525.1200 172.5200 530.3800 173.6000 ;
      RECT 7.4600 172.5200 522.9200 173.6000 ;
      RECT 0.0000 172.5200 5.2600 173.6000 ;
      RECT 0.0000 170.8800 530.3800 172.5200 ;
      RECT 527.7200 169.8000 530.3800 170.8800 ;
      RECT 4.8600 169.8000 525.5200 170.8800 ;
      RECT 0.0000 169.8000 2.6600 170.8800 ;
      RECT 0.0000 168.1600 530.3800 169.8000 ;
      RECT 525.1200 167.0800 530.3800 168.1600 ;
      RECT 7.4600 167.0800 522.9200 168.1600 ;
      RECT 0.0000 167.0800 5.2600 168.1600 ;
      RECT 0.0000 165.4400 530.3800 167.0800 ;
      RECT 527.7200 164.3600 530.3800 165.4400 ;
      RECT 4.8600 164.3600 525.5200 165.4400 ;
      RECT 0.0000 164.3600 2.6600 165.4400 ;
      RECT 0.0000 162.7200 530.3800 164.3600 ;
      RECT 525.1200 161.6400 530.3800 162.7200 ;
      RECT 7.4600 161.6400 522.9200 162.7200 ;
      RECT 0.0000 161.6400 5.2600 162.7200 ;
      RECT 0.0000 160.0000 530.3800 161.6400 ;
      RECT 527.7200 158.9200 530.3800 160.0000 ;
      RECT 4.8600 158.9200 525.5200 160.0000 ;
      RECT 0.0000 158.9200 2.6600 160.0000 ;
      RECT 0.0000 157.2800 530.3800 158.9200 ;
      RECT 525.1200 156.2000 530.3800 157.2800 ;
      RECT 7.4600 156.2000 522.9200 157.2800 ;
      RECT 0.0000 156.2000 5.2600 157.2800 ;
      RECT 0.0000 154.5600 530.3800 156.2000 ;
      RECT 527.7200 153.4800 530.3800 154.5600 ;
      RECT 4.8600 153.4800 525.5200 154.5600 ;
      RECT 0.0000 153.4800 2.6600 154.5600 ;
      RECT 0.0000 151.8400 530.3800 153.4800 ;
      RECT 525.1200 150.7600 530.3800 151.8400 ;
      RECT 7.4600 150.7600 522.9200 151.8400 ;
      RECT 0.0000 150.7600 5.2600 151.8400 ;
      RECT 0.0000 149.1200 530.3800 150.7600 ;
      RECT 527.7200 148.0400 530.3800 149.1200 ;
      RECT 4.8600 148.0400 525.5200 149.1200 ;
      RECT 0.0000 148.0400 2.6600 149.1200 ;
      RECT 0.0000 146.4000 530.3800 148.0400 ;
      RECT 525.1200 145.3200 530.3800 146.4000 ;
      RECT 7.4600 145.3200 522.9200 146.4000 ;
      RECT 0.0000 145.3200 5.2600 146.4000 ;
      RECT 0.0000 143.6800 530.3800 145.3200 ;
      RECT 527.7200 142.6000 530.3800 143.6800 ;
      RECT 4.8600 142.6000 525.5200 143.6800 ;
      RECT 0.0000 142.6000 2.6600 143.6800 ;
      RECT 0.0000 140.9600 530.3800 142.6000 ;
      RECT 525.1200 139.8800 530.3800 140.9600 ;
      RECT 7.4600 139.8800 522.9200 140.9600 ;
      RECT 0.0000 139.8800 5.2600 140.9600 ;
      RECT 0.0000 138.2400 530.3800 139.8800 ;
      RECT 527.7200 137.1600 530.3800 138.2400 ;
      RECT 4.8600 137.1600 525.5200 138.2400 ;
      RECT 0.0000 137.1600 2.6600 138.2400 ;
      RECT 0.0000 135.5200 530.3800 137.1600 ;
      RECT 525.1200 134.4400 530.3800 135.5200 ;
      RECT 7.4600 134.4400 522.9200 135.5200 ;
      RECT 0.0000 134.4400 5.2600 135.5200 ;
      RECT 0.0000 132.8000 530.3800 134.4400 ;
      RECT 527.7200 131.7200 530.3800 132.8000 ;
      RECT 4.8600 131.7200 525.5200 132.8000 ;
      RECT 0.0000 131.7200 2.6600 132.8000 ;
      RECT 0.0000 130.0800 530.3800 131.7200 ;
      RECT 525.1200 129.0000 530.3800 130.0800 ;
      RECT 7.4600 129.0000 522.9200 130.0800 ;
      RECT 0.0000 129.0000 5.2600 130.0800 ;
      RECT 0.0000 127.3600 530.3800 129.0000 ;
      RECT 527.7200 126.2800 530.3800 127.3600 ;
      RECT 4.8600 126.2800 525.5200 127.3600 ;
      RECT 0.0000 126.2800 2.6600 127.3600 ;
      RECT 0.0000 124.6400 530.3800 126.2800 ;
      RECT 525.1200 123.5600 530.3800 124.6400 ;
      RECT 7.4600 123.5600 522.9200 124.6400 ;
      RECT 0.0000 123.5600 5.2600 124.6400 ;
      RECT 0.0000 121.9200 530.3800 123.5600 ;
      RECT 527.7200 120.8400 530.3800 121.9200 ;
      RECT 4.8600 120.8400 525.5200 121.9200 ;
      RECT 0.0000 120.8400 2.6600 121.9200 ;
      RECT 0.0000 119.2000 530.3800 120.8400 ;
      RECT 525.1200 118.1200 530.3800 119.2000 ;
      RECT 7.4600 118.1200 522.9200 119.2000 ;
      RECT 0.0000 118.1200 5.2600 119.2000 ;
      RECT 0.0000 116.4800 530.3800 118.1200 ;
      RECT 527.7200 115.4000 530.3800 116.4800 ;
      RECT 4.8600 115.4000 525.5200 116.4800 ;
      RECT 0.0000 115.4000 2.6600 116.4800 ;
      RECT 0.0000 113.7600 530.3800 115.4000 ;
      RECT 525.1200 112.6800 530.3800 113.7600 ;
      RECT 7.4600 112.6800 522.9200 113.7600 ;
      RECT 0.0000 112.6800 5.2600 113.7600 ;
      RECT 0.0000 111.0400 530.3800 112.6800 ;
      RECT 527.7200 109.9600 530.3800 111.0400 ;
      RECT 4.8600 109.9600 525.5200 111.0400 ;
      RECT 0.0000 109.9600 2.6600 111.0400 ;
      RECT 0.0000 108.3200 530.3800 109.9600 ;
      RECT 525.1200 107.2400 530.3800 108.3200 ;
      RECT 7.4600 107.2400 522.9200 108.3200 ;
      RECT 0.0000 107.2400 5.2600 108.3200 ;
      RECT 0.0000 105.6000 530.3800 107.2400 ;
      RECT 527.7200 104.5200 530.3800 105.6000 ;
      RECT 4.8600 104.5200 525.5200 105.6000 ;
      RECT 0.0000 104.5200 2.6600 105.6000 ;
      RECT 0.0000 102.8800 530.3800 104.5200 ;
      RECT 525.1200 101.8000 530.3800 102.8800 ;
      RECT 7.4600 101.8000 522.9200 102.8800 ;
      RECT 0.0000 101.8000 5.2600 102.8800 ;
      RECT 0.0000 100.1600 530.3800 101.8000 ;
      RECT 527.7200 99.0800 530.3800 100.1600 ;
      RECT 4.8600 99.0800 525.5200 100.1600 ;
      RECT 0.0000 99.0800 2.6600 100.1600 ;
      RECT 0.0000 97.4400 530.3800 99.0800 ;
      RECT 525.1200 96.3600 530.3800 97.4400 ;
      RECT 7.4600 96.3600 522.9200 97.4400 ;
      RECT 0.0000 96.3600 5.2600 97.4400 ;
      RECT 0.0000 94.7200 530.3800 96.3600 ;
      RECT 527.7200 93.6400 530.3800 94.7200 ;
      RECT 4.8600 93.6400 525.5200 94.7200 ;
      RECT 0.0000 93.6400 2.6600 94.7200 ;
      RECT 0.0000 92.0000 530.3800 93.6400 ;
      RECT 525.1200 90.9200 530.3800 92.0000 ;
      RECT 7.4600 90.9200 522.9200 92.0000 ;
      RECT 0.0000 90.9200 5.2600 92.0000 ;
      RECT 0.0000 89.2800 530.3800 90.9200 ;
      RECT 527.7200 88.2000 530.3800 89.2800 ;
      RECT 4.8600 88.2000 525.5200 89.2800 ;
      RECT 0.0000 88.2000 2.6600 89.2800 ;
      RECT 0.0000 86.5600 530.3800 88.2000 ;
      RECT 525.1200 85.4800 530.3800 86.5600 ;
      RECT 7.4600 85.4800 522.9200 86.5600 ;
      RECT 0.0000 85.4800 5.2600 86.5600 ;
      RECT 0.0000 83.8400 530.3800 85.4800 ;
      RECT 527.7200 82.7600 530.3800 83.8400 ;
      RECT 4.8600 82.7600 525.5200 83.8400 ;
      RECT 0.0000 82.7600 2.6600 83.8400 ;
      RECT 0.0000 81.1200 530.3800 82.7600 ;
      RECT 525.1200 80.0400 530.3800 81.1200 ;
      RECT 7.4600 80.0400 522.9200 81.1200 ;
      RECT 0.0000 80.0400 5.2600 81.1200 ;
      RECT 0.0000 78.4000 530.3800 80.0400 ;
      RECT 527.7200 77.3200 530.3800 78.4000 ;
      RECT 4.8600 77.3200 525.5200 78.4000 ;
      RECT 0.0000 77.3200 2.6600 78.4000 ;
      RECT 0.0000 75.6800 530.3800 77.3200 ;
      RECT 525.1200 74.6000 530.3800 75.6800 ;
      RECT 7.4600 74.6000 522.9200 75.6800 ;
      RECT 0.0000 74.6000 5.2600 75.6800 ;
      RECT 0.0000 72.9600 530.3800 74.6000 ;
      RECT 527.7200 71.8800 530.3800 72.9600 ;
      RECT 4.8600 71.8800 525.5200 72.9600 ;
      RECT 0.0000 71.8800 2.6600 72.9600 ;
      RECT 0.0000 70.2400 530.3800 71.8800 ;
      RECT 525.1200 69.1600 530.3800 70.2400 ;
      RECT 7.4600 69.1600 522.9200 70.2400 ;
      RECT 0.0000 69.1600 5.2600 70.2400 ;
      RECT 0.0000 67.5200 530.3800 69.1600 ;
      RECT 527.7200 66.4400 530.3800 67.5200 ;
      RECT 4.8600 66.4400 525.5200 67.5200 ;
      RECT 0.0000 66.4400 2.6600 67.5200 ;
      RECT 0.0000 64.8000 530.3800 66.4400 ;
      RECT 525.1200 63.7200 530.3800 64.8000 ;
      RECT 7.4600 63.7200 522.9200 64.8000 ;
      RECT 0.0000 63.7200 5.2600 64.8000 ;
      RECT 0.0000 62.0800 530.3800 63.7200 ;
      RECT 527.7200 61.0000 530.3800 62.0800 ;
      RECT 4.8600 61.0000 525.5200 62.0800 ;
      RECT 0.0000 61.0000 2.6600 62.0800 ;
      RECT 0.0000 59.3600 530.3800 61.0000 ;
      RECT 525.1200 58.2800 530.3800 59.3600 ;
      RECT 7.4600 58.2800 522.9200 59.3600 ;
      RECT 0.0000 58.2800 5.2600 59.3600 ;
      RECT 0.0000 56.6400 530.3800 58.2800 ;
      RECT 527.7200 55.5600 530.3800 56.6400 ;
      RECT 4.8600 55.5600 525.5200 56.6400 ;
      RECT 0.0000 55.5600 2.6600 56.6400 ;
      RECT 0.0000 53.9200 530.3800 55.5600 ;
      RECT 525.1200 52.8400 530.3800 53.9200 ;
      RECT 7.4600 52.8400 522.9200 53.9200 ;
      RECT 0.0000 52.8400 5.2600 53.9200 ;
      RECT 0.0000 51.2000 530.3800 52.8400 ;
      RECT 527.7200 50.1200 530.3800 51.2000 ;
      RECT 4.8600 50.1200 525.5200 51.2000 ;
      RECT 0.0000 50.1200 2.6600 51.2000 ;
      RECT 0.0000 48.4800 530.3800 50.1200 ;
      RECT 525.1200 47.4000 530.3800 48.4800 ;
      RECT 7.4600 47.4000 522.9200 48.4800 ;
      RECT 0.0000 47.4000 5.2600 48.4800 ;
      RECT 0.0000 45.7600 530.3800 47.4000 ;
      RECT 527.7200 44.6800 530.3800 45.7600 ;
      RECT 4.8600 44.6800 525.5200 45.7600 ;
      RECT 0.0000 44.6800 2.6600 45.7600 ;
      RECT 0.0000 43.0400 530.3800 44.6800 ;
      RECT 525.1200 41.9600 530.3800 43.0400 ;
      RECT 7.4600 41.9600 522.9200 43.0400 ;
      RECT 0.0000 41.9600 5.2600 43.0400 ;
      RECT 0.0000 40.3200 530.3800 41.9600 ;
      RECT 527.7200 39.2400 530.3800 40.3200 ;
      RECT 4.8600 39.2400 525.5200 40.3200 ;
      RECT 0.0000 39.2400 2.6600 40.3200 ;
      RECT 0.0000 37.6000 530.3800 39.2400 ;
      RECT 525.1200 36.5200 530.3800 37.6000 ;
      RECT 7.4600 36.5200 522.9200 37.6000 ;
      RECT 0.0000 36.5200 5.2600 37.6000 ;
      RECT 0.0000 34.8800 530.3800 36.5200 ;
      RECT 527.7200 33.8000 530.3800 34.8800 ;
      RECT 4.8600 33.8000 525.5200 34.8800 ;
      RECT 0.0000 33.8000 2.6600 34.8800 ;
      RECT 0.0000 32.1600 530.3800 33.8000 ;
      RECT 525.1200 31.0800 530.3800 32.1600 ;
      RECT 7.4600 31.0800 522.9200 32.1600 ;
      RECT 0.0000 31.0800 5.2600 32.1600 ;
      RECT 0.0000 29.4400 530.3800 31.0800 ;
      RECT 527.7200 28.3600 530.3800 29.4400 ;
      RECT 4.8600 28.3600 525.5200 29.4400 ;
      RECT 0.0000 28.3600 2.6600 29.4400 ;
      RECT 0.0000 26.7200 530.3800 28.3600 ;
      RECT 525.1200 25.6400 530.3800 26.7200 ;
      RECT 7.4600 25.6400 522.9200 26.7200 ;
      RECT 0.0000 25.6400 5.2600 26.7200 ;
      RECT 0.0000 24.0000 530.3800 25.6400 ;
      RECT 527.7200 22.9200 530.3800 24.0000 ;
      RECT 4.8600 22.9200 525.5200 24.0000 ;
      RECT 0.0000 22.9200 2.6600 24.0000 ;
      RECT 0.0000 21.2800 530.3800 22.9200 ;
      RECT 525.1200 20.2000 530.3800 21.2800 ;
      RECT 7.4600 20.2000 522.9200 21.2800 ;
      RECT 0.0000 20.2000 5.2600 21.2800 ;
      RECT 0.0000 18.5600 530.3800 20.2000 ;
      RECT 527.7200 17.4800 530.3800 18.5600 ;
      RECT 4.8600 17.4800 525.5200 18.5600 ;
      RECT 0.0000 17.4800 2.6600 18.5600 ;
      RECT 0.0000 15.8400 530.3800 17.4800 ;
      RECT 525.1200 14.7600 530.3800 15.8400 ;
      RECT 7.4600 14.7600 522.9200 15.8400 ;
      RECT 0.0000 14.7600 5.2600 15.8400 ;
      RECT 0.0000 13.1200 530.3800 14.7600 ;
      RECT 527.7200 12.0400 530.3800 13.1200 ;
      RECT 4.8600 12.0400 525.5200 13.1200 ;
      RECT 0.0000 12.0400 2.6600 13.1200 ;
      RECT 0.0000 10.4000 530.3800 12.0400 ;
      RECT 525.1200 9.3200 530.3800 10.4000 ;
      RECT 7.4600 9.3200 522.9200 10.4000 ;
      RECT 0.0000 9.3200 5.2600 10.4000 ;
      RECT 0.0000 7.3300 530.3800 9.3200 ;
      RECT 0.0000 4.7300 530.3800 5.1300 ;
      RECT 0.0000 0.0000 530.3800 2.5300 ;
    LAYER met4 ;
      RECT 7.4600 434.9100 522.9200 470.9000 ;
      RECT 28.5450 432.7100 522.9200 434.9100 ;
      RECT 7.4600 432.7100 26.5250 434.9100 ;
      RECT 7.4600 431.5100 522.9200 432.7100 ;
      RECT 31.9450 429.3100 522.9200 431.5100 ;
      RECT 7.4600 429.3100 29.9250 431.5100 ;
      RECT 7.4600 1.0200 522.9200 429.3100 ;
      RECT 527.7200 0.0000 530.3800 470.9000 ;
      RECT 525.1200 0.0000 525.5200 470.9000 ;
      RECT 10.1500 0.0000 522.9200 1.0200 ;
      RECT 7.4600 0.0000 9.1700 1.0200 ;
      RECT 4.8600 0.0000 5.2600 470.9000 ;
      RECT 0.0000 0.0000 2.6600 470.9000 ;
  END
END BlockRAM_1KB
MACRO DSP
  CLASS BLOCK ;
  FOREIGN DSP ;
  ORIGIN 0.000 0.000 ;
  SIZE 223.275 BY 471.230 ;
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.400 463.720 204.540 471.230 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.640 0.000 201.780 11.940 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.080 458.280 208.220 471.230 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.380 461.340 210.520 471.230 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.480 0.000 203.620 36.760 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.320 0.000 205.460 1.090 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.160 0.000 207.300 17.410 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.000 0.000 209.140 14.660 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.220 425.980 212.360 471.230 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.590 13.890 462.890 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.840 0.000 210.980 18.400 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.280 0.000 194.420 9.560 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.120 0.000 196.260 6.500 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.830 6.990 458.130 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.190 6.990 459.490 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.960 0.000 198.100 15.000 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.240 452.840 206.380 471.230 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 203.690 459.190 223.275 459.490 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.230 7.450 461.530 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.800 0.000 199.940 17.380 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.680 0.000 212.820 5.820 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 468.030 15.730 468.330 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 464.630 223.275 464.930 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.730 466.670 223.275 466.970 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.870 468.030 223.275 468.330 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.200 0.000 218.340 8.880 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 470.070 17.110 470.370 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.040 458.960 220.180 471.230 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.390 470.070 223.275 470.370 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.040 0.000 220.180 14.320 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.880 0.000 222.020 13.980 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 464.630 19.410 464.930 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.060 465.390 214.200 471.230 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.410 461.230 223.275 461.530 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.900 456.580 216.040 471.230 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 466.670 20.330 466.970 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.200 462.020 218.340 471.230 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.520 0.000 214.660 19.760 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.360 0.000 216.500 25.200 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 200.930 462.590 223.275 462.890 ;
    END
  END FrameStrobe_O[9]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.880 424.960 222.020 471.230 ;
    END
  END UserCLK
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 5.200 99.440 465.360 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 5.200 22.640 465.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 5.200 176.240 465.360 ;
    END
  END VPWR
  PIN bot_E1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 86.550 223.275 86.850 ;
    END
  END bot_E1BEG[0]
  PIN bot_E1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 88.590 223.275 88.890 ;
    END
  END bot_E1BEG[1]
  PIN bot_E1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.210 89.950 223.275 90.250 ;
    END
  END bot_E1BEG[2]
  PIN bot_E1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 91.990 223.275 92.290 ;
    END
  END bot_E1BEG[3]
  PIN bot_E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.550 8.830 86.850 ;
    END
  END bot_E1END[0]
  PIN bot_E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.910 6.990 88.210 ;
    END
  END bot_E1END[1]
  PIN bot_E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.950 6.990 90.250 ;
    END
  END bot_E1END[2]
  PIN bot_E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.310 7.450 91.610 ;
    END
  END bot_E1END[3]
  PIN bot_E2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 94.030 223.275 94.330 ;
    END
  END bot_E2BEG[0]
  PIN bot_E2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.210 95.390 223.275 95.690 ;
    END
  END bot_E2BEG[1]
  PIN bot_E2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 97.430 223.275 97.730 ;
    END
  END bot_E2BEG[2]
  PIN bot_E2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.590 98.790 223.275 99.090 ;
    END
  END bot_E2BEG[3]
  PIN bot_E2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 100.830 223.275 101.130 ;
    END
  END bot_E2BEG[4]
  PIN bot_E2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 102.870 223.275 103.170 ;
    END
  END bot_E2BEG[5]
  PIN bot_E2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.590 104.230 223.275 104.530 ;
    END
  END bot_E2BEG[6]
  PIN bot_E2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 106.270 223.275 106.570 ;
    END
  END bot_E2BEG[7]
  PIN bot_E2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 108.310 223.275 108.610 ;
    END
  END bot_E2BEGb[0]
  PIN bot_E2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.590 109.670 223.275 109.970 ;
    END
  END bot_E2BEGb[1]
  PIN bot_E2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 111.710 223.275 112.010 ;
    END
  END bot_E2BEGb[2]
  PIN bot_E2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 113.750 223.275 114.050 ;
    END
  END bot_E2BEGb[3]
  PIN bot_E2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.590 115.110 223.275 115.410 ;
    END
  END bot_E2BEGb[4]
  PIN bot_E2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 117.150 223.275 117.450 ;
    END
  END bot_E2BEGb[5]
  PIN bot_E2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 220.710 118.510 223.275 118.810 ;
    END
  END bot_E2BEGb[6]
  PIN bot_E2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.590 120.550 223.275 120.850 ;
    END
  END bot_E2BEGb[7]
  PIN bot_E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.630 9.290 107.930 ;
    END
  END bot_E2END[0]
  PIN bot_E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.670 8.830 109.970 ;
    END
  END bot_E2END[1]
  PIN bot_E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.030 6.990 111.330 ;
    END
  END bot_E2END[2]
  PIN bot_E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.070 8.830 113.370 ;
    END
  END bot_E2END[3]
  PIN bot_E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.110 7.050 115.410 ;
    END
  END bot_E2END[4]
  PIN bot_E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.470 13.890 116.770 ;
    END
  END bot_E2END[5]
  PIN bot_E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.510 6.990 118.810 ;
    END
  END bot_E2END[6]
  PIN bot_E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.870 9.290 120.170 ;
    END
  END bot_E2END[7]
  PIN bot_E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.350 6.990 93.650 ;
    END
  END bot_E2MID[0]
  PIN bot_E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.390 6.070 95.690 ;
    END
  END bot_E2MID[1]
  PIN bot_E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.750 9.290 97.050 ;
    END
  END bot_E2MID[2]
  PIN bot_E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.790 12.050 99.090 ;
    END
  END bot_E2MID[3]
  PIN bot_E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.830 13.890 101.130 ;
    END
  END bot_E2MID[4]
  PIN bot_E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.190 19.410 102.490 ;
    END
  END bot_E2MID[5]
  PIN bot_E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.230 8.830 104.530 ;
    END
  END bot_E2MID[6]
  PIN bot_E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.590 13.890 105.890 ;
    END
  END bot_E2MID[7]
  PIN bot_E6BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 151.150 223.275 151.450 ;
    END
  END bot_E6BEG[0]
  PIN bot_E6BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 168.830 223.275 169.130 ;
    END
  END bot_E6BEG[10]
  PIN bot_E6BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 170.870 223.275 171.170 ;
    END
  END bot_E6BEG[11]
  PIN bot_E6BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 217.030 152.510 223.275 152.810 ;
    END
  END bot_E6BEG[1]
  PIN bot_E6BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 154.550 223.275 154.850 ;
    END
  END bot_E6BEG[2]
  PIN bot_E6BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 217.030 156.590 223.275 156.890 ;
    END
  END bot_E6BEG[3]
  PIN bot_E6BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 157.950 223.275 158.250 ;
    END
  END bot_E6BEG[4]
  PIN bot_E6BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.410 159.990 223.275 160.290 ;
    END
  END bot_E6BEG[5]
  PIN bot_E6BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 162.030 223.275 162.330 ;
    END
  END bot_E6BEG[6]
  PIN bot_E6BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.130 163.390 223.275 163.690 ;
    END
  END bot_E6BEG[7]
  PIN bot_E6BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.210 165.430 223.275 165.730 ;
    END
  END bot_E6BEG[8]
  PIN bot_E6BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.130 167.470 223.275 167.770 ;
    END
  END bot_E6BEG[9]
  PIN bot_E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 150.470 8.830 150.770 ;
    END
  END bot_E6END[0]
  PIN bot_E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.150 13.890 168.450 ;
    END
  END bot_E6END[10]
  PIN bot_E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.190 20.330 170.490 ;
    END
  END bot_E6END[11]
  PIN bot_E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.510 8.830 152.810 ;
    END
  END bot_E6END[1]
  PIN bot_E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.870 19.870 154.170 ;
    END
  END bot_E6END[2]
  PIN bot_E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.910 14.810 156.210 ;
    END
  END bot_E6END[3]
  PIN bot_E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.950 13.890 158.250 ;
    END
  END bot_E6END[4]
  PIN bot_E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.310 17.110 159.610 ;
    END
  END bot_E6END[5]
  PIN bot_E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.350 20.330 161.650 ;
    END
  END bot_E6END[6]
  PIN bot_E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.710 17.570 163.010 ;
    END
  END bot_E6END[7]
  PIN bot_E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.750 17.110 165.050 ;
    END
  END bot_E6END[8]
  PIN bot_E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.790 20.330 167.090 ;
    END
  END bot_E6END[9]
  PIN bot_EE4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 122.590 223.275 122.890 ;
    END
  END bot_EE4BEG[0]
  PIN bot_EE4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 140.270 223.275 140.570 ;
    END
  END bot_EE4BEG[10]
  PIN bot_EE4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.110 142.310 223.275 142.610 ;
    END
  END bot_EE4BEG[11]
  PIN bot_EE4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 143.670 223.275 143.970 ;
    END
  END bot_EE4BEG[12]
  PIN bot_EE4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 145.710 223.275 146.010 ;
    END
  END bot_EE4BEG[13]
  PIN bot_EE4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.590 147.750 223.275 148.050 ;
    END
  END bot_EE4BEG[14]
  PIN bot_EE4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.210 149.110 223.275 149.410 ;
    END
  END bot_EE4BEG[15]
  PIN bot_EE4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 123.950 223.275 124.250 ;
    END
  END bot_EE4BEG[1]
  PIN bot_EE4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.590 125.990 223.275 126.290 ;
    END
  END bot_EE4BEG[2]
  PIN bot_EE4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 128.030 223.275 128.330 ;
    END
  END bot_EE4BEG[3]
  PIN bot_EE4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 129.390 223.275 129.690 ;
    END
  END bot_EE4BEG[4]
  PIN bot_EE4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.590 131.430 223.275 131.730 ;
    END
  END bot_EE4BEG[5]
  PIN bot_EE4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 132.790 223.275 133.090 ;
    END
  END bot_EE4BEG[6]
  PIN bot_EE4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.130 134.830 223.275 135.130 ;
    END
  END bot_EE4BEG[7]
  PIN bot_EE4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.210 136.870 223.275 137.170 ;
    END
  END bot_EE4BEG[8]
  PIN bot_EE4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.210 138.230 223.275 138.530 ;
    END
  END bot_EE4BEG[9]
  PIN bot_EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.910 9.290 122.210 ;
    END
  END bot_EE4END[0]
  PIN bot_EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.590 13.890 139.890 ;
    END
  END bot_EE4END[10]
  PIN bot_EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.630 13.890 141.930 ;
    END
  END bot_EE4END[11]
  PIN bot_EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.670 14.350 143.970 ;
    END
  END bot_EE4END[12]
  PIN bot_EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.030 17.110 145.330 ;
    END
  END bot_EE4END[13]
  PIN bot_EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.070 16.650 147.370 ;
    END
  END bot_EE4END[14]
  PIN bot_EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.430 19.870 148.730 ;
    END
  END bot_EE4END[15]
  PIN bot_EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.950 6.990 124.250 ;
    END
  END bot_EE4END[1]
  PIN bot_EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.310 9.290 125.610 ;
    END
  END bot_EE4END[2]
  PIN bot_EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.350 17.110 127.650 ;
    END
  END bot_EE4END[3]
  PIN bot_EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.390 13.890 129.690 ;
    END
  END bot_EE4END[4]
  PIN bot_EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.750 20.330 131.050 ;
    END
  END bot_EE4END[5]
  PIN bot_EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.790 17.110 133.090 ;
    END
  END bot_EE4END[6]
  PIN bot_EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.150 20.330 134.450 ;
    END
  END bot_EE4END[7]
  PIN bot_EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.190 18.030 136.490 ;
    END
  END bot_EE4END[8]
  PIN bot_EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.230 17.110 138.530 ;
    END
  END bot_EE4END[9]
  PIN bot_FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.230 8.830 172.530 ;
    END
  END bot_FrameData[0]
  PIN bot_FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.910 16.190 190.210 ;
    END
  END bot_FrameData[10]
  PIN bot_FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.270 19.870 191.570 ;
    END
  END bot_FrameData[11]
  PIN bot_FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.310 13.890 193.610 ;
    END
  END bot_FrameData[12]
  PIN bot_FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.350 7.450 195.650 ;
    END
  END bot_FrameData[13]
  PIN bot_FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.710 8.830 197.010 ;
    END
  END bot_FrameData[14]
  PIN bot_FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.750 6.990 199.050 ;
    END
  END bot_FrameData[15]
  PIN bot_FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.790 6.990 201.090 ;
    END
  END bot_FrameData[16]
  PIN bot_FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.150 7.450 202.450 ;
    END
  END bot_FrameData[17]
  PIN bot_FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.190 14.350 204.490 ;
    END
  END bot_FrameData[18]
  PIN bot_FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.550 6.530 205.850 ;
    END
  END bot_FrameData[19]
  PIN bot_FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.590 7.450 173.890 ;
    END
  END bot_FrameData[1]
  PIN bot_FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.590 7.450 207.890 ;
    END
  END bot_FrameData[20]
  PIN bot_FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.630 6.990 209.930 ;
    END
  END bot_FrameData[21]
  PIN bot_FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.990 14.350 211.290 ;
    END
  END bot_FrameData[22]
  PIN bot_FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.030 16.650 213.330 ;
    END
  END bot_FrameData[23]
  PIN bot_FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.070 19.410 215.370 ;
    END
  END bot_FrameData[24]
  PIN bot_FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.430 20.330 216.730 ;
    END
  END bot_FrameData[25]
  PIN bot_FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 218.470 6.990 218.770 ;
    END
  END bot_FrameData[26]
  PIN bot_FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.830 6.530 220.130 ;
    END
  END bot_FrameData[27]
  PIN bot_FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.870 7.450 222.170 ;
    END
  END bot_FrameData[28]
  PIN bot_FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.910 8.830 224.210 ;
    END
  END bot_FrameData[29]
  PIN bot_FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.630 8.830 175.930 ;
    END
  END bot_FrameData[2]
  PIN bot_FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.270 6.990 225.570 ;
    END
  END bot_FrameData[30]
  PIN bot_FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.310 6.530 227.610 ;
    END
  END bot_FrameData[31]
  PIN bot_FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.990 7.450 177.290 ;
    END
  END bot_FrameData[3]
  PIN bot_FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.030 18.950 179.330 ;
    END
  END bot_FrameData[4]
  PIN bot_FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 181.070 6.990 181.370 ;
    END
  END bot_FrameData[5]
  PIN bot_FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.430 8.830 182.730 ;
    END
  END bot_FrameData[6]
  PIN bot_FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.470 7.450 184.770 ;
    END
  END bot_FrameData[7]
  PIN bot_FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.510 18.950 186.810 ;
    END
  END bot_FrameData[8]
  PIN bot_FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.870 17.570 188.170 ;
    END
  END bot_FrameData[9]
  PIN bot_FrameData_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 172.230 223.275 172.530 ;
    END
  END bot_FrameData_O[0]
  PIN bot_FrameData_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 190.590 223.275 190.890 ;
    END
  END bot_FrameData_O[10]
  PIN bot_FrameData_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 191.950 223.275 192.250 ;
    END
  END bot_FrameData_O[11]
  PIN bot_FrameData_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 193.990 223.275 194.290 ;
    END
  END bot_FrameData_O[12]
  PIN bot_FrameData_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.410 196.030 223.275 196.330 ;
    END
  END bot_FrameData_O[13]
  PIN bot_FrameData_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 197.390 223.275 197.690 ;
    END
  END bot_FrameData_O[14]
  PIN bot_FrameData_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 199.430 223.275 199.730 ;
    END
  END bot_FrameData_O[15]
  PIN bot_FrameData_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.130 201.470 223.275 201.770 ;
    END
  END bot_FrameData_O[16]
  PIN bot_FrameData_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 202.830 223.275 203.130 ;
    END
  END bot_FrameData_O[17]
  PIN bot_FrameData_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 204.870 223.275 205.170 ;
    END
  END bot_FrameData_O[18]
  PIN bot_FrameData_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 206.910 223.275 207.210 ;
    END
  END bot_FrameData_O[19]
  PIN bot_FrameData_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 174.270 223.275 174.570 ;
    END
  END bot_FrameData_O[1]
  PIN bot_FrameData_O[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.410 208.270 223.275 208.570 ;
    END
  END bot_FrameData_O[20]
  PIN bot_FrameData_O[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 210.310 223.275 210.610 ;
    END
  END bot_FrameData_O[21]
  PIN bot_FrameData_O[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 211.670 223.275 211.970 ;
    END
  END bot_FrameData_O[22]
  PIN bot_FrameData_O[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 213.710 223.275 214.010 ;
    END
  END bot_FrameData_O[23]
  PIN bot_FrameData_O[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 215.750 223.275 216.050 ;
    END
  END bot_FrameData_O[24]
  PIN bot_FrameData_O[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 217.110 223.275 217.410 ;
    END
  END bot_FrameData_O[25]
  PIN bot_FrameData_O[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 219.150 223.275 219.450 ;
    END
  END bot_FrameData_O[26]
  PIN bot_FrameData_O[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.410 221.190 223.275 221.490 ;
    END
  END bot_FrameData_O[27]
  PIN bot_FrameData_O[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.130 222.550 223.275 222.850 ;
    END
  END bot_FrameData_O[28]
  PIN bot_FrameData_O[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.210 224.590 223.275 224.890 ;
    END
  END bot_FrameData_O[29]
  PIN bot_FrameData_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 176.310 223.275 176.610 ;
    END
  END bot_FrameData_O[2]
  PIN bot_FrameData_O[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 226.630 223.275 226.930 ;
    END
  END bot_FrameData_O[30]
  PIN bot_FrameData_O[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.410 227.990 223.275 228.290 ;
    END
  END bot_FrameData_O[31]
  PIN bot_FrameData_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 177.670 223.275 177.970 ;
    END
  END bot_FrameData_O[3]
  PIN bot_FrameData_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 179.710 223.275 180.010 ;
    END
  END bot_FrameData_O[4]
  PIN bot_FrameData_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.410 181.750 223.275 182.050 ;
    END
  END bot_FrameData_O[5]
  PIN bot_FrameData_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 183.110 223.275 183.410 ;
    END
  END bot_FrameData_O[6]
  PIN bot_FrameData_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 185.150 223.275 185.450 ;
    END
  END bot_FrameData_O[7]
  PIN bot_FrameData_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.210 187.190 223.275 187.490 ;
    END
  END bot_FrameData_O[8]
  PIN bot_FrameData_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.130 188.550 223.275 188.850 ;
    END
  END bot_FrameData_O[9]
  PIN bot_N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.080 0.000 1.220 6.500 ;
    END
  END bot_N1END[0]
  PIN bot_N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.920 0.000 3.060 11.940 ;
    END
  END bot_N1END[1]
  PIN bot_N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.760 0.000 4.900 9.560 ;
    END
  END bot_N1END[2]
  PIN bot_N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.600 0.000 6.740 15.000 ;
    END
  END bot_N1END[3]
  PIN bot_N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.160 0.000 23.300 6.160 ;
    END
  END bot_N2END[0]
  PIN bot_N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.000 0.000 25.140 6.500 ;
    END
  END bot_N2END[1]
  PIN bot_N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.840 0.000 26.980 9.220 ;
    END
  END bot_N2END[2]
  PIN bot_N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.680 0.000 28.820 6.160 ;
    END
  END bot_N2END[3]
  PIN bot_N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.520 0.000 30.660 15.000 ;
    END
  END bot_N2END[4]
  PIN bot_N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.360 0.000 32.500 9.560 ;
    END
  END bot_N2END[5]
  PIN bot_N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.200 0.000 34.340 11.940 ;
    END
  END bot_N2END[6]
  PIN bot_N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.040 0.000 36.180 6.160 ;
    END
  END bot_N2END[7]
  PIN bot_N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.440 0.000 8.580 11.940 ;
    END
  END bot_N2MID[0]
  PIN bot_N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.280 0.000 10.420 3.780 ;
    END
  END bot_N2MID[1]
  PIN bot_N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.120 0.000 12.260 9.560 ;
    END
  END bot_N2MID[2]
  PIN bot_N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.960 0.000 14.100 15.000 ;
    END
  END bot_N2MID[3]
  PIN bot_N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.800 0.000 15.940 1.090 ;
    END
  END bot_N2MID[4]
  PIN bot_N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.640 0.000 17.780 1.090 ;
    END
  END bot_N2MID[5]
  PIN bot_N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.480 0.000 19.620 11.940 ;
    END
  END bot_N2MID[6]
  PIN bot_N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.320 0.000 21.460 6.840 ;
    END
  END bot_N2MID[7]
  PIN bot_N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.880 0.000 38.020 11.940 ;
    END
  END bot_N4END[0]
  PIN bot_N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.740 0.000 56.880 9.560 ;
    END
  END bot_N4END[10]
  PIN bot_N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.580 0.000 58.720 1.090 ;
    END
  END bot_N4END[11]
  PIN bot_N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.420 0.000 60.560 9.220 ;
    END
  END bot_N4END[12]
  PIN bot_N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.260 0.000 62.400 6.840 ;
    END
  END bot_N4END[13]
  PIN bot_N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.100 0.000 64.240 7.520 ;
    END
  END bot_N4END[14]
  PIN bot_N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.940 0.000 66.080 13.870 ;
    END
  END bot_N4END[15]
  PIN bot_N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.720 0.000 39.860 9.560 ;
    END
  END bot_N4END[1]
  PIN bot_N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.560 0.000 41.700 9.760 ;
    END
  END bot_N4END[2]
  PIN bot_N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.400 0.000 43.540 6.160 ;
    END
  END bot_N4END[3]
  PIN bot_N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.700 0.000 45.840 14.520 ;
    END
  END bot_N4END[4]
  PIN bot_N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.540 0.000 47.680 16.700 ;
    END
  END bot_N4END[5]
  PIN bot_N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.380 0.000 49.520 14.690 ;
    END
  END bot_N4END[6]
  PIN bot_N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.220 0.000 51.360 31.320 ;
    END
  END bot_N4END[7]
  PIN bot_N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.060 0.000 53.200 16.700 ;
    END
  END bot_N4END[8]
  PIN bot_N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.900 0.000 55.040 5.170 ;
    END
  END bot_N4END[9]
  PIN bot_NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.780 0.000 67.920 6.500 ;
    END
  END bot_NN4END[0]
  PIN bot_NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.180 0.000 86.320 25.540 ;
    END
  END bot_NN4END[10]
  PIN bot_NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.020 0.000 88.160 1.090 ;
    END
  END bot_NN4END[11]
  PIN bot_NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.320 0.000 90.460 39.140 ;
    END
  END bot_NN4END[12]
  PIN bot_NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.160 0.000 92.300 12.820 ;
    END
  END bot_NN4END[13]
  PIN bot_NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.000 0.000 94.140 1.090 ;
    END
  END bot_NN4END[14]
  PIN bot_NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.840 0.000 95.980 19.420 ;
    END
  END bot_NN4END[15]
  PIN bot_NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.620 0.000 69.760 5.820 ;
    END
  END bot_NN4END[1]
  PIN bot_NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.460 0.000 71.600 6.160 ;
    END
  END bot_NN4END[2]
  PIN bot_NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.300 0.000 73.440 6.500 ;
    END
  END bot_NN4END[3]
  PIN bot_NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.140 0.000 75.280 22.850 ;
    END
  END bot_NN4END[4]
  PIN bot_NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.980 0.000 77.120 13.870 ;
    END
  END bot_NN4END[5]
  PIN bot_NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.820 0.000 78.960 7.210 ;
    END
  END bot_NN4END[6]
  PIN bot_NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.660 0.000 80.800 42.200 ;
    END
  END bot_NN4END[7]
  PIN bot_NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.500 0.000 82.640 14.480 ;
    END
  END bot_NN4END[8]
  PIN bot_NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.340 0.000 84.480 6.020 ;
    END
  END bot_NN4END[9]
  PIN bot_S1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.680 0.000 97.820 1.400 ;
    END
  END bot_S1BEG[0]
  PIN bot_S1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.520 0.000 99.660 3.130 ;
    END
  END bot_S1BEG[1]
  PIN bot_S1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.360 0.000 101.500 1.090 ;
    END
  END bot_S1BEG[2]
  PIN bot_S1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.200 0.000 103.340 8.540 ;
    END
  END bot_S1BEG[3]
  PIN bot_S2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.760 0.000 119.900 5.820 ;
    END
  END bot_S2BEG[0]
  PIN bot_S2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.600 0.000 121.740 6.500 ;
    END
  END bot_S2BEG[1]
  PIN bot_S2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.440 0.000 123.580 8.540 ;
    END
  END bot_S2BEG[2]
  PIN bot_S2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.280 0.000 125.420 5.820 ;
    END
  END bot_S2BEG[3]
  PIN bot_S2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.120 0.000 127.260 8.540 ;
    END
  END bot_S2BEG[4]
  PIN bot_S2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.960 0.000 129.100 3.100 ;
    END
  END bot_S2BEG[5]
  PIN bot_S2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.800 0.000 130.940 8.880 ;
    END
  END bot_S2BEG[6]
  PIN bot_S2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.640 0.000 132.780 6.500 ;
    END
  END bot_S2BEG[7]
  PIN bot_S2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.040 0.000 105.180 2.080 ;
    END
  END bot_S2BEGb[0]
  PIN bot_S2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.880 0.000 107.020 4.460 ;
    END
  END bot_S2BEGb[1]
  PIN bot_S2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.720 0.000 108.860 13.980 ;
    END
  END bot_S2BEGb[2]
  PIN bot_S2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.560 0.000 110.700 13.800 ;
    END
  END bot_S2BEGb[3]
  PIN bot_S2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.400 0.000 112.540 3.780 ;
    END
  END bot_S2BEGb[4]
  PIN bot_S2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.240 0.000 114.380 15.840 ;
    END
  END bot_S2BEGb[5]
  PIN bot_S2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.080 0.000 116.220 13.800 ;
    END
  END bot_S2BEGb[6]
  PIN bot_S2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.920 0.000 118.060 13.980 ;
    END
  END bot_S2BEGb[7]
  PIN bot_S4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.940 0.000 135.080 8.540 ;
    END
  END bot_S4BEG[0]
  PIN bot_S4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.340 0.000 153.480 5.820 ;
    END
  END bot_S4BEG[10]
  PIN bot_S4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.180 0.000 155.320 8.540 ;
    END
  END bot_S4BEG[11]
  PIN bot_S4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.020 0.000 157.160 5.820 ;
    END
  END bot_S4BEG[12]
  PIN bot_S4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.860 0.000 159.000 8.540 ;
    END
  END bot_S4BEG[13]
  PIN bot_S4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.700 0.000 160.840 6.160 ;
    END
  END bot_S4BEG[14]
  PIN bot_S4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.540 0.000 162.680 8.880 ;
    END
  END bot_S4BEG[15]
  PIN bot_S4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.780 0.000 136.920 6.840 ;
    END
  END bot_S4BEG[1]
  PIN bot_S4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.620 0.000 138.760 8.880 ;
    END
  END bot_S4BEG[2]
  PIN bot_S4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.460 0.000 140.600 1.090 ;
    END
  END bot_S4BEG[3]
  PIN bot_S4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.300 0.000 142.440 11.260 ;
    END
  END bot_S4BEG[4]
  PIN bot_S4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.140 0.000 144.280 7.210 ;
    END
  END bot_S4BEG[5]
  PIN bot_S4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.980 0.000 146.120 4.460 ;
    END
  END bot_S4BEG[6]
  PIN bot_S4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.820 0.000 147.960 6.840 ;
    END
  END bot_S4BEG[7]
  PIN bot_S4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.660 0.000 149.800 3.100 ;
    END
  END bot_S4BEG[8]
  PIN bot_S4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.500 0.000 151.640 11.940 ;
    END
  END bot_S4BEG[9]
  PIN bot_SS4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.380 0.000 164.520 8.540 ;
    END
  END bot_SS4BEG[0]
  PIN bot_SS4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.240 0.000 183.380 5.820 ;
    END
  END bot_SS4BEG[10]
  PIN bot_SS4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.080 0.000 185.220 8.880 ;
    END
  END bot_SS4BEG[11]
  PIN bot_SS4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.920 0.000 187.060 6.160 ;
    END
  END bot_SS4BEG[12]
  PIN bot_SS4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.760 0.000 188.900 13.980 ;
    END
  END bot_SS4BEG[13]
  PIN bot_SS4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.600 0.000 190.740 5.850 ;
    END
  END bot_SS4BEG[14]
  PIN bot_SS4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.440 0.000 192.580 8.540 ;
    END
  END bot_SS4BEG[15]
  PIN bot_SS4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.220 0.000 166.360 13.980 ;
    END
  END bot_SS4BEG[1]
  PIN bot_SS4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.060 0.000 168.200 1.090 ;
    END
  END bot_SS4BEG[2]
  PIN bot_SS4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.900 0.000 170.040 8.880 ;
    END
  END bot_SS4BEG[3]
  PIN bot_SS4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.740 0.000 171.880 13.980 ;
    END
  END bot_SS4BEG[4]
  PIN bot_SS4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.580 0.000 173.720 12.280 ;
    END
  END bot_SS4BEG[5]
  PIN bot_SS4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.420 0.000 175.560 1.090 ;
    END
  END bot_SS4BEG[6]
  PIN bot_SS4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.260 0.000 177.400 14.320 ;
    END
  END bot_SS4BEG[7]
  PIN bot_SS4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.560 0.000 179.700 16.700 ;
    END
  END bot_SS4BEG[8]
  PIN bot_SS4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.400 0.000 181.540 16.700 ;
    END
  END bot_SS4BEG[9]
  PIN bot_W1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.870 15.270 1.170 ;
    END
  END bot_W1BEG[0]
  PIN bot_W1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.230 15.730 2.530 ;
    END
  END bot_W1BEG[1]
  PIN bot_W1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.270 14.810 4.570 ;
    END
  END bot_W1BEG[2]
  PIN bot_W1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.630 18.030 5.930 ;
    END
  END bot_W1BEG[3]
  PIN bot_W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.450 0.870 223.275 1.170 ;
    END
  END bot_W1END[0]
  PIN bot_W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.390 2.230 223.275 2.530 ;
    END
  END bot_W1END[1]
  PIN bot_W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.130 4.270 223.275 4.570 ;
    END
  END bot_W1END[2]
  PIN bot_W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 200.930 5.630 223.275 5.930 ;
    END
  END bot_W1END[3]
  PIN bot_W2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.670 19.870 7.970 ;
    END
  END bot_W2BEG[0]
  PIN bot_W2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.710 16.190 10.010 ;
    END
  END bot_W2BEG[1]
  PIN bot_W2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.070 16.650 11.370 ;
    END
  END bot_W2BEG[2]
  PIN bot_W2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.110 17.110 13.410 ;
    END
  END bot_W2BEG[3]
  PIN bot_W2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.150 20.330 15.450 ;
    END
  END bot_W2BEG[4]
  PIN bot_W2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.510 15.270 16.810 ;
    END
  END bot_W2BEG[5]
  PIN bot_W2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.550 6.530 18.850 ;
    END
  END bot_W2BEG[6]
  PIN bot_W2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.910 19.870 20.210 ;
    END
  END bot_W2BEG[7]
  PIN bot_W2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.950 6.990 22.250 ;
    END
  END bot_W2BEGb[0]
  PIN bot_W2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.990 13.890 24.290 ;
    END
  END bot_W2BEGb[1]
  PIN bot_W2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.350 17.110 25.650 ;
    END
  END bot_W2BEGb[2]
  PIN bot_W2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.390 9.750 27.690 ;
    END
  END bot_W2BEGb[3]
  PIN bot_W2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.430 6.990 29.730 ;
    END
  END bot_W2BEGb[4]
  PIN bot_W2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.790 13.890 31.090 ;
    END
  END bot_W2BEGb[5]
  PIN bot_W2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.830 9.750 33.130 ;
    END
  END bot_W2BEGb[6]
  PIN bot_W2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.190 6.990 34.490 ;
    END
  END bot_W2BEGb[7]
  PIN bot_W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 205.070 21.950 223.275 22.250 ;
    END
  END bot_W2END[0]
  PIN bot_W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.390 23.990 223.275 24.290 ;
    END
  END bot_W2END[1]
  PIN bot_W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 205.530 25.350 223.275 25.650 ;
    END
  END bot_W2END[2]
  PIN bot_W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 207.370 27.390 223.275 27.690 ;
    END
  END bot_W2END[3]
  PIN bot_W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 202.770 29.430 223.275 29.730 ;
    END
  END bot_W2END[4]
  PIN bot_W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 212.430 30.790 223.275 31.090 ;
    END
  END bot_W2END[5]
  PIN bot_W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 205.530 32.830 223.275 33.130 ;
    END
  END bot_W2END[6]
  PIN bot_W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 34.870 223.275 35.170 ;
    END
  END bot_W2END[7]
  PIN bot_W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 211.970 7.670 223.275 7.970 ;
    END
  END bot_W2MID[0]
  PIN bot_W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 200.930 9.710 223.275 10.010 ;
    END
  END bot_W2MID[1]
  PIN bot_W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 200.470 11.070 223.275 11.370 ;
    END
  END bot_W2MID[2]
  PIN bot_W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 200.470 13.110 223.275 13.410 ;
    END
  END bot_W2MID[3]
  PIN bot_W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 200.930 15.150 223.275 15.450 ;
    END
  END bot_W2MID[4]
  PIN bot_W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 202.770 16.510 223.275 16.810 ;
    END
  END bot_W2MID[5]
  PIN bot_W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.450 18.550 223.275 18.850 ;
    END
  END bot_W2MID[6]
  PIN bot_W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 19.910 223.275 20.210 ;
    END
  END bot_W2MID[7]
  PIN bot_W6BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.790 9.750 65.090 ;
    END
  END bot_W6BEG[0]
  PIN bot_W6BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.470 10.210 82.770 ;
    END
  END bot_W6BEG[10]
  PIN bot_W6BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.510 16.650 84.810 ;
    END
  END bot_W6BEG[11]
  PIN bot_W6BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.830 9.750 67.130 ;
    END
  END bot_W6BEG[1]
  PIN bot_W6BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.190 6.990 68.490 ;
    END
  END bot_W6BEG[2]
  PIN bot_W6BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.230 9.750 70.530 ;
    END
  END bot_W6BEG[3]
  PIN bot_W6BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.270 6.990 72.570 ;
    END
  END bot_W6BEG[4]
  PIN bot_W6BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.630 13.890 73.930 ;
    END
  END bot_W6BEG[5]
  PIN bot_W6BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.670 9.750 75.970 ;
    END
  END bot_W6BEG[6]
  PIN bot_W6BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.030 13.890 77.330 ;
    END
  END bot_W6BEG[7]
  PIN bot_W6BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.070 13.890 79.370 ;
    END
  END bot_W6BEG[8]
  PIN bot_W6BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.110 13.890 81.410 ;
    END
  END bot_W6BEG[9]
  PIN bot_W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 211.970 64.790 223.275 65.090 ;
    END
  END bot_W6END[0]
  PIN bot_W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 83.150 223.275 83.450 ;
    END
  END bot_W6END[10]
  PIN bot_W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.130 84.510 223.275 84.810 ;
    END
  END bot_W6END[11]
  PIN bot_W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 66.830 223.275 67.130 ;
    END
  END bot_W6END[1]
  PIN bot_W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 68.870 223.275 69.170 ;
    END
  END bot_W6END[2]
  PIN bot_W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.130 70.230 223.275 70.530 ;
    END
  END bot_W6END[3]
  PIN bot_W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.510 72.270 223.275 72.570 ;
    END
  END bot_W6END[4]
  PIN bot_W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.670 74.310 223.275 74.610 ;
    END
  END bot_W6END[5]
  PIN bot_W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.910 75.670 223.275 75.970 ;
    END
  END bot_W6END[6]
  PIN bot_W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 205.990 77.710 223.275 78.010 ;
    END
  END bot_W6END[7]
  PIN bot_W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.910 79.070 223.275 79.370 ;
    END
  END bot_W6END[8]
  PIN bot_W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 203.690 81.110 223.275 81.410 ;
    END
  END bot_W6END[9]
  PIN bot_WW4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.230 13.890 36.530 ;
    END
  END bot_WW4BEG[0]
  PIN bot_WW4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.910 10.210 54.210 ;
    END
  END bot_WW4BEG[10]
  PIN bot_WW4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.950 9.750 56.250 ;
    END
  END bot_WW4BEG[11]
  PIN bot_WW4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.990 9.750 58.290 ;
    END
  END bot_WW4BEG[12]
  PIN bot_WW4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.350 6.990 59.650 ;
    END
  END bot_WW4BEG[13]
  PIN bot_WW4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.390 13.890 61.690 ;
    END
  END bot_WW4BEG[14]
  PIN bot_WW4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.750 17.110 63.050 ;
    END
  END bot_WW4BEG[15]
  PIN bot_WW4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.270 10.210 38.570 ;
    END
  END bot_WW4BEG[1]
  PIN bot_WW4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.630 6.990 39.930 ;
    END
  END bot_WW4BEG[2]
  PIN bot_WW4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.670 13.890 41.970 ;
    END
  END bot_WW4BEG[3]
  PIN bot_WW4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.710 9.750 44.010 ;
    END
  END bot_WW4BEG[4]
  PIN bot_WW4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.070 6.990 45.370 ;
    END
  END bot_WW4BEG[5]
  PIN bot_WW4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.110 13.890 47.410 ;
    END
  END bot_WW4BEG[6]
  PIN bot_WW4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.470 9.750 48.770 ;
    END
  END bot_WW4BEG[7]
  PIN bot_WW4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.510 13.890 50.810 ;
    END
  END bot_WW4BEG[8]
  PIN bot_WW4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.550 17.110 52.850 ;
    END
  END bot_WW4BEG[9]
  PIN bot_WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.910 36.230 223.275 36.530 ;
    END
  END bot_WW4END[0]
  PIN bot_WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.450 54.590 223.275 54.890 ;
    END
  END bot_WW4END[10]
  PIN bot_WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.510 55.950 223.275 56.250 ;
    END
  END bot_WW4END[11]
  PIN bot_WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 205.990 57.990 223.275 58.290 ;
    END
  END bot_WW4END[12]
  PIN bot_WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 59.350 223.275 59.650 ;
    END
  END bot_WW4END[13]
  PIN bot_WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.450 61.390 223.275 61.690 ;
    END
  END bot_WW4END[14]
  PIN bot_WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.910 63.430 223.275 63.730 ;
    END
  END bot_WW4END[15]
  PIN bot_WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 208.290 38.270 223.275 38.570 ;
    END
  END bot_WW4END[1]
  PIN bot_WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 211.970 39.630 223.275 39.930 ;
    END
  END bot_WW4END[2]
  PIN bot_WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.910 41.670 223.275 41.970 ;
    END
  END bot_WW4END[3]
  PIN bot_WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 43.710 223.275 44.010 ;
    END
  END bot_WW4END[4]
  PIN bot_WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.130 45.070 223.275 45.370 ;
    END
  END bot_WW4END[5]
  PIN bot_WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.670 47.110 223.275 47.410 ;
    END
  END bot_WW4END[6]
  PIN bot_WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.910 49.150 223.275 49.450 ;
    END
  END bot_WW4END[7]
  PIN bot_WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 205.990 50.510 223.275 50.810 ;
    END
  END bot_WW4END[8]
  PIN bot_WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 212.830 52.550 223.275 52.850 ;
    END
  END bot_WW4END[9]
  PIN top_E1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 315.710 223.275 316.010 ;
    END
  END top_E1BEG[0]
  PIN top_E1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.870 317.750 223.275 318.050 ;
    END
  END top_E1BEG[1]
  PIN top_E1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 220.250 319.790 223.275 320.090 ;
    END
  END top_E1BEG[2]
  PIN top_E1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.130 321.150 223.275 321.450 ;
    END
  END top_E1BEG[3]
  PIN top_E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 315.030 7.450 315.330 ;
    END
  END top_E1END[0]
  PIN top_E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.390 8.830 316.690 ;
    END
  END top_E1END[1]
  PIN top_E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.430 6.990 318.730 ;
    END
  END top_E1END[2]
  PIN top_E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.790 6.530 320.090 ;
    END
  END top_E1END[3]
  PIN top_E2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 323.190 223.275 323.490 ;
    END
  END top_E2BEG[0]
  PIN top_E2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 324.550 223.275 324.850 ;
    END
  END top_E2BEG[1]
  PIN top_E2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.410 326.590 223.275 326.890 ;
    END
  END top_E2BEG[2]
  PIN top_E2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 328.630 223.275 328.930 ;
    END
  END top_E2BEG[3]
  PIN top_E2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 329.990 223.275 330.290 ;
    END
  END top_E2BEG[4]
  PIN top_E2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.410 332.030 223.275 332.330 ;
    END
  END top_E2BEG[5]
  PIN top_E2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 334.070 223.275 334.370 ;
    END
  END top_E2BEG[6]
  PIN top_E2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 335.430 223.275 335.730 ;
    END
  END top_E2BEG[7]
  PIN top_E2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 222.090 337.470 223.275 337.770 ;
    END
  END top_E2BEGb[0]
  PIN top_E2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.410 339.510 223.275 339.810 ;
    END
  END top_E2BEGb[1]
  PIN top_E2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 340.870 223.275 341.170 ;
    END
  END top_E2BEGb[2]
  PIN top_E2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 342.910 223.275 343.210 ;
    END
  END top_E2BEGb[3]
  PIN top_E2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.350 344.270 223.275 344.570 ;
    END
  END top_E2BEGb[4]
  PIN top_E2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 346.310 223.275 346.610 ;
    END
  END top_E2BEGb[5]
  PIN top_E2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 220.710 348.350 223.275 348.650 ;
    END
  END top_E2BEGb[6]
  PIN top_E2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 349.710 223.275 350.010 ;
    END
  END top_E2BEGb[7]
  PIN top_E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.110 6.990 336.410 ;
    END
  END top_E2END[0]
  PIN top_E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.150 11.590 338.450 ;
    END
  END top_E2END[1]
  PIN top_E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 339.510 6.990 339.810 ;
    END
  END top_E2END[2]
  PIN top_E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.550 6.530 341.850 ;
    END
  END top_E2END[3]
  PIN top_E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.590 11.590 343.890 ;
    END
  END top_E2END[4]
  PIN top_E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.950 9.290 345.250 ;
    END
  END top_E2END[5]
  PIN top_E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.990 6.990 347.290 ;
    END
  END top_E2END[6]
  PIN top_E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.350 9.290 348.650 ;
    END
  END top_E2END[7]
  PIN top_E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.830 8.830 322.130 ;
    END
  END top_E2MID[0]
  PIN top_E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.870 6.990 324.170 ;
    END
  END top_E2MID[1]
  PIN top_E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.230 19.410 325.530 ;
    END
  END top_E2MID[2]
  PIN top_E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.270 9.290 327.570 ;
    END
  END top_E2MID[3]
  PIN top_E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.310 6.990 329.610 ;
    END
  END top_E2MID[4]
  PIN top_E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 330.670 6.530 330.970 ;
    END
  END top_E2MID[5]
  PIN top_E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 332.710 13.890 333.010 ;
    END
  END top_E2MID[6]
  PIN top_E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.070 13.890 334.370 ;
    END
  END top_E2MID[7]
  PIN top_E6BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.410 380.310 223.275 380.610 ;
    END
  END top_E6BEG[0]
  PIN top_E6BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.410 397.990 223.275 398.290 ;
    END
  END top_E6BEG[10]
  PIN top_E6BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 400.030 223.275 400.330 ;
    END
  END top_E6BEG[11]
  PIN top_E6BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.410 382.350 223.275 382.650 ;
    END
  END top_E6BEG[1]
  PIN top_E6BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 383.710 223.275 384.010 ;
    END
  END top_E6BEG[2]
  PIN top_E6BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 212.890 385.750 223.275 386.050 ;
    END
  END top_E6BEG[3]
  PIN top_E6BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.410 387.790 223.275 388.090 ;
    END
  END top_E6BEG[4]
  PIN top_E6BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.210 389.150 223.275 389.450 ;
    END
  END top_E6BEG[5]
  PIN top_E6BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 391.190 223.275 391.490 ;
    END
  END top_E6BEG[6]
  PIN top_E6BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.210 393.230 223.275 393.530 ;
    END
  END top_E6BEG[7]
  PIN top_E6BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.590 394.590 223.275 394.890 ;
    END
  END top_E6BEG[8]
  PIN top_E6BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.130 396.630 223.275 396.930 ;
    END
  END top_E6BEG[9]
  PIN top_E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.950 7.450 379.250 ;
    END
  END top_E6END[0]
  PIN top_E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 396.630 13.890 396.930 ;
    END
  END top_E6END[10]
  PIN top_E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.670 13.890 398.970 ;
    END
  END top_E6END[11]
  PIN top_E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.990 8.830 381.290 ;
    END
  END top_E6END[1]
  PIN top_E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.350 13.890 382.650 ;
    END
  END top_E6END[2]
  PIN top_E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.390 15.730 384.690 ;
    END
  END top_E6END[3]
  PIN top_E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.430 17.570 386.730 ;
    END
  END top_E6END[4]
  PIN top_E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.790 14.350 388.090 ;
    END
  END top_E6END[5]
  PIN top_E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.830 17.110 390.130 ;
    END
  END top_E6END[6]
  PIN top_E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.190 20.330 391.490 ;
    END
  END top_E6END[7]
  PIN top_E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.230 20.330 393.530 ;
    END
  END top_E6END[8]
  PIN top_E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.270 7.280 395.570 ;
    END
  END top_E6END[9]
  PIN top_EE4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 351.750 223.275 352.050 ;
    END
  END top_EE4BEG[0]
  PIN top_EE4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.410 369.430 223.275 369.730 ;
    END
  END top_EE4BEG[10]
  PIN top_EE4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 371.470 223.275 371.770 ;
    END
  END top_EE4BEG[11]
  PIN top_EE4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.410 373.510 223.275 373.810 ;
    END
  END top_EE4BEG[12]
  PIN top_EE4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.870 374.870 223.275 375.170 ;
    END
  END top_EE4BEG[13]
  PIN top_EE4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.210 376.910 223.275 377.210 ;
    END
  END top_EE4BEG[14]
  PIN top_EE4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.130 378.270 223.275 378.570 ;
    END
  END top_EE4BEG[15]
  PIN top_EE4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.410 353.790 223.275 354.090 ;
    END
  END top_EE4BEG[1]
  PIN top_EE4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.350 355.150 223.275 355.450 ;
    END
  END top_EE4BEG[2]
  PIN top_EE4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 357.190 223.275 357.490 ;
    END
  END top_EE4BEG[3]
  PIN top_EE4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 358.550 223.275 358.850 ;
    END
  END top_EE4BEG[4]
  PIN top_EE4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 220.710 360.590 223.275 360.890 ;
    END
  END top_EE4BEG[5]
  PIN top_EE4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 362.630 223.275 362.930 ;
    END
  END top_EE4BEG[6]
  PIN top_EE4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 363.990 223.275 364.290 ;
    END
  END top_EE4BEG[7]
  PIN top_EE4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.210 366.030 223.275 366.330 ;
    END
  END top_EE4BEG[8]
  PIN top_EE4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.130 368.070 223.275 368.370 ;
    END
  END top_EE4BEG[9]
  PIN top_EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.390 6.990 350.690 ;
    END
  END top_EE4END[0]
  PIN top_EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.070 13.890 368.370 ;
    END
  END top_EE4END[10]
  PIN top_EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.110 14.350 370.410 ;
    END
  END top_EE4END[11]
  PIN top_EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.150 13.890 372.450 ;
    END
  END top_EE4END[12]
  PIN top_EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 373.510 17.110 373.810 ;
    END
  END top_EE4END[13]
  PIN top_EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 375.550 14.350 375.850 ;
    END
  END top_EE4END[14]
  PIN top_EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.910 17.110 377.210 ;
    END
  END top_EE4END[15]
  PIN top_EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.430 13.890 352.730 ;
    END
  END top_EE4END[1]
  PIN top_EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.790 9.290 354.090 ;
    END
  END top_EE4END[2]
  PIN top_EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.830 17.110 356.130 ;
    END
  END top_EE4END[3]
  PIN top_EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.870 13.890 358.170 ;
    END
  END top_EE4END[4]
  PIN top_EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.230 17.570 359.530 ;
    END
  END top_EE4END[5]
  PIN top_EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.270 17.110 361.570 ;
    END
  END top_EE4END[6]
  PIN top_EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 362.630 20.330 362.930 ;
    END
  END top_EE4END[7]
  PIN top_EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.670 17.570 364.970 ;
    END
  END top_EE4END[8]
  PIN top_EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 366.710 17.110 367.010 ;
    END
  END top_EE4END[9]
  PIN top_FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 400.710 7.450 401.010 ;
    END
  END top_FrameData[0]
  PIN top_FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.390 6.990 418.690 ;
    END
  END top_FrameData[10]
  PIN top_FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 419.750 7.450 420.050 ;
    END
  END top_FrameData[11]
  PIN top_FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.790 8.830 422.090 ;
    END
  END top_FrameData[12]
  PIN top_FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.830 7.450 424.130 ;
    END
  END top_FrameData[13]
  PIN top_FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.190 6.990 425.490 ;
    END
  END top_FrameData[14]
  PIN top_FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.230 8.830 427.530 ;
    END
  END top_FrameData[15]
  PIN top_FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.270 18.950 429.570 ;
    END
  END top_FrameData[16]
  PIN top_FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 430.630 16.190 430.930 ;
    END
  END top_FrameData[17]
  PIN top_FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 432.670 6.990 432.970 ;
    END
  END top_FrameData[18]
  PIN top_FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 434.030 6.530 434.330 ;
    END
  END top_FrameData[19]
  PIN top_FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 402.070 6.990 402.370 ;
    END
  END top_FrameData[1]
  PIN top_FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.070 7.450 436.370 ;
    END
  END top_FrameData[20]
  PIN top_FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 438.110 8.830 438.410 ;
    END
  END top_FrameData[21]
  PIN top_FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 439.470 18.950 439.770 ;
    END
  END top_FrameData[22]
  PIN top_FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 441.510 18.950 441.810 ;
    END
  END top_FrameData[23]
  PIN top_FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 443.550 8.830 443.850 ;
    END
  END top_FrameData[24]
  PIN top_FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.910 7.450 445.210 ;
    END
  END top_FrameData[25]
  PIN top_FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.950 19.870 447.250 ;
    END
  END top_FrameData[26]
  PIN top_FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.310 8.830 448.610 ;
    END
  END top_FrameData[27]
  PIN top_FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.350 6.990 450.650 ;
    END
  END top_FrameData[28]
  PIN top_FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.390 7.450 452.690 ;
    END
  END top_FrameData[29]
  PIN top_FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.110 6.990 404.410 ;
    END
  END top_FrameData[2]
  PIN top_FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 453.750 16.190 454.050 ;
    END
  END top_FrameData[30]
  PIN top_FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.790 18.950 456.090 ;
    END
  END top_FrameData[31]
  PIN top_FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.470 6.530 405.770 ;
    END
  END top_FrameData[3]
  PIN top_FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 407.510 6.990 407.810 ;
    END
  END top_FrameData[4]
  PIN top_FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 409.550 8.830 409.850 ;
    END
  END top_FrameData[5]
  PIN top_FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.910 14.350 411.210 ;
    END
  END top_FrameData[6]
  PIN top_FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.950 14.350 413.250 ;
    END
  END top_FrameData[7]
  PIN top_FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.990 19.410 415.290 ;
    END
  END top_FrameData[8]
  PIN top_FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.350 19.410 416.650 ;
    END
  END top_FrameData[9]
  PIN top_FrameData_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.410 402.070 223.275 402.370 ;
    END
  END top_FrameData_O[0]
  PIN top_FrameData_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.410 419.750 223.275 420.050 ;
    END
  END top_FrameData_O[10]
  PIN top_FrameData_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.410 421.790 223.275 422.090 ;
    END
  END top_FrameData_O[11]
  PIN top_FrameData_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.410 423.150 223.275 423.450 ;
    END
  END top_FrameData_O[12]
  PIN top_FrameData_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 425.190 223.275 425.490 ;
    END
  END top_FrameData_O[13]
  PIN top_FrameData_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 427.230 223.275 427.530 ;
    END
  END top_FrameData_O[14]
  PIN top_FrameData_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.410 428.590 223.275 428.890 ;
    END
  END top_FrameData_O[15]
  PIN top_FrameData_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.590 430.630 223.275 430.930 ;
    END
  END top_FrameData_O[16]
  PIN top_FrameData_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 432.670 223.275 432.970 ;
    END
  END top_FrameData_O[17]
  PIN top_FrameData_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 434.030 223.275 434.330 ;
    END
  END top_FrameData_O[18]
  PIN top_FrameData_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.590 436.070 223.275 436.370 ;
    END
  END top_FrameData_O[19]
  PIN top_FrameData_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.870 403.430 223.275 403.730 ;
    END
  END top_FrameData_O[1]
  PIN top_FrameData_O[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.410 437.430 223.275 437.730 ;
    END
  END top_FrameData_O[20]
  PIN top_FrameData_O[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 439.470 223.275 439.770 ;
    END
  END top_FrameData_O[21]
  PIN top_FrameData_O[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.590 441.510 223.275 441.810 ;
    END
  END top_FrameData_O[22]
  PIN top_FrameData_O[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 442.870 223.275 443.170 ;
    END
  END top_FrameData_O[23]
  PIN top_FrameData_O[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.130 444.910 223.275 445.210 ;
    END
  END top_FrameData_O[24]
  PIN top_FrameData_O[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 446.950 223.275 447.250 ;
    END
  END top_FrameData_O[25]
  PIN top_FrameData_O[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 205.990 448.310 223.275 448.610 ;
    END
  END top_FrameData_O[26]
  PIN top_FrameData_O[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 204.610 450.350 223.275 450.650 ;
    END
  END top_FrameData_O[27]
  PIN top_FrameData_O[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 200.930 452.390 223.275 452.690 ;
    END
  END top_FrameData_O[28]
  PIN top_FrameData_O[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.850 453.750 223.275 454.050 ;
    END
  END top_FrameData_O[29]
  PIN top_FrameData_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 405.470 223.275 405.770 ;
    END
  END top_FrameData_O[2]
  PIN top_FrameData_O[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.850 455.790 223.275 456.090 ;
    END
  END top_FrameData_O[30]
  PIN top_FrameData_O[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 199.550 457.150 223.275 457.450 ;
    END
  END top_FrameData_O[31]
  PIN top_FrameData_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.410 407.510 223.275 407.810 ;
    END
  END top_FrameData_O[3]
  PIN top_FrameData_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.590 408.870 223.275 409.170 ;
    END
  END top_FrameData_O[4]
  PIN top_FrameData_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 410.910 223.275 411.210 ;
    END
  END top_FrameData_O[5]
  PIN top_FrameData_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.730 412.950 223.275 413.250 ;
    END
  END top_FrameData_O[6]
  PIN top_FrameData_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.590 414.310 223.275 414.610 ;
    END
  END top_FrameData_O[7]
  PIN top_FrameData_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.210 416.350 223.275 416.650 ;
    END
  END top_FrameData_O[8]
  PIN top_FrameData_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.130 417.710 223.275 418.010 ;
    END
  END top_FrameData_O[9]
  PIN top_N1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.080 464.060 1.220 471.230 ;
    END
  END top_N1BEG[0]
  PIN top_N1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.920 467.120 3.060 471.230 ;
    END
  END top_N1BEG[1]
  PIN top_N1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.760 453.520 4.900 471.230 ;
    END
  END top_N1BEG[2]
  PIN top_N1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.600 453.180 6.740 471.230 ;
    END
  END top_N1BEG[3]
  PIN top_N2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.900 455.220 9.040 471.230 ;
    END
  END top_N2BEG[0]
  PIN top_N2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.740 454.880 10.880 471.230 ;
    END
  END top_N2BEG[1]
  PIN top_N2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.580 464.060 12.720 471.230 ;
    END
  END top_N2BEG[2]
  PIN top_N2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.420 460.660 14.560 471.230 ;
    END
  END top_N2BEG[3]
  PIN top_N2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.720 458.620 16.860 471.230 ;
    END
  END top_N2BEG[4]
  PIN top_N2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.560 461.480 18.700 471.230 ;
    END
  END top_N2BEG[5]
  PIN top_N2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.400 470.150 20.540 471.230 ;
    END
  END top_N2BEG[6]
  PIN top_N2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.240 470.150 22.380 471.230 ;
    END
  END top_N2BEG[7]
  PIN top_N2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.540 464.030 24.680 471.230 ;
    END
  END top_N2BEGb[0]
  PIN top_N2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.380 466.780 26.520 471.230 ;
    END
  END top_N2BEGb[1]
  PIN top_N2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.220 461.680 28.360 471.230 ;
    END
  END top_N2BEGb[2]
  PIN top_N2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.060 459.300 30.200 471.230 ;
    END
  END top_N2BEGb[3]
  PIN top_N2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.360 464.400 32.500 471.230 ;
    END
  END top_N2BEGb[4]
  PIN top_N2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.200 460.660 34.340 471.230 ;
    END
  END top_N2BEGb[5]
  PIN top_N2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.040 466.750 36.180 471.230 ;
    END
  END top_N2BEGb[6]
  PIN top_N2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.880 465.390 38.020 471.230 ;
    END
  END top_N2BEGb[7]
  PIN top_N4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.180 466.070 40.320 471.230 ;
    END
  END top_N4BEG[0]
  PIN top_N4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.500 464.740 59.640 471.230 ;
    END
  END top_N4BEG[10]
  PIN top_N4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.340 464.740 61.480 471.230 ;
    END
  END top_N4BEG[11]
  PIN top_N4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.640 461.680 63.780 471.230 ;
    END
  END top_N4BEG[12]
  PIN top_N4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.480 464.740 65.620 471.230 ;
    END
  END top_N4BEG[13]
  PIN top_N4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.320 462.020 67.460 471.230 ;
    END
  END top_N4BEG[14]
  PIN top_N4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.160 464.400 69.300 471.230 ;
    END
  END top_N4BEG[15]
  PIN top_N4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.020 460.320 42.160 471.230 ;
    END
  END top_N4BEG[1]
  PIN top_N4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.860 454.880 44.000 471.230 ;
    END
  END top_N4BEG[2]
  PIN top_N4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.700 456.580 45.840 471.230 ;
    END
  END top_N4BEG[3]
  PIN top_N4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.000 461.310 48.140 471.230 ;
    END
  END top_N4BEG[4]
  PIN top_N4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.840 466.750 49.980 471.230 ;
    END
  END top_N4BEG[5]
  PIN top_N4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.680 462.020 51.820 471.230 ;
    END
  END top_N4BEG[6]
  PIN top_N4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.520 470.150 53.660 471.230 ;
    END
  END top_N4BEG[7]
  PIN top_N4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.820 470.150 55.960 471.230 ;
    END
  END top_N4BEG[8]
  PIN top_N4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.660 462.020 57.800 471.230 ;
    END
  END top_N4BEG[9]
  PIN top_NN4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.460 462.020 71.600 471.230 ;
    END
  END top_NN4BEG[0]
  PIN top_NN4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.780 464.740 90.920 471.230 ;
    END
  END top_NN4BEG[10]
  PIN top_NN4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.620 462.020 92.760 471.230 ;
    END
  END top_NN4BEG[11]
  PIN top_NN4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.920 462.020 95.060 471.230 ;
    END
  END top_NN4BEG[12]
  PIN top_NN4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.760 461.680 96.900 471.230 ;
    END
  END top_NN4BEG[13]
  PIN top_NN4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.600 470.150 98.740 471.230 ;
    END
  END top_NN4BEG[14]
  PIN top_NN4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.440 464.740 100.580 471.230 ;
    END
  END top_NN4BEG[15]
  PIN top_NN4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.300 464.540 73.440 471.230 ;
    END
  END top_NN4BEG[1]
  PIN top_NN4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.140 462.020 75.280 471.230 ;
    END
  END top_NN4BEG[2]
  PIN top_NN4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.980 470.150 77.120 471.230 ;
    END
  END top_NN4BEG[3]
  PIN top_NN4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.280 462.020 79.420 471.230 ;
    END
  END top_NN4BEG[4]
  PIN top_NN4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.120 461.680 81.260 471.230 ;
    END
  END top_NN4BEG[5]
  PIN top_NN4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.960 457.600 83.100 471.230 ;
    END
  END top_NN4BEG[6]
  PIN top_NN4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.800 458.960 84.940 471.230 ;
    END
  END top_NN4BEG[7]
  PIN top_NN4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.100 470.150 87.240 471.230 ;
    END
  END top_NN4BEG[8]
  PIN top_NN4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.940 462.020 89.080 471.230 ;
    END
  END top_NN4BEG[9]
  PIN top_S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.740 463.720 102.880 471.230 ;
    END
  END top_S1END[0]
  PIN top_S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.580 461.340 104.720 471.230 ;
    END
  END top_S1END[1]
  PIN top_S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.420 463.720 106.560 471.230 ;
    END
  END top_S1END[2]
  PIN top_S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.260 464.400 108.400 471.230 ;
    END
  END top_S1END[3]
  PIN top_S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.560 463.720 110.700 471.230 ;
    END
  END top_S2END[0]
  PIN top_S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.400 461.680 112.540 471.230 ;
    END
  END top_S2END[1]
  PIN top_S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.240 458.280 114.380 471.230 ;
    END
  END top_S2END[2]
  PIN top_S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.540 461.680 116.680 471.230 ;
    END
  END top_S2END[3]
  PIN top_S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.380 464.060 118.520 471.230 ;
    END
  END top_S2END[4]
  PIN top_S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.220 462.840 120.360 471.230 ;
    END
  END top_S2END[5]
  PIN top_S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.060 461.340 122.200 471.230 ;
    END
  END top_S2END[6]
  PIN top_S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.360 464.710 124.500 471.230 ;
    END
  END top_S2END[7]
  PIN top_S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.200 461.680 126.340 471.230 ;
    END
  END top_S2MID[0]
  PIN top_S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.040 462.020 128.180 471.230 ;
    END
  END top_S2MID[1]
  PIN top_S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.880 458.280 130.020 471.230 ;
    END
  END top_S2MID[2]
  PIN top_S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.180 458.620 132.320 471.230 ;
    END
  END top_S2MID[3]
  PIN top_S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.020 463.720 134.160 471.230 ;
    END
  END top_S2MID[4]
  PIN top_S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.860 464.060 136.000 471.230 ;
    END
  END top_S2MID[5]
  PIN top_S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.700 463.040 137.840 471.230 ;
    END
  END top_S2MID[6]
  PIN top_S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.000 467.460 140.140 471.230 ;
    END
  END top_S2MID[7]
  PIN top_S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.840 470.150 141.980 471.230 ;
    END
  END top_S4END[0]
  PIN top_S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.160 462.020 161.300 471.230 ;
    END
  END top_S4END[10]
  PIN top_S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.460 459.950 163.600 471.230 ;
    END
  END top_S4END[11]
  PIN top_S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.300 467.430 165.440 471.230 ;
    END
  END top_S4END[12]
  PIN top_S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.140 461.310 167.280 471.230 ;
    END
  END top_S4END[13]
  PIN top_S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.980 455.400 169.120 471.230 ;
    END
  END top_S4END[14]
  PIN top_S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.280 455.220 171.420 471.230 ;
    END
  END top_S4END[15]
  PIN top_S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.680 467.120 143.820 471.230 ;
    END
  END top_S4END[1]
  PIN top_S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.520 467.800 145.660 471.230 ;
    END
  END top_S4END[2]
  PIN top_S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.820 455.220 147.960 471.230 ;
    END
  END top_S4END[3]
  PIN top_S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.660 453.860 149.800 471.230 ;
    END
  END top_S4END[4]
  PIN top_S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.500 442.270 151.640 471.230 ;
    END
  END top_S4END[5]
  PIN top_S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.340 461.990 153.480 471.230 ;
    END
  END top_S4END[6]
  PIN top_S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.640 461.820 155.780 471.230 ;
    END
  END top_S4END[7]
  PIN top_S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.480 453.520 157.620 471.230 ;
    END
  END top_S4END[8]
  PIN top_S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.320 453.660 159.460 471.230 ;
    END
  END top_S4END[9]
  PIN top_SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.120 461.340 173.260 471.230 ;
    END
  END top_SS4END[0]
  PIN top_SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.440 455.220 192.580 471.230 ;
    END
  END top_SS4END[10]
  PIN top_SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.740 459.480 194.880 471.230 ;
    END
  END top_SS4END[11]
  PIN top_SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.580 464.710 196.720 471.230 ;
    END
  END top_SS4END[12]
  PIN top_SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.420 428.700 198.560 471.230 ;
    END
  END top_SS4END[13]
  PIN top_SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.260 463.040 200.400 471.230 ;
    END
  END top_SS4END[14]
  PIN top_SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.560 455.220 202.700 471.230 ;
    END
  END top_SS4END[15]
  PIN top_SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.960 467.430 175.100 471.230 ;
    END
  END top_SS4END[1]
  PIN top_SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.800 461.340 176.940 471.230 ;
    END
  END top_SS4END[2]
  PIN top_SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.100 462.020 179.240 471.230 ;
    END
  END top_SS4END[3]
  PIN top_SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.940 434.140 181.080 471.230 ;
    END
  END top_SS4END[4]
  PIN top_SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.780 466.750 182.920 471.230 ;
    END
  END top_SS4END[5]
  PIN top_SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.620 431.080 184.760 471.230 ;
    END
  END top_SS4END[6]
  PIN top_SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.920 457.910 187.060 471.230 ;
    END
  END top_SS4END[7]
  PIN top_SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.760 459.100 188.900 471.230 ;
    END
  END top_SS4END[8]
  PIN top_SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.600 464.030 190.740 471.230 ;
    END
  END top_SS4END[9]
  PIN top_W1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.350 9.750 229.650 ;
    END
  END top_W1BEG[0]
  PIN top_W1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 230.710 10.210 231.010 ;
    END
  END top_W1BEG[1]
  PIN top_W1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.750 6.990 233.050 ;
    END
  END top_W1BEG[2]
  PIN top_W1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.110 13.890 234.410 ;
    END
  END top_W1BEG[3]
  PIN top_W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.130 230.030 223.275 230.330 ;
    END
  END top_W1END[0]
  PIN top_W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.450 231.390 223.275 231.690 ;
    END
  END top_W1END[1]
  PIN top_W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.130 233.430 223.275 233.730 ;
    END
  END top_W1END[2]
  PIN top_W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.910 235.470 223.275 235.770 ;
    END
  END top_W1END[3]
  PIN top_W2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.150 9.750 236.450 ;
    END
  END top_W2BEG[0]
  PIN top_W2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.190 6.990 238.490 ;
    END
  END top_W2BEG[1]
  PIN top_W2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.550 13.890 239.850 ;
    END
  END top_W2BEG[2]
  PIN top_W2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.590 9.750 241.890 ;
    END
  END top_W2BEG[3]
  PIN top_W2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.630 10.210 243.930 ;
    END
  END top_W2BEG[4]
  PIN top_W2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.990 13.890 245.290 ;
    END
  END top_W2BEG[5]
  PIN top_W2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.030 6.990 247.330 ;
    END
  END top_W2BEG[6]
  PIN top_W2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.390 13.890 248.690 ;
    END
  END top_W2BEG[7]
  PIN top_W2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.430 9.750 250.730 ;
    END
  END top_W2BEGb[0]
  PIN top_W2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 252.470 6.990 252.770 ;
    END
  END top_W2BEGb[1]
  PIN top_W2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.830 13.890 254.130 ;
    END
  END top_W2BEGb[2]
  PIN top_W2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.870 9.750 256.170 ;
    END
  END top_W2BEGb[3]
  PIN top_W2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.910 10.210 258.210 ;
    END
  END top_W2BEGb[4]
  PIN top_W2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.270 13.890 259.570 ;
    END
  END top_W2BEGb[5]
  PIN top_W2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.310 9.750 261.610 ;
    END
  END top_W2BEGb[6]
  PIN top_W2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.670 6.990 262.970 ;
    END
  END top_W2BEGb[7]
  PIN top_W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 205.530 251.110 223.275 251.410 ;
    END
  END top_W2END[0]
  PIN top_W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.910 253.150 223.275 253.450 ;
    END
  END top_W2END[1]
  PIN top_W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 205.070 255.190 223.275 255.490 ;
    END
  END top_W2END[2]
  PIN top_W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 256.550 223.275 256.850 ;
    END
  END top_W2END[3]
  PIN top_W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.910 258.590 223.275 258.890 ;
    END
  END top_W2END[4]
  PIN top_W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 205.530 260.630 223.275 260.930 ;
    END
  END top_W2END[5]
  PIN top_W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 207.830 261.990 223.275 262.290 ;
    END
  END top_W2END[6]
  PIN top_W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 264.030 223.275 264.330 ;
    END
  END top_W2END[7]
  PIN top_W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 207.830 236.830 223.275 237.130 ;
    END
  END top_W2MID[0]
  PIN top_W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 204.610 238.870 223.275 239.170 ;
    END
  END top_W2MID[1]
  PIN top_W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 240.910 223.275 241.210 ;
    END
  END top_W2MID[2]
  PIN top_W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 212.890 242.270 223.275 242.570 ;
    END
  END top_W2MID[3]
  PIN top_W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 202.770 244.310 223.275 244.610 ;
    END
  END top_W2MID[4]
  PIN top_W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 203.690 245.670 223.275 245.970 ;
    END
  END top_W2MID[5]
  PIN top_W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 211.050 247.710 223.275 248.010 ;
    END
  END top_W2MID[6]
  PIN top_W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 205.070 249.750 223.275 250.050 ;
    END
  END top_W2MID[7]
  PIN top_W6BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.270 9.750 293.570 ;
    END
  END top_W6BEG[0]
  PIN top_W6BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.950 10.210 311.250 ;
    END
  END top_W6BEG[10]
  PIN top_W6BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.990 13.890 313.290 ;
    END
  END top_W6BEG[11]
  PIN top_W6BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.310 9.750 295.610 ;
    END
  END top_W6BEG[1]
  PIN top_W6BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.670 6.990 296.970 ;
    END
  END top_W6BEG[2]
  PIN top_W6BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 298.710 9.750 299.010 ;
    END
  END top_W6BEG[3]
  PIN top_W6BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.750 6.990 301.050 ;
    END
  END top_W6BEG[4]
  PIN top_W6BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.110 13.890 302.410 ;
    END
  END top_W6BEG[5]
  PIN top_W6BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.150 9.750 304.450 ;
    END
  END top_W6BEG[6]
  PIN top_W6BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 305.510 13.890 305.810 ;
    END
  END top_W6BEG[7]
  PIN top_W6BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.550 13.890 307.850 ;
    END
  END top_W6BEG[8]
  PIN top_W6BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.590 13.890 309.890 ;
    END
  END top_W6BEG[9]
  PIN top_W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 294.630 223.275 294.930 ;
    END
  END top_W6END[0]
  PIN top_W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 312.310 223.275 312.610 ;
    END
  END top_W6END[10]
  PIN top_W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.130 314.350 223.275 314.650 ;
    END
  END top_W6END[11]
  PIN top_W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 295.990 223.275 296.290 ;
    END
  END top_W6END[1]
  PIN top_W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.910 298.030 223.275 298.330 ;
    END
  END top_W6END[2]
  PIN top_W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 300.070 223.275 300.370 ;
    END
  END top_W6END[3]
  PIN top_W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 205.990 301.430 223.275 301.730 ;
    END
  END top_W6END[4]
  PIN top_W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.910 303.470 223.275 303.770 ;
    END
  END top_W6END[5]
  PIN top_W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 211.510 304.830 223.275 305.130 ;
    END
  END top_W6END[6]
  PIN top_W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.910 306.870 223.275 307.170 ;
    END
  END top_W6END[7]
  PIN top_W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.450 308.910 223.275 309.210 ;
    END
  END top_W6END[8]
  PIN top_W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 205.990 310.270 223.275 310.570 ;
    END
  END top_W6END[9]
  PIN top_WW4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 264.710 13.890 265.010 ;
    END
  END top_WW4BEG[0]
  PIN top_WW4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.390 9.750 282.690 ;
    END
  END top_WW4BEG[10]
  PIN top_WW4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.430 9.750 284.730 ;
    END
  END top_WW4BEG[11]
  PIN top_WW4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 286.470 9.750 286.770 ;
    END
  END top_WW4BEG[12]
  PIN top_WW4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.830 6.990 288.130 ;
    END
  END top_WW4BEG[13]
  PIN top_WW4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.870 13.890 290.170 ;
    END
  END top_WW4BEG[14]
  PIN top_WW4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.230 17.110 291.530 ;
    END
  END top_WW4BEG[15]
  PIN top_WW4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.750 9.750 267.050 ;
    END
  END top_WW4BEG[1]
  PIN top_WW4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.110 6.990 268.410 ;
    END
  END top_WW4BEG[2]
  PIN top_WW4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.150 13.890 270.450 ;
    END
  END top_WW4BEG[3]
  PIN top_WW4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.190 9.750 272.490 ;
    END
  END top_WW4BEG[4]
  PIN top_WW4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.550 7.910 273.850 ;
    END
  END top_WW4BEG[5]
  PIN top_WW4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.590 13.890 275.890 ;
    END
  END top_WW4BEG[6]
  PIN top_WW4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.950 9.750 277.250 ;
    END
  END top_WW4BEG[7]
  PIN top_WW4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.990 13.890 279.290 ;
    END
  END top_WW4BEG[8]
  PIN top_WW4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.030 17.110 281.330 ;
    END
  END top_WW4BEG[9]
  PIN top_WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 212.430 265.390 223.275 265.690 ;
    END
  END top_WW4END[0]
  PIN top_WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 211.970 283.750 223.275 284.050 ;
    END
  END top_WW4END[10]
  PIN top_WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 285.110 223.275 285.410 ;
    END
  END top_WW4END[11]
  PIN top_WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.910 287.150 223.275 287.450 ;
    END
  END top_WW4END[12]
  PIN top_WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.450 289.190 223.275 289.490 ;
    END
  END top_WW4END[13]
  PIN top_WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.910 290.550 223.275 290.850 ;
    END
  END top_WW4END[14]
  PIN top_WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 204.150 292.590 223.275 292.890 ;
    END
  END top_WW4END[15]
  PIN top_WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.850 267.430 223.275 267.730 ;
    END
  END top_WW4END[1]
  PIN top_WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 269.470 223.275 269.770 ;
    END
  END top_WW4END[2]
  PIN top_WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 212.890 270.830 223.275 271.130 ;
    END
  END top_WW4END[3]
  PIN top_WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.670 272.870 223.275 273.170 ;
    END
  END top_WW4END[4]
  PIN top_WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.450 274.910 223.275 275.210 ;
    END
  END top_WW4END[5]
  PIN top_WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 205.530 276.270 223.275 276.570 ;
    END
  END top_WW4END[6]
  PIN top_WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 195.870 278.310 223.275 278.610 ;
    END
  END top_WW4END[7]
  PIN top_WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.790 280.350 223.275 280.650 ;
    END
  END top_WW4END[8]
  PIN top_WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.670 281.710 223.275 282.010 ;
    END
  END top_WW4END[9]
  OBS
      LAYER li1 ;
        RECT 5.520 2.465 222.955 468.095 ;
      LAYER met1 ;
        RECT 0.990 1.400 223.030 468.140 ;
      LAYER met2 ;
        RECT 1.500 466.840 2.640 470.970 ;
        RECT 3.340 466.840 4.480 470.970 ;
        RECT 1.500 463.780 4.480 466.840 ;
        RECT 1.020 453.240 4.480 463.780 ;
        RECT 5.180 453.240 6.320 470.970 ;
        RECT 1.020 452.900 6.320 453.240 ;
        RECT 7.020 454.940 8.620 470.970 ;
        RECT 9.320 454.940 10.460 470.970 ;
        RECT 7.020 454.600 10.460 454.940 ;
        RECT 11.160 463.780 12.300 470.970 ;
        RECT 13.000 463.780 14.140 470.970 ;
        RECT 11.160 460.380 14.140 463.780 ;
        RECT 14.840 460.380 16.440 470.970 ;
        RECT 11.160 458.340 16.440 460.380 ;
        RECT 17.140 461.200 18.280 470.970 ;
        RECT 18.980 469.870 20.120 470.970 ;
        RECT 20.820 469.870 21.960 470.970 ;
        RECT 22.660 469.870 24.260 470.970 ;
        RECT 18.980 463.750 24.260 469.870 ;
        RECT 24.960 466.500 26.100 470.970 ;
        RECT 26.800 466.500 27.940 470.970 ;
        RECT 24.960 463.750 27.940 466.500 ;
        RECT 18.980 461.400 27.940 463.750 ;
        RECT 28.640 461.400 29.780 470.970 ;
        RECT 18.980 461.200 29.780 461.400 ;
        RECT 17.140 459.020 29.780 461.200 ;
        RECT 30.480 464.120 32.080 470.970 ;
        RECT 32.780 464.120 33.920 470.970 ;
        RECT 30.480 460.380 33.920 464.120 ;
        RECT 34.620 466.470 35.760 470.970 ;
        RECT 36.460 466.470 37.600 470.970 ;
        RECT 34.620 465.110 37.600 466.470 ;
        RECT 38.300 465.790 39.900 470.970 ;
        RECT 40.600 465.790 41.740 470.970 ;
        RECT 38.300 465.110 41.740 465.790 ;
        RECT 34.620 460.380 41.740 465.110 ;
        RECT 30.480 460.040 41.740 460.380 ;
        RECT 42.440 460.040 43.580 470.970 ;
        RECT 30.480 459.020 43.580 460.040 ;
        RECT 17.140 458.340 43.580 459.020 ;
        RECT 11.160 454.600 43.580 458.340 ;
        RECT 44.280 456.300 45.420 470.970 ;
        RECT 46.120 461.030 47.720 470.970 ;
        RECT 48.420 466.470 49.560 470.970 ;
        RECT 50.260 466.470 51.400 470.970 ;
        RECT 48.420 461.740 51.400 466.470 ;
        RECT 52.100 469.870 53.240 470.970 ;
        RECT 53.940 469.870 55.540 470.970 ;
        RECT 56.240 469.870 57.380 470.970 ;
        RECT 52.100 461.740 57.380 469.870 ;
        RECT 58.080 464.460 59.220 470.970 ;
        RECT 59.920 464.460 61.060 470.970 ;
        RECT 61.760 464.460 63.360 470.970 ;
        RECT 58.080 461.740 63.360 464.460 ;
        RECT 48.420 461.400 63.360 461.740 ;
        RECT 64.060 464.460 65.200 470.970 ;
        RECT 65.900 464.460 67.040 470.970 ;
        RECT 64.060 461.740 67.040 464.460 ;
        RECT 67.740 464.120 68.880 470.970 ;
        RECT 69.580 464.120 71.180 470.970 ;
        RECT 67.740 461.740 71.180 464.120 ;
        RECT 71.880 464.260 73.020 470.970 ;
        RECT 73.720 464.260 74.860 470.970 ;
        RECT 71.880 461.740 74.860 464.260 ;
        RECT 75.560 469.870 76.700 470.970 ;
        RECT 77.400 469.870 79.000 470.970 ;
        RECT 75.560 461.740 79.000 469.870 ;
        RECT 79.700 461.740 80.840 470.970 ;
        RECT 64.060 461.400 80.840 461.740 ;
        RECT 81.540 461.400 82.680 470.970 ;
        RECT 48.420 461.030 82.680 461.400 ;
        RECT 46.120 457.320 82.680 461.030 ;
        RECT 83.380 458.680 84.520 470.970 ;
        RECT 85.220 469.870 86.820 470.970 ;
        RECT 87.520 469.870 88.660 470.970 ;
        RECT 85.220 461.740 88.660 469.870 ;
        RECT 89.360 464.460 90.500 470.970 ;
        RECT 91.200 464.460 92.340 470.970 ;
        RECT 89.360 461.740 92.340 464.460 ;
        RECT 93.040 461.740 94.640 470.970 ;
        RECT 95.340 461.740 96.480 470.970 ;
        RECT 85.220 461.400 96.480 461.740 ;
        RECT 97.180 469.870 98.320 470.970 ;
        RECT 99.020 469.870 100.160 470.970 ;
        RECT 97.180 464.460 100.160 469.870 ;
        RECT 100.860 464.460 102.460 470.970 ;
        RECT 97.180 463.440 102.460 464.460 ;
        RECT 103.160 463.440 104.300 470.970 ;
        RECT 97.180 461.400 104.300 463.440 ;
        RECT 85.220 461.060 104.300 461.400 ;
        RECT 105.000 463.440 106.140 470.970 ;
        RECT 106.840 464.120 107.980 470.970 ;
        RECT 108.680 464.120 110.280 470.970 ;
        RECT 106.840 463.440 110.280 464.120 ;
        RECT 110.980 463.440 112.120 470.970 ;
        RECT 105.000 461.400 112.120 463.440 ;
        RECT 112.820 461.400 113.960 470.970 ;
        RECT 105.000 461.060 113.960 461.400 ;
        RECT 85.220 458.680 113.960 461.060 ;
        RECT 83.380 458.000 113.960 458.680 ;
        RECT 114.660 461.400 116.260 470.970 ;
        RECT 116.960 463.780 118.100 470.970 ;
        RECT 118.800 463.780 119.940 470.970 ;
        RECT 116.960 462.560 119.940 463.780 ;
        RECT 120.640 462.560 121.780 470.970 ;
        RECT 116.960 461.400 121.780 462.560 ;
        RECT 114.660 461.060 121.780 461.400 ;
        RECT 122.480 464.430 124.080 470.970 ;
        RECT 124.780 464.430 125.920 470.970 ;
        RECT 122.480 461.400 125.920 464.430 ;
        RECT 126.620 461.740 127.760 470.970 ;
        RECT 128.460 461.740 129.600 470.970 ;
        RECT 126.620 461.400 129.600 461.740 ;
        RECT 122.480 461.060 129.600 461.400 ;
        RECT 114.660 458.000 129.600 461.060 ;
        RECT 130.300 458.340 131.900 470.970 ;
        RECT 132.600 463.440 133.740 470.970 ;
        RECT 134.440 463.780 135.580 470.970 ;
        RECT 136.280 463.780 137.420 470.970 ;
        RECT 134.440 463.440 137.420 463.780 ;
        RECT 132.600 462.760 137.420 463.440 ;
        RECT 138.120 467.180 139.720 470.970 ;
        RECT 140.420 469.870 141.560 470.970 ;
        RECT 142.260 469.870 143.400 470.970 ;
        RECT 140.420 467.180 143.400 469.870 ;
        RECT 138.120 466.840 143.400 467.180 ;
        RECT 144.100 467.520 145.240 470.970 ;
        RECT 145.940 467.520 147.540 470.970 ;
        RECT 144.100 466.840 147.540 467.520 ;
        RECT 138.120 462.760 147.540 466.840 ;
        RECT 132.600 458.340 147.540 462.760 ;
        RECT 130.300 458.000 147.540 458.340 ;
        RECT 83.380 457.320 147.540 458.000 ;
        RECT 46.120 456.300 147.540 457.320 ;
        RECT 44.280 454.940 147.540 456.300 ;
        RECT 148.240 454.940 149.380 470.970 ;
        RECT 44.280 454.600 149.380 454.940 ;
        RECT 7.020 453.580 149.380 454.600 ;
        RECT 150.080 453.580 151.220 470.970 ;
        RECT 7.020 452.900 151.220 453.580 ;
        RECT 1.020 441.990 151.220 452.900 ;
        RECT 151.920 461.710 153.060 470.970 ;
        RECT 153.760 461.710 155.360 470.970 ;
        RECT 151.920 461.540 155.360 461.710 ;
        RECT 156.060 461.540 157.200 470.970 ;
        RECT 151.920 453.240 157.200 461.540 ;
        RECT 157.900 453.380 159.040 470.970 ;
        RECT 159.740 461.740 160.880 470.970 ;
        RECT 161.580 461.740 163.180 470.970 ;
        RECT 159.740 459.670 163.180 461.740 ;
        RECT 163.880 467.150 165.020 470.970 ;
        RECT 165.720 467.150 166.860 470.970 ;
        RECT 163.880 461.030 166.860 467.150 ;
        RECT 167.560 461.030 168.700 470.970 ;
        RECT 163.880 459.670 168.700 461.030 ;
        RECT 159.740 455.120 168.700 459.670 ;
        RECT 169.400 455.120 171.000 470.970 ;
        RECT 159.740 454.940 171.000 455.120 ;
        RECT 171.700 461.060 172.840 470.970 ;
        RECT 173.540 467.150 174.680 470.970 ;
        RECT 175.380 467.150 176.520 470.970 ;
        RECT 173.540 461.060 176.520 467.150 ;
        RECT 177.220 461.740 178.820 470.970 ;
        RECT 179.520 461.740 180.660 470.970 ;
        RECT 177.220 461.060 180.660 461.740 ;
        RECT 171.700 454.940 180.660 461.060 ;
        RECT 159.740 453.380 180.660 454.940 ;
        RECT 157.900 453.240 180.660 453.380 ;
        RECT 151.920 441.990 180.660 453.240 ;
        RECT 1.020 433.860 180.660 441.990 ;
        RECT 181.360 466.470 182.500 470.970 ;
        RECT 183.200 466.470 184.340 470.970 ;
        RECT 181.360 433.860 184.340 466.470 ;
        RECT 1.020 430.800 184.340 433.860 ;
        RECT 185.040 457.630 186.640 470.970 ;
        RECT 187.340 458.820 188.480 470.970 ;
        RECT 189.180 463.750 190.320 470.970 ;
        RECT 191.020 463.750 192.160 470.970 ;
        RECT 189.180 458.820 192.160 463.750 ;
        RECT 187.340 457.630 192.160 458.820 ;
        RECT 185.040 454.940 192.160 457.630 ;
        RECT 192.860 459.200 194.460 470.970 ;
        RECT 195.160 464.430 196.300 470.970 ;
        RECT 197.000 464.430 198.140 470.970 ;
        RECT 195.160 459.200 198.140 464.430 ;
        RECT 192.860 454.940 198.140 459.200 ;
        RECT 185.040 430.800 198.140 454.940 ;
        RECT 1.020 428.420 198.140 430.800 ;
        RECT 198.840 462.760 199.980 470.970 ;
        RECT 200.680 462.760 202.280 470.970 ;
        RECT 198.840 454.940 202.280 462.760 ;
        RECT 202.980 463.440 204.120 470.970 ;
        RECT 204.820 463.440 205.960 470.970 ;
        RECT 202.980 454.940 205.960 463.440 ;
        RECT 198.840 452.560 205.960 454.940 ;
        RECT 206.660 458.000 207.800 470.970 ;
        RECT 208.500 461.060 210.100 470.970 ;
        RECT 210.800 461.060 211.940 470.970 ;
        RECT 208.500 458.000 211.940 461.060 ;
        RECT 206.660 452.560 211.940 458.000 ;
        RECT 198.840 428.420 211.940 452.560 ;
        RECT 1.020 425.700 211.940 428.420 ;
        RECT 212.640 465.110 213.780 470.970 ;
        RECT 214.480 465.110 215.620 470.970 ;
        RECT 212.640 456.300 215.620 465.110 ;
        RECT 216.320 461.740 217.920 470.970 ;
        RECT 218.620 461.740 219.760 470.970 ;
        RECT 216.320 458.680 219.760 461.740 ;
        RECT 220.460 458.680 221.600 470.970 ;
        RECT 216.320 456.300 221.600 458.680 ;
        RECT 212.640 425.700 221.600 456.300 ;
        RECT 1.020 424.680 221.600 425.700 ;
        RECT 222.300 424.680 223.000 470.970 ;
        RECT 1.020 42.480 223.000 424.680 ;
        RECT 1.020 31.600 80.380 42.480 ;
        RECT 1.020 16.980 50.940 31.600 ;
        RECT 1.020 15.280 47.260 16.980 ;
        RECT 1.020 12.220 6.320 15.280 ;
        RECT 1.020 6.780 2.640 12.220 ;
        RECT 1.500 0.270 2.640 6.780 ;
        RECT 3.340 9.840 6.320 12.220 ;
        RECT 3.340 0.270 4.480 9.840 ;
        RECT 5.180 0.270 6.320 9.840 ;
        RECT 7.020 12.220 13.680 15.280 ;
        RECT 7.020 0.270 8.160 12.220 ;
        RECT 8.860 9.840 13.680 12.220 ;
        RECT 8.860 4.060 11.840 9.840 ;
        RECT 8.860 0.270 10.000 4.060 ;
        RECT 10.700 0.270 11.840 4.060 ;
        RECT 12.540 0.270 13.680 9.840 ;
        RECT 14.380 12.220 30.240 15.280 ;
        RECT 14.380 1.370 19.200 12.220 ;
        RECT 14.380 0.270 15.520 1.370 ;
        RECT 16.220 0.270 17.360 1.370 ;
        RECT 18.060 0.270 19.200 1.370 ;
        RECT 19.900 9.500 30.240 12.220 ;
        RECT 19.900 7.120 26.560 9.500 ;
        RECT 19.900 0.270 21.040 7.120 ;
        RECT 21.740 6.780 26.560 7.120 ;
        RECT 21.740 6.440 24.720 6.780 ;
        RECT 21.740 0.270 22.880 6.440 ;
        RECT 23.580 0.270 24.720 6.440 ;
        RECT 25.420 0.270 26.560 6.780 ;
        RECT 27.260 6.440 30.240 9.500 ;
        RECT 27.260 0.270 28.400 6.440 ;
        RECT 29.100 0.270 30.240 6.440 ;
        RECT 30.940 14.800 47.260 15.280 ;
        RECT 30.940 12.220 45.420 14.800 ;
        RECT 30.940 9.840 33.920 12.220 ;
        RECT 30.940 0.270 32.080 9.840 ;
        RECT 32.780 0.270 33.920 9.840 ;
        RECT 34.620 6.440 37.600 12.220 ;
        RECT 34.620 0.270 35.760 6.440 ;
        RECT 36.460 0.270 37.600 6.440 ;
        RECT 38.300 10.040 45.420 12.220 ;
        RECT 38.300 9.840 41.280 10.040 ;
        RECT 38.300 0.270 39.440 9.840 ;
        RECT 40.140 0.270 41.280 9.840 ;
        RECT 41.980 6.440 45.420 10.040 ;
        RECT 41.980 0.270 43.120 6.440 ;
        RECT 43.820 0.270 45.420 6.440 ;
        RECT 46.120 0.270 47.260 14.800 ;
        RECT 47.960 14.970 50.940 16.980 ;
        RECT 47.960 0.270 49.100 14.970 ;
        RECT 49.800 0.270 50.940 14.970 ;
        RECT 51.640 23.130 80.380 31.600 ;
        RECT 51.640 16.980 74.860 23.130 ;
        RECT 51.640 0.270 52.780 16.980 ;
        RECT 53.480 14.150 74.860 16.980 ;
        RECT 53.480 9.840 65.660 14.150 ;
        RECT 53.480 5.450 56.460 9.840 ;
        RECT 53.480 0.270 54.620 5.450 ;
        RECT 55.320 0.270 56.460 5.450 ;
        RECT 57.160 9.500 65.660 9.840 ;
        RECT 57.160 1.370 60.140 9.500 ;
        RECT 57.160 0.270 58.300 1.370 ;
        RECT 59.000 0.270 60.140 1.370 ;
        RECT 60.840 7.800 65.660 9.500 ;
        RECT 60.840 7.120 63.820 7.800 ;
        RECT 60.840 0.270 61.980 7.120 ;
        RECT 62.680 0.270 63.820 7.120 ;
        RECT 64.520 0.270 65.660 7.800 ;
        RECT 66.360 6.780 74.860 14.150 ;
        RECT 66.360 0.270 67.500 6.780 ;
        RECT 68.200 6.440 73.020 6.780 ;
        RECT 68.200 6.100 71.180 6.440 ;
        RECT 68.200 0.270 69.340 6.100 ;
        RECT 70.040 0.270 71.180 6.100 ;
        RECT 71.880 0.270 73.020 6.440 ;
        RECT 73.720 0.270 74.860 6.780 ;
        RECT 75.560 14.150 80.380 23.130 ;
        RECT 75.560 0.270 76.700 14.150 ;
        RECT 77.400 7.490 80.380 14.150 ;
        RECT 77.400 0.270 78.540 7.490 ;
        RECT 79.240 0.270 80.380 7.490 ;
        RECT 81.080 39.420 223.000 42.480 ;
        RECT 81.080 25.820 90.040 39.420 ;
        RECT 81.080 14.760 85.900 25.820 ;
        RECT 81.080 0.270 82.220 14.760 ;
        RECT 82.920 6.300 85.900 14.760 ;
        RECT 82.920 0.270 84.060 6.300 ;
        RECT 84.760 0.270 85.900 6.300 ;
        RECT 86.600 1.370 90.040 25.820 ;
        RECT 86.600 0.270 87.740 1.370 ;
        RECT 88.440 0.270 90.040 1.370 ;
        RECT 90.740 37.040 223.000 39.420 ;
        RECT 90.740 19.700 203.200 37.040 ;
        RECT 90.740 13.100 95.560 19.700 ;
        RECT 90.740 0.270 91.880 13.100 ;
        RECT 92.580 1.370 95.560 13.100 ;
        RECT 92.580 0.270 93.720 1.370 ;
        RECT 94.420 0.270 95.560 1.370 ;
        RECT 96.260 17.660 203.200 19.700 ;
        RECT 96.260 16.980 199.520 17.660 ;
        RECT 96.260 16.120 179.280 16.980 ;
        RECT 96.260 14.260 113.960 16.120 ;
        RECT 96.260 8.820 108.440 14.260 ;
        RECT 96.260 3.410 102.920 8.820 ;
        RECT 96.260 1.680 99.240 3.410 ;
        RECT 96.260 0.270 97.400 1.680 ;
        RECT 98.100 0.270 99.240 1.680 ;
        RECT 99.940 1.370 102.920 3.410 ;
        RECT 99.940 0.270 101.080 1.370 ;
        RECT 101.780 0.270 102.920 1.370 ;
        RECT 103.620 4.740 108.440 8.820 ;
        RECT 103.620 2.360 106.600 4.740 ;
        RECT 103.620 0.270 104.760 2.360 ;
        RECT 105.460 0.270 106.600 2.360 ;
        RECT 107.300 0.270 108.440 4.740 ;
        RECT 109.140 14.080 113.960 14.260 ;
        RECT 109.140 0.270 110.280 14.080 ;
        RECT 110.980 4.060 113.960 14.080 ;
        RECT 110.980 0.270 112.120 4.060 ;
        RECT 112.820 0.270 113.960 4.060 ;
        RECT 114.660 14.600 179.280 16.120 ;
        RECT 114.660 14.260 176.980 14.600 ;
        RECT 114.660 14.080 117.640 14.260 ;
        RECT 114.660 0.270 115.800 14.080 ;
        RECT 116.500 0.270 117.640 14.080 ;
        RECT 118.340 12.220 165.940 14.260 ;
        RECT 118.340 11.540 151.220 12.220 ;
        RECT 118.340 9.160 142.020 11.540 ;
        RECT 118.340 8.820 130.520 9.160 ;
        RECT 118.340 6.780 123.160 8.820 ;
        RECT 118.340 6.100 121.320 6.780 ;
        RECT 118.340 0.270 119.480 6.100 ;
        RECT 120.180 0.270 121.320 6.100 ;
        RECT 122.020 0.270 123.160 6.780 ;
        RECT 123.860 6.100 126.840 8.820 ;
        RECT 123.860 0.270 125.000 6.100 ;
        RECT 125.700 0.270 126.840 6.100 ;
        RECT 127.540 3.380 130.520 8.820 ;
        RECT 127.540 0.270 128.680 3.380 ;
        RECT 129.380 0.270 130.520 3.380 ;
        RECT 131.220 8.820 138.340 9.160 ;
        RECT 131.220 6.780 134.660 8.820 ;
        RECT 131.220 0.270 132.360 6.780 ;
        RECT 133.060 0.270 134.660 6.780 ;
        RECT 135.360 7.120 138.340 8.820 ;
        RECT 135.360 0.270 136.500 7.120 ;
        RECT 137.200 0.270 138.340 7.120 ;
        RECT 139.040 1.370 142.020 9.160 ;
        RECT 139.040 0.270 140.180 1.370 ;
        RECT 140.880 0.270 142.020 1.370 ;
        RECT 142.720 7.490 151.220 11.540 ;
        RECT 142.720 0.270 143.860 7.490 ;
        RECT 144.560 7.120 151.220 7.490 ;
        RECT 144.560 4.740 147.540 7.120 ;
        RECT 144.560 0.270 145.700 4.740 ;
        RECT 146.400 0.270 147.540 4.740 ;
        RECT 148.240 3.380 151.220 7.120 ;
        RECT 148.240 0.270 149.380 3.380 ;
        RECT 150.080 0.270 151.220 3.380 ;
        RECT 151.920 9.160 165.940 12.220 ;
        RECT 151.920 8.820 162.260 9.160 ;
        RECT 151.920 6.100 154.900 8.820 ;
        RECT 151.920 0.270 153.060 6.100 ;
        RECT 153.760 0.270 154.900 6.100 ;
        RECT 155.600 6.100 158.580 8.820 ;
        RECT 155.600 0.270 156.740 6.100 ;
        RECT 157.440 0.270 158.580 6.100 ;
        RECT 159.280 6.440 162.260 8.820 ;
        RECT 159.280 0.270 160.420 6.440 ;
        RECT 161.120 0.270 162.260 6.440 ;
        RECT 162.960 8.820 165.940 9.160 ;
        RECT 162.960 0.270 164.100 8.820 ;
        RECT 164.800 0.270 165.940 8.820 ;
        RECT 166.640 9.160 171.460 14.260 ;
        RECT 166.640 1.370 169.620 9.160 ;
        RECT 166.640 0.270 167.780 1.370 ;
        RECT 168.480 0.270 169.620 1.370 ;
        RECT 170.320 0.270 171.460 9.160 ;
        RECT 172.160 12.560 176.980 14.260 ;
        RECT 172.160 0.270 173.300 12.560 ;
        RECT 174.000 1.370 176.980 12.560 ;
        RECT 174.000 0.270 175.140 1.370 ;
        RECT 175.840 0.270 176.980 1.370 ;
        RECT 177.680 0.270 179.280 14.600 ;
        RECT 179.980 0.270 181.120 16.980 ;
        RECT 181.820 15.280 199.520 16.980 ;
        RECT 181.820 14.260 197.680 15.280 ;
        RECT 181.820 9.160 188.480 14.260 ;
        RECT 181.820 6.100 184.800 9.160 ;
        RECT 181.820 0.270 182.960 6.100 ;
        RECT 183.660 0.270 184.800 6.100 ;
        RECT 185.500 6.440 188.480 9.160 ;
        RECT 185.500 0.270 186.640 6.440 ;
        RECT 187.340 0.270 188.480 6.440 ;
        RECT 189.180 9.840 197.680 14.260 ;
        RECT 189.180 8.820 194.000 9.840 ;
        RECT 189.180 6.130 192.160 8.820 ;
        RECT 189.180 0.270 190.320 6.130 ;
        RECT 191.020 0.270 192.160 6.130 ;
        RECT 192.860 0.270 194.000 8.820 ;
        RECT 194.700 6.780 197.680 9.840 ;
        RECT 194.700 0.270 195.840 6.780 ;
        RECT 196.540 0.270 197.680 6.780 ;
        RECT 198.380 0.270 199.520 15.280 ;
        RECT 200.220 12.220 203.200 17.660 ;
        RECT 200.220 0.270 201.360 12.220 ;
        RECT 202.060 0.270 203.200 12.220 ;
        RECT 203.900 25.480 223.000 37.040 ;
        RECT 203.900 20.040 216.080 25.480 ;
        RECT 203.900 18.680 214.240 20.040 ;
        RECT 203.900 17.690 210.560 18.680 ;
        RECT 203.900 1.370 206.880 17.690 ;
        RECT 203.900 0.270 205.040 1.370 ;
        RECT 205.740 0.270 206.880 1.370 ;
        RECT 207.580 14.940 210.560 17.690 ;
        RECT 207.580 0.270 208.720 14.940 ;
        RECT 209.420 0.270 210.560 14.940 ;
        RECT 211.260 6.100 214.240 18.680 ;
        RECT 211.260 0.270 212.400 6.100 ;
        RECT 213.100 0.270 214.240 6.100 ;
        RECT 214.940 0.270 216.080 20.040 ;
        RECT 216.780 14.600 223.000 25.480 ;
        RECT 216.780 9.160 219.760 14.600 ;
        RECT 216.780 0.270 217.920 9.160 ;
        RECT 218.620 0.270 219.760 9.160 ;
        RECT 220.460 14.260 223.000 14.600 ;
        RECT 220.460 0.270 221.600 14.260 ;
        RECT 222.300 0.270 223.000 14.260 ;
      LAYER met3 ;
        RECT 17.510 469.670 200.990 470.385 ;
        RECT 1.905 468.730 222.115 469.670 ;
        RECT 16.130 467.630 218.470 468.730 ;
        RECT 1.905 467.370 222.115 467.630 ;
        RECT 20.730 466.270 214.330 467.370 ;
        RECT 1.905 465.330 222.115 466.270 ;
        RECT 19.810 464.230 213.870 465.330 ;
        RECT 1.905 463.290 222.115 464.230 ;
        RECT 14.290 462.190 200.530 463.290 ;
        RECT 1.905 461.930 222.115 462.190 ;
        RECT 7.850 460.830 218.010 461.930 ;
        RECT 1.905 459.890 222.115 460.830 ;
        RECT 7.390 458.790 203.290 459.890 ;
        RECT 1.905 458.530 222.115 458.790 ;
        RECT 7.390 457.850 222.115 458.530 ;
        RECT 7.390 457.430 199.150 457.850 ;
        RECT 1.905 456.750 199.150 457.430 ;
        RECT 1.905 456.490 222.115 456.750 ;
        RECT 19.350 455.390 201.450 456.490 ;
        RECT 1.905 454.450 222.115 455.390 ;
        RECT 16.590 453.350 201.450 454.450 ;
        RECT 1.905 453.090 222.115 453.350 ;
        RECT 7.850 451.990 200.530 453.090 ;
        RECT 1.905 451.050 222.115 451.990 ;
        RECT 7.390 449.950 204.210 451.050 ;
        RECT 1.905 449.010 222.115 449.950 ;
        RECT 9.230 447.910 205.590 449.010 ;
        RECT 1.905 447.650 222.115 447.910 ;
        RECT 20.270 446.550 209.270 447.650 ;
        RECT 1.905 445.610 222.115 446.550 ;
        RECT 7.850 444.510 209.730 445.610 ;
        RECT 1.905 444.250 222.115 444.510 ;
        RECT 9.230 443.570 222.115 444.250 ;
        RECT 9.230 443.150 213.870 443.570 ;
        RECT 1.905 442.470 213.870 443.150 ;
        RECT 1.905 442.210 222.115 442.470 ;
        RECT 19.350 441.110 210.190 442.210 ;
        RECT 1.905 440.170 222.115 441.110 ;
        RECT 19.350 439.070 213.410 440.170 ;
        RECT 1.905 438.810 222.115 439.070 ;
        RECT 9.230 438.130 222.115 438.810 ;
        RECT 9.230 437.710 218.010 438.130 ;
        RECT 1.905 437.030 218.010 437.710 ;
        RECT 1.905 436.770 222.115 437.030 ;
        RECT 7.850 435.670 210.190 436.770 ;
        RECT 1.905 434.730 222.115 435.670 ;
        RECT 6.930 433.630 213.870 434.730 ;
        RECT 1.905 433.370 222.115 433.630 ;
        RECT 7.390 432.270 213.410 433.370 ;
        RECT 1.905 431.330 222.115 432.270 ;
        RECT 16.590 430.230 210.190 431.330 ;
        RECT 1.905 429.970 222.115 430.230 ;
        RECT 19.350 429.290 222.115 429.970 ;
        RECT 19.350 428.870 218.010 429.290 ;
        RECT 1.905 428.190 218.010 428.870 ;
        RECT 1.905 427.930 222.115 428.190 ;
        RECT 9.230 426.830 213.870 427.930 ;
        RECT 1.905 425.890 222.115 426.830 ;
        RECT 7.390 424.790 213.410 425.890 ;
        RECT 1.905 424.530 222.115 424.790 ;
        RECT 7.850 423.850 222.115 424.530 ;
        RECT 7.850 423.430 218.010 423.850 ;
        RECT 1.905 422.750 218.010 423.430 ;
        RECT 1.905 422.490 222.115 422.750 ;
        RECT 9.230 421.390 218.010 422.490 ;
        RECT 1.905 420.450 222.115 421.390 ;
        RECT 7.850 419.350 218.010 420.450 ;
        RECT 1.905 419.090 222.115 419.350 ;
        RECT 7.390 418.410 222.115 419.090 ;
        RECT 7.390 417.990 209.730 418.410 ;
        RECT 1.905 417.310 209.730 417.990 ;
        RECT 1.905 417.050 222.115 417.310 ;
        RECT 19.810 415.950 208.810 417.050 ;
        RECT 1.905 415.690 222.115 415.950 ;
        RECT 19.810 415.010 222.115 415.690 ;
        RECT 19.810 414.590 210.190 415.010 ;
        RECT 1.905 413.910 210.190 414.590 ;
        RECT 1.905 413.650 222.115 413.910 ;
        RECT 14.750 412.550 214.330 413.650 ;
        RECT 1.905 411.610 222.115 412.550 ;
        RECT 14.750 410.510 213.410 411.610 ;
        RECT 1.905 410.250 222.115 410.510 ;
        RECT 9.230 409.570 222.115 410.250 ;
        RECT 9.230 409.150 210.190 409.570 ;
        RECT 1.905 408.470 210.190 409.150 ;
        RECT 1.905 408.210 222.115 408.470 ;
        RECT 7.390 407.110 218.010 408.210 ;
        RECT 1.905 406.170 222.115 407.110 ;
        RECT 6.930 405.070 213.410 406.170 ;
        RECT 1.905 404.810 222.115 405.070 ;
        RECT 7.390 404.130 222.115 404.810 ;
        RECT 7.390 403.710 218.470 404.130 ;
        RECT 1.905 403.030 218.470 403.710 ;
        RECT 1.905 402.770 222.115 403.030 ;
        RECT 7.390 401.670 218.010 402.770 ;
        RECT 1.905 401.410 222.115 401.670 ;
        RECT 7.850 400.730 222.115 401.410 ;
        RECT 7.850 400.310 213.410 400.730 ;
        RECT 1.905 399.630 213.410 400.310 ;
        RECT 1.905 399.370 222.115 399.630 ;
        RECT 14.290 398.690 222.115 399.370 ;
        RECT 14.290 398.270 218.010 398.690 ;
        RECT 1.905 397.590 218.010 398.270 ;
        RECT 1.905 397.330 222.115 397.590 ;
        RECT 14.290 396.230 209.730 397.330 ;
        RECT 1.905 395.970 222.115 396.230 ;
        RECT 7.680 395.290 222.115 395.970 ;
        RECT 7.680 394.870 210.190 395.290 ;
        RECT 1.905 394.190 210.190 394.870 ;
        RECT 1.905 393.930 222.115 394.190 ;
        RECT 20.730 392.830 208.810 393.930 ;
        RECT 1.905 391.890 222.115 392.830 ;
        RECT 20.730 390.790 213.410 391.890 ;
        RECT 1.905 390.530 222.115 390.790 ;
        RECT 17.510 389.850 222.115 390.530 ;
        RECT 17.510 389.430 208.810 389.850 ;
        RECT 1.905 388.750 208.810 389.430 ;
        RECT 1.905 388.490 222.115 388.750 ;
        RECT 14.750 387.390 218.010 388.490 ;
        RECT 1.905 387.130 222.115 387.390 ;
        RECT 17.970 386.450 222.115 387.130 ;
        RECT 17.970 386.030 212.490 386.450 ;
        RECT 1.905 385.350 212.490 386.030 ;
        RECT 1.905 385.090 222.115 385.350 ;
        RECT 16.130 384.410 222.115 385.090 ;
        RECT 16.130 383.990 213.410 384.410 ;
        RECT 1.905 383.310 213.410 383.990 ;
        RECT 1.905 383.050 222.115 383.310 ;
        RECT 14.290 381.950 218.010 383.050 ;
        RECT 1.905 381.690 222.115 381.950 ;
        RECT 9.230 381.010 222.115 381.690 ;
        RECT 9.230 380.590 218.010 381.010 ;
        RECT 1.905 379.910 218.010 380.590 ;
        RECT 1.905 379.650 222.115 379.910 ;
        RECT 7.850 378.970 222.115 379.650 ;
        RECT 7.850 378.550 209.730 378.970 ;
        RECT 1.905 377.870 209.730 378.550 ;
        RECT 1.905 377.610 222.115 377.870 ;
        RECT 17.510 376.510 208.810 377.610 ;
        RECT 1.905 376.250 222.115 376.510 ;
        RECT 14.750 375.570 222.115 376.250 ;
        RECT 14.750 375.150 218.470 375.570 ;
        RECT 1.905 374.470 218.470 375.150 ;
        RECT 1.905 374.210 222.115 374.470 ;
        RECT 17.510 373.110 218.010 374.210 ;
        RECT 1.905 372.850 222.115 373.110 ;
        RECT 14.290 372.170 222.115 372.850 ;
        RECT 14.290 371.750 213.410 372.170 ;
        RECT 1.905 371.070 213.410 371.750 ;
        RECT 1.905 370.810 222.115 371.070 ;
        RECT 14.750 370.130 222.115 370.810 ;
        RECT 14.750 369.710 218.010 370.130 ;
        RECT 1.905 369.030 218.010 369.710 ;
        RECT 1.905 368.770 222.115 369.030 ;
        RECT 14.290 367.670 209.730 368.770 ;
        RECT 1.905 367.410 222.115 367.670 ;
        RECT 17.510 366.730 222.115 367.410 ;
        RECT 17.510 366.310 208.810 366.730 ;
        RECT 1.905 365.630 208.810 366.310 ;
        RECT 1.905 365.370 222.115 365.630 ;
        RECT 17.970 364.690 222.115 365.370 ;
        RECT 17.970 364.270 213.410 364.690 ;
        RECT 1.905 363.590 213.410 364.270 ;
        RECT 1.905 363.330 222.115 363.590 ;
        RECT 20.730 362.230 209.270 363.330 ;
        RECT 1.905 361.970 222.115 362.230 ;
        RECT 17.510 361.290 222.115 361.970 ;
        RECT 17.510 360.870 220.310 361.290 ;
        RECT 1.905 360.190 220.310 360.870 ;
        RECT 1.905 359.930 222.115 360.190 ;
        RECT 17.970 359.250 222.115 359.930 ;
        RECT 17.970 358.830 213.410 359.250 ;
        RECT 1.905 358.570 213.410 358.830 ;
        RECT 14.290 358.150 213.410 358.570 ;
        RECT 14.290 357.890 222.115 358.150 ;
        RECT 14.290 357.470 209.270 357.890 ;
        RECT 1.905 356.790 209.270 357.470 ;
        RECT 1.905 356.530 222.115 356.790 ;
        RECT 17.510 355.850 222.115 356.530 ;
        RECT 17.510 355.430 212.950 355.850 ;
        RECT 1.905 354.750 212.950 355.430 ;
        RECT 1.905 354.490 222.115 354.750 ;
        RECT 9.690 353.390 218.010 354.490 ;
        RECT 1.905 353.130 222.115 353.390 ;
        RECT 14.290 352.450 222.115 353.130 ;
        RECT 14.290 352.030 209.270 352.450 ;
        RECT 1.905 351.350 209.270 352.030 ;
        RECT 1.905 351.090 222.115 351.350 ;
        RECT 7.390 350.410 222.115 351.090 ;
        RECT 7.390 349.990 213.410 350.410 ;
        RECT 1.905 349.310 213.410 349.990 ;
        RECT 1.905 349.050 222.115 349.310 ;
        RECT 9.690 347.950 220.310 349.050 ;
        RECT 1.905 347.690 222.115 347.950 ;
        RECT 7.390 347.010 222.115 347.690 ;
        RECT 7.390 346.590 209.270 347.010 ;
        RECT 1.905 345.910 209.270 346.590 ;
        RECT 1.905 345.650 222.115 345.910 ;
        RECT 9.690 344.970 222.115 345.650 ;
        RECT 9.690 344.550 212.950 344.970 ;
        RECT 1.905 344.290 212.950 344.550 ;
        RECT 11.990 343.870 212.950 344.290 ;
        RECT 11.990 343.610 222.115 343.870 ;
        RECT 11.990 343.190 213.410 343.610 ;
        RECT 1.905 342.510 213.410 343.190 ;
        RECT 1.905 342.250 222.115 342.510 ;
        RECT 6.930 341.570 222.115 342.250 ;
        RECT 6.930 341.150 209.270 341.570 ;
        RECT 1.905 340.470 209.270 341.150 ;
        RECT 1.905 340.210 222.115 340.470 ;
        RECT 7.390 339.110 218.010 340.210 ;
        RECT 1.905 338.850 222.115 339.110 ;
        RECT 11.990 338.170 222.115 338.850 ;
        RECT 11.990 337.750 221.690 338.170 ;
        RECT 1.905 337.070 221.690 337.750 ;
        RECT 1.905 336.810 222.115 337.070 ;
        RECT 7.390 336.130 222.115 336.810 ;
        RECT 7.390 335.710 209.270 336.130 ;
        RECT 1.905 335.030 209.270 335.710 ;
        RECT 1.905 334.770 222.115 335.030 ;
        RECT 14.290 333.670 213.410 334.770 ;
        RECT 1.905 333.410 222.115 333.670 ;
        RECT 14.290 332.730 222.115 333.410 ;
        RECT 14.290 332.310 218.010 332.730 ;
        RECT 1.905 331.630 218.010 332.310 ;
        RECT 1.905 331.370 222.115 331.630 ;
        RECT 6.930 330.690 222.115 331.370 ;
        RECT 6.930 330.270 209.270 330.690 ;
        RECT 1.905 330.010 209.270 330.270 ;
        RECT 7.390 329.590 209.270 330.010 ;
        RECT 7.390 329.330 222.115 329.590 ;
        RECT 7.390 328.910 213.410 329.330 ;
        RECT 1.905 328.230 213.410 328.910 ;
        RECT 1.905 327.970 222.115 328.230 ;
        RECT 9.690 327.290 222.115 327.970 ;
        RECT 9.690 326.870 218.010 327.290 ;
        RECT 1.905 326.190 218.010 326.870 ;
        RECT 1.905 325.930 222.115 326.190 ;
        RECT 19.810 325.250 222.115 325.930 ;
        RECT 19.810 324.830 209.270 325.250 ;
        RECT 1.905 324.570 209.270 324.830 ;
        RECT 7.390 324.150 209.270 324.570 ;
        RECT 7.390 323.890 222.115 324.150 ;
        RECT 7.390 323.470 213.410 323.890 ;
        RECT 1.905 322.790 213.410 323.470 ;
        RECT 1.905 322.530 222.115 322.790 ;
        RECT 9.230 321.850 222.115 322.530 ;
        RECT 9.230 321.430 209.730 321.850 ;
        RECT 1.905 320.750 209.730 321.430 ;
        RECT 1.905 320.490 222.115 320.750 ;
        RECT 6.930 319.390 219.850 320.490 ;
        RECT 1.905 319.130 222.115 319.390 ;
        RECT 7.390 318.450 222.115 319.130 ;
        RECT 7.390 318.030 218.470 318.450 ;
        RECT 1.905 317.350 218.470 318.030 ;
        RECT 1.905 317.090 222.115 317.350 ;
        RECT 9.230 316.410 222.115 317.090 ;
        RECT 9.230 315.990 213.410 316.410 ;
        RECT 1.905 315.730 213.410 315.990 ;
        RECT 7.850 315.310 213.410 315.730 ;
        RECT 7.850 315.050 222.115 315.310 ;
        RECT 7.850 314.630 209.730 315.050 ;
        RECT 1.905 313.950 209.730 314.630 ;
        RECT 1.905 313.690 222.115 313.950 ;
        RECT 14.290 313.010 222.115 313.690 ;
        RECT 14.290 312.590 209.270 313.010 ;
        RECT 1.905 311.910 209.270 312.590 ;
        RECT 1.905 311.650 222.115 311.910 ;
        RECT 10.610 310.970 222.115 311.650 ;
        RECT 10.610 310.550 205.590 310.970 ;
        RECT 1.905 310.290 205.590 310.550 ;
        RECT 14.290 309.870 205.590 310.290 ;
        RECT 14.290 309.610 222.115 309.870 ;
        RECT 14.290 309.190 206.050 309.610 ;
        RECT 1.905 308.510 206.050 309.190 ;
        RECT 1.905 308.250 222.115 308.510 ;
        RECT 14.290 307.570 222.115 308.250 ;
        RECT 14.290 307.150 206.510 307.570 ;
        RECT 1.905 306.470 206.510 307.150 ;
        RECT 1.905 306.210 222.115 306.470 ;
        RECT 14.290 305.530 222.115 306.210 ;
        RECT 14.290 305.110 211.110 305.530 ;
        RECT 1.905 304.850 211.110 305.110 ;
        RECT 10.150 304.430 211.110 304.850 ;
        RECT 10.150 304.170 222.115 304.430 ;
        RECT 10.150 303.750 206.510 304.170 ;
        RECT 1.905 303.070 206.510 303.750 ;
        RECT 1.905 302.810 222.115 303.070 ;
        RECT 14.290 302.130 222.115 302.810 ;
        RECT 14.290 301.710 205.590 302.130 ;
        RECT 1.905 301.450 205.590 301.710 ;
        RECT 7.390 301.030 205.590 301.450 ;
        RECT 7.390 300.770 222.115 301.030 ;
        RECT 7.390 300.350 213.410 300.770 ;
        RECT 1.905 299.670 213.410 300.350 ;
        RECT 1.905 299.410 222.115 299.670 ;
        RECT 10.150 298.730 222.115 299.410 ;
        RECT 10.150 298.310 206.510 298.730 ;
        RECT 1.905 297.630 206.510 298.310 ;
        RECT 1.905 297.370 222.115 297.630 ;
        RECT 7.390 296.690 222.115 297.370 ;
        RECT 7.390 296.270 209.270 296.690 ;
        RECT 1.905 296.010 209.270 296.270 ;
        RECT 10.150 295.590 209.270 296.010 ;
        RECT 10.150 295.330 222.115 295.590 ;
        RECT 10.150 294.910 209.270 295.330 ;
        RECT 1.905 294.230 209.270 294.910 ;
        RECT 1.905 293.970 222.115 294.230 ;
        RECT 10.150 293.290 222.115 293.970 ;
        RECT 10.150 292.870 203.750 293.290 ;
        RECT 1.905 292.190 203.750 292.870 ;
        RECT 1.905 291.930 222.115 292.190 ;
        RECT 17.510 291.250 222.115 291.930 ;
        RECT 17.510 290.830 206.510 291.250 ;
        RECT 1.905 290.570 206.510 290.830 ;
        RECT 14.290 290.150 206.510 290.570 ;
        RECT 14.290 289.890 222.115 290.150 ;
        RECT 14.290 289.470 206.050 289.890 ;
        RECT 1.905 288.790 206.050 289.470 ;
        RECT 1.905 288.530 222.115 288.790 ;
        RECT 7.390 287.850 222.115 288.530 ;
        RECT 7.390 287.430 206.510 287.850 ;
        RECT 1.905 287.170 206.510 287.430 ;
        RECT 10.150 286.750 206.510 287.170 ;
        RECT 10.150 286.070 222.115 286.750 ;
        RECT 1.905 285.810 222.115 286.070 ;
        RECT 1.905 285.130 209.270 285.810 ;
        RECT 10.150 284.710 209.270 285.130 ;
        RECT 10.150 284.450 222.115 284.710 ;
        RECT 10.150 284.030 211.570 284.450 ;
        RECT 1.905 283.350 211.570 284.030 ;
        RECT 1.905 283.090 222.115 283.350 ;
        RECT 10.150 282.410 222.115 283.090 ;
        RECT 10.150 281.990 214.270 282.410 ;
        RECT 1.905 281.730 214.270 281.990 ;
        RECT 17.510 281.310 214.270 281.730 ;
        RECT 17.510 281.050 222.115 281.310 ;
        RECT 17.510 280.630 196.390 281.050 ;
        RECT 1.905 279.950 196.390 280.630 ;
        RECT 1.905 279.690 222.115 279.950 ;
        RECT 14.290 279.010 222.115 279.690 ;
        RECT 14.290 278.590 195.470 279.010 ;
        RECT 1.905 277.910 195.470 278.590 ;
        RECT 1.905 277.650 222.115 277.910 ;
        RECT 10.150 276.970 222.115 277.650 ;
        RECT 10.150 276.550 205.130 276.970 ;
        RECT 1.905 276.290 205.130 276.550 ;
        RECT 14.290 275.870 205.130 276.290 ;
        RECT 14.290 275.610 222.115 275.870 ;
        RECT 14.290 275.190 206.050 275.610 ;
        RECT 1.905 274.510 206.050 275.190 ;
        RECT 1.905 274.250 222.115 274.510 ;
        RECT 8.310 273.570 222.115 274.250 ;
        RECT 8.310 273.150 214.270 273.570 ;
        RECT 1.905 272.890 214.270 273.150 ;
        RECT 10.150 272.470 214.270 272.890 ;
        RECT 10.150 271.790 222.115 272.470 ;
        RECT 1.905 271.530 222.115 271.790 ;
        RECT 1.905 270.850 212.490 271.530 ;
        RECT 14.290 270.430 212.490 270.850 ;
        RECT 14.290 270.170 222.115 270.430 ;
        RECT 14.290 269.750 209.270 270.170 ;
        RECT 1.905 269.070 209.270 269.750 ;
        RECT 1.905 268.810 222.115 269.070 ;
        RECT 7.390 268.130 222.115 268.810 ;
        RECT 7.390 267.710 206.450 268.130 ;
        RECT 1.905 267.450 206.450 267.710 ;
        RECT 10.150 267.030 206.450 267.450 ;
        RECT 10.150 266.350 222.115 267.030 ;
        RECT 1.905 266.090 222.115 266.350 ;
        RECT 1.905 265.410 212.030 266.090 ;
        RECT 14.290 264.990 212.030 265.410 ;
        RECT 14.290 264.730 222.115 264.990 ;
        RECT 14.290 264.310 209.270 264.730 ;
        RECT 1.905 263.630 209.270 264.310 ;
        RECT 1.905 263.370 222.115 263.630 ;
        RECT 7.390 262.690 222.115 263.370 ;
        RECT 7.390 262.270 207.430 262.690 ;
        RECT 1.905 262.010 207.430 262.270 ;
        RECT 10.150 261.590 207.430 262.010 ;
        RECT 10.150 261.330 222.115 261.590 ;
        RECT 10.150 260.910 205.130 261.330 ;
        RECT 1.905 260.230 205.130 260.910 ;
        RECT 1.905 259.970 222.115 260.230 ;
        RECT 14.290 259.290 222.115 259.970 ;
        RECT 14.290 258.870 206.510 259.290 ;
        RECT 1.905 258.610 206.510 258.870 ;
        RECT 10.610 258.190 206.510 258.610 ;
        RECT 10.610 257.510 222.115 258.190 ;
        RECT 1.905 257.250 222.115 257.510 ;
        RECT 1.905 256.570 209.270 257.250 ;
        RECT 10.150 256.150 209.270 256.570 ;
        RECT 10.150 255.890 222.115 256.150 ;
        RECT 10.150 255.470 204.670 255.890 ;
        RECT 1.905 254.790 204.670 255.470 ;
        RECT 1.905 254.530 222.115 254.790 ;
        RECT 14.290 253.850 222.115 254.530 ;
        RECT 14.290 253.430 206.510 253.850 ;
        RECT 1.905 253.170 206.510 253.430 ;
        RECT 7.390 252.750 206.510 253.170 ;
        RECT 7.390 252.070 222.115 252.750 ;
        RECT 1.905 251.810 222.115 252.070 ;
        RECT 1.905 251.130 205.130 251.810 ;
        RECT 10.150 250.710 205.130 251.130 ;
        RECT 10.150 250.450 222.115 250.710 ;
        RECT 10.150 250.030 204.670 250.450 ;
        RECT 1.905 249.350 204.670 250.030 ;
        RECT 1.905 249.090 222.115 249.350 ;
        RECT 14.290 248.410 222.115 249.090 ;
        RECT 14.290 247.990 210.650 248.410 ;
        RECT 1.905 247.730 210.650 247.990 ;
        RECT 7.390 247.310 210.650 247.730 ;
        RECT 7.390 246.630 222.115 247.310 ;
        RECT 1.905 246.370 222.115 246.630 ;
        RECT 1.905 245.690 203.290 246.370 ;
        RECT 14.290 245.270 203.290 245.690 ;
        RECT 14.290 245.010 222.115 245.270 ;
        RECT 14.290 244.590 202.370 245.010 ;
        RECT 1.905 244.330 202.370 244.590 ;
        RECT 10.610 243.910 202.370 244.330 ;
        RECT 10.610 243.230 222.115 243.910 ;
        RECT 1.905 242.970 222.115 243.230 ;
        RECT 1.905 242.290 212.490 242.970 ;
        RECT 10.150 241.870 212.490 242.290 ;
        RECT 10.150 241.610 222.115 241.870 ;
        RECT 10.150 241.190 209.270 241.610 ;
        RECT 1.905 240.510 209.270 241.190 ;
        RECT 1.905 240.250 222.115 240.510 ;
        RECT 14.290 239.570 222.115 240.250 ;
        RECT 14.290 239.150 204.210 239.570 ;
        RECT 1.905 238.890 204.210 239.150 ;
        RECT 7.390 238.470 204.210 238.890 ;
        RECT 7.390 237.790 222.115 238.470 ;
        RECT 1.905 237.530 222.115 237.790 ;
        RECT 1.905 236.850 207.430 237.530 ;
        RECT 10.150 236.430 207.430 236.850 ;
        RECT 10.150 236.170 222.115 236.430 ;
        RECT 10.150 235.750 206.510 236.170 ;
        RECT 1.905 235.070 206.510 235.750 ;
        RECT 1.905 234.810 222.115 235.070 ;
        RECT 14.290 234.130 222.115 234.810 ;
        RECT 14.290 233.710 209.730 234.130 ;
        RECT 1.905 233.450 209.730 233.710 ;
        RECT 7.390 233.030 209.730 233.450 ;
        RECT 7.390 232.350 222.115 233.030 ;
        RECT 1.905 232.090 222.115 232.350 ;
        RECT 1.905 231.410 206.050 232.090 ;
        RECT 10.610 230.990 206.050 231.410 ;
        RECT 10.610 230.730 222.115 230.990 ;
        RECT 10.610 230.310 209.730 230.730 ;
        RECT 1.905 230.050 209.730 230.310 ;
        RECT 10.150 229.630 209.730 230.050 ;
        RECT 10.150 228.950 222.115 229.630 ;
        RECT 1.905 228.690 222.115 228.950 ;
        RECT 1.905 228.010 218.010 228.690 ;
        RECT 6.930 227.590 218.010 228.010 ;
        RECT 6.930 227.330 222.115 227.590 ;
        RECT 6.930 226.910 213.410 227.330 ;
        RECT 1.905 226.230 213.410 226.910 ;
        RECT 1.905 225.970 222.115 226.230 ;
        RECT 7.390 225.290 222.115 225.970 ;
        RECT 7.390 224.870 208.810 225.290 ;
        RECT 1.905 224.610 208.810 224.870 ;
        RECT 9.230 224.190 208.810 224.610 ;
        RECT 9.230 223.510 222.115 224.190 ;
        RECT 1.905 223.250 222.115 223.510 ;
        RECT 1.905 222.570 209.730 223.250 ;
        RECT 7.850 222.150 209.730 222.570 ;
        RECT 7.850 221.890 222.115 222.150 ;
        RECT 7.850 221.470 218.010 221.890 ;
        RECT 1.905 220.790 218.010 221.470 ;
        RECT 1.905 220.530 222.115 220.790 ;
        RECT 6.930 219.850 222.115 220.530 ;
        RECT 6.930 219.430 213.870 219.850 ;
        RECT 1.905 219.170 213.870 219.430 ;
        RECT 7.390 218.750 213.870 219.170 ;
        RECT 7.390 218.070 222.115 218.750 ;
        RECT 1.905 217.810 222.115 218.070 ;
        RECT 1.905 217.130 213.410 217.810 ;
        RECT 20.730 216.710 213.410 217.130 ;
        RECT 20.730 216.450 222.115 216.710 ;
        RECT 20.730 216.030 209.270 216.450 ;
        RECT 1.905 215.770 209.270 216.030 ;
        RECT 19.810 215.350 209.270 215.770 ;
        RECT 19.810 214.670 222.115 215.350 ;
        RECT 1.905 214.410 222.115 214.670 ;
        RECT 1.905 213.730 213.870 214.410 ;
        RECT 17.050 213.310 213.870 213.730 ;
        RECT 17.050 212.630 222.115 213.310 ;
        RECT 1.905 212.370 222.115 212.630 ;
        RECT 1.905 211.690 213.410 212.370 ;
        RECT 14.750 211.270 213.410 211.690 ;
        RECT 14.750 211.010 222.115 211.270 ;
        RECT 14.750 210.590 209.270 211.010 ;
        RECT 1.905 210.330 209.270 210.590 ;
        RECT 7.390 209.910 209.270 210.330 ;
        RECT 7.390 209.230 222.115 209.910 ;
        RECT 1.905 208.970 222.115 209.230 ;
        RECT 1.905 208.290 218.010 208.970 ;
        RECT 7.850 207.870 218.010 208.290 ;
        RECT 7.850 207.610 222.115 207.870 ;
        RECT 7.850 207.190 213.870 207.610 ;
        RECT 1.905 206.510 213.870 207.190 ;
        RECT 1.905 206.250 222.115 206.510 ;
        RECT 6.930 205.570 222.115 206.250 ;
        RECT 6.930 205.150 209.270 205.570 ;
        RECT 1.905 204.890 209.270 205.150 ;
        RECT 14.750 204.470 209.270 204.890 ;
        RECT 14.750 203.790 222.115 204.470 ;
        RECT 1.905 203.530 222.115 203.790 ;
        RECT 1.905 202.850 213.410 203.530 ;
        RECT 7.850 202.430 213.410 202.850 ;
        RECT 7.850 202.170 222.115 202.430 ;
        RECT 7.850 201.750 209.730 202.170 ;
        RECT 1.905 201.490 209.730 201.750 ;
        RECT 7.390 201.070 209.730 201.490 ;
        RECT 7.390 200.390 222.115 201.070 ;
        RECT 1.905 200.130 222.115 200.390 ;
        RECT 1.905 199.450 213.870 200.130 ;
        RECT 7.390 199.030 213.870 199.450 ;
        RECT 7.390 198.350 222.115 199.030 ;
        RECT 1.905 198.090 222.115 198.350 ;
        RECT 1.905 197.410 213.410 198.090 ;
        RECT 9.230 196.990 213.410 197.410 ;
        RECT 9.230 196.730 222.115 196.990 ;
        RECT 9.230 196.310 218.010 196.730 ;
        RECT 1.905 196.050 218.010 196.310 ;
        RECT 7.850 195.630 218.010 196.050 ;
        RECT 7.850 194.950 222.115 195.630 ;
        RECT 1.905 194.690 222.115 194.950 ;
        RECT 1.905 194.010 213.870 194.690 ;
        RECT 14.290 193.590 213.870 194.010 ;
        RECT 14.290 192.910 222.115 193.590 ;
        RECT 1.905 192.650 222.115 192.910 ;
        RECT 1.905 191.970 213.410 192.650 ;
        RECT 20.270 191.550 213.410 191.970 ;
        RECT 20.270 191.290 222.115 191.550 ;
        RECT 20.270 190.870 213.870 191.290 ;
        RECT 1.905 190.610 213.870 190.870 ;
        RECT 16.590 190.190 213.870 190.610 ;
        RECT 16.590 189.510 222.115 190.190 ;
        RECT 1.905 189.250 222.115 189.510 ;
        RECT 1.905 188.570 209.730 189.250 ;
        RECT 17.970 188.150 209.730 188.570 ;
        RECT 17.970 187.890 222.115 188.150 ;
        RECT 17.970 187.470 208.810 187.890 ;
        RECT 1.905 187.210 208.810 187.470 ;
        RECT 19.350 186.790 208.810 187.210 ;
        RECT 19.350 186.110 222.115 186.790 ;
        RECT 1.905 185.850 222.115 186.110 ;
        RECT 1.905 185.170 213.410 185.850 ;
        RECT 7.850 184.750 213.410 185.170 ;
        RECT 7.850 184.070 222.115 184.750 ;
        RECT 1.905 183.810 222.115 184.070 ;
        RECT 1.905 183.130 209.270 183.810 ;
        RECT 9.230 182.710 209.270 183.130 ;
        RECT 9.230 182.450 222.115 182.710 ;
        RECT 9.230 182.030 218.010 182.450 ;
        RECT 1.905 181.770 218.010 182.030 ;
        RECT 7.390 181.350 218.010 181.770 ;
        RECT 7.390 180.670 222.115 181.350 ;
        RECT 1.905 180.410 222.115 180.670 ;
        RECT 1.905 179.730 213.870 180.410 ;
        RECT 19.350 179.310 213.870 179.730 ;
        RECT 19.350 178.630 222.115 179.310 ;
        RECT 1.905 178.370 222.115 178.630 ;
        RECT 1.905 177.690 209.270 178.370 ;
        RECT 7.850 177.270 209.270 177.690 ;
        RECT 7.850 177.010 222.115 177.270 ;
        RECT 7.850 176.590 213.410 177.010 ;
        RECT 1.905 176.330 213.410 176.590 ;
        RECT 9.230 175.910 213.410 176.330 ;
        RECT 9.230 175.230 222.115 175.910 ;
        RECT 1.905 174.970 222.115 175.230 ;
        RECT 1.905 174.290 213.870 174.970 ;
        RECT 7.850 173.870 213.870 174.290 ;
        RECT 7.850 173.190 222.115 173.870 ;
        RECT 1.905 172.930 222.115 173.190 ;
        RECT 9.230 171.830 213.410 172.930 ;
        RECT 1.905 171.570 222.115 171.830 ;
        RECT 1.905 170.890 213.410 171.570 ;
        RECT 20.730 170.470 213.410 170.890 ;
        RECT 20.730 169.790 222.115 170.470 ;
        RECT 1.905 169.530 222.115 169.790 ;
        RECT 1.905 168.850 213.870 169.530 ;
        RECT 14.290 168.430 213.870 168.850 ;
        RECT 14.290 168.170 222.115 168.430 ;
        RECT 14.290 167.750 209.730 168.170 ;
        RECT 1.905 167.490 209.730 167.750 ;
        RECT 20.730 167.070 209.730 167.490 ;
        RECT 20.730 166.390 222.115 167.070 ;
        RECT 1.905 166.130 222.115 166.390 ;
        RECT 1.905 165.450 208.810 166.130 ;
        RECT 17.510 165.030 208.810 165.450 ;
        RECT 17.510 164.350 222.115 165.030 ;
        RECT 1.905 164.090 222.115 164.350 ;
        RECT 1.905 163.410 209.730 164.090 ;
        RECT 17.970 162.990 209.730 163.410 ;
        RECT 17.970 162.730 222.115 162.990 ;
        RECT 17.970 162.310 213.410 162.730 ;
        RECT 1.905 162.050 213.410 162.310 ;
        RECT 20.730 161.630 213.410 162.050 ;
        RECT 20.730 160.950 222.115 161.630 ;
        RECT 1.905 160.690 222.115 160.950 ;
        RECT 1.905 160.010 218.010 160.690 ;
        RECT 17.510 159.590 218.010 160.010 ;
        RECT 17.510 158.910 222.115 159.590 ;
        RECT 1.905 158.650 222.115 158.910 ;
        RECT 14.290 157.550 213.870 158.650 ;
        RECT 1.905 157.290 222.115 157.550 ;
        RECT 1.905 156.610 216.630 157.290 ;
        RECT 15.210 156.190 216.630 156.610 ;
        RECT 15.210 155.510 222.115 156.190 ;
        RECT 1.905 155.250 222.115 155.510 ;
        RECT 1.905 154.570 213.870 155.250 ;
        RECT 20.270 154.150 213.870 154.570 ;
        RECT 20.270 153.470 222.115 154.150 ;
        RECT 1.905 153.210 222.115 153.470 ;
        RECT 9.230 152.110 216.630 153.210 ;
        RECT 1.905 151.850 222.115 152.110 ;
        RECT 1.905 151.170 213.410 151.850 ;
        RECT 9.230 150.750 213.410 151.170 ;
        RECT 9.230 150.070 222.115 150.750 ;
        RECT 1.905 149.810 222.115 150.070 ;
        RECT 1.905 149.130 208.810 149.810 ;
        RECT 20.270 148.710 208.810 149.130 ;
        RECT 20.270 148.450 222.115 148.710 ;
        RECT 20.270 148.030 210.190 148.450 ;
        RECT 1.905 147.770 210.190 148.030 ;
        RECT 17.050 147.350 210.190 147.770 ;
        RECT 17.050 146.670 222.115 147.350 ;
        RECT 1.905 146.410 222.115 146.670 ;
        RECT 1.905 145.730 213.870 146.410 ;
        RECT 17.510 145.310 213.870 145.730 ;
        RECT 17.510 144.630 222.115 145.310 ;
        RECT 1.905 144.370 222.115 144.630 ;
        RECT 14.750 143.270 213.410 144.370 ;
        RECT 1.905 143.010 222.115 143.270 ;
        RECT 1.905 142.330 215.710 143.010 ;
        RECT 14.290 141.910 215.710 142.330 ;
        RECT 14.290 141.230 222.115 141.910 ;
        RECT 1.905 140.970 222.115 141.230 ;
        RECT 1.905 140.290 213.870 140.970 ;
        RECT 14.290 139.870 213.870 140.290 ;
        RECT 14.290 139.190 222.115 139.870 ;
        RECT 1.905 138.930 222.115 139.190 ;
        RECT 17.510 137.830 208.810 138.930 ;
        RECT 1.905 137.570 222.115 137.830 ;
        RECT 1.905 136.890 208.810 137.570 ;
        RECT 18.430 136.470 208.810 136.890 ;
        RECT 18.430 135.790 222.115 136.470 ;
        RECT 1.905 135.530 222.115 135.790 ;
        RECT 1.905 134.850 209.730 135.530 ;
        RECT 20.730 134.430 209.730 134.850 ;
        RECT 20.730 133.750 222.115 134.430 ;
        RECT 1.905 133.490 222.115 133.750 ;
        RECT 17.510 132.390 213.870 133.490 ;
        RECT 1.905 132.130 222.115 132.390 ;
        RECT 1.905 131.450 210.190 132.130 ;
        RECT 20.730 131.030 210.190 131.450 ;
        RECT 20.730 130.350 222.115 131.030 ;
        RECT 1.905 130.090 222.115 130.350 ;
        RECT 14.290 128.990 213.870 130.090 ;
        RECT 1.905 128.730 222.115 128.990 ;
        RECT 1.905 128.050 213.410 128.730 ;
        RECT 17.510 127.630 213.410 128.050 ;
        RECT 17.510 126.950 222.115 127.630 ;
        RECT 1.905 126.690 222.115 126.950 ;
        RECT 1.905 126.010 210.190 126.690 ;
        RECT 9.690 125.590 210.190 126.010 ;
        RECT 9.690 124.910 222.115 125.590 ;
        RECT 1.905 124.650 222.115 124.910 ;
        RECT 7.390 123.550 213.870 124.650 ;
        RECT 1.905 123.290 222.115 123.550 ;
        RECT 1.905 122.610 213.410 123.290 ;
        RECT 9.690 122.190 213.410 122.610 ;
        RECT 9.690 121.510 222.115 122.190 ;
        RECT 1.905 121.250 222.115 121.510 ;
        RECT 1.905 120.570 210.190 121.250 ;
        RECT 9.690 120.150 210.190 120.570 ;
        RECT 9.690 119.470 222.115 120.150 ;
        RECT 1.905 119.210 222.115 119.470 ;
        RECT 7.390 118.110 220.310 119.210 ;
        RECT 1.905 117.850 222.115 118.110 ;
        RECT 1.905 117.170 213.870 117.850 ;
        RECT 14.290 116.750 213.870 117.170 ;
        RECT 14.290 116.070 222.115 116.750 ;
        RECT 1.905 115.810 222.115 116.070 ;
        RECT 7.450 114.710 210.190 115.810 ;
        RECT 1.905 114.450 222.115 114.710 ;
        RECT 1.905 113.770 213.410 114.450 ;
        RECT 9.230 113.350 213.410 113.770 ;
        RECT 9.230 112.670 222.115 113.350 ;
        RECT 1.905 112.410 222.115 112.670 ;
        RECT 1.905 111.730 213.870 112.410 ;
        RECT 7.390 111.310 213.870 111.730 ;
        RECT 7.390 110.630 222.115 111.310 ;
        RECT 1.905 110.370 222.115 110.630 ;
        RECT 9.230 109.270 210.190 110.370 ;
        RECT 1.905 109.010 222.115 109.270 ;
        RECT 1.905 108.330 213.410 109.010 ;
        RECT 9.690 107.910 213.410 108.330 ;
        RECT 9.690 107.230 222.115 107.910 ;
        RECT 1.905 106.970 222.115 107.230 ;
        RECT 1.905 106.290 213.870 106.970 ;
        RECT 14.290 105.870 213.870 106.290 ;
        RECT 14.290 105.190 222.115 105.870 ;
        RECT 1.905 104.930 222.115 105.190 ;
        RECT 9.230 103.830 210.190 104.930 ;
        RECT 1.905 103.570 222.115 103.830 ;
        RECT 1.905 102.890 213.870 103.570 ;
        RECT 19.810 102.470 213.870 102.890 ;
        RECT 19.810 101.790 222.115 102.470 ;
        RECT 1.905 101.530 222.115 101.790 ;
        RECT 14.290 100.430 213.410 101.530 ;
        RECT 1.905 99.490 222.115 100.430 ;
        RECT 12.450 98.390 210.190 99.490 ;
        RECT 1.905 98.130 222.115 98.390 ;
        RECT 1.905 97.450 213.870 98.130 ;
        RECT 9.690 97.030 213.870 97.450 ;
        RECT 9.690 96.350 222.115 97.030 ;
        RECT 1.905 96.090 222.115 96.350 ;
        RECT 6.470 94.990 208.810 96.090 ;
        RECT 1.905 94.730 222.115 94.990 ;
        RECT 1.905 94.050 213.410 94.730 ;
        RECT 7.390 93.630 213.410 94.050 ;
        RECT 7.390 92.950 222.115 93.630 ;
        RECT 1.905 92.690 222.115 92.950 ;
        RECT 1.905 92.010 213.870 92.690 ;
        RECT 7.850 91.590 213.870 92.010 ;
        RECT 7.850 90.910 222.115 91.590 ;
        RECT 1.905 90.650 222.115 90.910 ;
        RECT 7.390 89.550 208.810 90.650 ;
        RECT 1.905 89.290 222.115 89.550 ;
        RECT 1.905 88.610 213.870 89.290 ;
        RECT 7.390 88.190 213.870 88.610 ;
        RECT 7.390 87.510 222.115 88.190 ;
        RECT 1.905 87.250 222.115 87.510 ;
        RECT 9.230 86.150 213.410 87.250 ;
        RECT 1.905 85.210 222.115 86.150 ;
        RECT 17.050 84.110 209.730 85.210 ;
        RECT 1.905 83.850 222.115 84.110 ;
        RECT 1.905 83.170 209.270 83.850 ;
        RECT 10.610 82.750 209.270 83.170 ;
        RECT 10.610 82.070 222.115 82.750 ;
        RECT 1.905 81.810 222.115 82.070 ;
        RECT 14.290 80.710 203.290 81.810 ;
        RECT 1.905 79.770 222.115 80.710 ;
        RECT 14.290 78.670 206.510 79.770 ;
        RECT 1.905 78.410 222.115 78.670 ;
        RECT 1.905 77.730 205.590 78.410 ;
        RECT 14.290 77.310 205.590 77.730 ;
        RECT 14.290 76.630 222.115 77.310 ;
        RECT 1.905 76.370 222.115 76.630 ;
        RECT 10.150 75.270 206.510 76.370 ;
        RECT 1.905 75.010 222.115 75.270 ;
        RECT 1.905 74.330 214.270 75.010 ;
        RECT 14.290 73.910 214.270 74.330 ;
        RECT 14.290 73.230 222.115 73.910 ;
        RECT 1.905 72.970 222.115 73.230 ;
        RECT 7.390 71.870 216.110 72.970 ;
        RECT 1.905 70.930 222.115 71.870 ;
        RECT 10.150 69.830 209.730 70.930 ;
        RECT 1.905 69.570 222.115 69.830 ;
        RECT 1.905 68.890 209.270 69.570 ;
        RECT 7.390 68.470 209.270 68.890 ;
        RECT 7.390 67.790 222.115 68.470 ;
        RECT 1.905 67.530 222.115 67.790 ;
        RECT 10.150 66.430 209.270 67.530 ;
        RECT 1.905 65.490 222.115 66.430 ;
        RECT 10.150 64.390 211.570 65.490 ;
        RECT 1.905 64.130 222.115 64.390 ;
        RECT 1.905 63.450 206.510 64.130 ;
        RECT 17.510 63.030 206.510 63.450 ;
        RECT 17.510 62.350 222.115 63.030 ;
        RECT 1.905 62.090 222.115 62.350 ;
        RECT 14.290 60.990 206.050 62.090 ;
        RECT 1.905 60.050 222.115 60.990 ;
        RECT 7.390 58.950 209.270 60.050 ;
        RECT 1.905 58.690 222.115 58.950 ;
        RECT 10.150 57.590 205.590 58.690 ;
        RECT 1.905 56.650 222.115 57.590 ;
        RECT 10.150 55.550 216.110 56.650 ;
        RECT 1.905 55.290 222.115 55.550 ;
        RECT 1.905 54.610 206.050 55.290 ;
        RECT 10.610 54.190 206.050 54.610 ;
        RECT 10.610 53.510 222.115 54.190 ;
        RECT 1.905 53.250 222.115 53.510 ;
        RECT 17.510 52.150 212.430 53.250 ;
        RECT 1.905 51.210 222.115 52.150 ;
        RECT 14.290 50.110 205.590 51.210 ;
        RECT 1.905 49.850 222.115 50.110 ;
        RECT 1.905 49.170 206.510 49.850 ;
        RECT 10.150 48.750 206.510 49.170 ;
        RECT 10.150 48.070 222.115 48.750 ;
        RECT 1.905 47.810 222.115 48.070 ;
        RECT 14.290 46.710 214.270 47.810 ;
        RECT 1.905 45.770 222.115 46.710 ;
        RECT 7.390 44.670 209.730 45.770 ;
        RECT 1.905 44.410 222.115 44.670 ;
        RECT 10.150 43.310 209.270 44.410 ;
        RECT 1.905 42.370 222.115 43.310 ;
        RECT 14.290 41.270 206.510 42.370 ;
        RECT 1.905 40.330 222.115 41.270 ;
        RECT 7.390 39.230 211.570 40.330 ;
        RECT 1.905 38.970 222.115 39.230 ;
        RECT 10.610 37.870 207.890 38.970 ;
        RECT 1.905 36.930 222.115 37.870 ;
        RECT 14.290 35.830 206.510 36.930 ;
        RECT 1.905 35.570 222.115 35.830 ;
        RECT 1.905 34.890 209.270 35.570 ;
        RECT 7.390 34.470 209.270 34.890 ;
        RECT 7.390 33.790 222.115 34.470 ;
        RECT 1.905 33.530 222.115 33.790 ;
        RECT 10.150 32.430 205.130 33.530 ;
        RECT 1.905 31.490 222.115 32.430 ;
        RECT 14.290 30.390 212.030 31.490 ;
        RECT 1.905 30.130 222.115 30.390 ;
        RECT 7.390 29.030 202.370 30.130 ;
        RECT 1.905 28.090 222.115 29.030 ;
        RECT 10.150 26.990 206.970 28.090 ;
        RECT 1.905 26.050 222.115 26.990 ;
        RECT 17.510 24.950 205.130 26.050 ;
        RECT 1.905 24.690 222.115 24.950 ;
        RECT 14.290 23.590 200.990 24.690 ;
        RECT 1.905 22.650 222.115 23.590 ;
        RECT 7.390 21.550 204.670 22.650 ;
        RECT 1.905 20.610 222.115 21.550 ;
        RECT 20.270 19.510 209.270 20.610 ;
        RECT 1.905 19.250 222.115 19.510 ;
        RECT 6.930 18.150 206.050 19.250 ;
        RECT 1.905 17.210 222.115 18.150 ;
        RECT 15.670 16.110 202.370 17.210 ;
        RECT 1.905 15.850 222.115 16.110 ;
        RECT 20.730 14.750 200.530 15.850 ;
        RECT 1.905 13.810 222.115 14.750 ;
        RECT 17.510 12.710 200.070 13.810 ;
        RECT 1.905 11.770 222.115 12.710 ;
        RECT 17.050 10.670 200.070 11.770 ;
        RECT 1.905 10.410 222.115 10.670 ;
        RECT 16.590 9.310 200.530 10.410 ;
        RECT 1.905 8.370 222.115 9.310 ;
        RECT 20.270 7.270 211.570 8.370 ;
        RECT 1.905 6.330 222.115 7.270 ;
        RECT 18.430 5.230 200.530 6.330 ;
        RECT 1.905 4.970 222.115 5.230 ;
        RECT 15.210 3.870 209.730 4.970 ;
        RECT 1.905 2.930 222.115 3.870 ;
        RECT 16.130 1.830 200.990 2.930 ;
        RECT 1.905 1.570 222.115 1.830 ;
        RECT 15.670 0.855 206.050 1.570 ;
      LAYER met4 ;
        RECT 5.815 4.935 20.640 460.185 ;
        RECT 23.040 4.935 97.440 460.185 ;
        RECT 99.840 4.935 174.240 460.185 ;
        RECT 176.640 4.935 209.465 460.185 ;
  END
END DSP
MACRO N_term_DSP
  CLASS BLOCK ;
  FOREIGN N_term_DSP ;
  ORIGIN 0.000 0.000 ;
  SIZE 223.275 BY 40.000 ;
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.380 0.000 187.520 6.500 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.320 0.000 205.460 6.500 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.160 0.000 207.300 9.560 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.000 0.000 209.140 7.890 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.840 0.000 210.980 17.380 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.680 0.000 212.820 1.770 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.520 0.000 214.660 15.340 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.360 0.000 216.500 22.820 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.200 0.000 218.340 15.680 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.040 0.000 220.180 17.040 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.880 0.000 222.020 17.720 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.220 0.000 189.360 6.500 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.060 0.000 191.200 9.220 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.900 0.000 193.040 6.160 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.740 0.000 194.880 9.560 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.580 0.000 196.720 9.220 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.420 0.000 198.560 11.600 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.260 0.000 200.400 5.850 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.100 0.000 202.240 11.940 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.480 0.000 203.620 6.160 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.680 39.030 5.820 40.000 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.000 31.920 117.140 40.000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.040 31.920 128.180 40.000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.540 31.920 139.680 40.000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.580 31.920 150.720 40.000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.620 31.920 161.760 40.000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.660 31.920 172.800 40.000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.160 31.920 184.300 40.000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.200 31.920 195.340 40.000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.240 31.920 206.380 40.000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.280 31.920 217.420 40.000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.720 31.920 16.860 40.000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.760 31.920 27.900 40.000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.800 31.920 38.940 40.000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.300 31.920 50.440 40.000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.340 31.920 61.480 40.000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.380 31.920 72.520 40.000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.420 31.920 83.560 40.000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.920 31.920 95.060 40.000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.960 31.920 106.100 40.000 ;
    END
  END FrameStrobe_O[9]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.620 0.000 0.760 6.500 ;
    END
  END N1END[0]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.000 0.000 2.140 15.000 ;
    END
  END N1END[1]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.840 0.000 3.980 17.380 ;
    END
  END N1END[2]
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.680 0.000 5.820 17.040 ;
    END
  END N1END[3]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.780 0.000 21.920 11.940 ;
    END
  END N2END[0]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.620 0.000 23.760 6.500 ;
    END
  END N2END[1]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.460 0.000 25.600 6.020 ;
    END
  END N2END[2]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.300 0.000 27.440 9.560 ;
    END
  END N2END[3]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.140 0.000 29.280 11.940 ;
    END
  END N2END[4]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.980 0.000 31.120 9.220 ;
    END
  END N2END[5]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.820 0.000 32.960 11.940 ;
    END
  END N2END[6]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.660 0.000 34.800 11.600 ;
    END
  END N2END[7]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.520 0.000 7.660 9.560 ;
    END
  END N2MID[0]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.360 0.000 9.500 11.600 ;
    END
  END N2MID[1]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.200 0.000 11.340 15.000 ;
    END
  END N2MID[2]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.040 0.000 13.180 15.000 ;
    END
  END N2MID[3]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.880 0.000 15.020 6.500 ;
    END
  END N2MID[4]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.720 0.000 16.860 9.220 ;
    END
  END N2MID[5]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.560 0.000 18.700 11.940 ;
    END
  END N2MID[6]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.400 0.000 20.540 9.220 ;
    END
  END N2MID[7]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.500 0.000 36.640 6.160 ;
    END
  END N4END[0]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.440 0.000 54.580 6.500 ;
    END
  END N4END[10]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.280 0.000 56.420 17.380 ;
    END
  END N4END[11]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.120 0.000 58.260 13.980 ;
    END
  END N4END[12]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.960 0.000 60.100 13.870 ;
    END
  END N4END[13]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.340 0.000 61.480 14.320 ;
    END
  END N4END[14]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.180 0.000 63.320 6.700 ;
    END
  END N4END[15]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.340 0.000 38.480 6.160 ;
    END
  END N4END[1]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.180 0.000 40.320 2.450 ;
    END
  END N4END[2]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.560 0.000 41.700 5.000 ;
    END
  END N4END[3]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.400 0.000 43.540 11.600 ;
    END
  END N4END[4]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.240 0.000 45.380 11.800 ;
    END
  END N4END[5]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.080 0.000 47.220 6.500 ;
    END
  END N4END[6]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.920 0.000 49.060 9.220 ;
    END
  END N4END[7]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.760 0.000 50.900 6.160 ;
    END
  END N4END[8]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.600 0.000 52.740 11.940 ;
    END
  END N4END[9]
  PIN NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.020 0.000 65.160 17.380 ;
    END
  END NN4END[0]
  PIN NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.960 0.000 83.100 11.940 ;
    END
  END NN4END[10]
  PIN NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.800 0.000 84.940 11.940 ;
    END
  END NN4END[11]
  PIN NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.640 0.000 86.780 15.000 ;
    END
  END NN4END[12]
  PIN NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.480 0.000 88.620 17.380 ;
    END
  END NN4END[13]
  PIN NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.320 0.000 90.460 17.380 ;
    END
  END NN4END[14]
  PIN NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.160 0.000 92.300 13.870 ;
    END
  END NN4END[15]
  PIN NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.860 0.000 67.000 5.850 ;
    END
  END NN4END[1]
  PIN NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.700 0.000 68.840 7.210 ;
    END
  END NN4END[2]
  PIN NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.540 0.000 70.680 7.680 ;
    END
  END NN4END[3]
  PIN NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.380 0.000 72.520 14.660 ;
    END
  END NN4END[4]
  PIN NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.220 0.000 74.360 17.380 ;
    END
  END NN4END[5]
  PIN NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.060 0.000 76.200 4.120 ;
    END
  END NN4END[6]
  PIN NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.900 0.000 78.040 17.380 ;
    END
  END NN4END[7]
  PIN NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.740 0.000 79.880 1.090 ;
    END
  END NN4END[8]
  PIN NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.580 0.000 81.720 7.210 ;
    END
  END NN4END[9]
  PIN S1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.000 0.000 94.140 6.160 ;
    END
  END S1BEG[0]
  PIN S1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.840 0.000 95.980 5.820 ;
    END
  END S1BEG[1]
  PIN S1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.680 0.000 97.820 8.880 ;
    END
  END S1BEG[2]
  PIN S1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.520 0.000 99.660 6.500 ;
    END
  END S1BEG[3]
  PIN S2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.620 0.000 115.760 6.160 ;
    END
  END S2BEG[0]
  PIN S2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.460 0.000 117.600 6.160 ;
    END
  END S2BEG[1]
  PIN S2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.300 0.000 119.440 8.880 ;
    END
  END S2BEG[2]
  PIN S2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.140 0.000 121.280 5.820 ;
    END
  END S2BEG[3]
  PIN S2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.520 0.000 122.660 8.880 ;
    END
  END S2BEG[4]
  PIN S2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.360 0.000 124.500 6.500 ;
    END
  END S2BEG[5]
  PIN S2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.200 0.000 126.340 8.880 ;
    END
  END S2BEG[6]
  PIN S2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.040 0.000 128.180 8.880 ;
    END
  END S2BEG[7]
  PIN S2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.360 0.000 101.500 8.880 ;
    END
  END S2BEGb[0]
  PIN S2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.740 0.000 102.880 5.820 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.580 0.000 104.720 1.060 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.420 0.000 106.560 11.600 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.260 0.000 108.400 2.420 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.100 0.000 110.240 11.600 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.940 0.000 112.080 5.850 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.780 0.000 113.920 11.260 ;
    END
  END S2BEGb[7]
  PIN S4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.880 0.000 130.020 5.820 ;
    END
  END S4BEG[0]
  PIN S4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.820 0.000 147.960 3.130 ;
    END
  END S4BEG[10]
  PIN S4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.660 0.000 149.800 6.160 ;
    END
  END S4BEG[11]
  PIN S4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.500 0.000 151.640 5.820 ;
    END
  END S4BEG[12]
  PIN S4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.340 0.000 153.480 8.880 ;
    END
  END S4BEG[13]
  PIN S4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.180 0.000 155.320 6.160 ;
    END
  END S4BEG[14]
  PIN S4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.020 0.000 157.160 8.880 ;
    END
  END S4BEG[15]
  PIN S4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.720 0.000 131.860 8.880 ;
    END
  END S4BEG[1]
  PIN S4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.560 0.000 133.700 6.500 ;
    END
  END S4BEG[2]
  PIN S4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.400 0.000 135.540 8.880 ;
    END
  END S4BEG[3]
  PIN S4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.240 0.000 137.380 5.820 ;
    END
  END S4BEG[4]
  PIN S4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.080 0.000 139.220 8.540 ;
    END
  END S4BEG[5]
  PIN S4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.920 0.000 141.060 11.600 ;
    END
  END S4BEG[6]
  PIN S4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.300 0.000 142.440 8.880 ;
    END
  END S4BEG[7]
  PIN S4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.140 0.000 144.280 8.540 ;
    END
  END S4BEG[8]
  PIN S4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.980 0.000 146.120 4.490 ;
    END
  END S4BEG[9]
  PIN SS4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.860 0.000 159.000 5.820 ;
    END
  END SS4BEG[0]
  PIN SS4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.800 0.000 176.940 6.160 ;
    END
  END SS4BEG[10]
  PIN SS4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.640 0.000 178.780 6.160 ;
    END
  END SS4BEG[11]
  PIN SS4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.480 0.000 180.620 8.880 ;
    END
  END SS4BEG[12]
  PIN SS4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.320 0.000 182.460 6.840 ;
    END
  END SS4BEG[13]
  PIN SS4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.700 0.000 183.840 11.600 ;
    END
  END SS4BEG[14]
  PIN SS4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.540 0.000 185.680 11.600 ;
    END
  END SS4BEG[15]
  PIN SS4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.700 0.000 160.840 9.560 ;
    END
  END SS4BEG[1]
  PIN SS4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.540 0.000 162.680 6.500 ;
    END
  END SS4BEG[2]
  PIN SS4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.920 0.000 164.060 8.540 ;
    END
  END SS4BEG[3]
  PIN SS4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.760 0.000 165.900 5.820 ;
    END
  END SS4BEG[4]
  PIN SS4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.600 0.000 167.740 8.880 ;
    END
  END SS4BEG[5]
  PIN SS4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.440 0.000 169.580 8.540 ;
    END
  END SS4BEG[6]
  PIN SS4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.280 0.000 171.420 11.600 ;
    END
  END SS4BEG[7]
  PIN SS4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.120 0.000 173.260 11.260 ;
    END
  END SS4BEG[8]
  PIN SS4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.960 0.000 175.100 14.320 ;
    END
  END SS4BEG[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 40.090 5.200 41.690 32.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 110.835 5.200 112.435 32.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 181.580 5.200 183.180 32.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 75.465 5.200 77.065 32.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 146.210 5.200 147.810 32.880 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 0.085 217.580 32.725 ;
      LAYER met1 ;
        RECT 0.530 0.040 222.110 32.880 ;
      LAYER met2 ;
        RECT 0.560 38.750 5.400 39.850 ;
        RECT 6.100 38.750 16.440 39.850 ;
        RECT 0.560 31.640 16.440 38.750 ;
        RECT 17.140 31.640 27.480 39.850 ;
        RECT 28.180 31.640 38.520 39.850 ;
        RECT 39.220 31.640 50.020 39.850 ;
        RECT 50.720 31.640 61.060 39.850 ;
        RECT 61.760 31.640 72.100 39.850 ;
        RECT 72.800 31.640 83.140 39.850 ;
        RECT 83.840 31.640 94.640 39.850 ;
        RECT 95.340 31.640 105.680 39.850 ;
        RECT 106.380 31.640 116.720 39.850 ;
        RECT 117.420 31.640 127.760 39.850 ;
        RECT 128.460 31.640 139.260 39.850 ;
        RECT 139.960 31.640 150.300 39.850 ;
        RECT 151.000 31.640 161.340 39.850 ;
        RECT 162.040 31.640 172.380 39.850 ;
        RECT 173.080 31.640 183.880 39.850 ;
        RECT 184.580 31.640 194.920 39.850 ;
        RECT 195.620 31.640 205.960 39.850 ;
        RECT 206.660 31.640 217.000 39.850 ;
        RECT 217.700 31.640 222.080 39.850 ;
        RECT 0.560 23.100 222.080 31.640 ;
        RECT 0.560 17.660 216.080 23.100 ;
        RECT 0.560 15.280 3.560 17.660 ;
        RECT 0.560 6.780 1.720 15.280 ;
        RECT 1.040 0.010 1.720 6.780 ;
        RECT 2.420 0.010 3.560 15.280 ;
        RECT 4.260 17.320 56.000 17.660 ;
        RECT 4.260 0.010 5.400 17.320 ;
        RECT 6.100 15.280 56.000 17.320 ;
        RECT 6.100 11.880 10.920 15.280 ;
        RECT 6.100 9.840 9.080 11.880 ;
        RECT 6.100 0.010 7.240 9.840 ;
        RECT 7.940 0.010 9.080 9.840 ;
        RECT 9.780 0.010 10.920 11.880 ;
        RECT 11.620 0.010 12.760 15.280 ;
        RECT 13.460 12.220 56.000 15.280 ;
        RECT 13.460 9.500 18.280 12.220 ;
        RECT 13.460 6.780 16.440 9.500 ;
        RECT 13.460 0.010 14.600 6.780 ;
        RECT 15.300 0.010 16.440 6.780 ;
        RECT 17.140 0.010 18.280 9.500 ;
        RECT 18.980 9.500 21.500 12.220 ;
        RECT 18.980 0.010 20.120 9.500 ;
        RECT 20.820 0.010 21.500 9.500 ;
        RECT 22.200 9.840 28.860 12.220 ;
        RECT 22.200 6.780 27.020 9.840 ;
        RECT 22.200 0.010 23.340 6.780 ;
        RECT 24.040 6.300 27.020 6.780 ;
        RECT 24.040 0.010 25.180 6.300 ;
        RECT 25.880 0.010 27.020 6.300 ;
        RECT 27.720 0.010 28.860 9.840 ;
        RECT 29.560 9.500 32.540 12.220 ;
        RECT 29.560 0.010 30.700 9.500 ;
        RECT 31.400 0.010 32.540 9.500 ;
        RECT 33.240 12.080 52.320 12.220 ;
        RECT 33.240 11.880 44.960 12.080 ;
        RECT 33.240 0.010 34.380 11.880 ;
        RECT 35.080 6.440 43.120 11.880 ;
        RECT 35.080 0.010 36.220 6.440 ;
        RECT 36.920 0.010 38.060 6.440 ;
        RECT 38.760 5.280 43.120 6.440 ;
        RECT 38.760 2.730 41.280 5.280 ;
        RECT 38.760 0.010 39.900 2.730 ;
        RECT 40.600 0.010 41.280 2.730 ;
        RECT 41.980 0.010 43.120 5.280 ;
        RECT 43.820 0.010 44.960 11.880 ;
        RECT 45.660 9.500 52.320 12.080 ;
        RECT 45.660 6.780 48.640 9.500 ;
        RECT 45.660 0.010 46.800 6.780 ;
        RECT 47.500 0.010 48.640 6.780 ;
        RECT 49.340 6.440 52.320 9.500 ;
        RECT 49.340 0.010 50.480 6.440 ;
        RECT 51.180 0.010 52.320 6.440 ;
        RECT 53.020 6.780 56.000 12.220 ;
        RECT 53.020 0.010 54.160 6.780 ;
        RECT 54.860 0.010 56.000 6.780 ;
        RECT 56.700 14.600 64.740 17.660 ;
        RECT 56.700 14.260 61.060 14.600 ;
        RECT 56.700 0.010 57.840 14.260 ;
        RECT 58.540 14.150 61.060 14.260 ;
        RECT 58.540 0.010 59.680 14.150 ;
        RECT 60.380 0.010 61.060 14.150 ;
        RECT 61.760 6.980 64.740 14.600 ;
        RECT 61.760 0.010 62.900 6.980 ;
        RECT 63.600 0.010 64.740 6.980 ;
        RECT 65.440 14.940 73.940 17.660 ;
        RECT 65.440 7.960 72.100 14.940 ;
        RECT 65.440 7.490 70.260 7.960 ;
        RECT 65.440 6.130 68.420 7.490 ;
        RECT 65.440 0.010 66.580 6.130 ;
        RECT 67.280 0.010 68.420 6.130 ;
        RECT 69.120 0.010 70.260 7.490 ;
        RECT 70.960 0.010 72.100 7.960 ;
        RECT 72.800 0.010 73.940 14.940 ;
        RECT 74.640 4.400 77.620 17.660 ;
        RECT 74.640 0.010 75.780 4.400 ;
        RECT 76.480 0.010 77.620 4.400 ;
        RECT 78.320 15.280 88.200 17.660 ;
        RECT 78.320 12.220 86.360 15.280 ;
        RECT 78.320 7.490 82.680 12.220 ;
        RECT 78.320 1.370 81.300 7.490 ;
        RECT 78.320 0.010 79.460 1.370 ;
        RECT 80.160 0.010 81.300 1.370 ;
        RECT 82.000 0.010 82.680 7.490 ;
        RECT 83.380 0.010 84.520 12.220 ;
        RECT 85.220 0.010 86.360 12.220 ;
        RECT 87.060 0.010 88.200 15.280 ;
        RECT 88.900 0.010 90.040 17.660 ;
        RECT 90.740 14.600 210.560 17.660 ;
        RECT 90.740 14.150 174.680 14.600 ;
        RECT 90.740 0.010 91.880 14.150 ;
        RECT 92.580 11.880 174.680 14.150 ;
        RECT 92.580 9.160 106.140 11.880 ;
        RECT 92.580 6.440 97.400 9.160 ;
        RECT 92.580 0.010 93.720 6.440 ;
        RECT 94.420 6.100 97.400 6.440 ;
        RECT 94.420 0.010 95.560 6.100 ;
        RECT 96.260 0.010 97.400 6.100 ;
        RECT 98.100 6.780 101.080 9.160 ;
        RECT 98.100 0.010 99.240 6.780 ;
        RECT 99.940 0.010 101.080 6.780 ;
        RECT 101.780 6.100 106.140 9.160 ;
        RECT 101.780 0.010 102.460 6.100 ;
        RECT 103.160 1.340 106.140 6.100 ;
        RECT 103.160 0.010 104.300 1.340 ;
        RECT 105.000 0.010 106.140 1.340 ;
        RECT 106.840 2.700 109.820 11.880 ;
        RECT 106.840 0.010 107.980 2.700 ;
        RECT 108.680 0.010 109.820 2.700 ;
        RECT 110.520 11.540 140.640 11.880 ;
        RECT 110.520 6.130 113.500 11.540 ;
        RECT 110.520 0.010 111.660 6.130 ;
        RECT 112.360 0.010 113.500 6.130 ;
        RECT 114.200 9.160 140.640 11.540 ;
        RECT 114.200 6.440 119.020 9.160 ;
        RECT 114.200 0.010 115.340 6.440 ;
        RECT 116.040 0.010 117.180 6.440 ;
        RECT 117.880 0.010 119.020 6.440 ;
        RECT 119.720 6.100 122.240 9.160 ;
        RECT 119.720 0.010 120.860 6.100 ;
        RECT 121.560 0.010 122.240 6.100 ;
        RECT 122.940 6.780 125.920 9.160 ;
        RECT 122.940 0.010 124.080 6.780 ;
        RECT 124.780 0.010 125.920 6.780 ;
        RECT 126.620 0.010 127.760 9.160 ;
        RECT 128.460 6.100 131.440 9.160 ;
        RECT 128.460 0.010 129.600 6.100 ;
        RECT 130.300 0.010 131.440 6.100 ;
        RECT 132.140 6.780 135.120 9.160 ;
        RECT 132.140 0.010 133.280 6.780 ;
        RECT 133.980 0.010 135.120 6.780 ;
        RECT 135.820 8.820 140.640 9.160 ;
        RECT 135.820 6.100 138.800 8.820 ;
        RECT 135.820 0.010 136.960 6.100 ;
        RECT 137.660 0.010 138.800 6.100 ;
        RECT 139.500 0.010 140.640 8.820 ;
        RECT 141.340 9.840 171.000 11.880 ;
        RECT 141.340 9.160 160.420 9.840 ;
        RECT 141.340 0.010 142.020 9.160 ;
        RECT 142.720 8.820 153.060 9.160 ;
        RECT 142.720 0.010 143.860 8.820 ;
        RECT 144.560 6.440 153.060 8.820 ;
        RECT 144.560 4.770 149.380 6.440 ;
        RECT 144.560 0.010 145.700 4.770 ;
        RECT 146.400 3.410 149.380 4.770 ;
        RECT 146.400 0.010 147.540 3.410 ;
        RECT 148.240 0.010 149.380 3.410 ;
        RECT 150.080 6.100 153.060 6.440 ;
        RECT 150.080 0.010 151.220 6.100 ;
        RECT 151.920 0.010 153.060 6.100 ;
        RECT 153.760 6.440 156.740 9.160 ;
        RECT 153.760 0.010 154.900 6.440 ;
        RECT 155.600 0.010 156.740 6.440 ;
        RECT 157.440 6.100 160.420 9.160 ;
        RECT 157.440 0.010 158.580 6.100 ;
        RECT 159.280 0.010 160.420 6.100 ;
        RECT 161.120 9.160 171.000 9.840 ;
        RECT 161.120 8.820 167.320 9.160 ;
        RECT 161.120 6.780 163.640 8.820 ;
        RECT 161.120 0.010 162.260 6.780 ;
        RECT 162.960 0.010 163.640 6.780 ;
        RECT 164.340 6.100 167.320 8.820 ;
        RECT 164.340 0.010 165.480 6.100 ;
        RECT 166.180 0.010 167.320 6.100 ;
        RECT 168.020 8.820 171.000 9.160 ;
        RECT 168.020 0.010 169.160 8.820 ;
        RECT 169.860 0.010 171.000 8.820 ;
        RECT 171.700 11.540 174.680 11.880 ;
        RECT 171.700 0.010 172.840 11.540 ;
        RECT 173.540 0.010 174.680 11.540 ;
        RECT 175.380 12.220 210.560 14.600 ;
        RECT 175.380 11.880 201.820 12.220 ;
        RECT 175.380 9.160 183.420 11.880 ;
        RECT 175.380 6.440 180.200 9.160 ;
        RECT 175.380 0.010 176.520 6.440 ;
        RECT 177.220 0.010 178.360 6.440 ;
        RECT 179.060 0.010 180.200 6.440 ;
        RECT 180.900 7.120 183.420 9.160 ;
        RECT 180.900 0.010 182.040 7.120 ;
        RECT 182.740 0.010 183.420 7.120 ;
        RECT 184.120 0.010 185.260 11.880 ;
        RECT 185.960 9.840 198.140 11.880 ;
        RECT 185.960 9.500 194.460 9.840 ;
        RECT 185.960 6.780 190.780 9.500 ;
        RECT 185.960 0.010 187.100 6.780 ;
        RECT 187.800 0.010 188.940 6.780 ;
        RECT 189.640 0.010 190.780 6.780 ;
        RECT 191.480 6.440 194.460 9.500 ;
        RECT 191.480 0.010 192.620 6.440 ;
        RECT 193.320 0.010 194.460 6.440 ;
        RECT 195.160 9.500 198.140 9.840 ;
        RECT 195.160 0.010 196.300 9.500 ;
        RECT 197.000 0.010 198.140 9.500 ;
        RECT 198.840 6.130 201.820 11.880 ;
        RECT 198.840 0.010 199.980 6.130 ;
        RECT 200.680 0.010 201.820 6.130 ;
        RECT 202.520 9.840 210.560 12.220 ;
        RECT 202.520 6.780 206.880 9.840 ;
        RECT 202.520 6.440 205.040 6.780 ;
        RECT 202.520 0.010 203.200 6.440 ;
        RECT 203.900 0.010 205.040 6.440 ;
        RECT 205.740 0.010 206.880 6.780 ;
        RECT 207.580 8.170 210.560 9.840 ;
        RECT 207.580 0.010 208.720 8.170 ;
        RECT 209.420 0.010 210.560 8.170 ;
        RECT 211.260 15.620 216.080 17.660 ;
        RECT 211.260 2.050 214.240 15.620 ;
        RECT 211.260 0.010 212.400 2.050 ;
        RECT 213.100 0.010 214.240 2.050 ;
        RECT 214.940 0.010 216.080 15.620 ;
        RECT 216.780 18.000 222.080 23.100 ;
        RECT 216.780 17.320 221.600 18.000 ;
        RECT 216.780 15.960 219.760 17.320 ;
        RECT 216.780 0.010 217.920 15.960 ;
        RECT 218.620 0.010 219.760 15.960 ;
        RECT 220.460 0.010 221.600 17.320 ;
      LAYER met3 ;
        RECT 13.405 3.575 200.035 32.805 ;
  END
END N_term_DSP
MACRO N_term_RAM_IO
  CLASS BLOCK ;
  FOREIGN N_term_RAM_IO ;
  ORIGIN 0.000 0.000 ;
  SIZE 125.000 BY 40.000 ;
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.140 0.000 98.280 7.890 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.940 0.000 112.080 9.560 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.320 0.000 113.460 11.940 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.700 0.000 114.840 9.220 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.080 0.000 116.220 15.000 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.460 0.000 117.600 11.600 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.840 0.000 118.980 14.660 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.220 0.000 120.360 12.280 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.600 0.000 121.740 11.260 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.980 0.000 123.120 17.040 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.360 0.000 124.500 14.320 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.520 0.000 99.660 7.210 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.900 0.000 101.040 7.210 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.280 0.000 102.420 17.040 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.660 0.000 103.800 6.700 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.040 0.000 105.180 6.500 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.420 0.000 106.560 10.610 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.800 0.000 107.940 20.440 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.180 0.000 109.320 9.930 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.560 0.000 110.700 2.450 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.920 31.920 3.060 40.000 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.480 31.920 65.620 40.000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.460 31.920 71.600 40.000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.900 31.920 78.040 40.000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.880 31.920 84.020 40.000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.320 31.920 90.460 40.000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.760 31.920 96.900 40.000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.740 31.920 102.880 40.000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.180 31.920 109.320 40.000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.160 32.260 115.300 40.000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.600 29.200 121.740 40.000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.900 31.920 9.040 40.000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.340 31.920 15.480 40.000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.320 31.920 21.460 40.000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.760 31.920 27.900 40.000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.200 31.920 34.340 40.000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.180 31.920 40.320 40.000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.620 31.920 46.760 40.000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.600 31.920 52.740 40.000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.040 31.920 59.180 40.000 ;
    END
  END FrameStrobe_O[9]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.620 0.000 0.760 9.560 ;
    END
  END N1END[0]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.540 0.000 1.680 11.940 ;
    END
  END N1END[1]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.920 0.000 3.060 9.220 ;
    END
  END N1END[2]
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.300 0.000 4.440 8.880 ;
    END
  END N1END[3]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.720 0.000 16.860 9.560 ;
    END
  END N2END[0]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.100 0.000 18.240 11.940 ;
    END
  END N2END[1]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.480 0.000 19.620 11.940 ;
    END
  END N2END[2]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.860 0.000 21.000 11.600 ;
    END
  END N2END[3]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.240 0.000 22.380 15.000 ;
    END
  END N2END[4]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.620 0.000 23.760 7.210 ;
    END
  END N2END[5]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.000 0.000 25.140 6.530 ;
    END
  END N2END[6]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.380 0.000 26.520 12.280 ;
    END
  END N2END[7]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.680 0.000 5.820 11.600 ;
    END
  END N2MID[0]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.060 0.000 7.200 15.000 ;
    END
  END N2MID[1]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.440 0.000 8.580 15.000 ;
    END
  END N2MID[2]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.820 0.000 9.960 11.600 ;
    END
  END N2MID[3]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.200 0.000 11.340 15.000 ;
    END
  END N2MID[4]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.580 0.000 12.720 14.660 ;
    END
  END N2MID[5]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.960 0.000 14.100 17.380 ;
    END
  END N2MID[6]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.340 0.000 15.480 17.380 ;
    END
  END N2MID[7]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.760 0.000 27.900 15.000 ;
    END
  END N4END[0]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.100 0.000 41.240 9.220 ;
    END
  END N4END[10]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.480 0.000 42.620 4.490 ;
    END
  END N4END[11]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.860 0.000 44.000 4.490 ;
    END
  END N4END[12]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.240 0.000 45.380 1.090 ;
    END
  END N4END[13]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.620 0.000 46.760 17.380 ;
    END
  END N4END[14]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.000 0.000 48.140 17.380 ;
    END
  END N4END[15]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.140 0.000 29.280 3.130 ;
    END
  END N4END[1]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.520 0.000 30.660 15.340 ;
    END
  END N4END[2]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.900 0.000 32.040 17.380 ;
    END
  END N4END[3]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.820 0.000 32.960 7.890 ;
    END
  END N4END[4]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.200 0.000 34.340 6.700 ;
    END
  END N4END[5]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.580 0.000 35.720 7.210 ;
    END
  END N4END[6]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.960 0.000 37.100 7.210 ;
    END
  END N4END[7]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.340 0.000 38.480 20.640 ;
    END
  END N4END[8]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.720 0.000 39.860 1.090 ;
    END
  END N4END[9]
  PIN S1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.380 0.000 49.520 6.160 ;
    END
  END S1BEG[0]
  PIN S1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.760 0.000 50.900 5.820 ;
    END
  END S1BEG[1]
  PIN S1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.140 0.000 52.280 8.880 ;
    END
  END S1BEG[2]
  PIN S1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.520 0.000 53.660 4.800 ;
    END
  END S1BEG[3]
  PIN S2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.480 0.000 65.620 6.160 ;
    END
  END S2BEG[0]
  PIN S2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.860 0.000 67.000 3.130 ;
    END
  END S2BEG[1]
  PIN S2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.240 0.000 68.380 8.880 ;
    END
  END S2BEG[2]
  PIN S2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.620 0.000 69.760 5.820 ;
    END
  END S2BEG[3]
  PIN S2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.000 0.000 71.140 4.490 ;
    END
  END S2BEG[4]
  PIN S2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.380 0.000 72.520 6.160 ;
    END
  END S2BEG[5]
  PIN S2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.760 0.000 73.900 4.490 ;
    END
  END S2BEG[6]
  PIN S2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.140 0.000 75.280 5.820 ;
    END
  END S2BEG[7]
  PIN S2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.900 0.000 55.040 8.880 ;
    END
  END S2BEGb[0]
  PIN S2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.280 0.000 56.420 5.820 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.660 0.000 57.800 4.490 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.040 0.000 59.180 11.600 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.420 0.000 60.560 8.540 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.800 0.000 61.940 5.850 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.180 0.000 63.320 7.210 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.100 0.000 64.240 7.210 ;
    END
  END S2BEGb[7]
  PIN S4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.520 0.000 76.660 11.600 ;
    END
  END S4BEG[0]
  PIN S4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.320 0.000 90.460 6.160 ;
    END
  END S4BEG[10]
  PIN S4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.700 0.000 91.840 3.130 ;
    END
  END S4BEG[11]
  PIN S4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.080 0.000 93.220 8.880 ;
    END
  END S4BEG[12]
  PIN S4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.460 0.000 94.600 8.880 ;
    END
  END S4BEG[13]
  PIN S4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.380 0.000 95.520 11.600 ;
    END
  END S4BEG[14]
  PIN S4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.760 0.000 96.900 8.540 ;
    END
  END S4BEG[15]
  PIN S4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.900 0.000 78.040 3.130 ;
    END
  END S4BEG[1]
  PIN S4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.280 0.000 79.420 8.880 ;
    END
  END S4BEG[2]
  PIN S4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.660 0.000 80.800 5.000 ;
    END
  END S4BEG[3]
  PIN S4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.040 0.000 82.180 4.490 ;
    END
  END S4BEG[4]
  PIN S4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.420 0.000 83.560 11.600 ;
    END
  END S4BEG[5]
  PIN S4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.800 0.000 84.940 5.850 ;
    END
  END S4BEG[6]
  PIN S4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.180 0.000 86.320 14.320 ;
    END
  END S4BEG[7]
  PIN S4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.560 0.000 87.700 12.280 ;
    END
  END S4BEG[8]
  PIN S4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.940 0.000 89.080 14.320 ;
    END
  END S4BEG[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 23.715 5.200 25.315 32.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 61.700 5.200 63.300 32.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 99.685 5.200 101.285 32.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 42.705 5.200 44.305 32.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 80.690 5.200 82.290 32.880 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 1.445 119.140 32.725 ;
      LAYER met1 ;
        RECT 0.530 1.400 124.590 34.300 ;
      LAYER met2 ;
        RECT 0.560 31.640 2.640 34.330 ;
        RECT 3.340 31.640 8.620 34.330 ;
        RECT 9.320 31.640 15.060 34.330 ;
        RECT 15.760 31.640 21.040 34.330 ;
        RECT 21.740 31.640 27.480 34.330 ;
        RECT 28.180 31.640 33.920 34.330 ;
        RECT 34.620 31.640 39.900 34.330 ;
        RECT 40.600 31.640 46.340 34.330 ;
        RECT 47.040 31.640 52.320 34.330 ;
        RECT 53.020 31.640 58.760 34.330 ;
        RECT 59.460 31.640 65.200 34.330 ;
        RECT 65.900 31.640 71.180 34.330 ;
        RECT 71.880 31.640 77.620 34.330 ;
        RECT 78.320 31.640 83.600 34.330 ;
        RECT 84.300 31.640 90.040 34.330 ;
        RECT 90.740 31.640 96.480 34.330 ;
        RECT 97.180 31.640 102.460 34.330 ;
        RECT 103.160 31.640 108.900 34.330 ;
        RECT 109.600 31.980 114.880 34.330 ;
        RECT 115.580 31.980 121.320 34.330 ;
        RECT 109.600 31.640 121.320 31.980 ;
        RECT 0.560 28.920 121.320 31.640 ;
        RECT 122.020 28.920 124.560 34.330 ;
        RECT 0.560 20.920 124.560 28.920 ;
        RECT 0.560 17.660 38.060 20.920 ;
        RECT 0.560 15.280 13.680 17.660 ;
        RECT 0.560 12.220 6.780 15.280 ;
        RECT 0.560 9.840 1.260 12.220 ;
        RECT 1.040 0.950 1.260 9.840 ;
        RECT 1.960 11.880 6.780 12.220 ;
        RECT 1.960 9.500 5.400 11.880 ;
        RECT 1.960 0.950 2.640 9.500 ;
        RECT 3.340 9.160 5.400 9.500 ;
        RECT 3.340 0.950 4.020 9.160 ;
        RECT 4.720 0.950 5.400 9.160 ;
        RECT 6.100 0.950 6.780 11.880 ;
        RECT 7.480 0.950 8.160 15.280 ;
        RECT 8.860 11.880 10.920 15.280 ;
        RECT 8.860 0.950 9.540 11.880 ;
        RECT 10.240 0.950 10.920 11.880 ;
        RECT 11.620 14.940 13.680 15.280 ;
        RECT 11.620 0.950 12.300 14.940 ;
        RECT 13.000 0.950 13.680 14.940 ;
        RECT 14.380 0.950 15.060 17.660 ;
        RECT 15.760 15.620 31.620 17.660 ;
        RECT 15.760 15.280 30.240 15.620 ;
        RECT 15.760 12.220 21.960 15.280 ;
        RECT 15.760 9.840 17.820 12.220 ;
        RECT 15.760 0.950 16.440 9.840 ;
        RECT 17.140 0.950 17.820 9.840 ;
        RECT 18.520 0.950 19.200 12.220 ;
        RECT 19.900 11.880 21.960 12.220 ;
        RECT 19.900 0.950 20.580 11.880 ;
        RECT 21.280 0.950 21.960 11.880 ;
        RECT 22.660 12.560 27.480 15.280 ;
        RECT 22.660 7.490 26.100 12.560 ;
        RECT 22.660 0.950 23.340 7.490 ;
        RECT 24.040 6.810 26.100 7.490 ;
        RECT 24.040 0.950 24.720 6.810 ;
        RECT 25.420 0.950 26.100 6.810 ;
        RECT 26.800 0.950 27.480 12.560 ;
        RECT 28.180 3.410 30.240 15.280 ;
        RECT 28.180 0.950 28.860 3.410 ;
        RECT 29.560 0.950 30.240 3.410 ;
        RECT 30.940 0.950 31.620 15.620 ;
        RECT 32.320 8.170 38.060 17.660 ;
        RECT 32.320 0.950 32.540 8.170 ;
        RECT 33.240 7.490 38.060 8.170 ;
        RECT 33.240 6.980 35.300 7.490 ;
        RECT 33.240 0.950 33.920 6.980 ;
        RECT 34.620 0.950 35.300 6.980 ;
        RECT 36.000 0.950 36.680 7.490 ;
        RECT 37.380 0.950 38.060 7.490 ;
        RECT 38.760 20.720 124.560 20.920 ;
        RECT 38.760 17.660 107.520 20.720 ;
        RECT 38.760 9.500 46.340 17.660 ;
        RECT 38.760 1.370 40.820 9.500 ;
        RECT 38.760 0.950 39.440 1.370 ;
        RECT 40.140 0.950 40.820 1.370 ;
        RECT 41.520 4.770 46.340 9.500 ;
        RECT 41.520 0.950 42.200 4.770 ;
        RECT 42.900 0.950 43.580 4.770 ;
        RECT 44.280 1.370 46.340 4.770 ;
        RECT 44.280 0.950 44.960 1.370 ;
        RECT 45.660 0.950 46.340 1.370 ;
        RECT 47.040 0.950 47.720 17.660 ;
        RECT 48.420 17.320 107.520 17.660 ;
        RECT 48.420 14.600 102.000 17.320 ;
        RECT 48.420 11.880 85.900 14.600 ;
        RECT 48.420 9.160 58.760 11.880 ;
        RECT 48.420 6.440 51.860 9.160 ;
        RECT 48.420 0.950 49.100 6.440 ;
        RECT 49.800 6.100 51.860 6.440 ;
        RECT 49.800 0.950 50.480 6.100 ;
        RECT 51.180 0.950 51.860 6.100 ;
        RECT 52.560 5.080 54.620 9.160 ;
        RECT 52.560 0.950 53.240 5.080 ;
        RECT 53.940 0.950 54.620 5.080 ;
        RECT 55.320 6.100 58.760 9.160 ;
        RECT 55.320 0.950 56.000 6.100 ;
        RECT 56.700 4.770 58.760 6.100 ;
        RECT 56.700 0.950 57.380 4.770 ;
        RECT 58.080 0.950 58.760 4.770 ;
        RECT 59.460 9.160 76.240 11.880 ;
        RECT 59.460 8.820 67.960 9.160 ;
        RECT 59.460 0.950 60.140 8.820 ;
        RECT 60.840 7.490 67.960 8.820 ;
        RECT 60.840 6.130 62.900 7.490 ;
        RECT 60.840 0.950 61.520 6.130 ;
        RECT 62.220 0.950 62.900 6.130 ;
        RECT 63.600 0.950 63.820 7.490 ;
        RECT 64.520 6.440 67.960 7.490 ;
        RECT 64.520 0.950 65.200 6.440 ;
        RECT 65.900 3.410 67.960 6.440 ;
        RECT 65.900 0.950 66.580 3.410 ;
        RECT 67.280 0.950 67.960 3.410 ;
        RECT 68.660 6.440 76.240 9.160 ;
        RECT 68.660 6.100 72.100 6.440 ;
        RECT 68.660 0.950 69.340 6.100 ;
        RECT 70.040 4.770 72.100 6.100 ;
        RECT 70.040 0.950 70.720 4.770 ;
        RECT 71.420 0.950 72.100 4.770 ;
        RECT 72.800 6.100 76.240 6.440 ;
        RECT 72.800 4.770 74.860 6.100 ;
        RECT 72.800 0.950 73.480 4.770 ;
        RECT 74.180 0.950 74.860 4.770 ;
        RECT 75.560 0.950 76.240 6.100 ;
        RECT 76.940 9.160 83.140 11.880 ;
        RECT 76.940 3.410 79.000 9.160 ;
        RECT 76.940 0.950 77.620 3.410 ;
        RECT 78.320 0.950 79.000 3.410 ;
        RECT 79.700 5.280 83.140 9.160 ;
        RECT 79.700 0.950 80.380 5.280 ;
        RECT 81.080 4.770 83.140 5.280 ;
        RECT 81.080 0.950 81.760 4.770 ;
        RECT 82.460 0.950 83.140 4.770 ;
        RECT 83.840 6.130 85.900 11.880 ;
        RECT 83.840 0.950 84.520 6.130 ;
        RECT 85.220 0.950 85.900 6.130 ;
        RECT 86.600 12.560 88.660 14.600 ;
        RECT 86.600 0.950 87.280 12.560 ;
        RECT 87.980 0.950 88.660 12.560 ;
        RECT 89.360 11.880 102.000 14.600 ;
        RECT 89.360 9.160 95.100 11.880 ;
        RECT 89.360 6.440 92.800 9.160 ;
        RECT 89.360 0.950 90.040 6.440 ;
        RECT 90.740 3.410 92.800 6.440 ;
        RECT 90.740 0.950 91.420 3.410 ;
        RECT 92.120 0.950 92.800 3.410 ;
        RECT 93.500 0.950 94.180 9.160 ;
        RECT 94.880 0.950 95.100 9.160 ;
        RECT 95.800 8.820 102.000 11.880 ;
        RECT 95.800 0.950 96.480 8.820 ;
        RECT 97.180 8.170 102.000 8.820 ;
        RECT 97.180 0.950 97.860 8.170 ;
        RECT 98.560 7.490 102.000 8.170 ;
        RECT 98.560 0.950 99.240 7.490 ;
        RECT 99.940 0.950 100.620 7.490 ;
        RECT 101.320 0.950 102.000 7.490 ;
        RECT 102.700 10.890 107.520 17.320 ;
        RECT 102.700 6.980 106.140 10.890 ;
        RECT 102.700 0.950 103.380 6.980 ;
        RECT 104.080 6.780 106.140 6.980 ;
        RECT 104.080 0.950 104.760 6.780 ;
        RECT 105.460 0.950 106.140 6.780 ;
        RECT 106.840 0.950 107.520 10.890 ;
        RECT 108.220 17.320 124.560 20.720 ;
        RECT 108.220 15.280 122.700 17.320 ;
        RECT 108.220 12.220 115.800 15.280 ;
        RECT 108.220 10.210 113.040 12.220 ;
        RECT 108.220 0.950 108.900 10.210 ;
        RECT 109.600 9.840 113.040 10.210 ;
        RECT 109.600 2.730 111.660 9.840 ;
        RECT 109.600 0.950 110.280 2.730 ;
        RECT 110.980 0.950 111.660 2.730 ;
        RECT 112.360 0.950 113.040 9.840 ;
        RECT 113.740 9.500 115.800 12.220 ;
        RECT 113.740 0.950 114.420 9.500 ;
        RECT 115.120 0.950 115.800 9.500 ;
        RECT 116.500 14.940 122.700 15.280 ;
        RECT 116.500 11.880 118.560 14.940 ;
        RECT 116.500 0.950 117.180 11.880 ;
        RECT 117.880 0.950 118.560 11.880 ;
        RECT 119.260 12.560 122.700 14.940 ;
        RECT 119.260 0.950 119.940 12.560 ;
        RECT 120.640 11.540 122.700 12.560 ;
        RECT 120.640 0.950 121.320 11.540 ;
        RECT 122.020 0.950 122.700 11.540 ;
        RECT 123.400 14.600 124.560 17.320 ;
        RECT 123.400 0.950 124.080 14.600 ;
      LAYER met3 ;
        RECT 14.325 5.275 101.285 32.805 ;
  END
END N_term_RAM_IO
MACRO N_term_single
  CLASS BLOCK ;
  FOREIGN N_term_single ;
  ORIGIN 0.000 0.000 ;
  SIZE 223.275 BY 40.000 ;
  PIN Ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.000 0.000 186.140 0.800 ;
    END
  END Ci
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.840 0.000 187.980 15.000 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.780 0.000 205.920 6.500 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.620 0.000 207.760 9.560 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.000 0.000 209.140 7.890 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.840 0.000 210.980 17.380 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.680 0.000 212.820 20.440 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.520 0.000 214.660 14.660 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.360 0.000 216.500 22.820 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.200 0.000 218.340 20.100 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.040 0.000 220.180 17.720 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.880 0.000 222.020 15.340 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.680 0.000 189.820 6.500 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.520 0.000 191.660 9.220 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.360 0.000 193.500 5.820 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.740 0.000 194.880 9.560 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.580 0.000 196.720 11.600 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.420 0.000 198.560 9.900 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.260 0.000 200.400 11.800 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.100 0.000 202.240 11.940 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.940 0.000 204.080 6.160 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.680 39.030 5.820 40.000 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.000 34.950 117.140 40.000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.040 31.920 128.180 40.000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.540 31.920 139.680 40.000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.580 31.920 150.720 40.000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.620 31.920 161.760 40.000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.660 31.920 172.800 40.000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.160 31.920 184.300 40.000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.200 31.920 195.340 40.000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.240 31.920 206.380 40.000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.280 31.920 217.420 40.000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.720 31.920 16.860 40.000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.760 31.920 27.900 40.000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.800 31.920 38.940 40.000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.300 31.920 50.440 40.000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.340 31.920 61.480 40.000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.380 31.920 72.520 40.000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.420 31.920 83.560 40.000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.920 31.920 95.060 40.000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.960 31.920 106.100 40.000 ;
    END
  END FrameStrobe_O[9]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.620 0.000 0.760 15.000 ;
    END
  END N1END[0]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.000 0.000 2.140 17.380 ;
    END
  END N1END[1]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.840 0.000 3.980 20.440 ;
    END
  END N1END[2]
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.680 0.000 5.820 17.040 ;
    END
  END N1END[3]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.780 0.000 21.920 11.940 ;
    END
  END N2END[0]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.620 0.000 23.760 3.440 ;
    END
  END N2END[1]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.460 0.000 25.600 12.140 ;
    END
  END N2END[2]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.300 0.000 27.440 9.560 ;
    END
  END N2END[3]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.140 0.000 29.280 11.940 ;
    END
  END N2END[4]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.520 0.000 30.660 9.220 ;
    END
  END N2END[5]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.360 0.000 32.500 1.090 ;
    END
  END N2END[6]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.200 0.000 34.340 11.600 ;
    END
  END N2END[7]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.520 0.000 7.660 9.560 ;
    END
  END N2MID[0]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.360 0.000 9.500 11.600 ;
    END
  END N2MID[1]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.200 0.000 11.340 5.850 ;
    END
  END N2MID[2]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.040 0.000 13.180 3.100 ;
    END
  END N2MID[3]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.880 0.000 15.020 6.500 ;
    END
  END N2MID[4]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.260 0.000 16.400 9.220 ;
    END
  END N2MID[5]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.100 0.000 18.240 11.940 ;
    END
  END N2MID[6]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.940 0.000 20.080 9.220 ;
    END
  END N2MID[7]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.040 0.000 36.180 6.160 ;
    END
  END N4END[0]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.980 0.000 54.120 11.940 ;
    END
  END N4END[10]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.820 0.000 55.960 11.940 ;
    END
  END N4END[11]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.660 0.000 57.800 15.000 ;
    END
  END N4END[12]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.500 0.000 59.640 9.900 ;
    END
  END N4END[13]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.880 0.000 61.020 15.200 ;
    END
  END N4END[14]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.720 0.000 62.860 17.380 ;
    END
  END N4END[15]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.880 0.000 38.020 6.160 ;
    END
  END N4END[1]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.720 0.000 39.860 9.560 ;
    END
  END N4END[2]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.560 0.000 41.700 5.170 ;
    END
  END N4END[3]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.400 0.000 43.540 11.600 ;
    END
  END N4END[4]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.240 0.000 45.380 6.020 ;
    END
  END N4END[5]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.620 0.000 46.760 6.500 ;
    END
  END N4END[6]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.460 0.000 48.600 9.220 ;
    END
  END N4END[7]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.300 0.000 50.440 3.440 ;
    END
  END N4END[8]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.140 0.000 52.280 15.000 ;
    END
  END N4END[9]
  PIN NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.560 0.000 64.700 17.380 ;
    END
  END NN4END[0]
  PIN NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.500 0.000 82.640 11.940 ;
    END
  END NN4END[10]
  PIN NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.340 0.000 84.480 15.000 ;
    END
  END NN4END[11]
  PIN NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.180 0.000 86.320 15.000 ;
    END
  END NN4END[12]
  PIN NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.020 0.000 88.160 7.210 ;
    END
  END NN4END[13]
  PIN NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.860 0.000 90.000 7.210 ;
    END
  END NN4END[14]
  PIN NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.240 0.000 91.380 5.850 ;
    END
  END NN4END[15]
  PIN NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.400 0.000 66.540 8.360 ;
    END
  END NN4END[1]
  PIN NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.240 0.000 68.380 13.870 ;
    END
  END NN4END[2]
  PIN NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.080 0.000 70.220 13.870 ;
    END
  END NN4END[3]
  PIN NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.920 0.000 72.060 15.680 ;
    END
  END NN4END[4]
  PIN NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.760 0.000 73.900 17.380 ;
    END
  END NN4END[5]
  PIN NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.140 0.000 75.280 15.680 ;
    END
  END NN4END[6]
  PIN NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.980 0.000 77.120 1.090 ;
    END
  END NN4END[7]
  PIN NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.820 0.000 78.960 7.210 ;
    END
  END NN4END[8]
  PIN NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.660 0.000 80.800 1.090 ;
    END
  END NN4END[9]
  PIN S1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.080 0.000 93.220 6.160 ;
    END
  END S1BEG[0]
  PIN S1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.920 0.000 95.060 4.490 ;
    END
  END S1BEG[1]
  PIN S1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.760 0.000 96.900 5.820 ;
    END
  END S1BEG[2]
  PIN S1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.600 0.000 98.740 8.880 ;
    END
  END S1BEG[3]
  PIN S2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.700 0.000 114.840 6.160 ;
    END
  END S2BEG[0]
  PIN S2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.540 0.000 116.680 8.880 ;
    END
  END S2BEG[1]
  PIN S2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.380 0.000 118.520 6.160 ;
    END
  END S2BEG[2]
  PIN S2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.760 0.000 119.900 8.880 ;
    END
  END S2BEG[3]
  PIN S2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.600 0.000 121.740 5.820 ;
    END
  END S2BEG[4]
  PIN S2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.440 0.000 123.580 8.880 ;
    END
  END S2BEG[5]
  PIN S2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.280 0.000 125.420 6.500 ;
    END
  END S2BEG[6]
  PIN S2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.120 0.000 127.260 8.880 ;
    END
  END S2BEG[7]
  PIN S2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.440 0.000 100.580 1.090 ;
    END
  END S2BEGb[0]
  PIN S2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.280 0.000 102.420 8.880 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.120 0.000 104.260 5.820 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.500 0.000 105.640 8.880 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.340 0.000 107.480 11.600 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.180 0.000 109.320 9.080 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.020 0.000 111.160 5.850 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.860 0.000 113.000 5.850 ;
    END
  END S2BEGb[7]
  PIN S4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.960 0.000 129.100 6.160 ;
    END
  END S4BEG[0]
  PIN S4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.900 0.000 147.040 1.090 ;
    END
  END S4BEG[10]
  PIN S4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.740 0.000 148.880 5.820 ;
    END
  END S4BEG[11]
  PIN S4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.120 0.000 150.260 8.880 ;
    END
  END S4BEG[12]
  PIN S4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.960 0.000 152.100 3.130 ;
    END
  END S4BEG[13]
  PIN S4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.800 0.000 153.940 8.880 ;
    END
  END S4BEG[14]
  PIN S4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.640 0.000 155.780 3.130 ;
    END
  END S4BEG[15]
  PIN S4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.800 0.000 130.940 8.880 ;
    END
  END S4BEG[1]
  PIN S4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.640 0.000 132.780 5.820 ;
    END
  END S4BEG[2]
  PIN S4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.480 0.000 134.620 8.540 ;
    END
  END S4BEG[3]
  PIN S4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.860 0.000 136.000 3.130 ;
    END
  END S4BEG[4]
  PIN S4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.700 0.000 137.840 9.220 ;
    END
  END S4BEG[5]
  PIN S4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.540 0.000 139.680 11.600 ;
    END
  END S4BEG[6]
  PIN S4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.380 0.000 141.520 8.880 ;
    END
  END S4BEG[7]
  PIN S4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.220 0.000 143.360 11.600 ;
    END
  END S4BEG[8]
  PIN S4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.060 0.000 145.200 11.600 ;
    END
  END S4BEG[9]
  PIN SS4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.480 0.000 157.620 4.490 ;
    END
  END SS4BEG[0]
  PIN SS4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.420 0.000 175.560 6.160 ;
    END
  END SS4BEG[10]
  PIN SS4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.260 0.000 177.400 6.160 ;
    END
  END SS4BEG[11]
  PIN SS4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.100 0.000 179.240 8.880 ;
    END
  END SS4BEG[12]
  PIN SS4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.480 0.000 180.620 6.360 ;
    END
  END SS4BEG[13]
  PIN SS4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.320 0.000 182.460 1.090 ;
    END
  END SS4BEG[14]
  PIN SS4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.160 0.000 184.300 11.600 ;
    END
  END SS4BEG[15]
  PIN SS4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.320 0.000 159.460 4.120 ;
    END
  END SS4BEG[1]
  PIN SS4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.160 0.000 161.300 1.090 ;
    END
  END SS4BEG[2]
  PIN SS4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.000 0.000 163.140 5.820 ;
    END
  END SS4BEG[3]
  PIN SS4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.380 0.000 164.520 8.740 ;
    END
  END SS4BEG[4]
  PIN SS4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.220 0.000 166.360 11.600 ;
    END
  END SS4BEG[5]
  PIN SS4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.060 0.000 168.200 9.220 ;
    END
  END SS4BEG[6]
  PIN SS4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.900 0.000 170.040 8.880 ;
    END
  END SS4BEG[7]
  PIN SS4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.740 0.000 171.880 11.600 ;
    END
  END SS4BEG[8]
  PIN SS4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.580 0.000 173.720 12.280 ;
    END
  END SS4BEG[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 40.090 5.200 41.690 32.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 110.835 5.200 112.435 32.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 181.580 5.200 183.180 32.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 75.465 5.200 77.065 32.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 146.210 5.200 147.810 32.880 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 0.085 217.580 32.725 ;
      LAYER met1 ;
        RECT 0.530 0.040 222.110 32.880 ;
      LAYER met2 ;
        RECT 0.560 38.750 5.400 39.850 ;
        RECT 6.100 38.750 16.440 39.850 ;
        RECT 0.560 31.640 16.440 38.750 ;
        RECT 17.140 31.640 27.480 39.850 ;
        RECT 28.180 31.640 38.520 39.850 ;
        RECT 39.220 31.640 50.020 39.850 ;
        RECT 50.720 31.640 61.060 39.850 ;
        RECT 61.760 31.640 72.100 39.850 ;
        RECT 72.800 31.640 83.140 39.850 ;
        RECT 83.840 31.640 94.640 39.850 ;
        RECT 95.340 31.640 105.680 39.850 ;
        RECT 106.380 34.670 116.720 39.850 ;
        RECT 117.420 34.670 127.760 39.850 ;
        RECT 106.380 31.640 127.760 34.670 ;
        RECT 128.460 31.640 139.260 39.850 ;
        RECT 139.960 31.640 150.300 39.850 ;
        RECT 151.000 31.640 161.340 39.850 ;
        RECT 162.040 31.640 172.380 39.850 ;
        RECT 173.080 31.640 183.880 39.850 ;
        RECT 184.580 31.640 194.920 39.850 ;
        RECT 195.620 31.640 205.960 39.850 ;
        RECT 206.660 31.640 217.000 39.850 ;
        RECT 217.700 31.640 222.080 39.850 ;
        RECT 0.560 23.100 222.080 31.640 ;
        RECT 0.560 20.720 216.080 23.100 ;
        RECT 0.560 17.660 3.560 20.720 ;
        RECT 0.560 15.280 1.720 17.660 ;
        RECT 1.040 0.010 1.720 15.280 ;
        RECT 2.420 0.010 3.560 17.660 ;
        RECT 4.260 17.660 212.400 20.720 ;
        RECT 4.260 17.320 62.440 17.660 ;
        RECT 4.260 0.010 5.400 17.320 ;
        RECT 6.100 15.480 62.440 17.320 ;
        RECT 6.100 15.280 60.600 15.480 ;
        RECT 6.100 12.420 51.860 15.280 ;
        RECT 6.100 12.220 25.180 12.420 ;
        RECT 6.100 11.880 17.820 12.220 ;
        RECT 6.100 9.840 9.080 11.880 ;
        RECT 6.100 0.010 7.240 9.840 ;
        RECT 7.940 0.010 9.080 9.840 ;
        RECT 9.780 9.500 17.820 11.880 ;
        RECT 9.780 6.780 15.980 9.500 ;
        RECT 9.780 6.130 14.600 6.780 ;
        RECT 9.780 0.010 10.920 6.130 ;
        RECT 11.620 3.380 14.600 6.130 ;
        RECT 11.620 0.010 12.760 3.380 ;
        RECT 13.460 0.010 14.600 3.380 ;
        RECT 15.300 0.010 15.980 6.780 ;
        RECT 16.680 0.010 17.820 9.500 ;
        RECT 18.520 9.500 21.500 12.220 ;
        RECT 18.520 0.010 19.660 9.500 ;
        RECT 20.360 0.010 21.500 9.500 ;
        RECT 22.200 3.720 25.180 12.220 ;
        RECT 22.200 0.010 23.340 3.720 ;
        RECT 24.040 0.010 25.180 3.720 ;
        RECT 25.880 12.220 51.860 12.420 ;
        RECT 25.880 9.840 28.860 12.220 ;
        RECT 25.880 0.010 27.020 9.840 ;
        RECT 27.720 0.010 28.860 9.840 ;
        RECT 29.560 11.880 51.860 12.220 ;
        RECT 29.560 9.500 33.920 11.880 ;
        RECT 29.560 0.010 30.240 9.500 ;
        RECT 30.940 1.370 33.920 9.500 ;
        RECT 30.940 0.010 32.080 1.370 ;
        RECT 32.780 0.010 33.920 1.370 ;
        RECT 34.620 9.840 43.120 11.880 ;
        RECT 34.620 6.440 39.440 9.840 ;
        RECT 34.620 0.010 35.760 6.440 ;
        RECT 36.460 0.010 37.600 6.440 ;
        RECT 38.300 0.010 39.440 6.440 ;
        RECT 40.140 5.450 43.120 9.840 ;
        RECT 40.140 0.010 41.280 5.450 ;
        RECT 41.980 0.010 43.120 5.450 ;
        RECT 43.820 9.500 51.860 11.880 ;
        RECT 43.820 6.780 48.180 9.500 ;
        RECT 43.820 6.300 46.340 6.780 ;
        RECT 43.820 0.010 44.960 6.300 ;
        RECT 45.660 0.010 46.340 6.300 ;
        RECT 47.040 0.010 48.180 6.780 ;
        RECT 48.880 3.720 51.860 9.500 ;
        RECT 48.880 0.010 50.020 3.720 ;
        RECT 50.720 0.010 51.860 3.720 ;
        RECT 52.560 12.220 57.380 15.280 ;
        RECT 52.560 0.010 53.700 12.220 ;
        RECT 54.400 0.010 55.540 12.220 ;
        RECT 56.240 0.010 57.380 12.220 ;
        RECT 58.080 10.180 60.600 15.280 ;
        RECT 58.080 0.010 59.220 10.180 ;
        RECT 59.920 0.010 60.600 10.180 ;
        RECT 61.300 0.010 62.440 15.480 ;
        RECT 63.140 0.010 64.280 17.660 ;
        RECT 64.980 15.960 73.480 17.660 ;
        RECT 64.980 14.150 71.640 15.960 ;
        RECT 64.980 8.640 67.960 14.150 ;
        RECT 64.980 0.010 66.120 8.640 ;
        RECT 66.820 0.010 67.960 8.640 ;
        RECT 68.660 0.010 69.800 14.150 ;
        RECT 70.500 0.010 71.640 14.150 ;
        RECT 72.340 0.010 73.480 15.960 ;
        RECT 74.180 15.960 210.560 17.660 ;
        RECT 74.180 0.010 74.860 15.960 ;
        RECT 75.560 15.280 210.560 15.960 ;
        RECT 75.560 12.220 84.060 15.280 ;
        RECT 75.560 7.490 82.220 12.220 ;
        RECT 75.560 1.370 78.540 7.490 ;
        RECT 75.560 0.010 76.700 1.370 ;
        RECT 77.400 0.010 78.540 1.370 ;
        RECT 79.240 1.370 82.220 7.490 ;
        RECT 79.240 0.010 80.380 1.370 ;
        RECT 81.080 0.010 82.220 1.370 ;
        RECT 82.920 0.010 84.060 12.220 ;
        RECT 84.760 0.010 85.900 15.280 ;
        RECT 86.600 12.560 187.560 15.280 ;
        RECT 86.600 11.880 173.300 12.560 ;
        RECT 86.600 9.160 107.060 11.880 ;
        RECT 86.600 7.490 98.320 9.160 ;
        RECT 86.600 0.010 87.740 7.490 ;
        RECT 88.440 0.010 89.580 7.490 ;
        RECT 90.280 6.440 98.320 7.490 ;
        RECT 90.280 6.130 92.800 6.440 ;
        RECT 90.280 0.010 90.960 6.130 ;
        RECT 91.660 0.010 92.800 6.130 ;
        RECT 93.500 6.100 98.320 6.440 ;
        RECT 93.500 4.770 96.480 6.100 ;
        RECT 93.500 0.010 94.640 4.770 ;
        RECT 95.340 0.010 96.480 4.770 ;
        RECT 97.180 0.010 98.320 6.100 ;
        RECT 99.020 1.370 102.000 9.160 ;
        RECT 99.020 0.010 100.160 1.370 ;
        RECT 100.860 0.010 102.000 1.370 ;
        RECT 102.700 6.100 105.220 9.160 ;
        RECT 102.700 0.010 103.840 6.100 ;
        RECT 104.540 0.010 105.220 6.100 ;
        RECT 105.920 0.010 107.060 9.160 ;
        RECT 107.760 9.500 139.260 11.880 ;
        RECT 107.760 9.360 137.420 9.500 ;
        RECT 107.760 0.010 108.900 9.360 ;
        RECT 109.600 9.160 137.420 9.360 ;
        RECT 109.600 6.440 116.260 9.160 ;
        RECT 109.600 6.130 114.420 6.440 ;
        RECT 109.600 0.010 110.740 6.130 ;
        RECT 111.440 0.010 112.580 6.130 ;
        RECT 113.280 0.010 114.420 6.130 ;
        RECT 115.120 0.010 116.260 6.440 ;
        RECT 116.960 6.440 119.480 9.160 ;
        RECT 116.960 0.010 118.100 6.440 ;
        RECT 118.800 0.010 119.480 6.440 ;
        RECT 120.180 6.100 123.160 9.160 ;
        RECT 120.180 0.010 121.320 6.100 ;
        RECT 122.020 0.010 123.160 6.100 ;
        RECT 123.860 6.780 126.840 9.160 ;
        RECT 123.860 0.010 125.000 6.780 ;
        RECT 125.700 0.010 126.840 6.780 ;
        RECT 127.540 6.440 130.520 9.160 ;
        RECT 127.540 0.010 128.680 6.440 ;
        RECT 129.380 0.010 130.520 6.440 ;
        RECT 131.220 8.820 137.420 9.160 ;
        RECT 131.220 6.100 134.200 8.820 ;
        RECT 131.220 0.010 132.360 6.100 ;
        RECT 133.060 0.010 134.200 6.100 ;
        RECT 134.900 3.410 137.420 8.820 ;
        RECT 134.900 0.010 135.580 3.410 ;
        RECT 136.280 0.010 137.420 3.410 ;
        RECT 138.120 0.010 139.260 9.500 ;
        RECT 139.960 9.160 142.940 11.880 ;
        RECT 139.960 0.010 141.100 9.160 ;
        RECT 141.800 0.010 142.940 9.160 ;
        RECT 143.640 0.010 144.780 11.880 ;
        RECT 145.480 9.160 165.940 11.880 ;
        RECT 145.480 6.100 149.840 9.160 ;
        RECT 145.480 1.370 148.460 6.100 ;
        RECT 145.480 0.010 146.620 1.370 ;
        RECT 147.320 0.010 148.460 1.370 ;
        RECT 149.160 0.010 149.840 6.100 ;
        RECT 150.540 3.410 153.520 9.160 ;
        RECT 150.540 0.010 151.680 3.410 ;
        RECT 152.380 0.010 153.520 3.410 ;
        RECT 154.220 9.020 165.940 9.160 ;
        RECT 154.220 6.100 164.100 9.020 ;
        RECT 154.220 4.770 162.720 6.100 ;
        RECT 154.220 3.410 157.200 4.770 ;
        RECT 154.220 0.010 155.360 3.410 ;
        RECT 156.060 0.010 157.200 3.410 ;
        RECT 157.900 4.400 162.720 4.770 ;
        RECT 157.900 0.010 159.040 4.400 ;
        RECT 159.740 1.370 162.720 4.400 ;
        RECT 159.740 0.010 160.880 1.370 ;
        RECT 161.580 0.010 162.720 1.370 ;
        RECT 163.420 0.010 164.100 6.100 ;
        RECT 164.800 0.010 165.940 9.020 ;
        RECT 166.640 9.500 171.460 11.880 ;
        RECT 166.640 0.010 167.780 9.500 ;
        RECT 168.480 9.160 171.460 9.500 ;
        RECT 168.480 0.010 169.620 9.160 ;
        RECT 170.320 0.010 171.460 9.160 ;
        RECT 172.160 0.010 173.300 11.880 ;
        RECT 174.000 11.880 187.560 12.560 ;
        RECT 174.000 9.160 183.880 11.880 ;
        RECT 174.000 6.440 178.820 9.160 ;
        RECT 174.000 0.010 175.140 6.440 ;
        RECT 175.840 0.010 176.980 6.440 ;
        RECT 177.680 0.010 178.820 6.440 ;
        RECT 179.520 6.640 183.880 9.160 ;
        RECT 179.520 0.010 180.200 6.640 ;
        RECT 180.900 1.370 183.880 6.640 ;
        RECT 180.900 0.010 182.040 1.370 ;
        RECT 182.740 0.010 183.880 1.370 ;
        RECT 184.580 1.080 187.560 11.880 ;
        RECT 184.580 0.010 185.720 1.080 ;
        RECT 186.420 0.010 187.560 1.080 ;
        RECT 188.260 12.220 210.560 15.280 ;
        RECT 188.260 12.080 201.820 12.220 ;
        RECT 188.260 11.880 199.980 12.080 ;
        RECT 188.260 9.840 196.300 11.880 ;
        RECT 188.260 9.500 194.460 9.840 ;
        RECT 188.260 6.780 191.240 9.500 ;
        RECT 188.260 0.010 189.400 6.780 ;
        RECT 190.100 0.010 191.240 6.780 ;
        RECT 191.940 6.100 194.460 9.500 ;
        RECT 191.940 0.010 193.080 6.100 ;
        RECT 193.780 0.010 194.460 6.100 ;
        RECT 195.160 0.010 196.300 9.840 ;
        RECT 197.000 10.180 199.980 11.880 ;
        RECT 197.000 0.010 198.140 10.180 ;
        RECT 198.840 0.010 199.980 10.180 ;
        RECT 200.680 0.010 201.820 12.080 ;
        RECT 202.520 9.840 210.560 12.220 ;
        RECT 202.520 6.780 207.340 9.840 ;
        RECT 202.520 6.440 205.500 6.780 ;
        RECT 202.520 0.010 203.660 6.440 ;
        RECT 204.360 0.010 205.500 6.440 ;
        RECT 206.200 0.010 207.340 6.780 ;
        RECT 208.040 8.170 210.560 9.840 ;
        RECT 208.040 0.010 208.720 8.170 ;
        RECT 209.420 0.010 210.560 8.170 ;
        RECT 211.260 0.010 212.400 17.660 ;
        RECT 213.100 14.940 216.080 20.720 ;
        RECT 213.100 0.010 214.240 14.940 ;
        RECT 214.940 0.010 216.080 14.940 ;
        RECT 216.780 20.380 222.080 23.100 ;
        RECT 216.780 0.010 217.920 20.380 ;
        RECT 218.620 18.000 222.080 20.380 ;
        RECT 218.620 0.010 219.760 18.000 ;
        RECT 220.460 15.620 222.080 18.000 ;
        RECT 220.460 0.010 221.600 15.620 ;
      LAYER met3 ;
        RECT 12.945 3.575 203.255 32.805 ;
  END
END N_term_single
MACRO N_term_single2
  CLASS BLOCK ;
  FOREIGN N_term_single2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 235.000 BY 40.000 ;
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.960 0.000 198.100 6.500 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.820 0.000 216.960 6.500 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.660 0.000 218.800 15.000 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.960 0.000 221.100 15.000 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.800 0.000 222.940 17.380 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.640 0.000 224.780 13.980 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.480 0.000 226.620 20.440 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.320 0.000 228.460 20.100 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.160 0.000 230.300 17.040 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.000 0.000 232.140 14.660 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.840 0.000 233.980 17.720 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.800 0.000 199.940 9.220 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.640 0.000 201.780 6.160 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.480 0.000 203.620 9.560 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.780 0.000 205.920 6.500 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.620 0.000 207.760 5.170 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.460 0.000 209.600 11.600 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.300 0.000 211.440 11.600 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.140 0.000 213.280 5.850 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.980 0.000 215.120 5.170 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.680 39.030 5.820 40.000 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.980 31.920 123.120 40.000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.940 31.920 135.080 40.000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.440 31.920 146.580 40.000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.400 31.920 158.540 40.000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.900 31.920 170.040 40.000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.860 31.920 182.000 40.000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.360 31.920 193.500 40.000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.320 31.920 205.460 40.000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.820 31.920 216.960 40.000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.780 31.920 228.920 40.000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.180 31.920 17.320 40.000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.140 31.920 29.280 40.000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.640 31.920 40.780 40.000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.600 31.920 52.740 40.000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.100 31.920 64.240 40.000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.060 31.920 76.200 40.000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.560 31.920 87.700 40.000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.520 29.200 99.660 40.000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.020 31.920 111.160 40.000 ;
    END
  END FrameStrobe_O[9]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.080 0.000 1.220 9.560 ;
    END
  END N1END[0]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.920 0.000 3.060 11.940 ;
    END
  END N1END[1]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.760 0.000 4.900 15.000 ;
    END
  END N1END[2]
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.600 0.000 6.740 14.660 ;
    END
  END N1END[3]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.620 0.000 23.760 6.500 ;
    END
  END N2END[0]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.460 0.000 25.600 3.810 ;
    END
  END N2END[1]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.300 0.000 27.440 9.560 ;
    END
  END N2END[2]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.140 0.000 29.280 3.100 ;
    END
  END N2END[3]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.980 0.000 31.120 9.220 ;
    END
  END N2END[4]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.280 0.000 33.420 11.940 ;
    END
  END N2END[5]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.120 0.000 35.260 5.000 ;
    END
  END N2END[6]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.960 0.000 37.100 11.940 ;
    END
  END N2END[7]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.440 0.000 8.580 6.160 ;
    END
  END N2MID[0]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.280 0.000 10.420 9.560 ;
    END
  END N2MID[1]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.120 0.000 12.260 11.600 ;
    END
  END N2MID[2]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.960 0.000 14.100 15.000 ;
    END
  END N2MID[3]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.800 0.000 15.940 15.000 ;
    END
  END N2MID[4]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.100 0.000 18.240 9.220 ;
    END
  END N2MID[5]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.940 0.000 20.080 11.940 ;
    END
  END N2MID[6]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.780 0.000 21.920 9.220 ;
    END
  END N2MID[7]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.800 0.000 38.940 6.160 ;
    END
  END N4END[0]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.660 0.000 57.800 6.500 ;
    END
  END N4END[10]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.500 0.000 59.640 15.000 ;
    END
  END N4END[11]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.340 0.000 61.480 15.000 ;
    END
  END N4END[12]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.180 0.000 63.320 13.870 ;
    END
  END N4END[13]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.480 0.000 65.620 11.600 ;
    END
  END N4END[14]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.320 0.000 67.460 15.000 ;
    END
  END N4END[15]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.640 0.000 40.780 6.160 ;
    END
  END N4END[1]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.480 0.000 42.620 1.090 ;
    END
  END N4END[2]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.320 0.000 44.460 9.560 ;
    END
  END N4END[3]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.160 0.000 46.300 9.900 ;
    END
  END N4END[4]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.460 0.000 48.600 11.600 ;
    END
  END N4END[5]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.300 0.000 50.440 11.600 ;
    END
  END N4END[6]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.140 0.000 52.280 6.160 ;
    END
  END N4END[7]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.980 0.000 54.120 9.420 ;
    END
  END N4END[8]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.820 0.000 55.960 11.940 ;
    END
  END N4END[9]
  PIN NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.160 0.000 69.300 7.210 ;
    END
  END NN4END[0]
  PIN NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.020 0.000 88.160 11.940 ;
    END
  END NN4END[10]
  PIN NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.860 0.000 90.000 15.000 ;
    END
  END NN4END[11]
  PIN NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.700 0.000 91.840 9.250 ;
    END
  END NN4END[12]
  PIN NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.540 0.000 93.680 7.210 ;
    END
  END NN4END[13]
  PIN NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.840 0.000 95.980 17.380 ;
    END
  END NN4END[14]
  PIN NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.680 0.000 97.820 5.640 ;
    END
  END NN4END[15]
  PIN NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.000 0.000 71.140 7.210 ;
    END
  END NN4END[1]
  PIN NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.840 0.000 72.980 14.320 ;
    END
  END NN4END[2]
  PIN NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.680 0.000 74.820 14.660 ;
    END
  END NN4END[3]
  PIN NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.520 0.000 76.660 5.820 ;
    END
  END NN4END[4]
  PIN NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.360 0.000 78.500 17.380 ;
    END
  END NN4END[5]
  PIN NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.660 0.000 80.800 4.490 ;
    END
  END NN4END[6]
  PIN NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.500 0.000 82.640 17.380 ;
    END
  END NN4END[7]
  PIN NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.340 0.000 84.480 17.380 ;
    END
  END NN4END[8]
  PIN NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.180 0.000 86.320 17.410 ;
    END
  END NN4END[9]
  PIN S1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.520 0.000 99.660 6.160 ;
    END
  END S1BEG[0]
  PIN S1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.360 0.000 101.500 6.160 ;
    END
  END S1BEG[1]
  PIN S1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.200 0.000 103.340 8.880 ;
    END
  END S1BEG[2]
  PIN S1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.040 0.000 105.180 6.160 ;
    END
  END S1BEG[3]
  PIN S2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.060 0.000 122.200 6.160 ;
    END
  END S2BEG[0]
  PIN S2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.900 0.000 124.040 6.160 ;
    END
  END S2BEG[1]
  PIN S2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.740 0.000 125.880 5.820 ;
    END
  END S2BEG[2]
  PIN S2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.040 0.000 128.180 8.880 ;
    END
  END S2BEG[3]
  PIN S2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.880 0.000 130.020 3.130 ;
    END
  END S2BEG[4]
  PIN S2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.720 0.000 131.860 8.880 ;
    END
  END S2BEG[5]
  PIN S2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.560 0.000 133.700 1.400 ;
    END
  END S2BEG[6]
  PIN S2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.400 0.000 135.540 8.880 ;
    END
  END S2BEG[7]
  PIN S2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.880 0.000 107.020 8.880 ;
    END
  END S2BEGb[0]
  PIN S2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.720 0.000 108.860 5.820 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.020 0.000 111.160 8.880 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.860 0.000 113.000 6.500 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.700 0.000 114.840 8.880 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.540 0.000 116.680 4.490 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.380 0.000 118.520 4.490 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.220 0.000 120.360 11.260 ;
    END
  END S2BEGb[7]
  PIN S4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.240 0.000 137.380 5.820 ;
    END
  END S4BEG[0]
  PIN S4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.100 0.000 156.240 6.160 ;
    END
  END S4BEG[10]
  PIN S4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.400 0.000 158.540 6.160 ;
    END
  END S4BEG[11]
  PIN S4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.240 0.000 160.380 5.820 ;
    END
  END S4BEG[12]
  PIN S4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.080 0.000 162.220 4.490 ;
    END
  END S4BEG[13]
  PIN S4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.920 0.000 164.060 6.160 ;
    END
  END S4BEG[14]
  PIN S4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.760 0.000 165.900 8.880 ;
    END
  END S4BEG[15]
  PIN S4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.080 0.000 139.220 9.560 ;
    END
  END S4BEG[1]
  PIN S4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.920 0.000 141.060 5.820 ;
    END
  END S4BEG[2]
  PIN S4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.220 0.000 143.360 8.880 ;
    END
  END S4BEG[3]
  PIN S4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.060 0.000 145.200 6.160 ;
    END
  END S4BEG[4]
  PIN S4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.900 0.000 147.040 8.880 ;
    END
  END S4BEG[5]
  PIN S4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.740 0.000 148.880 8.540 ;
    END
  END S4BEG[6]
  PIN S4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.580 0.000 150.720 11.600 ;
    END
  END S4BEG[7]
  PIN S4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.420 0.000 152.560 11.600 ;
    END
  END S4BEG[8]
  PIN S4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.260 0.000 154.400 4.660 ;
    END
  END S4BEG[9]
  PIN SS4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.600 0.000 167.740 8.880 ;
    END
  END SS4BEG[0]
  PIN SS4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.460 0.000 186.600 6.160 ;
    END
  END SS4BEG[10]
  PIN SS4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.300 0.000 188.440 6.160 ;
    END
  END SS4BEG[11]
  PIN SS4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.600 0.000 190.740 6.020 ;
    END
  END SS4BEG[12]
  PIN SS4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.440 0.000 192.580 1.090 ;
    END
  END SS4BEG[13]
  PIN SS4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.280 0.000 194.420 8.880 ;
    END
  END SS4BEG[14]
  PIN SS4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.120 0.000 196.260 11.600 ;
    END
  END SS4BEG[15]
  PIN SS4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.440 0.000 169.580 6.160 ;
    END
  END SS4BEG[1]
  PIN SS4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.280 0.000 171.420 9.900 ;
    END
  END SS4BEG[2]
  PIN SS4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.580 0.000 173.720 6.020 ;
    END
  END SS4BEG[3]
  PIN SS4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.420 0.000 175.560 8.880 ;
    END
  END SS4BEG[4]
  PIN SS4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.260 0.000 177.400 6.500 ;
    END
  END SS4BEG[5]
  PIN SS4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.100 0.000 179.240 8.880 ;
    END
  END SS4BEG[6]
  PIN SS4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.940 0.000 181.080 11.600 ;
    END
  END SS4BEG[7]
  PIN SS4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.780 0.000 182.920 8.880 ;
    END
  END SS4BEG[8]
  PIN SS4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.620 0.000 184.760 11.600 ;
    END
  END SS4BEG[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 42.045 5.200 43.645 32.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 116.695 5.200 118.295 32.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 191.350 5.200 192.950 32.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 79.370 5.200 80.970 32.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 154.025 5.200 155.625 32.880 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 0.085 229.080 32.725 ;
      LAYER met1 ;
        RECT 0.990 0.040 234.070 32.880 ;
      LAYER met2 ;
        RECT 1.020 38.750 5.400 39.850 ;
        RECT 6.100 38.750 16.900 39.850 ;
        RECT 1.020 31.640 16.900 38.750 ;
        RECT 17.600 31.640 28.860 39.850 ;
        RECT 29.560 31.640 40.360 39.850 ;
        RECT 41.060 31.640 52.320 39.850 ;
        RECT 53.020 31.640 63.820 39.850 ;
        RECT 64.520 31.640 75.780 39.850 ;
        RECT 76.480 31.640 87.280 39.850 ;
        RECT 87.980 31.640 99.240 39.850 ;
        RECT 1.020 28.920 99.240 31.640 ;
        RECT 99.940 31.640 110.740 39.850 ;
        RECT 111.440 31.640 122.700 39.850 ;
        RECT 123.400 31.640 134.660 39.850 ;
        RECT 135.360 31.640 146.160 39.850 ;
        RECT 146.860 31.640 158.120 39.850 ;
        RECT 158.820 31.640 169.620 39.850 ;
        RECT 170.320 31.640 181.580 39.850 ;
        RECT 182.280 31.640 193.080 39.850 ;
        RECT 193.780 31.640 205.040 39.850 ;
        RECT 205.740 31.640 216.540 39.850 ;
        RECT 217.240 31.640 228.500 39.850 ;
        RECT 229.200 31.640 234.040 39.850 ;
        RECT 99.940 28.920 234.040 31.640 ;
        RECT 1.020 20.720 234.040 28.920 ;
        RECT 1.020 17.690 226.200 20.720 ;
        RECT 1.020 17.660 85.900 17.690 ;
        RECT 1.020 15.280 78.080 17.660 ;
        RECT 1.020 12.220 4.480 15.280 ;
        RECT 1.020 9.840 2.640 12.220 ;
        RECT 1.500 0.010 2.640 9.840 ;
        RECT 3.340 0.010 4.480 12.220 ;
        RECT 5.180 14.940 13.680 15.280 ;
        RECT 5.180 0.010 6.320 14.940 ;
        RECT 7.020 11.880 13.680 14.940 ;
        RECT 7.020 9.840 11.840 11.880 ;
        RECT 7.020 6.440 10.000 9.840 ;
        RECT 7.020 0.010 8.160 6.440 ;
        RECT 8.860 0.010 10.000 6.440 ;
        RECT 10.700 0.010 11.840 9.840 ;
        RECT 12.540 0.010 13.680 11.880 ;
        RECT 14.380 0.010 15.520 15.280 ;
        RECT 16.220 12.220 59.220 15.280 ;
        RECT 16.220 9.500 19.660 12.220 ;
        RECT 16.220 0.010 17.820 9.500 ;
        RECT 18.520 0.010 19.660 9.500 ;
        RECT 20.360 9.840 33.000 12.220 ;
        RECT 20.360 9.500 27.020 9.840 ;
        RECT 20.360 0.010 21.500 9.500 ;
        RECT 22.200 6.780 27.020 9.500 ;
        RECT 22.200 0.010 23.340 6.780 ;
        RECT 24.040 4.090 27.020 6.780 ;
        RECT 24.040 0.010 25.180 4.090 ;
        RECT 25.880 0.010 27.020 4.090 ;
        RECT 27.720 9.500 33.000 9.840 ;
        RECT 27.720 3.380 30.700 9.500 ;
        RECT 27.720 0.010 28.860 3.380 ;
        RECT 29.560 0.010 30.700 3.380 ;
        RECT 31.400 0.010 33.000 9.500 ;
        RECT 33.700 5.280 36.680 12.220 ;
        RECT 33.700 0.010 34.840 5.280 ;
        RECT 35.540 0.010 36.680 5.280 ;
        RECT 37.380 11.880 55.540 12.220 ;
        RECT 37.380 10.180 48.180 11.880 ;
        RECT 37.380 9.840 45.880 10.180 ;
        RECT 37.380 6.440 44.040 9.840 ;
        RECT 37.380 0.010 38.520 6.440 ;
        RECT 39.220 0.010 40.360 6.440 ;
        RECT 41.060 1.370 44.040 6.440 ;
        RECT 41.060 0.010 42.200 1.370 ;
        RECT 42.900 0.010 44.040 1.370 ;
        RECT 44.740 0.010 45.880 9.840 ;
        RECT 46.580 0.010 48.180 10.180 ;
        RECT 48.880 0.010 50.020 11.880 ;
        RECT 50.720 9.700 55.540 11.880 ;
        RECT 50.720 6.440 53.700 9.700 ;
        RECT 50.720 0.010 51.860 6.440 ;
        RECT 52.560 0.010 53.700 6.440 ;
        RECT 54.400 0.010 55.540 9.700 ;
        RECT 56.240 6.780 59.220 12.220 ;
        RECT 56.240 0.010 57.380 6.780 ;
        RECT 58.080 0.010 59.220 6.780 ;
        RECT 59.920 0.010 61.060 15.280 ;
        RECT 61.760 14.150 67.040 15.280 ;
        RECT 61.760 0.010 62.900 14.150 ;
        RECT 63.600 11.880 67.040 14.150 ;
        RECT 63.600 0.010 65.200 11.880 ;
        RECT 65.900 0.010 67.040 11.880 ;
        RECT 67.740 14.940 78.080 15.280 ;
        RECT 67.740 14.600 74.400 14.940 ;
        RECT 67.740 7.490 72.560 14.600 ;
        RECT 67.740 0.010 68.880 7.490 ;
        RECT 69.580 0.010 70.720 7.490 ;
        RECT 71.420 0.010 72.560 7.490 ;
        RECT 73.260 0.010 74.400 14.600 ;
        RECT 75.100 6.100 78.080 14.940 ;
        RECT 75.100 0.010 76.240 6.100 ;
        RECT 76.940 0.010 78.080 6.100 ;
        RECT 78.780 4.770 82.220 17.660 ;
        RECT 78.780 0.010 80.380 4.770 ;
        RECT 81.080 0.010 82.220 4.770 ;
        RECT 82.920 0.010 84.060 17.660 ;
        RECT 84.760 0.010 85.900 17.660 ;
        RECT 86.600 17.660 226.200 17.690 ;
        RECT 86.600 15.280 95.560 17.660 ;
        RECT 86.600 12.220 89.580 15.280 ;
        RECT 86.600 0.010 87.740 12.220 ;
        RECT 88.440 0.010 89.580 12.220 ;
        RECT 90.280 9.530 95.560 15.280 ;
        RECT 90.280 0.010 91.420 9.530 ;
        RECT 92.120 7.490 95.560 9.530 ;
        RECT 92.120 0.010 93.260 7.490 ;
        RECT 93.960 0.010 95.560 7.490 ;
        RECT 96.260 15.280 222.520 17.660 ;
        RECT 96.260 11.880 218.380 15.280 ;
        RECT 96.260 11.540 150.300 11.880 ;
        RECT 96.260 9.160 119.940 11.540 ;
        RECT 96.260 6.440 102.920 9.160 ;
        RECT 96.260 5.920 99.240 6.440 ;
        RECT 96.260 0.010 97.400 5.920 ;
        RECT 98.100 0.010 99.240 5.920 ;
        RECT 99.940 0.010 101.080 6.440 ;
        RECT 101.780 0.010 102.920 6.440 ;
        RECT 103.620 6.440 106.600 9.160 ;
        RECT 103.620 0.010 104.760 6.440 ;
        RECT 105.460 0.010 106.600 6.440 ;
        RECT 107.300 6.100 110.740 9.160 ;
        RECT 107.300 0.010 108.440 6.100 ;
        RECT 109.140 0.010 110.740 6.100 ;
        RECT 111.440 6.780 114.420 9.160 ;
        RECT 111.440 0.010 112.580 6.780 ;
        RECT 113.280 0.010 114.420 6.780 ;
        RECT 115.120 4.770 119.940 9.160 ;
        RECT 115.120 0.010 116.260 4.770 ;
        RECT 116.960 0.010 118.100 4.770 ;
        RECT 118.800 0.010 119.940 4.770 ;
        RECT 120.640 9.840 150.300 11.540 ;
        RECT 120.640 9.160 138.800 9.840 ;
        RECT 120.640 6.440 127.760 9.160 ;
        RECT 120.640 0.010 121.780 6.440 ;
        RECT 122.480 0.010 123.620 6.440 ;
        RECT 124.320 6.100 127.760 6.440 ;
        RECT 124.320 0.010 125.460 6.100 ;
        RECT 126.160 0.010 127.760 6.100 ;
        RECT 128.460 3.410 131.440 9.160 ;
        RECT 128.460 0.010 129.600 3.410 ;
        RECT 130.300 0.010 131.440 3.410 ;
        RECT 132.140 1.680 135.120 9.160 ;
        RECT 132.140 0.010 133.280 1.680 ;
        RECT 133.980 0.010 135.120 1.680 ;
        RECT 135.820 6.100 138.800 9.160 ;
        RECT 135.820 0.010 136.960 6.100 ;
        RECT 137.660 0.010 138.800 6.100 ;
        RECT 139.500 9.160 150.300 9.840 ;
        RECT 139.500 6.100 142.940 9.160 ;
        RECT 139.500 0.010 140.640 6.100 ;
        RECT 141.340 0.010 142.940 6.100 ;
        RECT 143.640 6.440 146.620 9.160 ;
        RECT 143.640 0.010 144.780 6.440 ;
        RECT 145.480 0.010 146.620 6.440 ;
        RECT 147.320 8.820 150.300 9.160 ;
        RECT 147.320 0.010 148.460 8.820 ;
        RECT 149.160 0.010 150.300 8.820 ;
        RECT 151.000 0.010 152.140 11.880 ;
        RECT 152.840 10.180 180.660 11.880 ;
        RECT 152.840 9.160 171.000 10.180 ;
        RECT 152.840 6.440 165.480 9.160 ;
        RECT 152.840 4.940 155.820 6.440 ;
        RECT 152.840 0.010 153.980 4.940 ;
        RECT 154.680 0.010 155.820 4.940 ;
        RECT 156.520 0.010 158.120 6.440 ;
        RECT 158.820 6.100 163.640 6.440 ;
        RECT 158.820 0.010 159.960 6.100 ;
        RECT 160.660 4.770 163.640 6.100 ;
        RECT 160.660 0.010 161.800 4.770 ;
        RECT 162.500 0.010 163.640 4.770 ;
        RECT 164.340 0.010 165.480 6.440 ;
        RECT 166.180 0.010 167.320 9.160 ;
        RECT 168.020 6.440 171.000 9.160 ;
        RECT 168.020 0.010 169.160 6.440 ;
        RECT 169.860 0.010 171.000 6.440 ;
        RECT 171.700 9.160 180.660 10.180 ;
        RECT 171.700 6.300 175.140 9.160 ;
        RECT 171.700 0.010 173.300 6.300 ;
        RECT 174.000 0.010 175.140 6.300 ;
        RECT 175.840 6.780 178.820 9.160 ;
        RECT 175.840 0.010 176.980 6.780 ;
        RECT 177.680 0.010 178.820 6.780 ;
        RECT 179.520 0.010 180.660 9.160 ;
        RECT 181.360 9.160 184.340 11.880 ;
        RECT 181.360 0.010 182.500 9.160 ;
        RECT 183.200 0.010 184.340 9.160 ;
        RECT 185.040 9.160 195.840 11.880 ;
        RECT 185.040 6.440 194.000 9.160 ;
        RECT 185.040 0.010 186.180 6.440 ;
        RECT 186.880 0.010 188.020 6.440 ;
        RECT 188.720 6.300 194.000 6.440 ;
        RECT 188.720 0.010 190.320 6.300 ;
        RECT 191.020 1.370 194.000 6.300 ;
        RECT 191.020 0.010 192.160 1.370 ;
        RECT 192.860 0.010 194.000 1.370 ;
        RECT 194.700 0.010 195.840 9.160 ;
        RECT 196.540 9.840 209.180 11.880 ;
        RECT 196.540 9.500 203.200 9.840 ;
        RECT 196.540 6.780 199.520 9.500 ;
        RECT 196.540 0.010 197.680 6.780 ;
        RECT 198.380 0.010 199.520 6.780 ;
        RECT 200.220 6.440 203.200 9.500 ;
        RECT 200.220 0.010 201.360 6.440 ;
        RECT 202.060 0.010 203.200 6.440 ;
        RECT 203.900 6.780 209.180 9.840 ;
        RECT 203.900 0.010 205.500 6.780 ;
        RECT 206.200 5.450 209.180 6.780 ;
        RECT 206.200 0.010 207.340 5.450 ;
        RECT 208.040 0.010 209.180 5.450 ;
        RECT 209.880 0.010 211.020 11.880 ;
        RECT 211.720 6.780 218.380 11.880 ;
        RECT 211.720 6.130 216.540 6.780 ;
        RECT 211.720 0.010 212.860 6.130 ;
        RECT 213.560 5.450 216.540 6.130 ;
        RECT 213.560 0.010 214.700 5.450 ;
        RECT 215.400 0.010 216.540 5.450 ;
        RECT 217.240 0.010 218.380 6.780 ;
        RECT 219.080 0.010 220.680 15.280 ;
        RECT 221.380 0.010 222.520 15.280 ;
        RECT 223.220 14.260 226.200 17.660 ;
        RECT 223.220 0.010 224.360 14.260 ;
        RECT 225.060 0.010 226.200 14.260 ;
        RECT 226.900 20.380 234.040 20.720 ;
        RECT 226.900 0.010 228.040 20.380 ;
        RECT 228.740 18.000 234.040 20.380 ;
        RECT 228.740 17.320 233.560 18.000 ;
        RECT 228.740 0.010 229.880 17.320 ;
        RECT 230.580 14.940 233.560 17.320 ;
        RECT 230.580 0.010 231.720 14.940 ;
        RECT 232.420 0.010 233.560 14.940 ;
      LAYER met3 ;
        RECT 7.885 3.575 212.455 32.805 ;
      LAYER met4 ;
        RECT 96.895 5.200 116.295 32.880 ;
  END
END N_term_single2
MACRO RAM_IO
  CLASS BLOCK ;
  FOREIGN RAM_IO ;
  ORIGIN 0.000 0.000 ;
  SIZE 125.000 BY 223.115 ;
  PIN Config_accessC_bit0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.850 45.750 125.000 46.050 ;
    END
  END Config_accessC_bit0
  PIN Config_accessC_bit1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 115.830 48.470 125.000 48.770 ;
    END
  END Config_accessC_bit1
  PIN Config_accessC_bit2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 112.150 51.190 125.000 51.490 ;
    END
  END Config_accessC_bit2
  PIN Config_accessC_bit3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.290 53.910 125.000 54.210 ;
    END
  END Config_accessC_bit3
  PIN E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.510 7.910 84.810 ;
    END
  END E1END[0]
  PIN E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.870 20.330 86.170 ;
    END
  END E1END[1]
  PIN E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.910 20.790 88.210 ;
    END
  END E1END[2]
  PIN E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.270 14.350 89.570 ;
    END
  END E1END[3]
  PIN E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.910 19.410 105.210 ;
    END
  END E2END[0]
  PIN E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.950 15.730 107.250 ;
    END
  END E2END[1]
  PIN E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.310 20.790 108.610 ;
    END
  END E2END[2]
  PIN E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.350 7.050 110.650 ;
    END
  END E2END[3]
  PIN E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.390 8.370 112.690 ;
    END
  END E2END[4]
  PIN E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.750 13.950 114.050 ;
    END
  END E2END[5]
  PIN E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.790 18.030 116.090 ;
    END
  END E2END[6]
  PIN E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.150 19.870 117.450 ;
    END
  END E2END[7]
  PIN E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.310 17.570 91.610 ;
    END
  END E2MID[0]
  PIN E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.670 6.990 92.970 ;
    END
  END E2MID[1]
  PIN E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.710 20.330 95.010 ;
    END
  END E2MID[2]
  PIN E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.070 20.330 96.370 ;
    END
  END E2MID[3]
  PIN E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.110 19.410 98.410 ;
    END
  END E2MID[4]
  PIN E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.150 19.870 100.450 ;
    END
  END E2MID[5]
  PIN E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.510 17.570 101.810 ;
    END
  END E2MID[6]
  PIN E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.550 27.690 103.850 ;
    END
  END E2MID[7]
  PIN E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.070 6.990 147.370 ;
    END
  END E6END[0]
  PIN E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.070 6.990 164.370 ;
    END
  END E6END[10]
  PIN E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.110 16.190 166.410 ;
    END
  END E6END[11]
  PIN E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.430 11.130 148.730 ;
    END
  END E6END[1]
  PIN E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 150.470 13.430 150.770 ;
    END
  END E6END[2]
  PIN E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.830 13.890 152.130 ;
    END
  END E6END[3]
  PIN E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.870 2.390 154.170 ;
    END
  END E6END[4]
  PIN E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.910 19.240 156.210 ;
    END
  END E6END[5]
  PIN E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.270 19.870 157.570 ;
    END
  END E6END[6]
  PIN E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.310 20.330 159.610 ;
    END
  END E6END[7]
  PIN E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.670 19.870 160.970 ;
    END
  END E6END[8]
  PIN E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.710 17.110 163.010 ;
    END
  END E6END[9]
  PIN EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.190 6.990 119.490 ;
    END
  END EE4END[0]
  PIN EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.190 20.330 136.490 ;
    END
  END EE4END[10]
  PIN EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.230 6.990 138.530 ;
    END
  END EE4END[11]
  PIN EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.270 16.190 140.570 ;
    END
  END EE4END[12]
  PIN EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.630 20.330 141.930 ;
    END
  END EE4END[13]
  PIN EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.670 6.530 143.970 ;
    END
  END EE4END[14]
  PIN EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.030 14.350 145.330 ;
    END
  END EE4END[15]
  PIN EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.550 18.950 120.850 ;
    END
  END EE4END[1]
  PIN EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.590 20.330 122.890 ;
    END
  END EE4END[2]
  PIN EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.950 17.110 124.250 ;
    END
  END EE4END[3]
  PIN EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.990 20.330 126.290 ;
    END
  END EE4END[4]
  PIN EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.030 20.330 128.330 ;
    END
  END EE4END[5]
  PIN EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.390 13.950 129.690 ;
    END
  END EE4END[6]
  PIN EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.430 18.950 131.730 ;
    END
  END EE4END[7]
  PIN EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.790 20.330 133.090 ;
    END
  END EE4END[8]
  PIN EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.830 20.330 135.130 ;
    END
  END EE4END[9]
  PIN FAB2RAM_A0_O0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.850 79.070 125.000 79.370 ;
    END
  END FAB2RAM_A0_O0
  PIN FAB2RAM_A0_O1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.410 81.790 125.000 82.090 ;
    END
  END FAB2RAM_A0_O1
  PIN FAB2RAM_A0_O2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 113.530 85.190 125.000 85.490 ;
    END
  END FAB2RAM_A0_O2
  PIN FAB2RAM_A0_O3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 104.330 87.910 125.000 88.210 ;
    END
  END FAB2RAM_A0_O3
  PIN FAB2RAM_A1_O0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 115.370 68.190 125.000 68.490 ;
    END
  END FAB2RAM_A1_O0
  PIN FAB2RAM_A1_O1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 112.150 70.910 125.000 71.210 ;
    END
  END FAB2RAM_A1_O1
  PIN FAB2RAM_A1_O2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.630 73.630 125.000 73.930 ;
    END
  END FAB2RAM_A1_O2
  PIN FAB2RAM_A1_O3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 104.330 76.350 125.000 76.650 ;
    END
  END FAB2RAM_A1_O3
  PIN FAB2RAM_C_O0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.470 57.310 125.000 57.610 ;
    END
  END FAB2RAM_C_O0
  PIN FAB2RAM_C_O1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 117.150 60.030 125.000 60.330 ;
    END
  END FAB2RAM_C_O1
  PIN FAB2RAM_C_O2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.630 62.750 125.000 63.050 ;
    END
  END FAB2RAM_C_O2
  PIN FAB2RAM_C_O3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.630 65.470 125.000 65.770 ;
    END
  END FAB2RAM_C_O3
  PIN FAB2RAM_D0_O0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 115.370 123.950 125.000 124.250 ;
    END
  END FAB2RAM_D0_O0
  PIN FAB2RAM_D0_O1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.850 126.670 125.000 126.970 ;
    END
  END FAB2RAM_D0_O1
  PIN FAB2RAM_D0_O2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 110.310 129.390 125.000 129.690 ;
    END
  END FAB2RAM_D0_O2
  PIN FAB2RAM_D0_O3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.850 132.110 125.000 132.410 ;
    END
  END FAB2RAM_D0_O3
  PIN FAB2RAM_D1_O0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 110.770 113.070 125.000 113.370 ;
    END
  END FAB2RAM_D1_O0
  PIN FAB2RAM_D1_O1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.630 115.790 125.000 116.090 ;
    END
  END FAB2RAM_D1_O1
  PIN FAB2RAM_D1_O2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.870 118.510 125.000 118.810 ;
    END
  END FAB2RAM_D1_O2
  PIN FAB2RAM_D1_O3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.870 121.230 125.000 121.530 ;
    END
  END FAB2RAM_D1_O3
  PIN FAB2RAM_D2_O0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.870 101.510 125.000 101.810 ;
    END
  END FAB2RAM_D2_O0
  PIN FAB2RAM_D2_O1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.870 104.230 125.000 104.530 ;
    END
  END FAB2RAM_D2_O1
  PIN FAB2RAM_D2_O2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.410 106.950 125.000 107.250 ;
    END
  END FAB2RAM_D2_O2
  PIN FAB2RAM_D2_O3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 102.490 109.670 125.000 109.970 ;
    END
  END FAB2RAM_D2_O3
  PIN FAB2RAM_D3_O0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 104.330 90.630 125.000 90.930 ;
    END
  END FAB2RAM_D3_O0
  PIN FAB2RAM_D3_O1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.930 93.350 125.000 93.650 ;
    END
  END FAB2RAM_D3_O1
  PIN FAB2RAM_D3_O2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.410 96.070 125.000 96.370 ;
    END
  END FAB2RAM_D3_O2
  PIN FAB2RAM_D3_O3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.630 98.790 125.000 99.090 ;
    END
  END FAB2RAM_D3_O3
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.150 13.890 168.450 ;
    END
  END FrameData[0]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.150 8.830 185.450 ;
    END
  END FrameData[10]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.190 14.810 187.490 ;
    END
  END FrameData[11]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 188.550 14.350 188.850 ;
    END
  END FrameData[12]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.590 20.330 190.890 ;
    END
  END FrameData[13]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.950 16.190 192.250 ;
    END
  END FrameData[14]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.990 19.410 194.290 ;
    END
  END FrameData[15]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.030 14.410 196.330 ;
    END
  END FrameData[16]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.390 20.330 197.690 ;
    END
  END FrameData[17]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.430 20.850 199.730 ;
    END
  END FrameData[18]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.790 19.870 201.090 ;
    END
  END FrameData[19]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 169.510 14.350 169.810 ;
    END
  END FrameData[1]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.830 6.530 203.130 ;
    END
  END FrameData[20]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.190 7.450 204.490 ;
    END
  END FrameData[21]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.230 14.350 206.530 ;
    END
  END FrameData[22]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.590 20.330 207.890 ;
    END
  END FrameData[23]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.630 6.990 209.930 ;
    END
  END FrameData[24]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 211.670 18.950 211.970 ;
    END
  END FrameData[25]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.030 16.190 213.330 ;
    END
  END FrameData[26]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.070 15.270 215.370 ;
    END
  END FrameData[27]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.430 17.110 216.730 ;
    END
  END FrameData[28]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 218.470 19.870 218.770 ;
    END
  END FrameData[29]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.550 20.330 171.850 ;
    END
  END FrameData[2]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.830 20.330 220.130 ;
    END
  END FrameData[30]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.870 17.110 222.170 ;
    END
  END FrameData[31]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.910 28.610 173.210 ;
    END
  END FrameData[3]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.950 27.690 175.250 ;
    END
  END FrameData[4]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.310 19.870 176.610 ;
    END
  END FrameData[5]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.350 17.570 178.650 ;
    END
  END FrameData[6]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.710 17.570 180.010 ;
    END
  END FrameData[7]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 181.750 8.370 182.050 ;
    END
  END FrameData[8]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.790 20.790 184.090 ;
    END
  END FrameData[9]
  PIN FrameData_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.690 134.830 125.000 135.130 ;
    END
  END FrameData_O[0]
  PIN FrameData_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 115.370 162.710 125.000 163.010 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 115.830 165.430 125.000 165.730 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 112.150 168.830 125.000 169.130 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 117.210 171.550 125.000 171.850 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.850 174.270 125.000 174.570 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 115.830 176.990 125.000 177.290 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 115.370 179.710 125.000 180.010 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 115.830 182.430 125.000 182.730 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 115.370 185.150 125.000 185.450 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 117.210 187.870 125.000 188.170 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.630 137.550 125.000 137.850 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 115.830 190.590 125.000 190.890 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 115.370 193.310 125.000 193.610 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 115.370 196.710 125.000 197.010 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 115.830 199.430 125.000 199.730 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 115.370 202.150 125.000 202.450 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 115.830 204.870 125.000 205.170 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 115.370 207.590 125.000 207.890 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 115.370 210.310 125.000 210.610 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 115.830 213.030 125.000 213.330 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.230 215.750 125.000 216.050 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 110.770 140.950 125.000 141.250 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.930 218.470 125.000 218.770 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 107.090 221.190 125.000 221.490 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.630 143.670 125.000 143.970 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 115.830 146.390 125.000 146.690 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 117.210 149.110 125.000 149.410 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 113.990 151.830 125.000 152.130 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 117.840 154.550 125.000 154.850 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.470 157.270 125.000 157.570 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.470 159.990 125.000 160.290 ;
    END
  END FrameData_O[9]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.600 0.000 98.740 6.160 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.940 0.000 112.080 6.160 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.320 0.000 113.460 28.970 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.700 0.000 114.840 18.400 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.080 0.000 116.220 18.060 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.460 0.000 117.600 17.040 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.840 0.000 118.980 20.440 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.220 0.000 120.360 20.100 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.600 0.000 121.740 17.200 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.980 0.000 123.120 19.420 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.360 0.000 124.500 1.090 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.980 0.000 100.120 5.850 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.360 0.000 101.500 5.170 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.740 0.000 102.880 9.220 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.120 0.000 104.260 17.040 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.500 0.000 105.640 15.000 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.880 0.000 107.020 4.120 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.800 0.000 107.940 17.380 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.180 0.000 109.320 6.500 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.560 0.000 110.700 22.480 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.140 217.220 98.280 223.115 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.940 208.720 112.080 223.115 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.320 211.440 113.460 223.115 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.700 211.580 114.840 223.115 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.080 218.240 116.220 223.115 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.460 211.780 117.600 223.115 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.840 219.260 118.980 223.115 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.220 203.280 120.360 223.115 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.600 205.320 121.740 223.115 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.980 211.960 123.120 223.115 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.360 217.220 124.500 223.115 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.520 215.830 99.660 223.115 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.900 218.380 101.040 223.115 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.280 214.470 102.420 223.115 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.660 214.470 103.800 223.115 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.040 200.900 105.180 223.115 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.420 214.470 106.560 223.115 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.800 214.470 107.940 223.115 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.180 210.390 109.320 223.115 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.560 206.930 110.700 223.115 ;
    END
  END FrameStrobe_O[9]
  PIN N1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.620 217.220 0.760 223.115 ;
    END
  END N1BEG[0]
  PIN N1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.540 213.820 1.680 223.115 ;
    END
  END N1BEG[1]
  PIN N1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.920 219.600 3.060 223.115 ;
    END
  END N1BEG[2]
  PIN N1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.300 206.340 4.440 223.115 ;
    END
  END N1BEG[3]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.620 0.000 0.760 6.160 ;
    END
  END N1END[0]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.540 0.000 1.680 20.440 ;
    END
  END N1END[1]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.920 0.000 3.060 9.560 ;
    END
  END N1END[2]
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.300 0.000 4.440 6.500 ;
    END
  END N1END[3]
  PIN N2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.680 220.280 5.820 223.115 ;
    END
  END N2BEG[0]
  PIN N2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.060 220.620 7.200 223.115 ;
    END
  END N2BEG[1]
  PIN N2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.440 205.840 8.580 223.115 ;
    END
  END N2BEG[2]
  PIN N2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.820 210.600 9.960 223.115 ;
    END
  END N2BEG[3]
  PIN N2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.200 216.510 11.340 223.115 ;
    END
  END N2BEG[4]
  PIN N2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.580 209.060 12.720 223.115 ;
    END
  END N2BEG[5]
  PIN N2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.960 216.340 14.100 223.115 ;
    END
  END N2BEG[6]
  PIN N2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.340 218.240 15.480 223.115 ;
    END
  END N2BEG[7]
  PIN N2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.720 209.240 16.860 223.115 ;
    END
  END N2BEGb[0]
  PIN N2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.100 201.920 18.240 223.115 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.480 213.320 19.620 223.115 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.860 214.470 21.000 223.115 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.240 206.340 22.380 223.115 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.620 215.830 23.760 223.115 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.000 215.830 25.140 223.115 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.380 219.940 26.520 223.115 ;
    END
  END N2BEGb[7]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.720 0.000 16.860 6.160 ;
    END
  END N2END[0]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.100 0.000 18.240 2.420 ;
    END
  END N2END[1]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.020 0.000 19.160 3.780 ;
    END
  END N2END[2]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.400 0.000 20.540 15.000 ;
    END
  END N2END[3]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.780 0.000 21.920 13.870 ;
    END
  END N2END[4]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.160 0.000 23.300 14.320 ;
    END
  END N2END[5]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.540 0.000 24.680 6.160 ;
    END
  END N2END[6]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.920 0.000 26.060 9.560 ;
    END
  END N2END[7]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.680 0.000 5.820 9.900 ;
    END
  END N2MID[0]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.060 0.000 7.200 4.800 ;
    END
  END N2MID[1]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.440 0.000 8.580 8.880 ;
    END
  END N2MID[2]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.820 0.000 9.960 13.980 ;
    END
  END N2MID[3]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.200 0.000 11.340 2.760 ;
    END
  END N2MID[4]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.580 0.000 12.720 15.340 ;
    END
  END N2MID[5]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.960 0.000 14.100 3.440 ;
    END
  END N2MID[6]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.340 0.000 15.480 6.840 ;
    END
  END N2MID[7]
  PIN N4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.760 204.640 27.900 223.115 ;
    END
  END N4BEG[0]
  PIN N4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.100 216.510 41.240 223.115 ;
    END
  END N4BEG[10]
  PIN N4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.480 218.550 42.620 223.115 ;
    END
  END N4BEG[11]
  PIN N4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.860 218.550 44.000 223.115 ;
    END
  END N4BEG[12]
  PIN N4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.240 214.500 45.380 223.115 ;
    END
  END N4BEG[13]
  PIN N4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.620 209.240 46.760 223.115 ;
    END
  END N4BEG[14]
  PIN N4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.000 210.390 48.140 223.115 ;
    END
  END N4BEG[15]
  PIN N4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.140 206.340 29.280 223.115 ;
    END
  END N4BEG[1]
  PIN N4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.520 205.160 30.660 223.115 ;
    END
  END N4BEG[2]
  PIN N4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.900 202.600 32.040 223.115 ;
    END
  END N4BEG[3]
  PIN N4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.820 202.940 32.960 223.115 ;
    END
  END N4BEG[4]
  PIN N4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.200 206.930 34.340 223.115 ;
    END
  END N4BEG[5]
  PIN N4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.580 176.420 35.720 223.115 ;
    END
  END N4BEG[6]
  PIN N4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.960 173.700 37.100 223.115 ;
    END
  END N4BEG[7]
  PIN N4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.340 203.800 38.480 223.115 ;
    END
  END N4BEG[8]
  PIN N4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.720 211.960 39.860 223.115 ;
    END
  END N4BEG[9]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.300 0.000 27.440 3.810 ;
    END
  END N4END[0]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.640 0.000 40.780 24.210 ;
    END
  END N4END[10]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.020 0.000 42.160 3.780 ;
    END
  END N4END[11]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.400 0.000 43.540 4.660 ;
    END
  END N4END[12]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.780 0.000 44.920 12.280 ;
    END
  END N4END[13]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.160 0.000 46.300 13.870 ;
    END
  END N4END[14]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.540 0.000 47.680 16.700 ;
    END
  END N4END[15]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.680 0.000 28.820 7.210 ;
    END
  END N4END[1]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.060 0.000 30.200 13.980 ;
    END
  END N4END[2]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.440 0.000 31.580 15.340 ;
    END
  END N4END[3]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.820 0.000 32.960 13.870 ;
    END
  END N4END[4]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.200 0.000 34.340 7.210 ;
    END
  END N4END[5]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.580 0.000 35.720 36.620 ;
    END
  END N4END[6]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.500 0.000 36.640 15.000 ;
    END
  END N4END[7]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.880 0.000 38.020 13.870 ;
    END
  END N4END[8]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.260 0.000 39.400 18.770 ;
    END
  END N4END[9]
  PIN RAM2FAB_D0_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 107.550 34.870 125.000 35.170 ;
    END
  END RAM2FAB_D0_I0
  PIN RAM2FAB_D0_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.410 37.590 125.000 37.890 ;
    END
  END RAM2FAB_D0_I1
  PIN RAM2FAB_D0_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 110.310 40.310 125.000 40.610 ;
    END
  END RAM2FAB_D0_I2
  PIN RAM2FAB_D0_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.410 43.030 125.000 43.330 ;
    END
  END RAM2FAB_D0_I3
  PIN RAM2FAB_D1_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.390 23.310 125.000 23.610 ;
    END
  END RAM2FAB_D1_I0
  PIN RAM2FAB_D1_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 88.020 26.030 125.000 26.330 ;
    END
  END RAM2FAB_D1_I1
  PIN RAM2FAB_D1_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 113.070 29.430 125.000 29.730 ;
    END
  END RAM2FAB_D1_I2
  PIN RAM2FAB_D1_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 107.090 32.150 125.000 32.450 ;
    END
  END RAM2FAB_D1_I3
  PIN RAM2FAB_D2_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.970 12.430 125.000 12.730 ;
    END
  END RAM2FAB_D2_I0
  PIN RAM2FAB_D2_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 117.210 15.150 125.000 15.450 ;
    END
  END RAM2FAB_D2_I1
  PIN RAM2FAB_D2_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 123.590 17.870 125.000 18.170 ;
    END
  END RAM2FAB_D2_I2
  PIN RAM2FAB_D2_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 114.910 20.590 125.000 20.890 ;
    END
  END RAM2FAB_D2_I3
  PIN RAM2FAB_D3_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.870 1.550 125.000 1.850 ;
    END
  END RAM2FAB_D3_I0
  PIN RAM2FAB_D3_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 123.650 4.270 125.000 4.570 ;
    END
  END RAM2FAB_D3_I1
  PIN RAM2FAB_D3_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 123.650 6.990 125.000 7.290 ;
    END
  END RAM2FAB_D3_I2
  PIN RAM2FAB_D3_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 118.130 9.710 125.000 10.010 ;
    END
  END RAM2FAB_D3_I3
  PIN S1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.920 0.000 49.060 1.090 ;
    END
  END S1BEG[0]
  PIN S1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.300 0.000 50.440 7.520 ;
    END
  END S1BEG[1]
  PIN S1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.680 0.000 51.820 15.340 ;
    END
  END S1BEG[2]
  PIN S1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.060 0.000 53.200 2.080 ;
    END
  END S1BEG[3]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.380 216.880 49.520 223.115 ;
    END
  END S1END[0]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.760 213.480 50.900 223.115 ;
    END
  END S1END[1]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.140 216.880 52.280 223.115 ;
    END
  END S1END[2]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.520 213.480 53.660 223.115 ;
    END
  END S1END[3]
  PIN S2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.020 0.000 65.160 4.490 ;
    END
  END S2BEG[0]
  PIN S2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.400 0.000 66.540 16.700 ;
    END
  END S2BEG[1]
  PIN S2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.780 0.000 67.920 27.580 ;
    END
  END S2BEG[2]
  PIN S2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.160 0.000 69.300 19.760 ;
    END
  END S2BEG[3]
  PIN S2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.540 0.000 70.680 15.680 ;
    END
  END S2BEG[4]
  PIN S2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.920 0.000 72.060 13.980 ;
    END
  END S2BEG[5]
  PIN S2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.840 0.000 72.980 34.040 ;
    END
  END S2BEG[6]
  PIN S2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.220 0.000 74.360 9.420 ;
    END
  END S2BEG[7]
  PIN S2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.980 0.000 54.120 15.680 ;
    END
  END S2BEGb[0]
  PIN S2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.360 0.000 55.500 7.380 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.740 0.000 56.880 35.740 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.120 0.000 58.260 7.000 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.500 0.000 59.640 38.460 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.880 0.000 61.020 16.520 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.260 0.000 62.400 4.120 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.640 0.000 63.780 21.120 ;
    END
  END S2BEGb[7]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.900 206.930 55.040 223.115 ;
    END
  END S2END[0]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.280 153.640 56.420 223.115 ;
    END
  END S2END[1]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.660 191.380 57.800 223.115 ;
    END
  END S2END[2]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.040 200.700 59.180 223.115 ;
    END
  END S2END[3]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.420 213.480 60.560 223.115 ;
    END
  END S2END[4]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.800 216.040 61.940 223.115 ;
    END
  END S2END[5]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.180 216.540 63.320 223.115 ;
    END
  END S2END[6]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.100 220.590 64.240 223.115 ;
    END
  END S2END[7]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.480 216.880 65.620 223.115 ;
    END
  END S2MID[0]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.860 216.880 67.000 223.115 ;
    END
  END S2MID[1]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.240 213.480 68.380 223.115 ;
    END
  END S2MID[2]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.620 216.540 69.760 223.115 ;
    END
  END S2MID[3]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.000 213.140 71.140 223.115 ;
    END
  END S2MID[4]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.380 211.440 72.520 223.115 ;
    END
  END S2MID[5]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.760 213.480 73.900 223.115 ;
    END
  END S2MID[6]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.140 216.880 75.280 223.115 ;
    END
  END S2MID[7]
  PIN S4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.600 0.000 75.740 12.650 ;
    END
  END S4BEG[0]
  PIN S4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.400 0.000 89.540 35.740 ;
    END
  END S4BEG[10]
  PIN S4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.320 0.000 90.460 13.870 ;
    END
  END S4BEG[11]
  PIN S4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.700 0.000 91.840 18.400 ;
    END
  END S4BEG[12]
  PIN S4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.080 0.000 93.220 42.880 ;
    END
  END S4BEG[13]
  PIN S4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.460 0.000 94.600 44.920 ;
    END
  END S4BEG[14]
  PIN S4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.840 0.000 95.980 41.180 ;
    END
  END S4BEG[15]
  PIN S4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.980 0.000 77.120 15.000 ;
    END
  END S4BEG[1]
  PIN S4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.360 0.000 78.500 13.870 ;
    END
  END S4BEG[2]
  PIN S4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.740 0.000 79.880 11.290 ;
    END
  END S4BEG[3]
  PIN S4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.120 0.000 81.260 4.120 ;
    END
  END S4BEG[4]
  PIN S4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.500 0.000 82.640 18.400 ;
    END
  END S4BEG[5]
  PIN S4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.880 0.000 84.020 19.620 ;
    END
  END S4BEG[6]
  PIN S4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.260 0.000 85.400 15.680 ;
    END
  END S4BEG[7]
  PIN S4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.640 0.000 86.780 2.450 ;
    END
  END S4BEG[8]
  PIN S4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.020 0.000 88.160 2.450 ;
    END
  END S4BEG[9]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.520 211.440 76.660 223.115 ;
    END
  END S4END[0]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.320 201.760 90.460 223.115 ;
    END
  END S4END[10]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.700 201.920 91.840 223.115 ;
    END
  END S4END[11]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.080 216.510 93.220 223.115 ;
    END
  END S4END[12]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.460 206.930 94.600 223.115 ;
    END
  END S4END[13]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.380 214.470 95.520 223.115 ;
    END
  END S4END[14]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.760 214.470 96.900 223.115 ;
    END
  END S4END[15]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.900 212.940 78.040 223.115 ;
    END
  END S4END[1]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.280 216.540 79.420 223.115 ;
    END
  END S4END[2]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.660 218.380 80.800 223.115 ;
    END
  END S4END[3]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.040 219.260 82.180 223.115 ;
    END
  END S4END[4]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.420 204.950 83.560 223.115 ;
    END
  END S4END[5]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.800 212.800 84.940 223.115 ;
    END
  END S4END[6]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.180 216.510 86.320 223.115 ;
    END
  END S4END[7]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.560 192.540 87.700 223.115 ;
    END
  END S4END[8]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.940 214.470 89.080 223.115 ;
    END
  END S4END[9]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.220 0.000 97.360 19.420 ;
    END
  END UserCLK
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 42.705 5.200 44.305 217.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 80.690 5.200 82.290 217.840 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 23.715 5.200 25.315 217.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 61.700 5.200 63.300 217.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 99.685 5.200 101.285 217.840 ;
    END
  END VPWR
  PIN W1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.870 14.810 1.170 ;
    END
  END W1BEG[0]
  PIN W1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.230 7.450 2.530 ;
    END
  END W1BEG[1]
  PIN W1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.270 17.570 4.570 ;
    END
  END W1BEG[2]
  PIN W1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.630 26.770 5.930 ;
    END
  END W1BEG[3]
  PIN W2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.670 13.890 7.970 ;
    END
  END W2BEG[0]
  PIN W2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.030 3.310 9.330 ;
    END
  END W2BEG[1]
  PIN W2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.070 19.870 11.370 ;
    END
  END W2BEG[2]
  PIN W2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.430 18.950 12.730 ;
    END
  END W2BEG[3]
  PIN W2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.470 15.730 14.770 ;
    END
  END W2BEG[4]
  PIN W2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.510 18.490 16.810 ;
    END
  END W2BEG[5]
  PIN W2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.870 16.650 18.170 ;
    END
  END W2BEG[6]
  PIN W2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.910 22.630 20.210 ;
    END
  END W2BEG[7]
  PIN W2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.270 20.330 21.570 ;
    END
  END W2BEGb[0]
  PIN W2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.310 17.110 23.610 ;
    END
  END W2BEGb[1]
  PIN W2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.670 19.870 24.970 ;
    END
  END W2BEGb[2]
  PIN W2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.710 20.330 27.010 ;
    END
  END W2BEGb[3]
  PIN W2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.750 7.910 29.050 ;
    END
  END W2BEGb[4]
  PIN W2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.110 22.000 30.410 ;
    END
  END W2BEGb[5]
  PIN W2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.150 15.270 32.450 ;
    END
  END W2BEGb[6]
  PIN W2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.510 22.630 33.810 ;
    END
  END W2BEGb[7]
  PIN W6BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.430 7.910 63.730 ;
    END
  END W6BEG[0]
  PIN W6BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.430 9.290 80.730 ;
    END
  END W6BEG[10]
  PIN W6BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.470 16.650 82.770 ;
    END
  END W6BEG[11]
  PIN W6BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.790 17.570 65.090 ;
    END
  END W6BEG[1]
  PIN W6BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.830 19.870 67.130 ;
    END
  END W6BEG[2]
  PIN W6BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.190 20.330 68.490 ;
    END
  END W6BEG[3]
  PIN W6BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.230 20.330 70.530 ;
    END
  END W6BEG[4]
  PIN W6BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.270 18.490 72.570 ;
    END
  END W6BEG[5]
  PIN W6BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.630 17.860 73.930 ;
    END
  END W6BEG[6]
  PIN W6BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.670 20.330 75.970 ;
    END
  END W6BEG[7]
  PIN W6BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.030 20.330 77.330 ;
    END
  END W6BEG[8]
  PIN W6BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.070 19.870 79.370 ;
    END
  END W6BEG[9]
  PIN WW4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.550 19.870 35.850 ;
    END
  END WW4BEG[0]
  PIN WW4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.550 19.870 52.850 ;
    END
  END WW4BEG[10]
  PIN WW4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.590 20.330 54.890 ;
    END
  END WW4BEG[11]
  PIN WW4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.630 19.870 56.930 ;
    END
  END WW4BEG[12]
  PIN WW4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.990 21.080 58.290 ;
    END
  END WW4BEG[13]
  PIN WW4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.030 19.870 60.330 ;
    END
  END WW4BEG[14]
  PIN WW4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.390 20.330 61.690 ;
    END
  END WW4BEG[15]
  PIN WW4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.910 20.330 37.210 ;
    END
  END WW4BEG[1]
  PIN WW4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.950 17.570 39.250 ;
    END
  END WW4BEG[2]
  PIN WW4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.310 20.330 40.610 ;
    END
  END WW4BEG[3]
  PIN WW4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.350 19.870 42.650 ;
    END
  END WW4BEG[4]
  PIN WW4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.390 40.110 44.690 ;
    END
  END WW4BEG[5]
  PIN WW4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.750 23.380 46.050 ;
    END
  END WW4BEG[6]
  PIN WW4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.790 40.110 48.090 ;
    END
  END WW4BEG[7]
  PIN WW4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.150 20.330 49.450 ;
    END
  END WW4BEG[8]
  PIN WW4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.190 18.950 51.490 ;
    END
  END WW4BEG[9]
  OBS
      LAYER li1 ;
        RECT 4.285 1.445 124.975 217.685 ;
      LAYER met1 ;
        RECT 0.530 0.720 124.590 220.620 ;
      LAYER met2 ;
        RECT 1.040 216.940 1.260 222.205 ;
        RECT 0.560 213.540 1.260 216.940 ;
        RECT 1.960 219.320 2.640 222.205 ;
        RECT 3.340 219.320 4.020 222.205 ;
        RECT 1.960 213.540 4.020 219.320 ;
        RECT 0.560 206.060 4.020 213.540 ;
        RECT 4.720 220.000 5.400 222.205 ;
        RECT 6.100 220.340 6.780 222.205 ;
        RECT 7.480 220.340 8.160 222.205 ;
        RECT 6.100 220.000 8.160 220.340 ;
        RECT 4.720 206.060 8.160 220.000 ;
        RECT 0.560 205.560 8.160 206.060 ;
        RECT 8.860 210.320 9.540 222.205 ;
        RECT 10.240 216.230 10.920 222.205 ;
        RECT 11.620 216.230 12.300 222.205 ;
        RECT 10.240 210.320 12.300 216.230 ;
        RECT 8.860 208.780 12.300 210.320 ;
        RECT 13.000 216.060 13.680 222.205 ;
        RECT 14.380 217.960 15.060 222.205 ;
        RECT 15.760 217.960 16.440 222.205 ;
        RECT 14.380 216.060 16.440 217.960 ;
        RECT 13.000 208.960 16.440 216.060 ;
        RECT 17.140 208.960 17.820 222.205 ;
        RECT 13.000 208.780 17.820 208.960 ;
        RECT 8.860 205.560 17.820 208.780 ;
        RECT 0.560 201.640 17.820 205.560 ;
        RECT 18.520 213.040 19.200 222.205 ;
        RECT 19.900 214.190 20.580 222.205 ;
        RECT 21.280 214.190 21.960 222.205 ;
        RECT 19.900 213.040 21.960 214.190 ;
        RECT 18.520 206.060 21.960 213.040 ;
        RECT 22.660 215.550 23.340 222.205 ;
        RECT 24.040 215.550 24.720 222.205 ;
        RECT 25.420 219.660 26.100 222.205 ;
        RECT 26.800 219.660 27.480 222.205 ;
        RECT 25.420 215.550 27.480 219.660 ;
        RECT 22.660 206.060 27.480 215.550 ;
        RECT 18.520 204.360 27.480 206.060 ;
        RECT 28.180 206.060 28.860 222.205 ;
        RECT 29.560 206.060 30.240 222.205 ;
        RECT 28.180 204.880 30.240 206.060 ;
        RECT 30.940 204.880 31.620 222.205 ;
        RECT 28.180 204.360 31.620 204.880 ;
        RECT 18.520 202.320 31.620 204.360 ;
        RECT 32.320 202.660 32.540 222.205 ;
        RECT 33.240 206.650 33.920 222.205 ;
        RECT 34.620 206.650 35.300 222.205 ;
        RECT 33.240 202.660 35.300 206.650 ;
        RECT 32.320 202.320 35.300 202.660 ;
        RECT 18.520 201.640 35.300 202.320 ;
        RECT 0.560 176.140 35.300 201.640 ;
        RECT 36.000 176.140 36.680 222.205 ;
        RECT 0.560 173.420 36.680 176.140 ;
        RECT 37.380 203.520 38.060 222.205 ;
        RECT 38.760 211.680 39.440 222.205 ;
        RECT 40.140 216.230 40.820 222.205 ;
        RECT 41.520 218.270 42.200 222.205 ;
        RECT 42.900 218.270 43.580 222.205 ;
        RECT 44.280 218.270 44.960 222.205 ;
        RECT 41.520 216.230 44.960 218.270 ;
        RECT 40.140 214.220 44.960 216.230 ;
        RECT 45.660 214.220 46.340 222.205 ;
        RECT 40.140 211.680 46.340 214.220 ;
        RECT 38.760 208.960 46.340 211.680 ;
        RECT 47.040 210.110 47.720 222.205 ;
        RECT 48.420 216.600 49.100 222.205 ;
        RECT 49.800 216.600 50.480 222.205 ;
        RECT 48.420 213.200 50.480 216.600 ;
        RECT 51.180 216.600 51.860 222.205 ;
        RECT 52.560 216.600 53.240 222.205 ;
        RECT 51.180 213.200 53.240 216.600 ;
        RECT 53.940 213.200 54.620 222.205 ;
        RECT 48.420 210.110 54.620 213.200 ;
        RECT 47.040 208.960 54.620 210.110 ;
        RECT 38.760 206.650 54.620 208.960 ;
        RECT 55.320 206.650 56.000 222.205 ;
        RECT 38.760 203.520 56.000 206.650 ;
        RECT 37.380 173.420 56.000 203.520 ;
        RECT 0.560 153.360 56.000 173.420 ;
        RECT 56.700 191.100 57.380 222.205 ;
        RECT 58.080 200.420 58.760 222.205 ;
        RECT 59.460 213.200 60.140 222.205 ;
        RECT 60.840 215.760 61.520 222.205 ;
        RECT 62.220 216.260 62.900 222.205 ;
        RECT 63.600 220.310 63.820 222.205 ;
        RECT 64.520 220.310 65.200 222.205 ;
        RECT 63.600 216.600 65.200 220.310 ;
        RECT 65.900 216.600 66.580 222.205 ;
        RECT 67.280 216.600 67.960 222.205 ;
        RECT 63.600 216.260 67.960 216.600 ;
        RECT 62.220 215.760 67.960 216.260 ;
        RECT 60.840 213.200 67.960 215.760 ;
        RECT 68.660 216.260 69.340 222.205 ;
        RECT 70.040 216.260 70.720 222.205 ;
        RECT 68.660 213.200 70.720 216.260 ;
        RECT 59.460 212.860 70.720 213.200 ;
        RECT 71.420 212.860 72.100 222.205 ;
        RECT 59.460 211.160 72.100 212.860 ;
        RECT 72.800 213.200 73.480 222.205 ;
        RECT 74.180 216.600 74.860 222.205 ;
        RECT 75.560 216.600 76.240 222.205 ;
        RECT 74.180 213.200 76.240 216.600 ;
        RECT 72.800 211.160 76.240 213.200 ;
        RECT 76.940 212.660 77.620 222.205 ;
        RECT 78.320 216.260 79.000 222.205 ;
        RECT 79.700 218.100 80.380 222.205 ;
        RECT 81.080 218.980 81.760 222.205 ;
        RECT 82.460 218.980 83.140 222.205 ;
        RECT 81.080 218.100 83.140 218.980 ;
        RECT 79.700 216.260 83.140 218.100 ;
        RECT 78.320 212.660 83.140 216.260 ;
        RECT 76.940 211.160 83.140 212.660 ;
        RECT 59.460 204.670 83.140 211.160 ;
        RECT 83.840 212.520 84.520 222.205 ;
        RECT 85.220 216.230 85.900 222.205 ;
        RECT 86.600 216.230 87.280 222.205 ;
        RECT 85.220 212.520 87.280 216.230 ;
        RECT 83.840 204.670 87.280 212.520 ;
        RECT 59.460 200.420 87.280 204.670 ;
        RECT 58.080 192.260 87.280 200.420 ;
        RECT 87.980 214.190 88.660 222.205 ;
        RECT 89.360 214.190 90.040 222.205 ;
        RECT 87.980 201.480 90.040 214.190 ;
        RECT 90.740 201.640 91.420 222.205 ;
        RECT 92.120 216.230 92.800 222.205 ;
        RECT 93.500 216.230 94.180 222.205 ;
        RECT 92.120 206.650 94.180 216.230 ;
        RECT 94.880 214.190 95.100 222.205 ;
        RECT 95.800 214.190 96.480 222.205 ;
        RECT 97.180 216.940 97.860 222.205 ;
        RECT 98.560 216.940 99.240 222.205 ;
        RECT 97.180 215.550 99.240 216.940 ;
        RECT 99.940 218.100 100.620 222.205 ;
        RECT 101.320 218.100 102.000 222.205 ;
        RECT 99.940 215.550 102.000 218.100 ;
        RECT 97.180 214.190 102.000 215.550 ;
        RECT 102.700 214.190 103.380 222.205 ;
        RECT 104.080 214.190 104.760 222.205 ;
        RECT 94.880 206.650 104.760 214.190 ;
        RECT 92.120 201.640 104.760 206.650 ;
        RECT 90.740 201.480 104.760 201.640 ;
        RECT 87.980 200.620 104.760 201.480 ;
        RECT 105.460 214.190 106.140 222.205 ;
        RECT 106.840 214.190 107.520 222.205 ;
        RECT 108.220 214.190 108.900 222.205 ;
        RECT 105.460 210.110 108.900 214.190 ;
        RECT 109.600 210.110 110.280 222.205 ;
        RECT 105.460 206.650 110.280 210.110 ;
        RECT 110.980 208.440 111.660 222.205 ;
        RECT 112.360 211.160 113.040 222.205 ;
        RECT 113.740 211.300 114.420 222.205 ;
        RECT 115.120 217.960 115.800 222.205 ;
        RECT 116.500 217.960 117.180 222.205 ;
        RECT 115.120 211.500 117.180 217.960 ;
        RECT 117.880 218.980 118.560 222.205 ;
        RECT 119.260 218.980 119.940 222.205 ;
        RECT 117.880 211.500 119.940 218.980 ;
        RECT 115.120 211.300 119.940 211.500 ;
        RECT 113.740 211.160 119.940 211.300 ;
        RECT 112.360 208.440 119.940 211.160 ;
        RECT 110.980 206.650 119.940 208.440 ;
        RECT 105.460 203.000 119.940 206.650 ;
        RECT 120.640 205.040 121.320 222.205 ;
        RECT 122.020 211.680 122.700 222.205 ;
        RECT 123.400 216.940 124.080 222.205 ;
        RECT 124.780 216.940 124.960 222.205 ;
        RECT 123.400 211.680 124.960 216.940 ;
        RECT 122.020 205.040 124.960 211.680 ;
        RECT 120.640 203.000 124.960 205.040 ;
        RECT 105.460 200.620 124.960 203.000 ;
        RECT 87.980 192.260 124.960 200.620 ;
        RECT 58.080 191.100 124.960 192.260 ;
        RECT 56.700 153.360 124.960 191.100 ;
        RECT 0.560 45.200 124.960 153.360 ;
        RECT 0.560 43.160 94.180 45.200 ;
        RECT 0.560 38.740 92.800 43.160 ;
        RECT 0.560 36.900 59.220 38.740 ;
        RECT 0.560 20.720 35.300 36.900 ;
        RECT 0.560 6.440 1.260 20.720 ;
        RECT 1.040 0.690 1.260 6.440 ;
        RECT 1.960 15.620 35.300 20.720 ;
        RECT 1.960 14.260 12.300 15.620 ;
        RECT 1.960 10.180 9.540 14.260 ;
        RECT 1.960 9.840 5.400 10.180 ;
        RECT 1.960 0.690 2.640 9.840 ;
        RECT 3.340 6.780 5.400 9.840 ;
        RECT 3.340 0.690 4.020 6.780 ;
        RECT 4.720 0.690 5.400 6.780 ;
        RECT 6.100 9.160 9.540 10.180 ;
        RECT 6.100 5.080 8.160 9.160 ;
        RECT 6.100 0.690 6.780 5.080 ;
        RECT 7.480 0.690 8.160 5.080 ;
        RECT 8.860 0.690 9.540 9.160 ;
        RECT 10.240 3.040 12.300 14.260 ;
        RECT 10.240 0.690 10.920 3.040 ;
        RECT 11.620 0.690 12.300 3.040 ;
        RECT 13.000 15.280 31.160 15.620 ;
        RECT 13.000 7.120 20.120 15.280 ;
        RECT 13.000 3.720 15.060 7.120 ;
        RECT 13.000 0.690 13.680 3.720 ;
        RECT 14.380 0.690 15.060 3.720 ;
        RECT 15.760 6.440 20.120 7.120 ;
        RECT 15.760 0.690 16.440 6.440 ;
        RECT 17.140 4.060 20.120 6.440 ;
        RECT 17.140 2.700 18.740 4.060 ;
        RECT 17.140 0.690 17.820 2.700 ;
        RECT 18.520 0.690 18.740 2.700 ;
        RECT 19.440 0.690 20.120 4.060 ;
        RECT 20.820 14.600 31.160 15.280 ;
        RECT 20.820 14.150 22.880 14.600 ;
        RECT 20.820 0.690 21.500 14.150 ;
        RECT 22.200 0.690 22.880 14.150 ;
        RECT 23.580 14.260 31.160 14.600 ;
        RECT 23.580 9.840 29.780 14.260 ;
        RECT 23.580 6.440 25.640 9.840 ;
        RECT 23.580 0.690 24.260 6.440 ;
        RECT 24.960 0.690 25.640 6.440 ;
        RECT 26.340 7.490 29.780 9.840 ;
        RECT 26.340 4.090 28.400 7.490 ;
        RECT 26.340 0.690 27.020 4.090 ;
        RECT 27.720 0.690 28.400 4.090 ;
        RECT 29.100 0.690 29.780 7.490 ;
        RECT 30.480 0.690 31.160 14.260 ;
        RECT 31.860 14.150 35.300 15.620 ;
        RECT 31.860 0.690 32.540 14.150 ;
        RECT 33.240 7.490 35.300 14.150 ;
        RECT 33.240 0.690 33.920 7.490 ;
        RECT 34.620 0.690 35.300 7.490 ;
        RECT 36.000 36.020 59.220 36.900 ;
        RECT 36.000 24.490 56.460 36.020 ;
        RECT 36.000 19.050 40.360 24.490 ;
        RECT 36.000 15.280 38.980 19.050 ;
        RECT 36.000 0.690 36.220 15.280 ;
        RECT 36.920 14.150 38.980 15.280 ;
        RECT 36.920 0.690 37.600 14.150 ;
        RECT 38.300 0.690 38.980 14.150 ;
        RECT 39.680 0.690 40.360 19.050 ;
        RECT 41.060 16.980 56.460 24.490 ;
        RECT 41.060 14.150 47.260 16.980 ;
        RECT 41.060 12.560 45.880 14.150 ;
        RECT 41.060 4.940 44.500 12.560 ;
        RECT 41.060 4.060 43.120 4.940 ;
        RECT 41.060 0.690 41.740 4.060 ;
        RECT 42.440 0.690 43.120 4.060 ;
        RECT 43.820 0.690 44.500 4.940 ;
        RECT 45.200 0.690 45.880 12.560 ;
        RECT 46.580 0.690 47.260 14.150 ;
        RECT 47.960 15.960 56.460 16.980 ;
        RECT 47.960 15.620 53.700 15.960 ;
        RECT 47.960 7.800 51.400 15.620 ;
        RECT 47.960 1.370 50.020 7.800 ;
        RECT 47.960 0.690 48.640 1.370 ;
        RECT 49.340 0.690 50.020 1.370 ;
        RECT 50.720 0.690 51.400 7.800 ;
        RECT 52.100 2.360 53.700 15.620 ;
        RECT 52.100 0.690 52.780 2.360 ;
        RECT 53.480 0.690 53.700 2.360 ;
        RECT 54.400 7.660 56.460 15.960 ;
        RECT 54.400 0.690 55.080 7.660 ;
        RECT 55.780 0.690 56.460 7.660 ;
        RECT 57.160 7.280 59.220 36.020 ;
        RECT 57.160 0.690 57.840 7.280 ;
        RECT 58.540 0.690 59.220 7.280 ;
        RECT 59.920 36.020 92.800 38.740 ;
        RECT 59.920 34.320 89.120 36.020 ;
        RECT 59.920 27.860 72.560 34.320 ;
        RECT 59.920 21.400 67.500 27.860 ;
        RECT 59.920 16.800 63.360 21.400 ;
        RECT 59.920 0.690 60.600 16.800 ;
        RECT 61.300 4.400 63.360 16.800 ;
        RECT 61.300 0.690 61.980 4.400 ;
        RECT 62.680 0.690 63.360 4.400 ;
        RECT 64.060 16.980 67.500 21.400 ;
        RECT 64.060 4.770 66.120 16.980 ;
        RECT 64.060 0.690 64.740 4.770 ;
        RECT 65.440 0.690 66.120 4.770 ;
        RECT 66.820 0.690 67.500 16.980 ;
        RECT 68.200 20.040 72.560 27.860 ;
        RECT 68.200 0.690 68.880 20.040 ;
        RECT 69.580 15.960 72.560 20.040 ;
        RECT 69.580 0.690 70.260 15.960 ;
        RECT 70.960 14.260 72.560 15.960 ;
        RECT 70.960 0.690 71.640 14.260 ;
        RECT 72.340 0.690 72.560 14.260 ;
        RECT 73.260 19.900 89.120 34.320 ;
        RECT 73.260 18.680 83.600 19.900 ;
        RECT 73.260 15.280 82.220 18.680 ;
        RECT 73.260 12.930 76.700 15.280 ;
        RECT 73.260 9.700 75.320 12.930 ;
        RECT 73.260 0.690 73.940 9.700 ;
        RECT 74.640 0.690 75.320 9.700 ;
        RECT 76.020 0.690 76.700 12.930 ;
        RECT 77.400 14.150 82.220 15.280 ;
        RECT 77.400 0.690 78.080 14.150 ;
        RECT 78.780 11.570 82.220 14.150 ;
        RECT 78.780 0.690 79.460 11.570 ;
        RECT 80.160 4.400 82.220 11.570 ;
        RECT 80.160 0.690 80.840 4.400 ;
        RECT 81.540 0.690 82.220 4.400 ;
        RECT 82.920 0.690 83.600 18.680 ;
        RECT 84.300 15.960 89.120 19.900 ;
        RECT 84.300 0.690 84.980 15.960 ;
        RECT 85.680 2.730 89.120 15.960 ;
        RECT 85.680 0.690 86.360 2.730 ;
        RECT 87.060 0.690 87.740 2.730 ;
        RECT 88.440 0.690 89.120 2.730 ;
        RECT 89.820 18.680 92.800 36.020 ;
        RECT 89.820 14.150 91.420 18.680 ;
        RECT 89.820 0.690 90.040 14.150 ;
        RECT 90.740 0.690 91.420 14.150 ;
        RECT 92.120 0.690 92.800 18.680 ;
        RECT 93.500 0.690 94.180 43.160 ;
        RECT 94.880 41.460 124.960 45.200 ;
        RECT 94.880 0.690 95.560 41.460 ;
        RECT 96.260 29.250 124.960 41.460 ;
        RECT 96.260 22.760 113.040 29.250 ;
        RECT 96.260 19.700 110.280 22.760 ;
        RECT 96.260 0.690 96.940 19.700 ;
        RECT 97.640 17.660 110.280 19.700 ;
        RECT 97.640 17.320 107.520 17.660 ;
        RECT 97.640 9.500 103.840 17.320 ;
        RECT 97.640 6.440 102.460 9.500 ;
        RECT 97.640 0.690 98.320 6.440 ;
        RECT 99.020 6.130 102.460 6.440 ;
        RECT 99.020 0.690 99.700 6.130 ;
        RECT 100.400 5.450 102.460 6.130 ;
        RECT 100.400 0.690 101.080 5.450 ;
        RECT 101.780 0.690 102.460 5.450 ;
        RECT 103.160 0.690 103.840 9.500 ;
        RECT 104.540 15.280 107.520 17.320 ;
        RECT 104.540 0.690 105.220 15.280 ;
        RECT 105.920 4.400 107.520 15.280 ;
        RECT 105.920 0.690 106.600 4.400 ;
        RECT 107.300 0.690 107.520 4.400 ;
        RECT 108.220 6.780 110.280 17.660 ;
        RECT 108.220 0.690 108.900 6.780 ;
        RECT 109.600 0.690 110.280 6.780 ;
        RECT 110.980 6.440 113.040 22.760 ;
        RECT 110.980 0.690 111.660 6.440 ;
        RECT 112.360 0.690 113.040 6.440 ;
        RECT 113.740 20.720 124.960 29.250 ;
        RECT 113.740 18.680 118.560 20.720 ;
        RECT 113.740 0.690 114.420 18.680 ;
        RECT 115.120 18.340 118.560 18.680 ;
        RECT 115.120 0.690 115.800 18.340 ;
        RECT 116.500 17.320 118.560 18.340 ;
        RECT 116.500 0.690 117.180 17.320 ;
        RECT 117.880 0.690 118.560 17.320 ;
        RECT 119.260 20.380 124.960 20.720 ;
        RECT 119.260 0.690 119.940 20.380 ;
        RECT 120.640 19.700 124.960 20.380 ;
        RECT 120.640 17.480 122.700 19.700 ;
        RECT 120.640 0.690 121.320 17.480 ;
        RECT 122.020 0.690 122.700 17.480 ;
        RECT 123.400 1.370 124.960 19.700 ;
        RECT 123.400 0.690 124.080 1.370 ;
        RECT 124.780 0.690 124.960 1.370 ;
      LAYER met3 ;
        RECT 17.510 221.890 124.810 222.185 ;
        RECT 17.510 221.470 106.690 221.890 ;
        RECT 2.365 220.790 106.690 221.470 ;
        RECT 2.365 220.530 124.810 220.790 ;
        RECT 20.730 219.430 124.810 220.530 ;
        RECT 2.365 219.170 124.810 219.430 ;
        RECT 20.270 218.070 108.530 219.170 ;
        RECT 2.365 217.130 124.810 218.070 ;
        RECT 17.510 216.450 124.810 217.130 ;
        RECT 17.510 216.030 110.830 216.450 ;
        RECT 2.365 215.770 110.830 216.030 ;
        RECT 15.670 215.350 110.830 215.770 ;
        RECT 15.670 214.670 124.810 215.350 ;
        RECT 2.365 213.730 124.810 214.670 ;
        RECT 16.590 212.630 115.430 213.730 ;
        RECT 2.365 212.370 124.810 212.630 ;
        RECT 19.350 211.270 124.810 212.370 ;
        RECT 2.365 211.010 124.810 211.270 ;
        RECT 2.365 210.330 114.970 211.010 ;
        RECT 7.390 209.910 114.970 210.330 ;
        RECT 7.390 209.230 124.810 209.910 ;
        RECT 2.365 208.290 124.810 209.230 ;
        RECT 20.730 207.190 114.970 208.290 ;
        RECT 2.365 206.930 124.810 207.190 ;
        RECT 14.750 205.830 124.810 206.930 ;
        RECT 2.365 205.570 124.810 205.830 ;
        RECT 2.365 204.890 115.430 205.570 ;
        RECT 7.850 204.470 115.430 204.890 ;
        RECT 7.850 203.790 124.810 204.470 ;
        RECT 2.365 203.530 124.810 203.790 ;
        RECT 6.930 202.850 124.810 203.530 ;
        RECT 6.930 202.430 114.970 202.850 ;
        RECT 2.365 201.750 114.970 202.430 ;
        RECT 2.365 201.490 124.810 201.750 ;
        RECT 20.270 200.390 124.810 201.490 ;
        RECT 2.365 200.130 124.810 200.390 ;
        RECT 21.250 199.030 115.430 200.130 ;
        RECT 2.365 198.090 124.810 199.030 ;
        RECT 20.730 197.410 124.810 198.090 ;
        RECT 20.730 196.990 114.970 197.410 ;
        RECT 2.365 196.730 114.970 196.990 ;
        RECT 14.810 196.310 114.970 196.730 ;
        RECT 14.810 195.630 124.810 196.310 ;
        RECT 2.365 194.690 124.810 195.630 ;
        RECT 19.810 194.010 124.810 194.690 ;
        RECT 19.810 193.590 114.970 194.010 ;
        RECT 2.365 192.910 114.970 193.590 ;
        RECT 2.365 192.650 124.810 192.910 ;
        RECT 16.590 191.550 124.810 192.650 ;
        RECT 2.365 191.290 124.810 191.550 ;
        RECT 20.730 190.190 115.430 191.290 ;
        RECT 2.365 189.250 124.810 190.190 ;
        RECT 14.750 188.570 124.810 189.250 ;
        RECT 14.750 188.150 116.810 188.570 ;
        RECT 2.365 187.890 116.810 188.150 ;
        RECT 15.210 187.470 116.810 187.890 ;
        RECT 15.210 186.790 124.810 187.470 ;
        RECT 2.365 185.850 124.810 186.790 ;
        RECT 9.230 184.750 114.970 185.850 ;
        RECT 2.365 184.490 124.810 184.750 ;
        RECT 21.190 183.390 124.810 184.490 ;
        RECT 2.365 183.130 124.810 183.390 ;
        RECT 2.365 182.450 115.430 183.130 ;
        RECT 8.770 182.030 115.430 182.450 ;
        RECT 8.770 181.350 124.810 182.030 ;
        RECT 2.365 180.410 124.810 181.350 ;
        RECT 17.970 179.310 114.970 180.410 ;
        RECT 2.365 179.050 124.810 179.310 ;
        RECT 17.970 177.950 124.810 179.050 ;
        RECT 2.365 177.690 124.810 177.950 ;
        RECT 2.365 177.010 115.430 177.690 ;
        RECT 20.270 176.590 115.430 177.010 ;
        RECT 20.270 175.910 124.810 176.590 ;
        RECT 2.365 175.650 124.810 175.910 ;
        RECT 28.090 174.970 124.810 175.650 ;
        RECT 28.090 174.550 109.450 174.970 ;
        RECT 2.365 173.870 109.450 174.550 ;
        RECT 2.365 173.610 124.810 173.870 ;
        RECT 29.010 172.510 124.810 173.610 ;
        RECT 2.365 172.250 124.810 172.510 ;
        RECT 20.730 171.150 116.810 172.250 ;
        RECT 2.365 170.210 124.810 171.150 ;
        RECT 14.750 169.530 124.810 170.210 ;
        RECT 14.750 169.110 111.750 169.530 ;
        RECT 2.365 168.850 111.750 169.110 ;
        RECT 14.290 168.430 111.750 168.850 ;
        RECT 14.290 167.750 124.810 168.430 ;
        RECT 2.365 166.810 124.810 167.750 ;
        RECT 16.590 166.130 124.810 166.810 ;
        RECT 16.590 165.710 115.430 166.130 ;
        RECT 2.365 165.030 115.430 165.710 ;
        RECT 2.365 164.770 124.810 165.030 ;
        RECT 7.390 163.670 124.810 164.770 ;
        RECT 2.365 163.410 124.810 163.670 ;
        RECT 17.510 162.310 114.970 163.410 ;
        RECT 2.365 161.370 124.810 162.310 ;
        RECT 20.270 160.690 124.810 161.370 ;
        RECT 20.270 160.270 108.070 160.690 ;
        RECT 2.365 160.010 108.070 160.270 ;
        RECT 20.730 159.590 108.070 160.010 ;
        RECT 20.730 158.910 124.810 159.590 ;
        RECT 2.365 157.970 124.810 158.910 ;
        RECT 20.270 156.870 108.070 157.970 ;
        RECT 2.365 156.610 124.810 156.870 ;
        RECT 19.640 155.510 124.810 156.610 ;
        RECT 2.365 155.250 124.810 155.510 ;
        RECT 2.365 154.570 117.440 155.250 ;
        RECT 2.790 154.150 117.440 154.570 ;
        RECT 2.790 153.470 124.810 154.150 ;
        RECT 2.365 152.530 124.810 153.470 ;
        RECT 14.290 151.430 113.590 152.530 ;
        RECT 2.365 151.170 124.810 151.430 ;
        RECT 13.830 150.070 124.810 151.170 ;
        RECT 2.365 149.810 124.810 150.070 ;
        RECT 2.365 149.130 116.810 149.810 ;
        RECT 11.530 148.710 116.810 149.130 ;
        RECT 11.530 148.030 124.810 148.710 ;
        RECT 2.365 147.770 124.810 148.030 ;
        RECT 7.390 147.090 124.810 147.770 ;
        RECT 7.390 146.670 115.430 147.090 ;
        RECT 2.365 145.990 115.430 146.670 ;
        RECT 2.365 145.730 124.810 145.990 ;
        RECT 14.750 144.630 124.810 145.730 ;
        RECT 2.365 144.370 124.810 144.630 ;
        RECT 6.930 143.270 106.230 144.370 ;
        RECT 2.365 142.330 124.810 143.270 ;
        RECT 20.730 141.650 124.810 142.330 ;
        RECT 20.730 141.230 110.370 141.650 ;
        RECT 2.365 140.970 110.370 141.230 ;
        RECT 16.590 140.550 110.370 140.970 ;
        RECT 16.590 139.870 124.810 140.550 ;
        RECT 2.365 138.930 124.810 139.870 ;
        RECT 7.390 138.250 124.810 138.930 ;
        RECT 7.390 137.830 106.230 138.250 ;
        RECT 2.365 137.150 106.230 137.830 ;
        RECT 2.365 136.890 124.810 137.150 ;
        RECT 20.730 135.790 124.810 136.890 ;
        RECT 2.365 135.530 124.810 135.790 ;
        RECT 20.730 134.430 111.290 135.530 ;
        RECT 2.365 133.490 124.810 134.430 ;
        RECT 20.730 132.810 124.810 133.490 ;
        RECT 20.730 132.390 109.450 132.810 ;
        RECT 2.365 132.130 109.450 132.390 ;
        RECT 19.350 131.710 109.450 132.130 ;
        RECT 19.350 131.030 124.810 131.710 ;
        RECT 2.365 130.090 124.810 131.030 ;
        RECT 14.350 128.990 109.910 130.090 ;
        RECT 2.365 128.730 124.810 128.990 ;
        RECT 20.730 127.630 124.810 128.730 ;
        RECT 2.365 127.370 124.810 127.630 ;
        RECT 2.365 126.690 109.450 127.370 ;
        RECT 20.730 126.270 109.450 126.690 ;
        RECT 20.730 125.590 124.810 126.270 ;
        RECT 2.365 124.650 124.810 125.590 ;
        RECT 17.510 123.550 114.970 124.650 ;
        RECT 2.365 123.290 124.810 123.550 ;
        RECT 20.730 122.190 124.810 123.290 ;
        RECT 2.365 121.930 124.810 122.190 ;
        RECT 2.365 121.250 103.470 121.930 ;
        RECT 19.350 120.830 103.470 121.250 ;
        RECT 19.350 120.150 124.810 120.830 ;
        RECT 2.365 119.890 124.810 120.150 ;
        RECT 7.390 119.210 124.810 119.890 ;
        RECT 7.390 118.790 103.470 119.210 ;
        RECT 2.365 118.110 103.470 118.790 ;
        RECT 2.365 117.850 124.810 118.110 ;
        RECT 20.270 116.750 124.810 117.850 ;
        RECT 2.365 116.490 124.810 116.750 ;
        RECT 18.430 115.390 106.230 116.490 ;
        RECT 2.365 114.450 124.810 115.390 ;
        RECT 14.350 113.770 124.810 114.450 ;
        RECT 14.350 113.350 110.370 113.770 ;
        RECT 2.365 113.090 110.370 113.350 ;
        RECT 8.770 112.670 110.370 113.090 ;
        RECT 8.770 111.990 124.810 112.670 ;
        RECT 2.365 111.050 124.810 111.990 ;
        RECT 7.450 110.370 124.810 111.050 ;
        RECT 7.450 109.950 102.090 110.370 ;
        RECT 2.365 109.270 102.090 109.950 ;
        RECT 2.365 109.010 124.810 109.270 ;
        RECT 21.190 107.910 124.810 109.010 ;
        RECT 2.365 107.650 124.810 107.910 ;
        RECT 16.130 106.550 103.010 107.650 ;
        RECT 2.365 105.610 124.810 106.550 ;
        RECT 19.810 104.930 124.810 105.610 ;
        RECT 19.810 104.510 103.470 104.930 ;
        RECT 2.365 104.250 103.470 104.510 ;
        RECT 28.090 103.830 103.470 104.250 ;
        RECT 28.090 103.150 124.810 103.830 ;
        RECT 2.365 102.210 124.810 103.150 ;
        RECT 17.970 101.110 103.470 102.210 ;
        RECT 2.365 100.850 124.810 101.110 ;
        RECT 20.270 99.750 124.810 100.850 ;
        RECT 2.365 99.490 124.810 99.750 ;
        RECT 2.365 98.810 106.230 99.490 ;
        RECT 19.810 98.390 106.230 98.810 ;
        RECT 19.810 97.710 124.810 98.390 ;
        RECT 2.365 96.770 124.810 97.710 ;
        RECT 20.730 95.670 103.010 96.770 ;
        RECT 2.365 95.410 124.810 95.670 ;
        RECT 20.730 94.310 124.810 95.410 ;
        RECT 2.365 94.050 124.810 94.310 ;
        RECT 2.365 93.370 108.530 94.050 ;
        RECT 7.390 92.950 108.530 93.370 ;
        RECT 7.390 92.270 124.810 92.950 ;
        RECT 2.365 92.010 124.810 92.270 ;
        RECT 17.970 91.330 124.810 92.010 ;
        RECT 17.970 90.910 103.930 91.330 ;
        RECT 2.365 90.230 103.930 90.910 ;
        RECT 2.365 89.970 124.810 90.230 ;
        RECT 14.750 88.870 124.810 89.970 ;
        RECT 2.365 88.610 124.810 88.870 ;
        RECT 21.190 87.510 103.930 88.610 ;
        RECT 2.365 86.570 124.810 87.510 ;
        RECT 20.730 85.890 124.810 86.570 ;
        RECT 20.730 85.470 113.130 85.890 ;
        RECT 2.365 85.210 113.130 85.470 ;
        RECT 8.310 84.790 113.130 85.210 ;
        RECT 8.310 84.110 124.810 84.790 ;
        RECT 2.365 83.170 124.810 84.110 ;
        RECT 17.050 82.490 124.810 83.170 ;
        RECT 17.050 82.070 103.010 82.490 ;
        RECT 2.365 81.390 103.010 82.070 ;
        RECT 2.365 81.130 124.810 81.390 ;
        RECT 9.690 80.030 124.810 81.130 ;
        RECT 2.365 79.770 124.810 80.030 ;
        RECT 20.270 78.670 109.450 79.770 ;
        RECT 2.365 77.730 124.810 78.670 ;
        RECT 20.730 77.050 124.810 77.730 ;
        RECT 20.730 76.630 103.930 77.050 ;
        RECT 2.365 76.370 103.930 76.630 ;
        RECT 20.730 75.950 103.930 76.370 ;
        RECT 20.730 75.270 124.810 75.950 ;
        RECT 2.365 74.330 124.810 75.270 ;
        RECT 18.260 73.230 106.230 74.330 ;
        RECT 2.365 72.970 124.810 73.230 ;
        RECT 18.890 71.870 124.810 72.970 ;
        RECT 2.365 71.610 124.810 71.870 ;
        RECT 2.365 70.930 111.750 71.610 ;
        RECT 20.730 70.510 111.750 70.930 ;
        RECT 20.730 69.830 124.810 70.510 ;
        RECT 2.365 68.890 124.810 69.830 ;
        RECT 20.730 67.790 114.970 68.890 ;
        RECT 2.365 67.530 124.810 67.790 ;
        RECT 20.270 66.430 124.810 67.530 ;
        RECT 2.365 66.170 124.810 66.430 ;
        RECT 2.365 65.490 106.230 66.170 ;
        RECT 17.970 65.070 106.230 65.490 ;
        RECT 17.970 64.390 124.810 65.070 ;
        RECT 2.365 64.130 124.810 64.390 ;
        RECT 8.310 63.450 124.810 64.130 ;
        RECT 8.310 63.030 106.230 63.450 ;
        RECT 2.365 62.350 106.230 63.030 ;
        RECT 2.365 62.090 124.810 62.350 ;
        RECT 20.730 60.990 124.810 62.090 ;
        RECT 2.365 60.730 124.810 60.990 ;
        RECT 20.270 59.630 116.750 60.730 ;
        RECT 2.365 58.690 124.810 59.630 ;
        RECT 21.480 58.010 124.810 58.690 ;
        RECT 21.480 57.590 108.070 58.010 ;
        RECT 2.365 57.330 108.070 57.590 ;
        RECT 20.270 56.910 108.070 57.330 ;
        RECT 20.270 56.230 124.810 56.910 ;
        RECT 2.365 55.290 124.810 56.230 ;
        RECT 20.730 54.610 124.810 55.290 ;
        RECT 20.730 54.190 115.890 54.610 ;
        RECT 2.365 53.510 115.890 54.190 ;
        RECT 2.365 53.250 124.810 53.510 ;
        RECT 20.270 52.150 124.810 53.250 ;
        RECT 2.365 51.890 124.810 52.150 ;
        RECT 19.350 50.790 111.750 51.890 ;
        RECT 2.365 49.850 124.810 50.790 ;
        RECT 20.730 49.170 124.810 49.850 ;
        RECT 20.730 48.750 115.430 49.170 ;
        RECT 2.365 48.490 115.430 48.750 ;
        RECT 40.510 48.070 115.430 48.490 ;
        RECT 40.510 47.390 124.810 48.070 ;
        RECT 2.365 46.450 124.810 47.390 ;
        RECT 23.780 45.350 109.450 46.450 ;
        RECT 2.365 45.090 124.810 45.350 ;
        RECT 40.510 43.990 124.810 45.090 ;
        RECT 2.365 43.730 124.810 43.990 ;
        RECT 2.365 43.050 103.010 43.730 ;
        RECT 20.270 42.630 103.010 43.050 ;
        RECT 20.270 41.950 124.810 42.630 ;
        RECT 2.365 41.010 124.810 41.950 ;
        RECT 20.730 39.910 109.910 41.010 ;
        RECT 2.365 39.650 124.810 39.910 ;
        RECT 17.970 38.550 124.810 39.650 ;
        RECT 2.365 38.290 124.810 38.550 ;
        RECT 2.365 37.610 103.010 38.290 ;
        RECT 20.730 37.190 103.010 37.610 ;
        RECT 20.730 36.510 124.810 37.190 ;
        RECT 2.365 36.250 124.810 36.510 ;
        RECT 20.270 35.570 124.810 36.250 ;
        RECT 20.270 35.150 107.150 35.570 ;
        RECT 2.365 34.470 107.150 35.150 ;
        RECT 2.365 34.210 124.810 34.470 ;
        RECT 23.030 33.110 124.810 34.210 ;
        RECT 2.365 32.850 124.810 33.110 ;
        RECT 15.670 31.750 106.690 32.850 ;
        RECT 2.365 30.810 124.810 31.750 ;
        RECT 22.400 30.130 124.810 30.810 ;
        RECT 22.400 29.710 112.670 30.130 ;
        RECT 2.365 29.450 112.670 29.710 ;
        RECT 8.310 29.030 112.670 29.450 ;
        RECT 8.310 28.350 124.810 29.030 ;
        RECT 2.365 27.410 124.810 28.350 ;
        RECT 20.730 26.730 124.810 27.410 ;
        RECT 20.730 26.310 87.620 26.730 ;
        RECT 2.365 25.630 87.620 26.310 ;
        RECT 2.365 25.370 124.810 25.630 ;
        RECT 20.270 24.270 124.810 25.370 ;
        RECT 2.365 24.010 124.810 24.270 ;
        RECT 17.510 22.910 108.990 24.010 ;
        RECT 2.365 21.970 124.810 22.910 ;
        RECT 20.730 21.290 124.810 21.970 ;
        RECT 20.730 20.870 114.510 21.290 ;
        RECT 2.365 20.610 114.510 20.870 ;
        RECT 23.030 20.190 114.510 20.610 ;
        RECT 23.030 19.510 124.810 20.190 ;
        RECT 2.365 18.570 124.810 19.510 ;
        RECT 17.050 17.470 123.190 18.570 ;
        RECT 2.365 17.210 124.810 17.470 ;
        RECT 18.890 16.110 124.810 17.210 ;
        RECT 2.365 15.850 124.810 16.110 ;
        RECT 2.365 15.170 116.810 15.850 ;
        RECT 16.130 14.750 116.810 15.170 ;
        RECT 16.130 14.070 124.810 14.750 ;
        RECT 2.365 13.130 124.810 14.070 ;
        RECT 19.350 12.030 119.570 13.130 ;
        RECT 2.365 11.770 124.810 12.030 ;
        RECT 20.270 10.670 124.810 11.770 ;
        RECT 2.365 10.410 124.810 10.670 ;
        RECT 2.365 9.730 117.730 10.410 ;
        RECT 3.710 9.310 117.730 9.730 ;
        RECT 3.710 8.630 124.810 9.310 ;
        RECT 2.365 8.370 124.810 8.630 ;
        RECT 14.290 7.690 124.810 8.370 ;
        RECT 14.290 7.270 123.250 7.690 ;
        RECT 2.365 6.590 123.250 7.270 ;
        RECT 2.365 6.330 124.810 6.590 ;
        RECT 27.170 5.230 124.810 6.330 ;
        RECT 2.365 4.970 124.810 5.230 ;
        RECT 17.970 3.870 123.250 4.970 ;
        RECT 2.365 2.930 124.810 3.870 ;
        RECT 7.850 2.250 124.810 2.930 ;
        RECT 7.850 1.830 103.470 2.250 ;
        RECT 2.365 1.570 103.470 1.830 ;
        RECT 15.210 1.150 103.470 1.570 ;
        RECT 15.210 0.855 124.810 1.150 ;
      LAYER met4 ;
        RECT 3.055 218.240 122.985 218.785 ;
        RECT 3.055 4.800 23.315 218.240 ;
        RECT 25.715 4.800 42.305 218.240 ;
        RECT 44.705 4.800 61.300 218.240 ;
        RECT 63.700 4.800 80.290 218.240 ;
        RECT 82.690 4.800 99.285 218.240 ;
        RECT 101.685 4.800 122.985 218.240 ;
        RECT 3.055 2.215 122.985 4.800 ;
  END
END RAM_IO
MACRO RegFile
  CLASS BLOCK ;
  FOREIGN RegFile ;
  ORIGIN 0.000 0.000 ;
  SIZE 235.000 BY 223.115 ;
  PIN E1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 222.550 84.510 235.000 84.810 ;
    END
  END E1BEG[0]
  PIN E1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 225.770 85.870 235.000 86.170 ;
    END
  END E1BEG[1]
  PIN E1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 220.250 87.910 235.000 88.210 ;
    END
  END E1BEG[2]
  PIN E1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 217.490 89.270 235.000 89.570 ;
    END
  END E1BEG[3]
  PIN E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.510 8.830 84.810 ;
    END
  END E1END[0]
  PIN E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.870 19.410 86.170 ;
    END
  END E1END[1]
  PIN E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.910 8.830 88.210 ;
    END
  END E1END[2]
  PIN E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.270 7.450 89.570 ;
    END
  END E1END[3]
  PIN E2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 219.330 91.310 235.000 91.610 ;
    END
  END E2BEG[0]
  PIN E2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.410 92.670 235.000 92.970 ;
    END
  END E2BEG[1]
  PIN E2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 219.790 94.710 235.000 95.010 ;
    END
  END E2BEG[2]
  PIN E2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 215.650 96.070 235.000 96.370 ;
    END
  END E2BEG[3]
  PIN E2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 220.710 98.110 235.000 98.410 ;
    END
  END E2BEG[4]
  PIN E2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 217.030 100.150 235.000 100.450 ;
    END
  END E2BEG[5]
  PIN E2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 220.250 101.510 235.000 101.810 ;
    END
  END E2BEG[6]
  PIN E2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 219.790 103.550 235.000 103.850 ;
    END
  END E2BEG[7]
  PIN E2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 232.670 104.910 235.000 105.210 ;
    END
  END E2BEGb[0]
  PIN E2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 212.890 106.950 235.000 107.250 ;
    END
  END E2BEGb[1]
  PIN E2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.570 108.310 235.000 108.610 ;
    END
  END E2BEGb[2]
  PIN E2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 217.490 110.350 235.000 110.650 ;
    END
  END E2BEGb[3]
  PIN E2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.980 112.390 235.000 112.690 ;
    END
  END E2BEGb[4]
  PIN E2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 217.490 113.750 235.000 114.050 ;
    END
  END E2BEGb[5]
  PIN E2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 225.770 115.790 235.000 116.090 ;
    END
  END E2BEGb[6]
  PIN E2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 222.550 117.150 235.000 117.450 ;
    END
  END E2BEGb[7]
  PIN E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.910 7.910 105.210 ;
    END
  END E2END[0]
  PIN E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.950 13.890 107.250 ;
    END
  END E2END[1]
  PIN E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.310 16.190 108.610 ;
    END
  END E2END[2]
  PIN E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.350 8.830 110.650 ;
    END
  END E2END[3]
  PIN E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.390 6.990 112.690 ;
    END
  END E2END[4]
  PIN E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.750 17.570 114.050 ;
    END
  END E2END[5]
  PIN E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.790 9.290 116.090 ;
    END
  END E2END[6]
  PIN E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.150 14.350 117.450 ;
    END
  END E2END[7]
  PIN E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.310 20.330 91.610 ;
    END
  END E2MID[0]
  PIN E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.670 17.110 92.970 ;
    END
  END E2MID[1]
  PIN E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.710 18.030 95.010 ;
    END
  END E2MID[2]
  PIN E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.070 19.870 96.370 ;
    END
  END E2MID[3]
  PIN E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.110 18.490 98.410 ;
    END
  END E2MID[4]
  PIN E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.150 19.870 100.450 ;
    END
  END E2MID[5]
  PIN E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.510 20.330 101.810 ;
    END
  END E2MID[6]
  PIN E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.550 8.890 103.850 ;
    END
  END E2MID[7]
  PIN E6BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 225.310 147.070 235.000 147.370 ;
    END
  END E6BEG[0]
  PIN E6BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 225.310 164.070 235.000 164.370 ;
    END
  END E6BEG[10]
  PIN E6BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 225.310 166.110 235.000 166.410 ;
    END
  END E6BEG[11]
  PIN E6BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 220.710 148.430 235.000 148.730 ;
    END
  END E6BEG[1]
  PIN E6BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 225.770 150.470 235.000 150.770 ;
    END
  END E6BEG[2]
  PIN E6BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 219.790 151.830 235.000 152.130 ;
    END
  END E6BEG[3]
  PIN E6BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 223.930 153.870 235.000 154.170 ;
    END
  END E6BEG[4]
  PIN E6BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 224.790 155.910 235.000 156.210 ;
    END
  END E6BEG[5]
  PIN E6BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 228.470 157.270 235.000 157.570 ;
    END
  END E6BEG[6]
  PIN E6BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.870 159.310 235.000 159.610 ;
    END
  END E6BEG[7]
  PIN E6BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 220.250 160.670 235.000 160.970 ;
    END
  END E6BEG[8]
  PIN E6BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 220.710 162.710 235.000 163.010 ;
    END
  END E6BEG[9]
  PIN E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.070 7.450 147.370 ;
    END
  END E6END[0]
  PIN E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.070 19.410 164.370 ;
    END
  END E6END[10]
  PIN E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.110 14.350 166.410 ;
    END
  END E6END[11]
  PIN E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.430 6.990 148.730 ;
    END
  END E6END[1]
  PIN E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 150.470 20.330 150.770 ;
    END
  END E6END[2]
  PIN E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.830 18.950 152.130 ;
    END
  END E6END[3]
  PIN E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.870 18.030 154.170 ;
    END
  END E6END[4]
  PIN E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.910 19.870 156.210 ;
    END
  END E6END[5]
  PIN E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.270 18.950 157.570 ;
    END
  END E6END[6]
  PIN E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.310 20.330 159.610 ;
    END
  END E6END[7]
  PIN E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.670 18.030 160.970 ;
    END
  END E6END[8]
  PIN E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.710 3.770 163.010 ;
    END
  END E6END[9]
  PIN EE4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.570 119.190 235.000 119.490 ;
    END
  END EE4BEG[0]
  PIN EE4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 217.490 136.190 235.000 136.490 ;
    END
  END EE4BEG[10]
  PIN EE4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 220.710 138.230 235.000 138.530 ;
    END
  END EE4BEG[11]
  PIN EE4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.730 140.270 235.000 140.570 ;
    END
  END EE4BEG[12]
  PIN EE4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 217.950 141.630 235.000 141.930 ;
    END
  END EE4BEG[13]
  PIN EE4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 219.330 143.670 235.000 143.970 ;
    END
  END EE4BEG[14]
  PIN EE4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 219.790 145.030 235.000 145.330 ;
    END
  END EE4BEG[15]
  PIN EE4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 233.990 120.550 235.000 120.850 ;
    END
  END EE4BEG[1]
  PIN EE4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 224.850 122.590 235.000 122.890 ;
    END
  END EE4BEG[2]
  PIN EE4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 207.830 123.950 235.000 124.250 ;
    END
  END EE4BEG[3]
  PIN EE4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 212.140 125.990 235.000 126.290 ;
    END
  END EE4BEG[4]
  PIN EE4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 225.310 128.030 235.000 128.330 ;
    END
  END EE4BEG[5]
  PIN EE4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 211.510 129.390 235.000 129.690 ;
    END
  END EE4BEG[6]
  PIN EE4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 220.250 131.430 235.000 131.730 ;
    END
  END EE4BEG[7]
  PIN EE4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 212.430 132.790 235.000 133.090 ;
    END
  END EE4BEG[8]
  PIN EE4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.570 134.830 235.000 135.130 ;
    END
  END EE4BEG[9]
  PIN EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.190 19.870 119.490 ;
    END
  END EE4END[0]
  PIN EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.190 6.130 136.490 ;
    END
  END EE4END[10]
  PIN EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.230 19.870 138.530 ;
    END
  END EE4END[11]
  PIN EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.270 21.250 140.570 ;
    END
  END EE4END[12]
  PIN EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.630 13.890 141.930 ;
    END
  END EE4END[13]
  PIN EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.670 20.330 143.970 ;
    END
  END EE4END[14]
  PIN EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.030 13.950 145.330 ;
    END
  END EE4END[15]
  PIN EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.550 18.950 120.850 ;
    END
  END EE4END[1]
  PIN EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.590 13.890 122.890 ;
    END
  END EE4END[2]
  PIN EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.950 12.970 124.250 ;
    END
  END EE4END[3]
  PIN EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.990 19.870 126.290 ;
    END
  END EE4END[4]
  PIN EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.030 18.490 128.330 ;
    END
  END EE4END[5]
  PIN EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.390 18.950 129.690 ;
    END
  END EE4END[6]
  PIN EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.430 16.190 131.730 ;
    END
  END EE4END[7]
  PIN EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.790 20.620 133.090 ;
    END
  END EE4END[8]
  PIN EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.830 42.870 135.130 ;
    END
  END EE4END[9]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.150 13.890 168.450 ;
    END
  END FrameData[0]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.150 20.330 185.450 ;
    END
  END FrameData[10]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.190 19.870 187.490 ;
    END
  END FrameData[11]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 188.550 6.990 188.850 ;
    END
  END FrameData[12]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.590 6.990 190.890 ;
    END
  END FrameData[13]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.950 7.450 192.250 ;
    END
  END FrameData[14]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.990 9.750 194.290 ;
    END
  END FrameData[15]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.030 34.590 196.330 ;
    END
  END FrameData[16]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.390 18.030 197.690 ;
    END
  END FrameData[17]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.430 28.150 199.730 ;
    END
  END FrameData[18]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.790 21.080 201.090 ;
    END
  END FrameData[19]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 169.510 14.810 169.810 ;
    END
  END FrameData[1]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.830 16.650 203.130 ;
    END
  END FrameData[20]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.190 20.330 204.490 ;
    END
  END FrameData[21]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.230 26.770 206.530 ;
    END
  END FrameData[22]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.590 18.950 207.890 ;
    END
  END FrameData[23]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.630 20.330 209.930 ;
    END
  END FrameData[24]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 211.670 37.350 211.970 ;
    END
  END FrameData[25]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.030 6.990 213.330 ;
    END
  END FrameData[26]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.070 18.950 215.370 ;
    END
  END FrameData[27]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.430 16.190 216.730 ;
    END
  END FrameData[28]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 218.470 7.450 218.770 ;
    END
  END FrameData[29]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.550 18.950 171.850 ;
    END
  END FrameData[2]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.830 6.530 220.130 ;
    END
  END FrameData[30]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.870 14.350 222.170 ;
    END
  END FrameData[31]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.910 6.990 173.210 ;
    END
  END FrameData[3]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.950 7.450 175.250 ;
    END
  END FrameData[4]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.310 7.450 176.610 ;
    END
  END FrameData[5]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.350 6.530 178.650 ;
    END
  END FrameData[6]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.710 18.950 180.010 ;
    END
  END FrameData[7]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 181.750 20.330 182.050 ;
    END
  END FrameData[8]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.790 7.450 184.090 ;
    END
  END FrameData[9]
  PIN FrameData_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 227.610 168.150 235.000 168.450 ;
    END
  END FrameData_O[0]
  PIN FrameData_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 225.310 185.150 235.000 185.450 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 225.310 187.190 235.000 187.490 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 222.090 188.550 235.000 188.850 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 225.770 190.590 235.000 190.890 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 227.610 191.950 235.000 192.250 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 222.550 193.990 235.000 194.290 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 222.090 196.030 235.000 196.330 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 225.770 197.390 235.000 197.690 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 222.550 199.430 235.000 199.730 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 220.710 200.790 235.000 201.090 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.630 169.510 235.000 169.810 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 226.690 202.830 235.000 203.130 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 222.090 204.190 235.000 204.490 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 224.390 206.230 235.000 206.530 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.870 207.590 235.000 207.890 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 220.710 209.630 235.000 209.930 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 222.550 211.670 235.000 211.970 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.870 213.030 235.000 213.330 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.870 215.070 235.000 215.370 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 215.650 216.430 235.000 216.730 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.110 218.470 235.000 218.770 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.870 171.550 235.000 171.850 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 219.330 219.830 235.000 220.130 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 221.870 235.000 222.170 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 215.190 172.910 235.000 173.210 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 222.550 174.950 235.000 175.250 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.410 176.310 235.000 176.610 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 227.610 178.350 235.000 178.650 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 220.710 179.710 235.000 180.010 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 219.790 181.750 235.000 182.050 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 220.250 183.790 235.000 184.090 ;
    END
  END FrameData_O[9]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.420 0.000 198.560 6.500 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.280 0.000 217.420 6.500 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.120 0.000 219.260 11.940 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.960 0.000 221.100 4.800 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.800 0.000 222.940 18.560 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.640 0.000 224.780 15.680 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.480 0.000 226.620 14.480 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.320 0.000 228.460 15.160 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.160 0.000 230.300 15.840 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.000 0.000 232.140 18.400 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.840 0.000 233.980 13.800 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.260 0.000 200.400 20.440 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.100 0.000 202.240 1.400 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.940 0.000 204.080 7.210 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.780 0.000 205.920 1.090 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.620 0.000 207.760 25.880 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.460 0.000 209.600 15.680 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.300 0.000 211.440 6.700 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.140 0.000 213.280 2.420 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.440 0.000 215.580 4.120 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.960 212.600 198.100 223.115 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.820 208.720 216.960 223.115 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.660 216.510 218.800 223.115 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.960 203.280 221.100 223.115 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.800 218.240 222.940 223.115 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.640 209.060 224.780 223.115 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.480 211.780 226.620 223.115 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.320 206.340 228.460 223.115 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.160 211.440 230.300 223.115 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.000 202.940 232.140 223.115 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.840 202.600 233.980 223.115 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.800 209.060 199.940 223.115 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.640 206.340 201.780 223.115 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.480 206.000 203.620 223.115 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.780 206.930 205.920 223.115 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.620 199.880 207.760 223.115 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.460 207.840 209.600 223.115 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.300 193.760 211.440 223.115 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.140 204.980 213.280 223.115 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.980 214.470 215.120 223.115 ;
    END
  END FrameStrobe_O[9]
  PIN N1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.080 199.880 1.220 223.115 ;
    END
  END N1BEG[0]
  PIN N1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.920 211.780 3.060 223.115 ;
    END
  END N1BEG[1]
  PIN N1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.760 206.340 4.900 223.115 ;
    END
  END N1BEG[2]
  PIN N1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.600 220.590 6.740 223.115 ;
    END
  END N1BEG[3]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.080 0.000 1.220 10.240 ;
    END
  END N1END[0]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.920 0.000 3.060 6.500 ;
    END
  END N1END[1]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.760 0.000 4.900 9.560 ;
    END
  END N1END[2]
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.600 0.000 6.740 17.380 ;
    END
  END N1END[3]
  PIN N2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.440 206.930 8.580 223.115 ;
    END
  END N2BEG[0]
  PIN N2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.280 202.440 10.420 223.115 ;
    END
  END N2BEG[1]
  PIN N2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.120 201.920 12.260 223.115 ;
    END
  END N2BEG[2]
  PIN N2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.960 216.880 14.100 223.115 ;
    END
  END N2BEG[3]
  PIN N2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.800 221.950 15.940 223.115 ;
    END
  END N2BEG[4]
  PIN N2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.100 221.950 18.240 223.115 ;
    END
  END N2BEG[5]
  PIN N2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.940 221.270 20.080 223.115 ;
    END
  END N2BEG[6]
  PIN N2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.780 215.860 21.920 223.115 ;
    END
  END N2BEG[7]
  PIN N2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.620 202.600 23.760 223.115 ;
    END
  END N2BEGb[0]
  PIN N2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.460 201.920 25.600 223.115 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.300 218.580 27.440 223.115 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.140 217.020 29.280 223.115 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.980 206.930 31.120 223.115 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.280 206.930 33.420 223.115 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.120 221.950 35.260 223.115 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.960 218.240 37.100 223.115 ;
    END
  END N2BEGb[7]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.620 0.000 23.760 11.940 ;
    END
  END N2END[0]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.460 0.000 25.600 3.780 ;
    END
  END N2END[1]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.300 0.000 27.440 7.210 ;
    END
  END N2END[2]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.140 0.000 29.280 20.440 ;
    END
  END N2END[3]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.980 0.000 31.120 6.160 ;
    END
  END N2END[4]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.820 0.000 32.960 13.980 ;
    END
  END N2END[5]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.660 0.000 34.800 3.440 ;
    END
  END N2END[6]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.500 0.000 36.640 1.740 ;
    END
  END N2END[7]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.440 0.000 8.580 5.850 ;
    END
  END N2MID[0]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.280 0.000 10.420 7.890 ;
    END
  END N2MID[1]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.120 0.000 12.260 28.260 ;
    END
  END N2MID[2]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.960 0.000 14.100 28.600 ;
    END
  END N2MID[3]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.800 0.000 15.940 5.170 ;
    END
  END N2MID[4]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.640 0.000 17.780 14.660 ;
    END
  END N2MID[5]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.480 0.000 19.620 4.120 ;
    END
  END N2MID[6]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.320 0.000 21.460 7.180 ;
    END
  END N2MID[7]
  PIN N4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.800 213.110 38.940 223.115 ;
    END
  END N4BEG[0]
  PIN N4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.660 203.620 57.800 223.115 ;
    END
  END N4BEG[10]
  PIN N4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.500 204.980 59.640 223.115 ;
    END
  END N4BEG[11]
  PIN N4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.340 206.340 61.480 223.115 ;
    END
  END N4BEG[12]
  PIN N4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.180 214.500 63.320 223.115 ;
    END
  END N4BEG[13]
  PIN N4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.480 206.930 65.620 223.115 ;
    END
  END N4BEG[14]
  PIN N4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.320 221.980 67.460 223.115 ;
    END
  END N4BEG[15]
  PIN N4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.640 189.680 40.780 223.115 ;
    END
  END N4BEG[1]
  PIN N4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.480 214.470 42.620 223.115 ;
    END
  END N4BEG[2]
  PIN N4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.320 211.960 44.460 223.115 ;
    END
  END N4BEG[3]
  PIN N4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.160 214.470 46.300 223.115 ;
    END
  END N4BEG[4]
  PIN N4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.460 215.360 48.600 223.115 ;
    END
  END N4BEG[5]
  PIN N4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.300 221.950 50.440 223.115 ;
    END
  END N4BEG[6]
  PIN N4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.140 214.470 52.280 223.115 ;
    END
  END N4BEG[7]
  PIN N4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.980 206.000 54.120 223.115 ;
    END
  END N4BEG[8]
  PIN N4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.820 214.470 55.960 223.115 ;
    END
  END N4BEG[9]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.340 0.000 38.480 3.100 ;
    END
  END N4END[0]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.200 0.000 57.340 9.560 ;
    END
  END N4END[10]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.040 0.000 59.180 31.320 ;
    END
  END N4END[11]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.880 0.000 61.020 18.560 ;
    END
  END N4END[12]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.720 0.000 62.860 5.170 ;
    END
  END N4END[13]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.560 0.000 64.700 7.210 ;
    END
  END N4END[14]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.860 0.000 67.000 1.090 ;
    END
  END N4END[15]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.180 0.000 40.320 19.420 ;
    END
  END N4END[1]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.020 0.000 42.160 10.400 ;
    END
  END N4END[2]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.320 0.000 44.460 17.380 ;
    END
  END N4END[3]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.160 0.000 46.300 31.320 ;
    END
  END N4END[4]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.000 0.000 48.140 14.480 ;
    END
  END N4END[5]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.840 0.000 49.980 9.420 ;
    END
  END N4END[6]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.680 0.000 51.820 21.120 ;
    END
  END N4END[7]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.520 0.000 53.660 11.760 ;
    END
  END N4END[8]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.360 0.000 55.500 2.420 ;
    END
  END N4END[9]
  PIN NN4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.160 203.280 69.300 223.115 ;
    END
  END NN4BEG[0]
  PIN NN4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.020 203.620 88.160 223.115 ;
    END
  END NN4BEG[10]
  PIN NN4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.860 206.520 90.000 223.115 ;
    END
  END NN4BEG[11]
  PIN NN4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.700 214.470 91.840 223.115 ;
    END
  END NN4BEG[12]
  PIN NN4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.540 208.380 93.680 223.115 ;
    END
  END NN4BEG[13]
  PIN NN4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.840 214.470 95.980 223.115 ;
    END
  END NN4BEG[14]
  PIN NN4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.680 218.550 97.820 223.115 ;
    END
  END NN4BEG[15]
  PIN NN4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.000 221.950 71.140 223.115 ;
    END
  END NN4BEG[1]
  PIN NN4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.840 209.060 72.980 223.115 ;
    END
  END NN4BEG[2]
  PIN NN4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.680 205.160 74.820 223.115 ;
    END
  END NN4BEG[3]
  PIN NN4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.520 190.020 76.660 223.115 ;
    END
  END NN4BEG[4]
  PIN NN4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.360 214.470 78.500 223.115 ;
    END
  END NN4BEG[5]
  PIN NN4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.660 205.320 80.800 223.115 ;
    END
  END NN4BEG[6]
  PIN NN4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.500 206.000 82.640 223.115 ;
    END
  END NN4BEG[7]
  PIN NN4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.340 186.960 84.480 223.115 ;
    END
  END NN4BEG[8]
  PIN NN4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.180 206.930 86.320 223.115 ;
    END
  END NN4BEG[9]
  PIN NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.700 0.000 68.840 13.330 ;
    END
  END NN4END[0]
  PIN NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.560 0.000 87.700 15.880 ;
    END
  END NN4END[10]
  PIN NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.400 0.000 89.540 11.080 ;
    END
  END NN4END[11]
  PIN NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.240 0.000 91.380 39.140 ;
    END
  END NN4END[12]
  PIN NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.080 0.000 93.220 15.160 ;
    END
  END NN4END[13]
  PIN NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.920 0.000 95.060 17.240 ;
    END
  END NN4END[14]
  PIN NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.760 0.000 96.900 16.700 ;
    END
  END NN4END[15]
  PIN NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.540 0.000 70.680 1.090 ;
    END
  END NN4END[1]
  PIN NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.380 0.000 72.520 9.560 ;
    END
  END NN4END[2]
  PIN NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.220 0.000 74.360 6.160 ;
    END
  END NN4END[3]
  PIN NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.060 0.000 76.200 14.180 ;
    END
  END NN4END[4]
  PIN NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.900 0.000 78.040 42.200 ;
    END
  END NN4END[5]
  PIN NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.740 0.000 79.880 39.820 ;
    END
  END NN4END[6]
  PIN NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.580 0.000 81.720 20.100 ;
    END
  END NN4END[7]
  PIN NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.420 0.000 83.560 44.580 ;
    END
  END NN4END[8]
  PIN NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.260 0.000 85.400 15.680 ;
    END
  END NN4END[9]
  PIN S1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.600 0.000 98.740 3.100 ;
    END
  END S1BEG[0]
  PIN S1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.440 0.000 100.580 7.210 ;
    END
  END S1BEG[1]
  PIN S1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.280 0.000 102.420 1.740 ;
    END
  END S1BEG[2]
  PIN S1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.120 0.000 104.260 8.540 ;
    END
  END S1BEG[3]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.520 219.230 99.660 223.115 ;
    END
  END S1END[0]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.360 216.880 101.500 223.115 ;
    END
  END S1END[1]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.200 214.500 103.340 223.115 ;
    END
  END S1END[2]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.040 211.440 105.180 223.115 ;
    END
  END S1END[3]
  PIN S2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.140 0.000 121.280 6.500 ;
    END
  END S2BEG[0]
  PIN S2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.980 0.000 123.120 6.020 ;
    END
  END S2BEG[1]
  PIN S2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.820 0.000 124.960 2.760 ;
    END
  END S2BEG[2]
  PIN S2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.660 0.000 126.800 1.090 ;
    END
  END S2BEG[3]
  PIN S2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.500 0.000 128.640 3.100 ;
    END
  END S2BEG[4]
  PIN S2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.800 0.000 130.940 1.740 ;
    END
  END S2BEG[5]
  PIN S2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.640 0.000 132.780 13.980 ;
    END
  END S2BEG[6]
  PIN S2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.480 0.000 134.620 8.540 ;
    END
  END S2BEG[7]
  PIN S2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.960 0.000 106.100 13.980 ;
    END
  END S2BEGb[0]
  PIN S2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.260 0.000 108.400 11.260 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.100 0.000 110.240 3.810 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.940 0.000 112.080 15.680 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.780 0.000 113.920 5.170 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.620 0.000 115.760 11.290 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.460 0.000 117.600 1.940 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.300 0.000 119.440 18.060 ;
    END
  END S2BEGb[7]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.880 216.540 107.020 223.115 ;
    END
  END S2END[0]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.720 221.640 108.860 223.115 ;
    END
  END S2END[1]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.020 221.980 111.160 223.115 ;
    END
  END S2END[2]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.860 221.950 113.000 223.115 ;
    END
  END S2END[3]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.700 206.340 114.840 223.115 ;
    END
  END S2END[4]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.540 221.300 116.680 223.115 ;
    END
  END S2END[5]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.380 208.040 118.520 223.115 ;
    END
  END S2END[6]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.220 200.560 120.360 223.115 ;
    END
  END S2END[7]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.060 207.200 122.200 223.115 ;
    END
  END S2MID[0]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.900 202.910 124.040 223.115 ;
    END
  END S2MID[1]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.740 214.470 125.880 223.115 ;
    END
  END S2MID[2]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.040 215.660 128.180 223.115 ;
    END
  END S2MID[3]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.880 201.920 130.020 223.115 ;
    END
  END S2MID[4]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.720 206.930 131.860 223.115 ;
    END
  END S2MID[5]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.560 204.980 133.700 223.115 ;
    END
  END S2MID[6]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.400 201.920 135.540 223.115 ;
    END
  END S2MID[7]
  PIN S4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.320 0.000 136.460 2.080 ;
    END
  END S4BEG[0]
  PIN S4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.180 0.000 155.320 5.850 ;
    END
  END S4BEG[10]
  PIN S4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.020 0.000 157.160 4.120 ;
    END
  END S4BEG[11]
  PIN S4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.860 0.000 159.000 7.210 ;
    END
  END S4BEG[12]
  PIN S4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.700 0.000 160.840 24.860 ;
    END
  END S4BEG[13]
  PIN S4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.540 0.000 162.680 27.580 ;
    END
  END S4BEG[14]
  PIN S4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.380 0.000 164.520 3.810 ;
    END
  END S4BEG[15]
  PIN S4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.160 0.000 138.300 13.870 ;
    END
  END S4BEG[1]
  PIN S4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.000 0.000 140.140 19.760 ;
    END
  END S4BEG[2]
  PIN S4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.840 0.000 141.980 20.100 ;
    END
  END S4BEG[3]
  PIN S4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.680 0.000 143.820 7.210 ;
    END
  END S4BEG[4]
  PIN S4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.520 0.000 145.660 13.870 ;
    END
  END S4BEG[5]
  PIN S4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.360 0.000 147.500 4.460 ;
    END
  END S4BEG[6]
  PIN S4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.200 0.000 149.340 30.300 ;
    END
  END S4BEG[7]
  PIN S4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.500 0.000 151.640 28.260 ;
    END
  END S4BEG[8]
  PIN S4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.340 0.000 153.480 1.090 ;
    END
  END S4BEG[9]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.240 203.280 137.380 223.115 ;
    END
  END S4END[0]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.100 216.720 156.240 223.115 ;
    END
  END S4END[10]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.400 212.430 158.540 223.115 ;
    END
  END S4END[11]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.240 196.790 160.380 223.115 ;
    END
  END S4END[12]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.080 151.260 162.220 223.115 ;
    END
  END S4END[13]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.920 206.930 164.060 223.115 ;
    END
  END S4END[14]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.760 202.740 165.900 223.115 ;
    END
  END S4END[15]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.080 216.880 139.220 223.115 ;
    END
  END S4END[1]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.920 219.230 141.060 223.115 ;
    END
  END S4END[2]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.220 207.670 143.360 223.115 ;
    END
  END S4END[3]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.060 179.320 145.200 223.115 ;
    END
  END S4END[4]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.900 216.720 147.040 223.115 ;
    END
  END S4END[5]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.740 207.200 148.880 223.115 ;
    END
  END S4END[6]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.580 214.500 150.720 223.115 ;
    END
  END S4END[7]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.420 206.930 152.560 223.115 ;
    END
  END S4END[8]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.260 221.950 154.400 223.115 ;
    END
  END S4END[9]
  PIN SS4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.220 0.000 166.360 41.520 ;
    END
  END SS4BEG[0]
  PIN SS4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.080 0.000 185.220 3.810 ;
    END
  END SS4BEG[10]
  PIN SS4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.920 0.000 187.060 9.040 ;
    END
  END SS4BEG[11]
  PIN SS4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.760 0.000 188.900 3.100 ;
    END
  END SS4BEG[12]
  PIN SS4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.600 0.000 190.740 1.090 ;
    END
  END SS4BEG[13]
  PIN SS4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.440 0.000 192.580 1.090 ;
    END
  END SS4BEG[14]
  PIN SS4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.740 0.000 194.880 13.870 ;
    END
  END SS4BEG[15]
  PIN SS4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.060 0.000 168.200 3.440 ;
    END
  END SS4BEG[1]
  PIN SS4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.900 0.000 170.040 1.090 ;
    END
  END SS4BEG[2]
  PIN SS4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.200 0.000 172.340 9.040 ;
    END
  END SS4BEG[3]
  PIN SS4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.040 0.000 174.180 13.120 ;
    END
  END SS4BEG[4]
  PIN SS4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.880 0.000 176.020 5.820 ;
    END
  END SS4BEG[5]
  PIN SS4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.720 0.000 177.860 17.410 ;
    END
  END SS4BEG[6]
  PIN SS4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.560 0.000 179.700 11.080 ;
    END
  END SS4BEG[7]
  PIN SS4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.400 0.000 181.540 1.740 ;
    END
  END SS4BEG[8]
  PIN SS4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.240 0.000 183.380 15.370 ;
    END
  END SS4BEG[9]
  PIN SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.600 220.960 167.740 223.115 ;
    END
  END SS4END[0]
  PIN SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.460 218.920 186.600 223.115 ;
    END
  END SS4END[10]
  PIN SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.300 194.100 188.440 223.115 ;
    END
  END SS4END[11]
  PIN SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.600 214.470 190.740 223.115 ;
    END
  END SS4END[12]
  PIN SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.440 216.040 192.580 223.115 ;
    END
  END SS4END[13]
  PIN SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.280 202.940 194.420 223.115 ;
    END
  END SS4END[14]
  PIN SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.120 211.580 196.260 223.115 ;
    END
  END SS4END[15]
  PIN SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.440 200.560 169.580 223.115 ;
    END
  END SS4END[1]
  PIN SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.280 218.240 171.420 223.115 ;
    END
  END SS4END[2]
  PIN SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.580 217.220 173.720 223.115 ;
    END
  END SS4END[3]
  PIN SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.420 221.950 175.560 223.115 ;
    END
  END SS4END[4]
  PIN SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.260 206.930 177.400 223.115 ;
    END
  END SS4END[5]
  PIN SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.100 216.720 179.240 223.115 ;
    END
  END SS4END[6]
  PIN SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.940 214.470 181.080 223.115 ;
    END
  END SS4END[7]
  PIN SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.780 206.000 182.920 223.115 ;
    END
  END SS4END[8]
  PIN SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.620 166.400 184.760 223.115 ;
    END
  END SS4END[9]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.580 0.000 196.720 17.200 ;
    END
  END UserCLK
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 5.200 99.440 217.840 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 5.200 22.640 217.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 5.200 176.240 217.840 ;
    END
  END VPWR
  PIN W1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.870 14.810 1.170 ;
    END
  END W1BEG[0]
  PIN W1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.230 15.270 2.530 ;
    END
  END W1BEG[1]
  PIN W1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.270 6.990 4.570 ;
    END
  END W1BEG[2]
  PIN W1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.630 5.150 5.930 ;
    END
  END W1BEG[3]
  PIN W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 222.550 0.870 235.000 1.170 ;
    END
  END W1END[0]
  PIN W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 219.790 2.230 235.000 2.530 ;
    END
  END W1END[1]
  PIN W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 198.170 4.270 235.000 4.570 ;
    END
  END W1END[2]
  PIN W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 5.630 235.000 5.930 ;
    END
  END W1END[3]
  PIN W2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.670 7.450 7.970 ;
    END
  END W2BEG[0]
  PIN W2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.030 20.330 9.330 ;
    END
  END W2BEG[1]
  PIN W2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.070 7.910 11.370 ;
    END
  END W2BEG[2]
  PIN W2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.430 4.230 12.730 ;
    END
  END W2BEG[3]
  PIN W2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.470 14.350 14.770 ;
    END
  END W2BEG[4]
  PIN W2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.510 20.330 16.810 ;
    END
  END W2BEG[5]
  PIN W2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.870 9.750 18.170 ;
    END
  END W2BEG[6]
  PIN W2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.910 15.730 20.210 ;
    END
  END W2BEG[7]
  PIN W2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.270 17.570 21.570 ;
    END
  END W2BEGb[0]
  PIN W2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.310 11.590 23.610 ;
    END
  END W2BEGb[1]
  PIN W2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.670 3.310 24.970 ;
    END
  END W2BEGb[2]
  PIN W2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.710 24.470 27.010 ;
    END
  END W2BEGb[3]
  PIN W2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.750 23.090 29.050 ;
    END
  END W2BEGb[4]
  PIN W2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.110 13.950 30.410 ;
    END
  END W2BEGb[5]
  PIN W2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.150 20.330 32.450 ;
    END
  END W2BEGb[6]
  PIN W2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.510 29.530 33.810 ;
    END
  END W2BEGb[7]
  PIN W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 220.710 21.270 235.000 21.570 ;
    END
  END W2END[0]
  PIN W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 220.710 23.310 235.000 23.610 ;
    END
  END W2END[1]
  PIN W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 220.710 24.670 235.000 24.970 ;
    END
  END W2END[2]
  PIN W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 222.550 26.710 235.000 27.010 ;
    END
  END W2END[3]
  PIN W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 227.150 28.750 235.000 29.050 ;
    END
  END W2END[4]
  PIN W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 184.830 30.110 235.000 30.410 ;
    END
  END W2END[5]
  PIN W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 220.710 32.150 235.000 32.450 ;
    END
  END W2END[6]
  PIN W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 182.530 33.510 235.000 33.810 ;
    END
  END W2END[7]
  PIN W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.110 7.670 235.000 7.970 ;
    END
  END W2MID[0]
  PIN W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 9.030 235.000 9.330 ;
    END
  END W2MID[1]
  PIN W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 215.190 11.070 235.000 11.370 ;
    END
  END W2MID[2]
  PIN W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 215.190 12.430 235.000 12.730 ;
    END
  END W2MID[3]
  PIN W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 227.610 14.470 235.000 14.770 ;
    END
  END W2MID[4]
  PIN W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 229.910 16.510 235.000 16.810 ;
    END
  END W2MID[5]
  PIN W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.570 17.870 235.000 18.170 ;
    END
  END W2MID[6]
  PIN W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 224.850 19.910 235.000 20.210 ;
    END
  END W2MID[7]
  PIN W6BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.430 9.750 63.730 ;
    END
  END W6BEG[0]
  PIN W6BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.430 6.990 80.730 ;
    END
  END W6BEG[10]
  PIN W6BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.470 20.330 82.770 ;
    END
  END W6BEG[11]
  PIN W6BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.790 9.750 65.090 ;
    END
  END W6BEG[1]
  PIN W6BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.830 9.750 67.130 ;
    END
  END W6BEG[2]
  PIN W6BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.190 13.890 68.490 ;
    END
  END W6BEG[3]
  PIN W6BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.230 17.110 70.530 ;
    END
  END W6BEG[4]
  PIN W6BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.270 13.890 72.570 ;
    END
  END W6BEG[5]
  PIN W6BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.630 17.570 73.930 ;
    END
  END W6BEG[6]
  PIN W6BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.670 11.130 75.970 ;
    END
  END W6BEG[7]
  PIN W6BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.030 14.350 77.330 ;
    END
  END W6BEG[8]
  PIN W6BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.070 20.330 79.370 ;
    END
  END W6BEG[9]
  PIN W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 215.190 63.430 235.000 63.730 ;
    END
  END W6END[0]
  PIN W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.350 80.430 235.000 80.730 ;
    END
  END W6END[10]
  PIN W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 233.990 82.470 235.000 82.770 ;
    END
  END W6END[11]
  PIN W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 220.710 64.790 235.000 65.090 ;
    END
  END W6END[1]
  PIN W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 183.450 66.830 235.000 67.130 ;
    END
  END W6END[2]
  PIN W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 68.190 235.000 68.490 ;
    END
  END W6END[3]
  PIN W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 233.990 70.230 235.000 70.530 ;
    END
  END W6END[4]
  PIN W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.590 72.270 235.000 72.570 ;
    END
  END W6END[5]
  PIN W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 220.250 73.630 235.000 73.930 ;
    END
  END W6END[6]
  PIN W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 217.950 75.670 235.000 75.970 ;
    END
  END W6END[7]
  PIN W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 233.990 77.030 235.000 77.330 ;
    END
  END W6END[8]
  PIN W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.730 79.070 235.000 79.370 ;
    END
  END W6END[9]
  PIN WW4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.550 19.410 35.850 ;
    END
  END WW4BEG[0]
  PIN WW4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.550 10.210 52.850 ;
    END
  END WW4BEG[10]
  PIN WW4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.590 9.750 54.890 ;
    END
  END WW4BEG[11]
  PIN WW4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.630 13.890 56.930 ;
    END
  END WW4BEG[12]
  PIN WW4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.990 19.870 58.290 ;
    END
  END WW4BEG[13]
  PIN WW4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.030 13.890 60.330 ;
    END
  END WW4BEG[14]
  PIN WW4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.390 19.870 61.690 ;
    END
  END WW4BEG[15]
  PIN WW4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.910 19.870 37.210 ;
    END
  END WW4BEG[1]
  PIN WW4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.950 19.870 39.250 ;
    END
  END WW4BEG[2]
  PIN WW4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.310 20.330 40.610 ;
    END
  END WW4BEG[3]
  PIN WW4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.350 13.950 42.650 ;
    END
  END WW4BEG[4]
  PIN WW4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.390 18.490 44.690 ;
    END
  END WW4BEG[5]
  PIN WW4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.750 20.330 46.050 ;
    END
  END WW4BEG[6]
  PIN WW4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.790 18.950 48.090 ;
    END
  END WW4BEG[7]
  PIN WW4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.150 15.730 49.450 ;
    END
  END WW4BEG[8]
  PIN WW4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.190 18.030 51.490 ;
    END
  END WW4BEG[9]
  PIN WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 212.890 35.550 235.000 35.850 ;
    END
  END WW4END[0]
  PIN WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 233.990 52.550 235.000 52.850 ;
    END
  END WW4END[10]
  PIN WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 220.710 54.590 235.000 54.890 ;
    END
  END WW4END[11]
  PIN WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.110 56.630 235.000 56.930 ;
    END
  END WW4END[12]
  PIN WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 233.990 57.990 235.000 58.290 ;
    END
  END WW4END[13]
  PIN WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 215.650 60.030 235.000 60.330 ;
    END
  END WW4END[14]
  PIN WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 187.590 61.390 235.000 61.690 ;
    END
  END WW4END[15]
  PIN WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 215.650 36.910 235.000 37.210 ;
    END
  END WW4END[1]
  PIN WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 220.250 38.950 235.000 39.250 ;
    END
  END WW4END[2]
  PIN WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 211.970 40.310 235.000 40.610 ;
    END
  END WW4END[3]
  PIN WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 217.490 42.350 235.000 42.650 ;
    END
  END WW4END[4]
  PIN WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 233.990 44.390 235.000 44.690 ;
    END
  END WW4END[5]
  PIN WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 229.390 45.750 235.000 46.050 ;
    END
  END WW4END[6]
  PIN WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 233.990 47.790 235.000 48.090 ;
    END
  END WW4END[7]
  PIN WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 220.710 49.150 235.000 49.450 ;
    END
  END WW4END[8]
  PIN WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 233.990 51.190 235.000 51.490 ;
    END
  END WW4END[9]
  OBS
      LAYER li1 ;
        RECT 4.745 2.805 233.075 221.255 ;
      LAYER met1 ;
        RECT 0.990 1.400 234.530 221.980 ;
      LAYER met2 ;
        RECT 1.500 211.500 2.640 222.770 ;
        RECT 3.340 211.500 4.480 222.770 ;
        RECT 1.500 206.060 4.480 211.500 ;
        RECT 5.180 220.310 6.320 222.770 ;
        RECT 7.020 220.310 8.160 222.770 ;
        RECT 5.180 206.650 8.160 220.310 ;
        RECT 8.860 206.650 10.000 222.770 ;
        RECT 5.180 206.060 10.000 206.650 ;
        RECT 1.500 202.160 10.000 206.060 ;
        RECT 10.700 202.160 11.840 222.770 ;
        RECT 1.500 201.640 11.840 202.160 ;
        RECT 12.540 216.600 13.680 222.770 ;
        RECT 14.380 221.670 15.520 222.770 ;
        RECT 16.220 221.670 17.820 222.770 ;
        RECT 18.520 221.670 19.660 222.770 ;
        RECT 14.380 220.990 19.660 221.670 ;
        RECT 20.360 220.990 21.500 222.770 ;
        RECT 14.380 216.600 21.500 220.990 ;
        RECT 12.540 215.580 21.500 216.600 ;
        RECT 22.200 215.580 23.340 222.770 ;
        RECT 12.540 202.320 23.340 215.580 ;
        RECT 24.040 202.320 25.180 222.770 ;
        RECT 12.540 201.640 25.180 202.320 ;
        RECT 25.880 218.300 27.020 222.770 ;
        RECT 27.720 218.300 28.860 222.770 ;
        RECT 25.880 216.740 28.860 218.300 ;
        RECT 29.560 216.740 30.700 222.770 ;
        RECT 25.880 206.650 30.700 216.740 ;
        RECT 31.400 206.650 33.000 222.770 ;
        RECT 33.700 221.670 34.840 222.770 ;
        RECT 35.540 221.670 36.680 222.770 ;
        RECT 33.700 217.960 36.680 221.670 ;
        RECT 37.380 217.960 38.520 222.770 ;
        RECT 33.700 212.830 38.520 217.960 ;
        RECT 39.220 212.830 40.360 222.770 ;
        RECT 33.700 206.650 40.360 212.830 ;
        RECT 25.880 201.640 40.360 206.650 ;
        RECT 1.500 199.600 40.360 201.640 ;
        RECT 1.020 189.400 40.360 199.600 ;
        RECT 41.060 214.190 42.200 222.770 ;
        RECT 42.900 214.190 44.040 222.770 ;
        RECT 41.060 211.680 44.040 214.190 ;
        RECT 44.740 214.190 45.880 222.770 ;
        RECT 46.580 215.080 48.180 222.770 ;
        RECT 48.880 221.670 50.020 222.770 ;
        RECT 50.720 221.670 51.860 222.770 ;
        RECT 48.880 215.080 51.860 221.670 ;
        RECT 46.580 214.190 51.860 215.080 ;
        RECT 52.560 214.190 53.700 222.770 ;
        RECT 44.740 211.680 53.700 214.190 ;
        RECT 41.060 205.720 53.700 211.680 ;
        RECT 54.400 214.190 55.540 222.770 ;
        RECT 56.240 214.190 57.380 222.770 ;
        RECT 54.400 205.720 57.380 214.190 ;
        RECT 41.060 203.340 57.380 205.720 ;
        RECT 58.080 204.700 59.220 222.770 ;
        RECT 59.920 206.060 61.060 222.770 ;
        RECT 61.760 214.220 62.900 222.770 ;
        RECT 63.600 214.220 65.200 222.770 ;
        RECT 61.760 206.650 65.200 214.220 ;
        RECT 65.900 221.700 67.040 222.770 ;
        RECT 67.740 221.700 68.880 222.770 ;
        RECT 65.900 206.650 68.880 221.700 ;
        RECT 61.760 206.060 68.880 206.650 ;
        RECT 59.920 204.700 68.880 206.060 ;
        RECT 58.080 203.340 68.880 204.700 ;
        RECT 41.060 203.000 68.880 203.340 ;
        RECT 69.580 221.670 70.720 222.770 ;
        RECT 71.420 221.670 72.560 222.770 ;
        RECT 69.580 208.780 72.560 221.670 ;
        RECT 73.260 208.780 74.400 222.770 ;
        RECT 69.580 204.880 74.400 208.780 ;
        RECT 75.100 204.880 76.240 222.770 ;
        RECT 69.580 203.000 76.240 204.880 ;
        RECT 41.060 189.740 76.240 203.000 ;
        RECT 76.940 214.190 78.080 222.770 ;
        RECT 78.780 214.190 80.380 222.770 ;
        RECT 76.940 205.040 80.380 214.190 ;
        RECT 81.080 205.720 82.220 222.770 ;
        RECT 82.920 205.720 84.060 222.770 ;
        RECT 81.080 205.040 84.060 205.720 ;
        RECT 76.940 189.740 84.060 205.040 ;
        RECT 41.060 189.400 84.060 189.740 ;
        RECT 1.020 186.680 84.060 189.400 ;
        RECT 84.760 206.650 85.900 222.770 ;
        RECT 86.600 206.650 87.740 222.770 ;
        RECT 84.760 203.340 87.740 206.650 ;
        RECT 88.440 206.240 89.580 222.770 ;
        RECT 90.280 214.190 91.420 222.770 ;
        RECT 92.120 214.190 93.260 222.770 ;
        RECT 90.280 208.100 93.260 214.190 ;
        RECT 93.960 214.190 95.560 222.770 ;
        RECT 96.260 218.270 97.400 222.770 ;
        RECT 98.100 218.950 99.240 222.770 ;
        RECT 99.940 218.950 101.080 222.770 ;
        RECT 98.100 218.270 101.080 218.950 ;
        RECT 96.260 216.600 101.080 218.270 ;
        RECT 101.780 216.600 102.920 222.770 ;
        RECT 96.260 214.220 102.920 216.600 ;
        RECT 103.620 214.220 104.760 222.770 ;
        RECT 96.260 214.190 104.760 214.220 ;
        RECT 93.960 211.160 104.760 214.190 ;
        RECT 105.460 216.260 106.600 222.770 ;
        RECT 107.300 221.360 108.440 222.770 ;
        RECT 109.140 221.700 110.740 222.770 ;
        RECT 111.440 221.700 112.580 222.770 ;
        RECT 109.140 221.670 112.580 221.700 ;
        RECT 113.280 221.670 114.420 222.770 ;
        RECT 109.140 221.360 114.420 221.670 ;
        RECT 107.300 216.260 114.420 221.360 ;
        RECT 105.460 211.160 114.420 216.260 ;
        RECT 93.960 208.100 114.420 211.160 ;
        RECT 90.280 206.240 114.420 208.100 ;
        RECT 88.440 206.060 114.420 206.240 ;
        RECT 115.120 221.020 116.260 222.770 ;
        RECT 116.960 221.020 118.100 222.770 ;
        RECT 115.120 207.760 118.100 221.020 ;
        RECT 118.800 207.760 119.940 222.770 ;
        RECT 115.120 206.060 119.940 207.760 ;
        RECT 88.440 203.340 119.940 206.060 ;
        RECT 84.760 200.280 119.940 203.340 ;
        RECT 120.640 206.920 121.780 222.770 ;
        RECT 122.480 206.920 123.620 222.770 ;
        RECT 120.640 202.630 123.620 206.920 ;
        RECT 124.320 214.190 125.460 222.770 ;
        RECT 126.160 215.380 127.760 222.770 ;
        RECT 128.460 215.380 129.600 222.770 ;
        RECT 126.160 214.190 129.600 215.380 ;
        RECT 124.320 202.630 129.600 214.190 ;
        RECT 120.640 201.640 129.600 202.630 ;
        RECT 130.300 206.650 131.440 222.770 ;
        RECT 132.140 206.650 133.280 222.770 ;
        RECT 130.300 204.700 133.280 206.650 ;
        RECT 133.980 204.700 135.120 222.770 ;
        RECT 130.300 201.640 135.120 204.700 ;
        RECT 135.820 203.000 136.960 222.770 ;
        RECT 137.660 216.600 138.800 222.770 ;
        RECT 139.500 218.950 140.640 222.770 ;
        RECT 141.340 218.950 142.940 222.770 ;
        RECT 139.500 216.600 142.940 218.950 ;
        RECT 137.660 207.390 142.940 216.600 ;
        RECT 143.640 207.390 144.780 222.770 ;
        RECT 137.660 203.000 144.780 207.390 ;
        RECT 135.820 201.640 144.780 203.000 ;
        RECT 120.640 200.280 144.780 201.640 ;
        RECT 84.760 186.680 144.780 200.280 ;
        RECT 1.020 179.040 144.780 186.680 ;
        RECT 145.480 216.440 146.620 222.770 ;
        RECT 147.320 216.440 148.460 222.770 ;
        RECT 145.480 206.920 148.460 216.440 ;
        RECT 149.160 214.220 150.300 222.770 ;
        RECT 151.000 214.220 152.140 222.770 ;
        RECT 149.160 206.920 152.140 214.220 ;
        RECT 145.480 206.650 152.140 206.920 ;
        RECT 152.840 221.670 153.980 222.770 ;
        RECT 154.680 221.670 155.820 222.770 ;
        RECT 152.840 216.440 155.820 221.670 ;
        RECT 156.520 216.440 158.120 222.770 ;
        RECT 152.840 212.150 158.120 216.440 ;
        RECT 158.820 212.150 159.960 222.770 ;
        RECT 152.840 206.650 159.960 212.150 ;
        RECT 145.480 196.510 159.960 206.650 ;
        RECT 160.660 196.510 161.800 222.770 ;
        RECT 145.480 179.040 161.800 196.510 ;
        RECT 1.020 150.980 161.800 179.040 ;
        RECT 162.500 206.650 163.640 222.770 ;
        RECT 164.340 206.650 165.480 222.770 ;
        RECT 162.500 202.460 165.480 206.650 ;
        RECT 166.180 220.680 167.320 222.770 ;
        RECT 168.020 220.680 169.160 222.770 ;
        RECT 166.180 202.460 169.160 220.680 ;
        RECT 162.500 200.280 169.160 202.460 ;
        RECT 169.860 217.960 171.000 222.770 ;
        RECT 171.700 217.960 173.300 222.770 ;
        RECT 169.860 216.940 173.300 217.960 ;
        RECT 174.000 221.670 175.140 222.770 ;
        RECT 175.840 221.670 176.980 222.770 ;
        RECT 174.000 216.940 176.980 221.670 ;
        RECT 169.860 206.650 176.980 216.940 ;
        RECT 177.680 216.440 178.820 222.770 ;
        RECT 179.520 216.440 180.660 222.770 ;
        RECT 177.680 214.190 180.660 216.440 ;
        RECT 181.360 214.190 182.500 222.770 ;
        RECT 177.680 206.650 182.500 214.190 ;
        RECT 169.860 205.720 182.500 206.650 ;
        RECT 183.200 205.720 184.340 222.770 ;
        RECT 169.860 200.280 184.340 205.720 ;
        RECT 162.500 166.120 184.340 200.280 ;
        RECT 185.040 218.640 186.180 222.770 ;
        RECT 186.880 218.640 188.020 222.770 ;
        RECT 185.040 193.820 188.020 218.640 ;
        RECT 188.720 214.190 190.320 222.770 ;
        RECT 191.020 215.760 192.160 222.770 ;
        RECT 192.860 215.760 194.000 222.770 ;
        RECT 191.020 214.190 194.000 215.760 ;
        RECT 188.720 202.660 194.000 214.190 ;
        RECT 194.700 211.300 195.840 222.770 ;
        RECT 196.540 212.320 197.680 222.770 ;
        RECT 198.380 212.320 199.520 222.770 ;
        RECT 196.540 211.300 199.520 212.320 ;
        RECT 194.700 208.780 199.520 211.300 ;
        RECT 200.220 208.780 201.360 222.770 ;
        RECT 194.700 206.060 201.360 208.780 ;
        RECT 202.060 206.060 203.200 222.770 ;
        RECT 194.700 205.720 203.200 206.060 ;
        RECT 203.900 206.650 205.500 222.770 ;
        RECT 206.200 206.650 207.340 222.770 ;
        RECT 203.900 205.720 207.340 206.650 ;
        RECT 194.700 202.660 207.340 205.720 ;
        RECT 188.720 199.600 207.340 202.660 ;
        RECT 208.040 207.560 209.180 222.770 ;
        RECT 209.880 207.560 211.020 222.770 ;
        RECT 208.040 199.600 211.020 207.560 ;
        RECT 188.720 193.820 211.020 199.600 ;
        RECT 185.040 193.480 211.020 193.820 ;
        RECT 211.720 204.700 212.860 222.770 ;
        RECT 213.560 214.190 214.700 222.770 ;
        RECT 215.400 214.190 216.540 222.770 ;
        RECT 213.560 208.440 216.540 214.190 ;
        RECT 217.240 216.230 218.380 222.770 ;
        RECT 219.080 216.230 220.680 222.770 ;
        RECT 217.240 208.440 220.680 216.230 ;
        RECT 213.560 204.700 220.680 208.440 ;
        RECT 211.720 203.000 220.680 204.700 ;
        RECT 221.380 217.960 222.520 222.770 ;
        RECT 223.220 217.960 224.360 222.770 ;
        RECT 221.380 208.780 224.360 217.960 ;
        RECT 225.060 211.500 226.200 222.770 ;
        RECT 226.900 211.500 228.040 222.770 ;
        RECT 225.060 208.780 228.040 211.500 ;
        RECT 221.380 206.060 228.040 208.780 ;
        RECT 228.740 211.160 229.880 222.770 ;
        RECT 230.580 211.160 231.720 222.770 ;
        RECT 228.740 206.060 231.720 211.160 ;
        RECT 221.380 203.000 231.720 206.060 ;
        RECT 211.720 202.660 231.720 203.000 ;
        RECT 232.420 202.660 233.560 222.770 ;
        RECT 211.720 202.320 233.560 202.660 ;
        RECT 234.260 202.320 234.500 222.770 ;
        RECT 211.720 193.480 234.500 202.320 ;
        RECT 185.040 166.120 234.500 193.480 ;
        RECT 162.500 150.980 234.500 166.120 ;
        RECT 1.020 44.860 234.500 150.980 ;
        RECT 1.020 42.480 83.140 44.860 ;
        RECT 1.020 31.600 77.620 42.480 ;
        RECT 1.020 28.880 45.880 31.600 ;
        RECT 1.020 28.540 13.680 28.880 ;
        RECT 1.020 17.660 11.840 28.540 ;
        RECT 1.020 10.520 6.320 17.660 ;
        RECT 1.500 9.840 6.320 10.520 ;
        RECT 1.500 6.780 4.480 9.840 ;
        RECT 1.500 0.270 2.640 6.780 ;
        RECT 3.340 0.270 4.480 6.780 ;
        RECT 5.180 0.270 6.320 9.840 ;
        RECT 7.020 8.170 11.840 17.660 ;
        RECT 7.020 6.130 10.000 8.170 ;
        RECT 7.020 0.270 8.160 6.130 ;
        RECT 8.860 0.270 10.000 6.130 ;
        RECT 10.700 0.270 11.840 8.170 ;
        RECT 12.540 0.270 13.680 28.540 ;
        RECT 14.380 20.720 45.880 28.880 ;
        RECT 14.380 14.940 28.860 20.720 ;
        RECT 14.380 5.450 17.360 14.940 ;
        RECT 14.380 0.270 15.520 5.450 ;
        RECT 16.220 0.270 17.360 5.450 ;
        RECT 18.060 12.220 28.860 14.940 ;
        RECT 18.060 7.460 23.340 12.220 ;
        RECT 18.060 4.400 21.040 7.460 ;
        RECT 18.060 0.270 19.200 4.400 ;
        RECT 19.900 0.270 21.040 4.400 ;
        RECT 21.740 0.270 23.340 7.460 ;
        RECT 24.040 7.490 28.860 12.220 ;
        RECT 24.040 4.060 27.020 7.490 ;
        RECT 24.040 0.270 25.180 4.060 ;
        RECT 25.880 0.270 27.020 4.060 ;
        RECT 27.720 0.270 28.860 7.490 ;
        RECT 29.560 19.700 45.880 20.720 ;
        RECT 29.560 14.260 39.900 19.700 ;
        RECT 29.560 6.440 32.540 14.260 ;
        RECT 29.560 0.270 30.700 6.440 ;
        RECT 31.400 0.270 32.540 6.440 ;
        RECT 33.240 3.720 39.900 14.260 ;
        RECT 33.240 0.270 34.380 3.720 ;
        RECT 35.080 3.380 39.900 3.720 ;
        RECT 35.080 2.020 38.060 3.380 ;
        RECT 35.080 0.270 36.220 2.020 ;
        RECT 36.920 0.270 38.060 2.020 ;
        RECT 38.760 0.270 39.900 3.380 ;
        RECT 40.600 17.660 45.880 19.700 ;
        RECT 40.600 10.680 44.040 17.660 ;
        RECT 40.600 0.270 41.740 10.680 ;
        RECT 42.440 0.270 44.040 10.680 ;
        RECT 44.740 0.270 45.880 17.660 ;
        RECT 46.580 21.400 58.760 31.600 ;
        RECT 46.580 14.760 51.400 21.400 ;
        RECT 46.580 0.270 47.720 14.760 ;
        RECT 48.420 9.700 51.400 14.760 ;
        RECT 48.420 0.270 49.560 9.700 ;
        RECT 50.260 0.270 51.400 9.700 ;
        RECT 52.100 12.040 58.760 21.400 ;
        RECT 52.100 0.270 53.240 12.040 ;
        RECT 53.940 9.840 58.760 12.040 ;
        RECT 53.940 2.700 56.920 9.840 ;
        RECT 53.940 0.270 55.080 2.700 ;
        RECT 55.780 0.270 56.920 2.700 ;
        RECT 57.620 0.270 58.760 9.840 ;
        RECT 59.460 18.840 77.620 31.600 ;
        RECT 59.460 0.270 60.600 18.840 ;
        RECT 61.300 14.460 77.620 18.840 ;
        RECT 61.300 13.610 75.780 14.460 ;
        RECT 61.300 7.490 68.420 13.610 ;
        RECT 61.300 5.450 64.280 7.490 ;
        RECT 61.300 0.270 62.440 5.450 ;
        RECT 63.140 0.270 64.280 5.450 ;
        RECT 64.980 1.370 68.420 7.490 ;
        RECT 64.980 0.270 66.580 1.370 ;
        RECT 67.280 0.270 68.420 1.370 ;
        RECT 69.120 9.840 75.780 13.610 ;
        RECT 69.120 1.370 72.100 9.840 ;
        RECT 69.120 0.270 70.260 1.370 ;
        RECT 70.960 0.270 72.100 1.370 ;
        RECT 72.800 6.440 75.780 9.840 ;
        RECT 72.800 0.270 73.940 6.440 ;
        RECT 74.640 0.270 75.780 6.440 ;
        RECT 76.480 0.270 77.620 14.460 ;
        RECT 78.320 40.100 83.140 42.480 ;
        RECT 78.320 0.270 79.460 40.100 ;
        RECT 80.160 20.380 83.140 40.100 ;
        RECT 80.160 0.270 81.300 20.380 ;
        RECT 82.000 0.270 83.140 20.380 ;
        RECT 83.840 41.800 234.500 44.860 ;
        RECT 83.840 39.420 165.940 41.800 ;
        RECT 83.840 16.160 90.960 39.420 ;
        RECT 83.840 15.960 87.280 16.160 ;
        RECT 83.840 0.270 84.980 15.960 ;
        RECT 85.680 0.270 87.280 15.960 ;
        RECT 87.980 11.360 90.960 16.160 ;
        RECT 87.980 0.270 89.120 11.360 ;
        RECT 89.820 0.270 90.960 11.360 ;
        RECT 91.660 30.580 165.940 39.420 ;
        RECT 91.660 20.380 148.920 30.580 ;
        RECT 91.660 20.040 141.560 20.380 ;
        RECT 91.660 18.340 139.720 20.040 ;
        RECT 91.660 17.520 119.020 18.340 ;
        RECT 91.660 15.440 94.640 17.520 ;
        RECT 91.660 0.270 92.800 15.440 ;
        RECT 93.500 0.270 94.640 15.440 ;
        RECT 95.340 16.980 119.020 17.520 ;
        RECT 95.340 0.270 96.480 16.980 ;
        RECT 97.180 15.960 119.020 16.980 ;
        RECT 97.180 14.260 111.660 15.960 ;
        RECT 97.180 8.820 105.680 14.260 ;
        RECT 97.180 7.490 103.840 8.820 ;
        RECT 97.180 3.380 100.160 7.490 ;
        RECT 97.180 0.270 98.320 3.380 ;
        RECT 99.020 0.270 100.160 3.380 ;
        RECT 100.860 2.020 103.840 7.490 ;
        RECT 100.860 0.270 102.000 2.020 ;
        RECT 102.700 0.270 103.840 2.020 ;
        RECT 104.540 0.270 105.680 8.820 ;
        RECT 106.380 11.540 111.660 14.260 ;
        RECT 106.380 0.270 107.980 11.540 ;
        RECT 108.680 4.090 111.660 11.540 ;
        RECT 108.680 0.270 109.820 4.090 ;
        RECT 110.520 0.270 111.660 4.090 ;
        RECT 112.360 11.570 119.020 15.960 ;
        RECT 112.360 5.450 115.340 11.570 ;
        RECT 112.360 0.270 113.500 5.450 ;
        RECT 114.200 0.270 115.340 5.450 ;
        RECT 116.040 2.220 119.020 11.570 ;
        RECT 116.040 0.270 117.180 2.220 ;
        RECT 117.880 0.270 119.020 2.220 ;
        RECT 119.720 14.260 139.720 18.340 ;
        RECT 119.720 6.780 132.360 14.260 ;
        RECT 119.720 0.270 120.860 6.780 ;
        RECT 121.560 6.300 132.360 6.780 ;
        RECT 121.560 0.270 122.700 6.300 ;
        RECT 123.400 3.380 132.360 6.300 ;
        RECT 123.400 3.040 128.220 3.380 ;
        RECT 123.400 0.270 124.540 3.040 ;
        RECT 125.240 1.370 128.220 3.040 ;
        RECT 125.240 0.270 126.380 1.370 ;
        RECT 127.080 0.270 128.220 1.370 ;
        RECT 128.920 2.020 132.360 3.380 ;
        RECT 128.920 0.270 130.520 2.020 ;
        RECT 131.220 0.270 132.360 2.020 ;
        RECT 133.060 14.150 139.720 14.260 ;
        RECT 133.060 8.820 137.880 14.150 ;
        RECT 133.060 0.270 134.200 8.820 ;
        RECT 134.900 2.360 137.880 8.820 ;
        RECT 134.900 0.270 136.040 2.360 ;
        RECT 136.740 0.270 137.880 2.360 ;
        RECT 138.580 0.270 139.720 14.150 ;
        RECT 140.420 0.270 141.560 20.040 ;
        RECT 142.260 14.150 148.920 20.380 ;
        RECT 142.260 7.490 145.240 14.150 ;
        RECT 142.260 0.270 143.400 7.490 ;
        RECT 144.100 0.270 145.240 7.490 ;
        RECT 145.940 4.740 148.920 14.150 ;
        RECT 145.940 0.270 147.080 4.740 ;
        RECT 147.780 0.270 148.920 4.740 ;
        RECT 149.620 28.540 165.940 30.580 ;
        RECT 149.620 0.270 151.220 28.540 ;
        RECT 151.920 27.860 165.940 28.540 ;
        RECT 151.920 25.140 162.260 27.860 ;
        RECT 151.920 7.490 160.420 25.140 ;
        RECT 151.920 6.130 158.580 7.490 ;
        RECT 151.920 1.370 154.900 6.130 ;
        RECT 151.920 0.270 153.060 1.370 ;
        RECT 153.760 0.270 154.900 1.370 ;
        RECT 155.600 4.400 158.580 6.130 ;
        RECT 155.600 0.270 156.740 4.400 ;
        RECT 157.440 0.270 158.580 4.400 ;
        RECT 159.280 0.270 160.420 7.490 ;
        RECT 161.120 0.270 162.260 25.140 ;
        RECT 162.960 4.090 165.940 27.860 ;
        RECT 162.960 0.270 164.100 4.090 ;
        RECT 164.800 0.270 165.940 4.090 ;
        RECT 166.640 26.160 234.500 41.800 ;
        RECT 166.640 20.720 207.340 26.160 ;
        RECT 166.640 17.690 199.980 20.720 ;
        RECT 166.640 13.400 177.440 17.690 ;
        RECT 166.640 9.320 173.760 13.400 ;
        RECT 166.640 3.720 171.920 9.320 ;
        RECT 166.640 0.270 167.780 3.720 ;
        RECT 168.480 1.370 171.920 3.720 ;
        RECT 168.480 0.270 169.620 1.370 ;
        RECT 170.320 0.270 171.920 1.370 ;
        RECT 172.620 0.270 173.760 9.320 ;
        RECT 174.460 6.100 177.440 13.400 ;
        RECT 174.460 0.270 175.600 6.100 ;
        RECT 176.300 0.270 177.440 6.100 ;
        RECT 178.140 17.480 199.980 17.690 ;
        RECT 178.140 15.650 196.300 17.480 ;
        RECT 178.140 11.360 182.960 15.650 ;
        RECT 178.140 0.270 179.280 11.360 ;
        RECT 179.980 2.020 182.960 11.360 ;
        RECT 179.980 0.270 181.120 2.020 ;
        RECT 181.820 0.270 182.960 2.020 ;
        RECT 183.660 14.150 196.300 15.650 ;
        RECT 183.660 9.320 194.460 14.150 ;
        RECT 183.660 4.090 186.640 9.320 ;
        RECT 183.660 0.270 184.800 4.090 ;
        RECT 185.500 0.270 186.640 4.090 ;
        RECT 187.340 3.380 194.460 9.320 ;
        RECT 187.340 0.270 188.480 3.380 ;
        RECT 189.180 1.370 194.460 3.380 ;
        RECT 189.180 0.270 190.320 1.370 ;
        RECT 191.020 0.270 192.160 1.370 ;
        RECT 192.860 0.270 194.460 1.370 ;
        RECT 195.160 0.270 196.300 14.150 ;
        RECT 197.000 6.780 199.980 17.480 ;
        RECT 197.000 0.270 198.140 6.780 ;
        RECT 198.840 0.270 199.980 6.780 ;
        RECT 200.680 7.490 207.340 20.720 ;
        RECT 200.680 1.680 203.660 7.490 ;
        RECT 200.680 0.270 201.820 1.680 ;
        RECT 202.520 0.270 203.660 1.680 ;
        RECT 204.360 1.370 207.340 7.490 ;
        RECT 204.360 0.270 205.500 1.370 ;
        RECT 206.200 0.270 207.340 1.370 ;
        RECT 208.040 18.840 234.500 26.160 ;
        RECT 208.040 15.960 222.520 18.840 ;
        RECT 208.040 0.270 209.180 15.960 ;
        RECT 209.880 12.220 222.520 15.960 ;
        RECT 209.880 6.980 218.840 12.220 ;
        RECT 209.880 0.270 211.020 6.980 ;
        RECT 211.720 6.780 218.840 6.980 ;
        RECT 211.720 4.400 217.000 6.780 ;
        RECT 211.720 2.700 215.160 4.400 ;
        RECT 211.720 0.270 212.860 2.700 ;
        RECT 213.560 0.270 215.160 2.700 ;
        RECT 215.860 0.270 217.000 4.400 ;
        RECT 217.700 0.270 218.840 6.780 ;
        RECT 219.540 5.080 222.520 12.220 ;
        RECT 219.540 0.270 220.680 5.080 ;
        RECT 221.380 0.270 222.520 5.080 ;
        RECT 223.220 18.680 234.500 18.840 ;
        RECT 223.220 16.120 231.720 18.680 ;
        RECT 223.220 15.960 229.880 16.120 ;
        RECT 223.220 0.270 224.360 15.960 ;
        RECT 225.060 15.440 229.880 15.960 ;
        RECT 225.060 14.760 228.040 15.440 ;
        RECT 225.060 0.270 226.200 14.760 ;
        RECT 226.900 0.270 228.040 14.760 ;
        RECT 228.740 0.270 229.880 15.440 ;
        RECT 230.580 0.270 231.720 16.120 ;
        RECT 232.420 14.080 234.500 18.680 ;
        RECT 232.420 0.270 233.560 14.080 ;
        RECT 234.260 0.270 234.500 14.080 ;
      LAYER met3 ;
        RECT 14.750 221.470 213.870 222.185 ;
        RECT 3.285 220.530 234.750 221.470 ;
        RECT 6.930 219.430 218.930 220.530 ;
        RECT 3.285 219.170 234.750 219.430 ;
        RECT 7.850 218.070 215.710 219.170 ;
        RECT 3.285 217.130 234.750 218.070 ;
        RECT 16.590 216.030 215.250 217.130 ;
        RECT 3.285 215.770 234.750 216.030 ;
        RECT 19.350 214.670 218.470 215.770 ;
        RECT 3.285 213.730 234.750 214.670 ;
        RECT 7.390 212.630 218.470 213.730 ;
        RECT 3.285 212.370 234.750 212.630 ;
        RECT 37.750 211.270 222.150 212.370 ;
        RECT 3.285 210.330 234.750 211.270 ;
        RECT 20.730 209.230 220.310 210.330 ;
        RECT 3.285 208.290 234.750 209.230 ;
        RECT 19.350 207.190 218.470 208.290 ;
        RECT 3.285 206.930 234.750 207.190 ;
        RECT 27.170 205.830 223.990 206.930 ;
        RECT 3.285 204.890 234.750 205.830 ;
        RECT 20.730 203.790 221.690 204.890 ;
        RECT 3.285 203.530 234.750 203.790 ;
        RECT 17.050 202.430 226.290 203.530 ;
        RECT 3.285 201.490 234.750 202.430 ;
        RECT 21.480 200.390 220.310 201.490 ;
        RECT 3.285 200.130 234.750 200.390 ;
        RECT 28.550 199.030 222.150 200.130 ;
        RECT 3.285 198.090 234.750 199.030 ;
        RECT 18.430 196.990 225.370 198.090 ;
        RECT 3.285 196.730 234.750 196.990 ;
        RECT 34.990 195.630 221.690 196.730 ;
        RECT 3.285 194.690 234.750 195.630 ;
        RECT 10.150 193.590 222.150 194.690 ;
        RECT 3.285 192.650 234.750 193.590 ;
        RECT 7.850 191.550 227.210 192.650 ;
        RECT 3.285 191.290 234.750 191.550 ;
        RECT 7.390 190.190 225.370 191.290 ;
        RECT 3.285 189.250 234.750 190.190 ;
        RECT 7.390 188.150 221.690 189.250 ;
        RECT 3.285 187.890 234.750 188.150 ;
        RECT 20.270 186.790 224.910 187.890 ;
        RECT 3.285 185.850 234.750 186.790 ;
        RECT 20.730 184.750 224.910 185.850 ;
        RECT 3.285 184.490 234.750 184.750 ;
        RECT 7.850 183.390 219.850 184.490 ;
        RECT 3.285 182.450 234.750 183.390 ;
        RECT 20.730 181.350 219.390 182.450 ;
        RECT 3.285 180.410 234.750 181.350 ;
        RECT 19.350 179.310 220.310 180.410 ;
        RECT 3.285 179.050 234.750 179.310 ;
        RECT 6.930 177.950 227.210 179.050 ;
        RECT 3.285 177.010 234.750 177.950 ;
        RECT 7.850 175.910 218.010 177.010 ;
        RECT 3.285 175.650 234.750 175.910 ;
        RECT 7.850 174.550 222.150 175.650 ;
        RECT 3.285 173.610 234.750 174.550 ;
        RECT 7.390 172.510 214.790 173.610 ;
        RECT 3.285 172.250 234.750 172.510 ;
        RECT 19.350 171.150 218.470 172.250 ;
        RECT 3.285 170.210 234.750 171.150 ;
        RECT 15.210 169.110 221.230 170.210 ;
        RECT 3.285 168.850 234.750 169.110 ;
        RECT 14.290 167.750 227.210 168.850 ;
        RECT 3.285 166.810 234.750 167.750 ;
        RECT 14.750 165.710 224.910 166.810 ;
        RECT 3.285 164.770 234.750 165.710 ;
        RECT 19.810 163.670 224.910 164.770 ;
        RECT 3.285 163.410 234.750 163.670 ;
        RECT 4.170 162.310 220.310 163.410 ;
        RECT 3.285 161.370 234.750 162.310 ;
        RECT 18.430 160.270 219.850 161.370 ;
        RECT 3.285 160.010 234.750 160.270 ;
        RECT 20.730 158.910 218.470 160.010 ;
        RECT 3.285 157.970 234.750 158.910 ;
        RECT 19.350 156.870 228.070 157.970 ;
        RECT 3.285 156.610 234.750 156.870 ;
        RECT 20.270 155.510 224.390 156.610 ;
        RECT 3.285 154.570 234.750 155.510 ;
        RECT 18.430 153.470 223.530 154.570 ;
        RECT 3.285 152.530 234.750 153.470 ;
        RECT 19.350 151.430 219.390 152.530 ;
        RECT 3.285 151.170 234.750 151.430 ;
        RECT 20.730 150.070 225.370 151.170 ;
        RECT 3.285 149.130 234.750 150.070 ;
        RECT 7.390 148.030 220.310 149.130 ;
        RECT 3.285 147.770 234.750 148.030 ;
        RECT 7.850 146.670 224.910 147.770 ;
        RECT 3.285 145.730 234.750 146.670 ;
        RECT 14.350 144.630 219.390 145.730 ;
        RECT 3.285 144.370 234.750 144.630 ;
        RECT 20.730 143.270 218.930 144.370 ;
        RECT 3.285 142.330 234.750 143.270 ;
        RECT 14.290 141.230 217.550 142.330 ;
        RECT 3.285 140.970 234.750 141.230 ;
        RECT 21.650 139.870 214.330 140.970 ;
        RECT 3.285 138.930 234.750 139.870 ;
        RECT 20.270 137.830 220.310 138.930 ;
        RECT 3.285 136.890 234.750 137.830 ;
        RECT 6.530 135.790 217.090 136.890 ;
        RECT 3.285 135.530 234.750 135.790 ;
        RECT 43.270 134.430 216.170 135.530 ;
        RECT 3.285 133.490 234.750 134.430 ;
        RECT 21.020 132.390 212.030 133.490 ;
        RECT 3.285 132.130 234.750 132.390 ;
        RECT 16.590 131.030 219.850 132.130 ;
        RECT 3.285 130.090 234.750 131.030 ;
        RECT 19.350 128.990 211.110 130.090 ;
        RECT 3.285 128.730 234.750 128.990 ;
        RECT 18.890 127.630 224.910 128.730 ;
        RECT 3.285 126.690 234.750 127.630 ;
        RECT 20.270 125.590 211.740 126.690 ;
        RECT 3.285 124.650 234.750 125.590 ;
        RECT 13.370 123.550 207.430 124.650 ;
        RECT 3.285 123.290 234.750 123.550 ;
        RECT 14.290 122.190 224.450 123.290 ;
        RECT 3.285 121.250 234.750 122.190 ;
        RECT 19.350 120.150 233.590 121.250 ;
        RECT 3.285 119.890 234.750 120.150 ;
        RECT 20.270 118.790 216.170 119.890 ;
        RECT 3.285 117.850 234.750 118.790 ;
        RECT 14.750 116.750 222.150 117.850 ;
        RECT 3.285 116.490 234.750 116.750 ;
        RECT 9.690 115.390 225.370 116.490 ;
        RECT 3.285 114.450 234.750 115.390 ;
        RECT 17.970 113.350 217.090 114.450 ;
        RECT 3.285 113.090 234.750 113.350 ;
        RECT 7.390 111.990 213.580 113.090 ;
        RECT 3.285 111.050 234.750 111.990 ;
        RECT 9.230 109.950 217.090 111.050 ;
        RECT 3.285 109.010 234.750 109.950 ;
        RECT 16.590 107.910 216.170 109.010 ;
        RECT 3.285 107.650 234.750 107.910 ;
        RECT 14.290 106.550 212.490 107.650 ;
        RECT 3.285 105.610 234.750 106.550 ;
        RECT 8.310 104.510 232.270 105.610 ;
        RECT 3.285 104.250 234.750 104.510 ;
        RECT 9.290 103.150 219.390 104.250 ;
        RECT 3.285 102.210 234.750 103.150 ;
        RECT 20.730 101.110 219.850 102.210 ;
        RECT 3.285 100.850 234.750 101.110 ;
        RECT 20.270 99.750 216.630 100.850 ;
        RECT 3.285 98.810 234.750 99.750 ;
        RECT 18.890 97.710 220.310 98.810 ;
        RECT 3.285 96.770 234.750 97.710 ;
        RECT 20.270 95.670 215.250 96.770 ;
        RECT 3.285 95.410 234.750 95.670 ;
        RECT 18.430 94.310 219.390 95.410 ;
        RECT 3.285 93.370 234.750 94.310 ;
        RECT 17.510 92.270 218.010 93.370 ;
        RECT 3.285 92.010 234.750 92.270 ;
        RECT 20.730 90.910 218.930 92.010 ;
        RECT 3.285 89.970 234.750 90.910 ;
        RECT 7.850 88.870 217.090 89.970 ;
        RECT 3.285 88.610 234.750 88.870 ;
        RECT 9.230 87.510 219.850 88.610 ;
        RECT 3.285 86.570 234.750 87.510 ;
        RECT 19.810 85.470 225.370 86.570 ;
        RECT 3.285 85.210 234.750 85.470 ;
        RECT 9.230 84.110 222.150 85.210 ;
        RECT 3.285 83.170 234.750 84.110 ;
        RECT 20.730 82.070 233.590 83.170 ;
        RECT 3.285 81.130 234.750 82.070 ;
        RECT 7.390 80.030 212.950 81.130 ;
        RECT 3.285 79.770 234.750 80.030 ;
        RECT 20.730 78.670 214.330 79.770 ;
        RECT 3.285 77.730 234.750 78.670 ;
        RECT 14.750 76.630 233.590 77.730 ;
        RECT 3.285 76.370 234.750 76.630 ;
        RECT 11.530 75.270 217.550 76.370 ;
        RECT 3.285 74.330 234.750 75.270 ;
        RECT 17.970 73.230 219.850 74.330 ;
        RECT 3.285 72.970 234.750 73.230 ;
        RECT 14.290 71.870 210.190 72.970 ;
        RECT 3.285 70.930 234.750 71.870 ;
        RECT 17.510 69.830 233.590 70.930 ;
        RECT 3.285 68.890 234.750 69.830 ;
        RECT 14.290 67.790 209.270 68.890 ;
        RECT 3.285 67.530 234.750 67.790 ;
        RECT 10.150 66.430 183.050 67.530 ;
        RECT 3.285 65.490 234.750 66.430 ;
        RECT 10.150 64.390 220.310 65.490 ;
        RECT 3.285 64.130 234.750 64.390 ;
        RECT 10.150 63.030 214.790 64.130 ;
        RECT 3.285 62.090 234.750 63.030 ;
        RECT 20.270 60.990 187.190 62.090 ;
        RECT 3.285 60.730 234.750 60.990 ;
        RECT 14.290 59.630 215.250 60.730 ;
        RECT 3.285 58.690 234.750 59.630 ;
        RECT 20.270 57.590 233.590 58.690 ;
        RECT 3.285 57.330 234.750 57.590 ;
        RECT 14.290 56.230 215.710 57.330 ;
        RECT 3.285 55.290 234.750 56.230 ;
        RECT 10.150 54.190 220.310 55.290 ;
        RECT 3.285 53.250 234.750 54.190 ;
        RECT 10.610 52.150 233.590 53.250 ;
        RECT 3.285 51.890 234.750 52.150 ;
        RECT 18.430 50.790 233.590 51.890 ;
        RECT 3.285 49.850 234.750 50.790 ;
        RECT 16.130 48.750 220.310 49.850 ;
        RECT 3.285 48.490 234.750 48.750 ;
        RECT 19.350 47.390 233.590 48.490 ;
        RECT 3.285 46.450 234.750 47.390 ;
        RECT 20.730 45.350 228.990 46.450 ;
        RECT 3.285 45.090 234.750 45.350 ;
        RECT 18.890 43.990 233.590 45.090 ;
        RECT 3.285 43.050 234.750 43.990 ;
        RECT 14.350 41.950 217.090 43.050 ;
        RECT 3.285 41.010 234.750 41.950 ;
        RECT 20.730 39.910 211.570 41.010 ;
        RECT 3.285 39.650 234.750 39.910 ;
        RECT 20.270 38.550 219.850 39.650 ;
        RECT 3.285 37.610 234.750 38.550 ;
        RECT 20.270 36.510 215.250 37.610 ;
        RECT 3.285 36.250 234.750 36.510 ;
        RECT 19.810 35.150 212.490 36.250 ;
        RECT 3.285 34.210 234.750 35.150 ;
        RECT 29.930 33.110 182.130 34.210 ;
        RECT 3.285 32.850 234.750 33.110 ;
        RECT 20.730 31.750 220.310 32.850 ;
        RECT 3.285 30.810 234.750 31.750 ;
        RECT 14.350 29.710 184.430 30.810 ;
        RECT 3.285 29.450 234.750 29.710 ;
        RECT 23.490 28.350 226.750 29.450 ;
        RECT 3.285 27.410 234.750 28.350 ;
        RECT 24.870 26.310 222.150 27.410 ;
        RECT 3.285 25.370 234.750 26.310 ;
        RECT 3.710 24.270 220.310 25.370 ;
        RECT 3.285 24.010 234.750 24.270 ;
        RECT 11.990 22.910 220.310 24.010 ;
        RECT 3.285 21.970 234.750 22.910 ;
        RECT 17.970 20.870 220.310 21.970 ;
        RECT 3.285 20.610 234.750 20.870 ;
        RECT 16.130 19.510 224.450 20.610 ;
        RECT 3.285 18.570 234.750 19.510 ;
        RECT 10.150 17.470 216.170 18.570 ;
        RECT 3.285 17.210 234.750 17.470 ;
        RECT 20.730 16.110 229.510 17.210 ;
        RECT 3.285 15.170 234.750 16.110 ;
        RECT 14.750 14.070 227.210 15.170 ;
        RECT 3.285 13.130 234.750 14.070 ;
        RECT 4.630 12.030 214.790 13.130 ;
        RECT 3.285 11.770 234.750 12.030 ;
        RECT 8.310 10.670 214.790 11.770 ;
        RECT 3.285 9.730 234.750 10.670 ;
        RECT 20.730 8.630 213.870 9.730 ;
        RECT 3.285 8.370 234.750 8.630 ;
        RECT 7.850 7.270 215.710 8.370 ;
        RECT 3.285 6.330 234.750 7.270 ;
        RECT 5.550 5.230 213.870 6.330 ;
        RECT 3.285 4.970 234.750 5.230 ;
        RECT 7.390 3.870 197.770 4.970 ;
        RECT 3.285 2.930 234.750 3.870 ;
        RECT 15.670 1.830 219.390 2.930 ;
        RECT 3.285 1.570 234.750 1.830 ;
        RECT 15.210 0.855 222.150 1.570 ;
      LAYER met4 ;
        RECT 10.415 4.800 20.640 216.745 ;
        RECT 23.040 4.800 97.440 216.745 ;
        RECT 99.840 4.800 174.240 216.745 ;
        RECT 176.640 4.800 224.185 216.745 ;
        RECT 10.415 3.575 224.185 4.800 ;
  END
END RegFile
MACRO S_term_DSP
  CLASS BLOCK ;
  FOREIGN S_term_DSP ;
  ORIGIN 0.000 0.000 ;
  SIZE 223.275 BY 40.000 ;
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.680 0.000 5.820 6.160 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.000 0.000 117.140 6.500 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.040 0.000 128.180 6.500 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.540 0.000 139.680 6.500 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.580 0.000 150.720 6.500 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.620 0.000 161.760 6.500 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.660 0.000 172.800 6.500 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.160 0.000 184.300 6.500 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.200 0.000 195.340 6.500 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.240 0.000 206.380 6.500 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.280 0.000 217.420 6.500 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.720 0.000 16.860 6.160 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.760 0.000 27.900 6.500 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.800 0.000 38.940 6.500 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.300 0.000 50.440 6.500 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.340 0.000 61.480 6.700 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.380 0.000 72.520 6.500 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.420 0.000 83.560 6.500 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.920 0.000 95.060 6.500 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.960 0.000 106.100 6.500 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.380 29.540 187.520 40.000 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.320 32.260 205.460 40.000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.160 29.540 207.300 40.000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.000 32.260 209.140 40.000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.840 29.540 210.980 40.000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.680 26.820 212.820 40.000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.520 31.920 214.660 40.000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.360 23.760 216.500 40.000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.200 26.480 218.340 40.000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.040 29.200 220.180 40.000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.880 20.700 222.020 40.000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.220 32.260 189.360 40.000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.060 29.200 191.200 40.000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.900 26.820 193.040 40.000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.740 29.540 194.880 40.000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.580 26.820 196.720 40.000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.420 26.820 198.560 40.000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.260 26.480 200.400 40.000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.100 24.100 202.240 40.000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.480 30.870 203.620 40.000 ;
    END
  END FrameStrobe_O[9]
  PIN N1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.620 32.260 0.760 40.000 ;
    END
  END N1BEG[0]
  PIN N1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.000 29.540 2.140 40.000 ;
    END
  END N1BEG[1]
  PIN N1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.840 31.920 3.980 40.000 ;
    END
  END N1BEG[2]
  PIN N1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.680 31.240 5.820 40.000 ;
    END
  END N1BEG[3]
  PIN N2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.520 33.590 7.660 40.000 ;
    END
  END N2BEG[0]
  PIN N2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.360 26.820 9.500 40.000 ;
    END
  END N2BEG[1]
  PIN N2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.200 39.030 11.340 40.000 ;
    END
  END N2BEG[2]
  PIN N2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.040 32.260 13.180 40.000 ;
    END
  END N2BEG[3]
  PIN N2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.880 29.200 15.020 40.000 ;
    END
  END N2BEG[4]
  PIN N2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.720 31.920 16.860 40.000 ;
    END
  END N2BEG[5]
  PIN N2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.560 29.540 18.700 40.000 ;
    END
  END N2BEG[6]
  PIN N2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.400 32.260 20.540 40.000 ;
    END
  END N2BEG[7]
  PIN N2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.780 29.200 21.920 40.000 ;
    END
  END N2BEGb[0]
  PIN N2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.620 30.560 23.760 40.000 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.460 29.540 25.600 40.000 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.300 31.240 27.440 40.000 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.140 29.200 29.280 40.000 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.980 32.260 31.120 40.000 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.820 29.540 32.960 40.000 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.660 26.820 34.800 40.000 ;
    END
  END N2BEGb[7]
  PIN N4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.500 31.580 36.640 40.000 ;
    END
  END N4BEG[0]
  PIN N4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.440 32.260 54.580 40.000 ;
    END
  END N4BEG[10]
  PIN N4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.280 39.030 56.420 40.000 ;
    END
  END N4BEG[11]
  PIN N4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.120 34.950 58.260 40.000 ;
    END
  END N4BEG[12]
  PIN N4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.960 29.540 60.100 40.000 ;
    END
  END N4BEG[13]
  PIN N4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.340 31.920 61.480 40.000 ;
    END
  END N4BEG[14]
  PIN N4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.180 29.340 63.320 40.000 ;
    END
  END N4BEG[15]
  PIN N4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.340 26.820 38.480 40.000 ;
    END
  END N4BEG[1]
  PIN N4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.180 33.590 40.320 40.000 ;
    END
  END N4BEG[2]
  PIN N4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.560 32.260 41.700 40.000 ;
    END
  END N4BEG[3]
  PIN N4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.400 26.820 43.540 40.000 ;
    END
  END N4BEG[4]
  PIN N4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.240 29.200 45.380 40.000 ;
    END
  END N4BEG[5]
  PIN N4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.080 26.820 47.220 40.000 ;
    END
  END N4BEG[6]
  PIN N4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.920 29.540 49.060 40.000 ;
    END
  END N4BEG[7]
  PIN N4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.760 26.820 50.900 40.000 ;
    END
  END N4BEG[8]
  PIN N4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.600 24.100 52.740 40.000 ;
    END
  END N4BEG[9]
  PIN NN4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.020 31.240 65.160 40.000 ;
    END
  END NN4BEG[0]
  PIN NN4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.960 32.260 83.100 40.000 ;
    END
  END NN4BEG[10]
  PIN NN4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.800 32.260 84.940 40.000 ;
    END
  END NN4BEG[11]
  PIN NN4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.640 31.240 86.780 40.000 ;
    END
  END NN4BEG[12]
  PIN NN4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.480 29.540 88.620 40.000 ;
    END
  END NN4BEG[13]
  PIN NN4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.320 26.820 90.460 40.000 ;
    END
  END NN4BEG[14]
  PIN NN4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.160 29.540 92.300 40.000 ;
    END
  END NN4BEG[15]
  PIN NN4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.860 29.340 67.000 40.000 ;
    END
  END NN4BEG[1]
  PIN NN4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.700 31.920 68.840 40.000 ;
    END
  END NN4BEG[2]
  PIN NN4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.540 29.200 70.680 40.000 ;
    END
  END NN4BEG[3]
  PIN NN4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.380 31.240 72.520 40.000 ;
    END
  END NN4BEG[4]
  PIN NN4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.220 29.540 74.360 40.000 ;
    END
  END NN4BEG[5]
  PIN NN4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.060 39.030 76.200 40.000 ;
    END
  END NN4BEG[6]
  PIN NN4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.900 26.820 78.040 40.000 ;
    END
  END NN4BEG[7]
  PIN NN4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.740 23.080 79.880 40.000 ;
    END
  END NN4BEG[8]
  PIN NN4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.580 26.480 81.720 40.000 ;
    END
  END NN4BEG[9]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.000 20.700 94.140 40.000 ;
    END
  END S1END[0]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.840 23.080 95.980 40.000 ;
    END
  END S1END[1]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.680 21.040 97.820 40.000 ;
    END
  END S1END[2]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.520 31.240 99.660 40.000 ;
    END
  END S1END[3]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.360 30.870 101.500 40.000 ;
    END
  END S2END[0]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.740 17.640 102.880 40.000 ;
    END
  END S2END[1]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.580 20.700 104.720 40.000 ;
    END
  END S2END[2]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.420 38.350 106.560 40.000 ;
    END
  END S2END[3]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.260 39.030 108.400 40.000 ;
    END
  END S2END[4]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.100 22.880 110.240 40.000 ;
    END
  END S2END[5]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.940 39.030 112.080 40.000 ;
    END
  END S2END[6]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.780 39.030 113.920 40.000 ;
    END
  END S2END[7]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.620 32.230 115.760 40.000 ;
    END
  END S2MID[0]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.460 20.020 117.600 40.000 ;
    END
  END S2MID[1]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.300 22.740 119.440 40.000 ;
    END
  END S2MID[2]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.140 20.360 121.280 40.000 ;
    END
  END S2MID[3]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.520 22.400 122.660 40.000 ;
    END
  END S2MID[4]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.360 20.360 124.500 40.000 ;
    END
  END S2MID[5]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.200 26.820 126.340 40.000 ;
    END
  END S2MID[6]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.040 36.340 128.180 40.000 ;
    END
  END S2MID[7]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.880 31.550 130.020 40.000 ;
    END
  END S4END[0]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.820 33.590 147.960 40.000 ;
    END
  END S4END[10]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.660 26.140 149.800 40.000 ;
    END
  END S4END[11]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.500 28.830 151.640 40.000 ;
    END
  END S4END[12]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.340 32.230 153.480 40.000 ;
    END
  END S4END[13]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.180 23.080 155.320 40.000 ;
    END
  END S4END[14]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.020 26.140 157.160 40.000 ;
    END
  END S4END[15]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.720 34.980 131.860 40.000 ;
    END
  END S4END[1]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.560 25.800 133.700 40.000 ;
    END
  END S4END[2]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.400 26.820 135.540 40.000 ;
    END
  END S4END[3]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.240 20.020 137.380 40.000 ;
    END
  END S4END[4]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.080 31.550 139.220 40.000 ;
    END
  END S4END[5]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.920 17.640 141.060 40.000 ;
    END
  END S4END[6]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.300 20.360 142.440 40.000 ;
    END
  END S4END[7]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.140 28.830 144.280 40.000 ;
    END
  END S4END[8]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.980 33.620 146.120 40.000 ;
    END
  END S4END[9]
  PIN SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.860 28.520 159.000 40.000 ;
    END
  END SS4END[0]
  PIN SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.800 31.920 176.940 40.000 ;
    END
  END SS4END[10]
  PIN SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.640 28.520 178.780 40.000 ;
    END
  END SS4END[11]
  PIN SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.480 28.320 180.620 40.000 ;
    END
  END SS4END[12]
  PIN SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.320 31.920 182.460 40.000 ;
    END
  END SS4END[13]
  PIN SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.700 28.180 183.840 40.000 ;
    END
  END SS4END[14]
  PIN SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.540 31.580 185.680 40.000 ;
    END
  END SS4END[15]
  PIN SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.700 25.800 160.840 40.000 ;
    END
  END SS4END[1]
  PIN SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.540 28.860 162.680 40.000 ;
    END
  END SS4END[2]
  PIN SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.920 25.940 164.060 40.000 ;
    END
  END SS4END[3]
  PIN SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.760 25.800 165.900 40.000 ;
    END
  END SS4END[4]
  PIN SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.600 31.580 167.740 40.000 ;
    END
  END SS4END[5]
  PIN SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.440 31.580 169.580 40.000 ;
    END
  END SS4END[6]
  PIN SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.280 28.860 171.420 40.000 ;
    END
  END SS4END[7]
  PIN SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.120 26.140 173.260 40.000 ;
    END
  END SS4END[8]
  PIN SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.960 26.140 175.100 40.000 ;
    END
  END SS4END[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 40.090 5.200 41.690 32.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 110.835 5.200 112.435 32.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 181.580 5.200 183.180 32.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 75.465 5.200 77.065 32.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 146.210 5.200 147.810 32.880 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 217.580 39.355 ;
      LAYER met1 ;
        RECT 0.530 4.120 222.110 39.400 ;
      LAYER met2 ;
        RECT 1.040 31.980 1.720 39.850 ;
        RECT 0.560 29.260 1.720 31.980 ;
        RECT 2.420 31.640 3.560 39.850 ;
        RECT 4.260 31.640 5.400 39.850 ;
        RECT 2.420 30.960 5.400 31.640 ;
        RECT 6.100 33.310 7.240 39.850 ;
        RECT 7.940 33.310 9.080 39.850 ;
        RECT 6.100 30.960 9.080 33.310 ;
        RECT 2.420 29.260 9.080 30.960 ;
        RECT 0.560 26.540 9.080 29.260 ;
        RECT 9.780 38.750 10.920 39.850 ;
        RECT 11.620 38.750 12.760 39.850 ;
        RECT 9.780 31.980 12.760 38.750 ;
        RECT 13.460 31.980 14.600 39.850 ;
        RECT 9.780 28.920 14.600 31.980 ;
        RECT 15.300 31.640 16.440 39.850 ;
        RECT 17.140 31.640 18.280 39.850 ;
        RECT 15.300 29.260 18.280 31.640 ;
        RECT 18.980 31.980 20.120 39.850 ;
        RECT 20.820 31.980 21.500 39.850 ;
        RECT 18.980 29.260 21.500 31.980 ;
        RECT 15.300 28.920 21.500 29.260 ;
        RECT 22.200 30.280 23.340 39.850 ;
        RECT 24.040 30.280 25.180 39.850 ;
        RECT 22.200 29.260 25.180 30.280 ;
        RECT 25.880 30.960 27.020 39.850 ;
        RECT 27.720 30.960 28.860 39.850 ;
        RECT 25.880 29.260 28.860 30.960 ;
        RECT 22.200 28.920 28.860 29.260 ;
        RECT 29.560 31.980 30.700 39.850 ;
        RECT 31.400 31.980 32.540 39.850 ;
        RECT 29.560 29.260 32.540 31.980 ;
        RECT 33.240 29.260 34.380 39.850 ;
        RECT 29.560 28.920 34.380 29.260 ;
        RECT 9.780 26.540 34.380 28.920 ;
        RECT 35.080 31.300 36.220 39.850 ;
        RECT 36.920 31.300 38.060 39.850 ;
        RECT 35.080 26.540 38.060 31.300 ;
        RECT 38.760 33.310 39.900 39.850 ;
        RECT 40.600 33.310 41.280 39.850 ;
        RECT 38.760 31.980 41.280 33.310 ;
        RECT 41.980 31.980 43.120 39.850 ;
        RECT 38.760 26.540 43.120 31.980 ;
        RECT 43.820 28.920 44.960 39.850 ;
        RECT 45.660 28.920 46.800 39.850 ;
        RECT 43.820 26.540 46.800 28.920 ;
        RECT 47.500 29.260 48.640 39.850 ;
        RECT 49.340 29.260 50.480 39.850 ;
        RECT 47.500 26.540 50.480 29.260 ;
        RECT 51.180 26.540 52.320 39.850 ;
        RECT 0.560 23.820 52.320 26.540 ;
        RECT 53.020 31.980 54.160 39.850 ;
        RECT 54.860 38.750 56.000 39.850 ;
        RECT 56.700 38.750 57.840 39.850 ;
        RECT 54.860 34.670 57.840 38.750 ;
        RECT 58.540 34.670 59.680 39.850 ;
        RECT 54.860 31.980 59.680 34.670 ;
        RECT 53.020 29.260 59.680 31.980 ;
        RECT 60.380 31.640 61.060 39.850 ;
        RECT 61.760 31.640 62.900 39.850 ;
        RECT 60.380 29.260 62.900 31.640 ;
        RECT 53.020 29.060 62.900 29.260 ;
        RECT 63.600 30.960 64.740 39.850 ;
        RECT 65.440 30.960 66.580 39.850 ;
        RECT 63.600 29.060 66.580 30.960 ;
        RECT 67.280 31.640 68.420 39.850 ;
        RECT 69.120 31.640 70.260 39.850 ;
        RECT 67.280 29.060 70.260 31.640 ;
        RECT 53.020 28.920 70.260 29.060 ;
        RECT 70.960 30.960 72.100 39.850 ;
        RECT 72.800 30.960 73.940 39.850 ;
        RECT 70.960 29.260 73.940 30.960 ;
        RECT 74.640 38.750 75.780 39.850 ;
        RECT 76.480 38.750 77.620 39.850 ;
        RECT 74.640 29.260 77.620 38.750 ;
        RECT 70.960 28.920 77.620 29.260 ;
        RECT 53.020 26.540 77.620 28.920 ;
        RECT 78.320 26.540 79.460 39.850 ;
        RECT 53.020 23.820 79.460 26.540 ;
        RECT 0.560 22.800 79.460 23.820 ;
        RECT 80.160 26.200 81.300 39.850 ;
        RECT 82.000 31.980 82.680 39.850 ;
        RECT 83.380 31.980 84.520 39.850 ;
        RECT 85.220 31.980 86.360 39.850 ;
        RECT 82.000 30.960 86.360 31.980 ;
        RECT 87.060 30.960 88.200 39.850 ;
        RECT 82.000 29.260 88.200 30.960 ;
        RECT 88.900 29.260 90.040 39.850 ;
        RECT 82.000 26.540 90.040 29.260 ;
        RECT 90.740 29.260 91.880 39.850 ;
        RECT 92.580 29.260 93.720 39.850 ;
        RECT 90.740 26.540 93.720 29.260 ;
        RECT 82.000 26.200 93.720 26.540 ;
        RECT 80.160 22.800 93.720 26.200 ;
        RECT 0.560 20.420 93.720 22.800 ;
        RECT 94.420 22.800 95.560 39.850 ;
        RECT 96.260 22.800 97.400 39.850 ;
        RECT 94.420 20.760 97.400 22.800 ;
        RECT 98.100 30.960 99.240 39.850 ;
        RECT 99.940 30.960 101.080 39.850 ;
        RECT 98.100 30.590 101.080 30.960 ;
        RECT 101.780 30.590 102.460 39.850 ;
        RECT 98.100 20.760 102.460 30.590 ;
        RECT 94.420 20.420 102.460 20.760 ;
        RECT 0.560 17.360 102.460 20.420 ;
        RECT 103.160 20.420 104.300 39.850 ;
        RECT 105.000 38.070 106.140 39.850 ;
        RECT 106.840 38.750 107.980 39.850 ;
        RECT 108.680 38.750 109.820 39.850 ;
        RECT 106.840 38.070 109.820 38.750 ;
        RECT 105.000 22.600 109.820 38.070 ;
        RECT 110.520 38.750 111.660 39.850 ;
        RECT 112.360 38.750 113.500 39.850 ;
        RECT 114.200 38.750 115.340 39.850 ;
        RECT 110.520 31.950 115.340 38.750 ;
        RECT 116.040 31.950 117.180 39.850 ;
        RECT 110.520 22.600 117.180 31.950 ;
        RECT 105.000 20.420 117.180 22.600 ;
        RECT 103.160 19.740 117.180 20.420 ;
        RECT 117.880 22.460 119.020 39.850 ;
        RECT 119.720 22.460 120.860 39.850 ;
        RECT 117.880 20.080 120.860 22.460 ;
        RECT 121.560 22.120 122.240 39.850 ;
        RECT 122.940 22.120 124.080 39.850 ;
        RECT 121.560 20.080 124.080 22.120 ;
        RECT 124.780 26.540 125.920 39.850 ;
        RECT 126.620 36.060 127.760 39.850 ;
        RECT 128.460 36.060 129.600 39.850 ;
        RECT 126.620 31.270 129.600 36.060 ;
        RECT 130.300 34.700 131.440 39.850 ;
        RECT 132.140 34.700 133.280 39.850 ;
        RECT 130.300 31.270 133.280 34.700 ;
        RECT 126.620 26.540 133.280 31.270 ;
        RECT 124.780 25.520 133.280 26.540 ;
        RECT 133.980 26.540 135.120 39.850 ;
        RECT 135.820 26.540 136.960 39.850 ;
        RECT 133.980 25.520 136.960 26.540 ;
        RECT 124.780 20.080 136.960 25.520 ;
        RECT 117.880 19.740 136.960 20.080 ;
        RECT 137.660 31.270 138.800 39.850 ;
        RECT 139.500 31.270 140.640 39.850 ;
        RECT 137.660 19.740 140.640 31.270 ;
        RECT 103.160 17.360 140.640 19.740 ;
        RECT 141.340 20.080 142.020 39.850 ;
        RECT 142.720 28.550 143.860 39.850 ;
        RECT 144.560 33.340 145.700 39.850 ;
        RECT 146.400 33.340 147.540 39.850 ;
        RECT 144.560 33.310 147.540 33.340 ;
        RECT 148.240 33.310 149.380 39.850 ;
        RECT 144.560 28.550 149.380 33.310 ;
        RECT 142.720 25.860 149.380 28.550 ;
        RECT 150.080 28.550 151.220 39.850 ;
        RECT 151.920 31.950 153.060 39.850 ;
        RECT 153.760 31.950 154.900 39.850 ;
        RECT 151.920 28.550 154.900 31.950 ;
        RECT 150.080 25.860 154.900 28.550 ;
        RECT 142.720 22.800 154.900 25.860 ;
        RECT 155.600 25.860 156.740 39.850 ;
        RECT 157.440 28.240 158.580 39.850 ;
        RECT 159.280 28.240 160.420 39.850 ;
        RECT 157.440 25.860 160.420 28.240 ;
        RECT 155.600 25.520 160.420 25.860 ;
        RECT 161.120 28.580 162.260 39.850 ;
        RECT 162.960 28.580 163.640 39.850 ;
        RECT 161.120 25.660 163.640 28.580 ;
        RECT 164.340 25.660 165.480 39.850 ;
        RECT 161.120 25.520 165.480 25.660 ;
        RECT 166.180 31.300 167.320 39.850 ;
        RECT 168.020 31.300 169.160 39.850 ;
        RECT 169.860 31.300 171.000 39.850 ;
        RECT 166.180 28.580 171.000 31.300 ;
        RECT 171.700 28.580 172.840 39.850 ;
        RECT 166.180 25.860 172.840 28.580 ;
        RECT 173.540 25.860 174.680 39.850 ;
        RECT 175.380 31.640 176.520 39.850 ;
        RECT 177.220 31.640 178.360 39.850 ;
        RECT 175.380 28.240 178.360 31.640 ;
        RECT 179.060 28.240 180.200 39.850 ;
        RECT 175.380 28.040 180.200 28.240 ;
        RECT 180.900 31.640 182.040 39.850 ;
        RECT 182.740 31.640 183.420 39.850 ;
        RECT 180.900 28.040 183.420 31.640 ;
        RECT 175.380 27.900 183.420 28.040 ;
        RECT 184.120 31.300 185.260 39.850 ;
        RECT 185.960 31.300 187.100 39.850 ;
        RECT 184.120 29.260 187.100 31.300 ;
        RECT 187.800 31.980 188.940 39.850 ;
        RECT 189.640 31.980 190.780 39.850 ;
        RECT 187.800 29.260 190.780 31.980 ;
        RECT 184.120 28.920 190.780 29.260 ;
        RECT 191.480 28.920 192.620 39.850 ;
        RECT 184.120 27.900 192.620 28.920 ;
        RECT 175.380 26.540 192.620 27.900 ;
        RECT 193.320 29.260 194.460 39.850 ;
        RECT 195.160 29.260 196.300 39.850 ;
        RECT 193.320 26.540 196.300 29.260 ;
        RECT 197.000 26.540 198.140 39.850 ;
        RECT 198.840 26.540 199.980 39.850 ;
        RECT 175.380 26.200 199.980 26.540 ;
        RECT 200.680 26.200 201.820 39.850 ;
        RECT 175.380 25.860 201.820 26.200 ;
        RECT 166.180 25.520 201.820 25.860 ;
        RECT 155.600 23.820 201.820 25.520 ;
        RECT 202.520 30.590 203.200 39.850 ;
        RECT 203.900 31.980 205.040 39.850 ;
        RECT 205.740 31.980 206.880 39.850 ;
        RECT 203.900 30.590 206.880 31.980 ;
        RECT 202.520 29.260 206.880 30.590 ;
        RECT 207.580 31.980 208.720 39.850 ;
        RECT 209.420 31.980 210.560 39.850 ;
        RECT 207.580 29.260 210.560 31.980 ;
        RECT 211.260 29.260 212.400 39.850 ;
        RECT 202.520 26.540 212.400 29.260 ;
        RECT 213.100 31.640 214.240 39.850 ;
        RECT 214.940 31.640 216.080 39.850 ;
        RECT 213.100 26.540 216.080 31.640 ;
        RECT 202.520 23.820 216.080 26.540 ;
        RECT 155.600 23.480 216.080 23.820 ;
        RECT 216.780 26.200 217.920 39.850 ;
        RECT 218.620 28.920 219.760 39.850 ;
        RECT 220.460 28.920 221.600 39.850 ;
        RECT 218.620 26.200 221.600 28.920 ;
        RECT 216.780 23.480 221.600 26.200 ;
        RECT 155.600 22.800 221.600 23.480 ;
        RECT 142.720 20.420 221.600 22.800 ;
        RECT 142.720 20.080 222.080 20.420 ;
        RECT 141.340 17.360 222.080 20.080 ;
        RECT 0.560 6.980 222.080 17.360 ;
        RECT 0.560 6.780 61.060 6.980 ;
        RECT 0.560 6.440 27.480 6.780 ;
        RECT 0.560 4.090 5.400 6.440 ;
        RECT 6.100 4.090 16.440 6.440 ;
        RECT 17.140 4.090 27.480 6.440 ;
        RECT 28.180 4.090 38.520 6.780 ;
        RECT 39.220 4.090 50.020 6.780 ;
        RECT 50.720 4.090 61.060 6.780 ;
        RECT 61.760 6.780 222.080 6.980 ;
        RECT 61.760 4.090 72.100 6.780 ;
        RECT 72.800 4.090 83.140 6.780 ;
        RECT 83.840 4.090 94.640 6.780 ;
        RECT 95.340 4.090 105.680 6.780 ;
        RECT 106.380 4.090 116.720 6.780 ;
        RECT 117.420 4.090 127.760 6.780 ;
        RECT 128.460 4.090 139.260 6.780 ;
        RECT 139.960 4.090 150.300 6.780 ;
        RECT 151.000 4.090 161.340 6.780 ;
        RECT 162.040 4.090 172.380 6.780 ;
        RECT 173.080 4.090 183.880 6.780 ;
        RECT 184.580 4.090 194.920 6.780 ;
        RECT 195.620 4.090 205.960 6.780 ;
        RECT 206.660 4.090 217.000 6.780 ;
        RECT 217.700 4.090 222.080 6.780 ;
      LAYER met3 ;
        RECT 40.090 5.275 183.180 32.805 ;
  END
END S_term_DSP
MACRO S_term_RAM_IO
  CLASS BLOCK ;
  FOREIGN S_term_RAM_IO ;
  ORIGIN 0.000 0.000 ;
  SIZE 125.000 BY 40.000 ;
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.920 0.000 3.060 6.500 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.480 0.000 65.620 6.500 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.460 0.000 71.600 6.160 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.900 0.000 78.040 9.560 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.880 0.000 84.020 11.940 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.320 0.000 90.460 11.940 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.760 0.000 96.900 11.940 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.740 0.000 102.880 11.940 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.180 0.000 109.320 7.210 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.160 0.000 115.300 11.600 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.600 0.000 121.740 14.660 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.900 0.000 9.040 6.500 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.340 0.000 15.480 6.500 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.320 0.000 21.460 6.500 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.760 0.000 27.900 6.500 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.200 0.000 34.340 9.560 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.180 0.000 40.320 6.500 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.620 0.000 46.760 11.940 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.600 0.000 52.740 11.940 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.040 0.000 59.180 11.940 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.140 31.920 98.280 40.000 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.940 31.920 112.080 40.000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.320 29.200 113.460 40.000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.700 26.820 114.840 40.000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.080 29.540 116.220 40.000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.460 32.260 117.600 40.000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.840 23.760 118.980 40.000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.220 26.480 120.360 40.000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.600 28.860 121.740 40.000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.980 20.700 123.120 40.000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.360 24.100 124.500 40.000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.520 30.870 99.660 40.000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.900 32.230 101.040 40.000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.280 26.820 102.420 40.000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.660 23.760 103.800 40.000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.040 29.540 105.180 40.000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.420 20.700 106.560 40.000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.800 18.320 107.940 40.000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.180 20.020 109.320 40.000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.560 18.320 110.700 40.000 ;
    END
  END FrameStrobe_O[9]
  PIN N1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.620 31.920 0.760 40.000 ;
    END
  END N1BEG[0]
  PIN N1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.540 29.200 1.680 40.000 ;
    END
  END N1BEG[1]
  PIN N1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.920 32.260 3.060 40.000 ;
    END
  END N1BEG[2]
  PIN N1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.300 30.560 4.440 40.000 ;
    END
  END N1BEG[3]
  PIN N2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.680 26.480 5.820 40.000 ;
    END
  END N2BEG[0]
  PIN N2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.060 28.520 7.200 40.000 ;
    END
  END N2BEG[1]
  PIN N2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.440 26.480 8.580 40.000 ;
    END
  END N2BEG[2]
  PIN N2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.820 29.200 9.960 40.000 ;
    END
  END N2BEG[3]
  PIN N2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.200 32.230 11.340 40.000 ;
    END
  END N2BEG[4]
  PIN N2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.580 26.480 12.720 40.000 ;
    END
  END N2BEG[5]
  PIN N2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.960 32.260 14.100 40.000 ;
    END
  END N2BEG[6]
  PIN N2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.340 29.200 15.480 40.000 ;
    END
  END N2BEG[7]
  PIN N2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.720 26.480 16.860 40.000 ;
    END
  END N2BEGb[0]
  PIN N2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.100 28.860 18.240 40.000 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.480 31.920 19.620 40.000 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.860 26.480 21.000 40.000 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.240 29.540 22.380 40.000 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.620 32.260 23.760 40.000 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.000 32.230 25.140 40.000 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.380 29.200 26.520 40.000 ;
    END
  END N2BEGb[7]
  PIN N4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.760 31.920 27.900 40.000 ;
    END
  END N4BEG[0]
  PIN N4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.100 32.260 41.240 40.000 ;
    END
  END N4BEG[10]
  PIN N4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.480 34.950 42.620 40.000 ;
    END
  END N4BEG[11]
  PIN N4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.860 33.960 44.000 40.000 ;
    END
  END N4BEG[12]
  PIN N4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.240 28.860 45.380 40.000 ;
    END
  END N4BEG[13]
  PIN N4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.620 29.200 46.760 40.000 ;
    END
  END N4BEG[14]
  PIN N4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.000 31.920 48.140 40.000 ;
    END
  END N4BEG[15]
  PIN N4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.140 29.540 29.280 40.000 ;
    END
  END N4BEG[1]
  PIN N4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.520 26.480 30.660 40.000 ;
    END
  END N4BEG[2]
  PIN N4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.900 29.200 32.040 40.000 ;
    END
  END N4BEG[3]
  PIN N4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.820 26.820 32.960 40.000 ;
    END
  END N4BEG[4]
  PIN N4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.200 22.710 34.340 40.000 ;
    END
  END N4BEG[5]
  PIN N4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.580 26.480 35.720 40.000 ;
    END
  END N4BEG[6]
  PIN N4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.960 23.760 37.100 40.000 ;
    END
  END N4BEG[7]
  PIN N4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.340 26.820 38.480 40.000 ;
    END
  END N4BEG[8]
  PIN N4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.720 26.480 39.860 40.000 ;
    END
  END N4BEG[9]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.380 32.230 49.520 40.000 ;
    END
  END S1END[0]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.760 31.720 50.900 40.000 ;
    END
  END S1END[1]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.140 29.040 52.280 40.000 ;
    END
  END S1END[2]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.520 31.380 53.660 40.000 ;
    END
  END S1END[3]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.900 31.720 55.040 40.000 ;
    END
  END S2END[0]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.280 26.820 56.420 40.000 ;
    END
  END S2END[1]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.660 27.680 57.800 40.000 ;
    END
  END S2END[2]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.040 20.700 59.180 40.000 ;
    END
  END S2END[3]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.420 31.550 60.560 40.000 ;
    END
  END S2END[4]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.800 32.260 61.940 40.000 ;
    END
  END S2END[5]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.180 32.230 63.320 40.000 ;
    END
  END S2END[6]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.100 32.910 64.240 40.000 ;
    END
  END S2END[7]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.480 20.700 65.620 40.000 ;
    END
  END S2MID[0]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.860 23.080 67.000 40.000 ;
    END
  END S2MID[1]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.240 26.480 68.380 40.000 ;
    END
  END S2MID[2]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.620 23.420 69.760 40.000 ;
    END
  END S2MID[3]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.000 25.120 71.140 40.000 ;
    END
  END S2MID[4]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.380 23.760 72.520 40.000 ;
    END
  END S2MID[5]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.760 28.180 73.900 40.000 ;
    END
  END S2MID[6]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.140 25.460 75.280 40.000 ;
    END
  END S2MID[7]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.520 31.380 76.660 40.000 ;
    END
  END S4END[0]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.320 26.140 90.460 40.000 ;
    END
  END S4END[10]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.700 23.080 91.840 40.000 ;
    END
  END S4END[11]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.080 28.860 93.220 40.000 ;
    END
  END S4END[12]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.460 23.080 94.600 40.000 ;
    END
  END S4END[13]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.380 31.240 95.520 40.000 ;
    END
  END S4END[14]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.760 22.740 96.900 40.000 ;
    END
  END S4END[15]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.900 32.910 78.040 40.000 ;
    END
  END S4END[1]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.280 31.240 79.420 40.000 ;
    END
  END S4END[2]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.660 33.590 80.800 40.000 ;
    END
  END S4END[3]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.040 34.270 82.180 40.000 ;
    END
  END S4END[4]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.420 28.830 83.560 40.000 ;
    END
  END S4END[5]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.800 17.640 84.940 40.000 ;
    END
  END S4END[6]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.180 20.360 86.320 40.000 ;
    END
  END S4END[7]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.560 17.640 87.700 40.000 ;
    END
  END S4END[8]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.940 20.360 89.080 40.000 ;
    END
  END S4END[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 23.715 5.200 25.315 32.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 61.700 5.200 63.300 32.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 99.685 5.200 101.285 32.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 42.705 5.200 44.305 32.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 80.690 5.200 82.290 32.880 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 119.140 32.725 ;
      LAYER met1 ;
        RECT 0.530 4.120 124.590 36.340 ;
      LAYER met2 ;
        RECT 1.040 31.640 1.260 36.370 ;
        RECT 0.560 28.920 1.260 31.640 ;
        RECT 1.960 31.980 2.640 36.370 ;
        RECT 3.340 31.980 4.020 36.370 ;
        RECT 1.960 30.280 4.020 31.980 ;
        RECT 4.720 30.280 5.400 36.370 ;
        RECT 1.960 28.920 5.400 30.280 ;
        RECT 0.560 26.200 5.400 28.920 ;
        RECT 6.100 28.240 6.780 36.370 ;
        RECT 7.480 28.240 8.160 36.370 ;
        RECT 6.100 26.200 8.160 28.240 ;
        RECT 8.860 28.920 9.540 36.370 ;
        RECT 10.240 31.950 10.920 36.370 ;
        RECT 11.620 31.950 12.300 36.370 ;
        RECT 10.240 28.920 12.300 31.950 ;
        RECT 8.860 26.200 12.300 28.920 ;
        RECT 13.000 31.980 13.680 36.370 ;
        RECT 14.380 31.980 15.060 36.370 ;
        RECT 13.000 28.920 15.060 31.980 ;
        RECT 15.760 28.920 16.440 36.370 ;
        RECT 13.000 26.200 16.440 28.920 ;
        RECT 17.140 28.580 17.820 36.370 ;
        RECT 18.520 31.640 19.200 36.370 ;
        RECT 19.900 31.640 20.580 36.370 ;
        RECT 18.520 28.580 20.580 31.640 ;
        RECT 17.140 26.200 20.580 28.580 ;
        RECT 21.280 29.260 21.960 36.370 ;
        RECT 22.660 31.980 23.340 36.370 ;
        RECT 24.040 31.980 24.720 36.370 ;
        RECT 22.660 31.950 24.720 31.980 ;
        RECT 25.420 31.950 26.100 36.370 ;
        RECT 22.660 29.260 26.100 31.950 ;
        RECT 21.280 28.920 26.100 29.260 ;
        RECT 26.800 31.640 27.480 36.370 ;
        RECT 28.180 31.640 28.860 36.370 ;
        RECT 26.800 29.260 28.860 31.640 ;
        RECT 29.560 29.260 30.240 36.370 ;
        RECT 26.800 28.920 30.240 29.260 ;
        RECT 21.280 26.200 30.240 28.920 ;
        RECT 30.940 28.920 31.620 36.370 ;
        RECT 32.320 28.920 32.540 36.370 ;
        RECT 30.940 26.540 32.540 28.920 ;
        RECT 33.240 26.540 33.920 36.370 ;
        RECT 30.940 26.200 33.920 26.540 ;
        RECT 0.560 22.430 33.920 26.200 ;
        RECT 34.620 26.200 35.300 36.370 ;
        RECT 36.000 26.200 36.680 36.370 ;
        RECT 34.620 23.480 36.680 26.200 ;
        RECT 37.380 26.540 38.060 36.370 ;
        RECT 38.760 26.540 39.440 36.370 ;
        RECT 37.380 26.200 39.440 26.540 ;
        RECT 40.140 31.980 40.820 36.370 ;
        RECT 41.520 34.670 42.200 36.370 ;
        RECT 42.900 34.670 43.580 36.370 ;
        RECT 41.520 33.680 43.580 34.670 ;
        RECT 44.280 33.680 44.960 36.370 ;
        RECT 41.520 31.980 44.960 33.680 ;
        RECT 40.140 28.580 44.960 31.980 ;
        RECT 45.660 28.920 46.340 36.370 ;
        RECT 47.040 31.640 47.720 36.370 ;
        RECT 48.420 31.950 49.100 36.370 ;
        RECT 49.800 31.950 50.480 36.370 ;
        RECT 48.420 31.640 50.480 31.950 ;
        RECT 47.040 31.440 50.480 31.640 ;
        RECT 51.180 31.440 51.860 36.370 ;
        RECT 47.040 28.920 51.860 31.440 ;
        RECT 45.660 28.760 51.860 28.920 ;
        RECT 52.560 31.100 53.240 36.370 ;
        RECT 53.940 31.440 54.620 36.370 ;
        RECT 55.320 31.440 56.000 36.370 ;
        RECT 53.940 31.100 56.000 31.440 ;
        RECT 52.560 28.760 56.000 31.100 ;
        RECT 45.660 28.580 56.000 28.760 ;
        RECT 40.140 26.540 56.000 28.580 ;
        RECT 56.700 27.400 57.380 36.370 ;
        RECT 58.080 27.400 58.760 36.370 ;
        RECT 56.700 26.540 58.760 27.400 ;
        RECT 40.140 26.200 58.760 26.540 ;
        RECT 37.380 23.480 58.760 26.200 ;
        RECT 34.620 22.430 58.760 23.480 ;
        RECT 0.560 20.420 58.760 22.430 ;
        RECT 59.460 31.270 60.140 36.370 ;
        RECT 60.840 31.980 61.520 36.370 ;
        RECT 62.220 31.980 62.900 36.370 ;
        RECT 60.840 31.950 62.900 31.980 ;
        RECT 63.600 32.630 63.820 36.370 ;
        RECT 64.520 32.630 65.200 36.370 ;
        RECT 63.600 31.950 65.200 32.630 ;
        RECT 60.840 31.270 65.200 31.950 ;
        RECT 59.460 20.420 65.200 31.270 ;
        RECT 65.900 22.800 66.580 36.370 ;
        RECT 67.280 26.200 67.960 36.370 ;
        RECT 68.660 26.200 69.340 36.370 ;
        RECT 67.280 23.140 69.340 26.200 ;
        RECT 70.040 24.840 70.720 36.370 ;
        RECT 71.420 24.840 72.100 36.370 ;
        RECT 70.040 23.480 72.100 24.840 ;
        RECT 72.800 27.900 73.480 36.370 ;
        RECT 74.180 27.900 74.860 36.370 ;
        RECT 72.800 25.180 74.860 27.900 ;
        RECT 75.560 31.100 76.240 36.370 ;
        RECT 76.940 32.630 77.620 36.370 ;
        RECT 78.320 32.630 79.000 36.370 ;
        RECT 76.940 31.100 79.000 32.630 ;
        RECT 75.560 30.960 79.000 31.100 ;
        RECT 79.700 33.310 80.380 36.370 ;
        RECT 81.080 33.990 81.760 36.370 ;
        RECT 82.460 33.990 83.140 36.370 ;
        RECT 81.080 33.310 83.140 33.990 ;
        RECT 79.700 30.960 83.140 33.310 ;
        RECT 75.560 28.550 83.140 30.960 ;
        RECT 83.840 28.550 84.520 36.370 ;
        RECT 75.560 25.180 84.520 28.550 ;
        RECT 72.800 23.480 84.520 25.180 ;
        RECT 70.040 23.140 84.520 23.480 ;
        RECT 67.280 22.800 84.520 23.140 ;
        RECT 65.900 20.420 84.520 22.800 ;
        RECT 0.560 17.360 84.520 20.420 ;
        RECT 85.220 20.080 85.900 36.370 ;
        RECT 86.600 20.080 87.280 36.370 ;
        RECT 85.220 17.360 87.280 20.080 ;
        RECT 87.980 20.080 88.660 36.370 ;
        RECT 89.360 25.860 90.040 36.370 ;
        RECT 90.740 25.860 91.420 36.370 ;
        RECT 89.360 22.800 91.420 25.860 ;
        RECT 92.120 28.580 92.800 36.370 ;
        RECT 93.500 28.580 94.180 36.370 ;
        RECT 92.120 22.800 94.180 28.580 ;
        RECT 94.880 30.960 95.100 36.370 ;
        RECT 95.800 30.960 96.480 36.370 ;
        RECT 94.880 22.800 96.480 30.960 ;
        RECT 89.360 22.460 96.480 22.800 ;
        RECT 97.180 31.640 97.860 36.370 ;
        RECT 98.560 31.640 99.240 36.370 ;
        RECT 97.180 30.590 99.240 31.640 ;
        RECT 99.940 31.950 100.620 36.370 ;
        RECT 101.320 31.950 102.000 36.370 ;
        RECT 99.940 30.590 102.000 31.950 ;
        RECT 97.180 26.540 102.000 30.590 ;
        RECT 102.700 26.540 103.380 36.370 ;
        RECT 97.180 23.480 103.380 26.540 ;
        RECT 104.080 29.260 104.760 36.370 ;
        RECT 105.460 29.260 106.140 36.370 ;
        RECT 104.080 23.480 106.140 29.260 ;
        RECT 97.180 22.460 106.140 23.480 ;
        RECT 89.360 20.420 106.140 22.460 ;
        RECT 106.840 20.420 107.520 36.370 ;
        RECT 89.360 20.080 107.520 20.420 ;
        RECT 87.980 18.040 107.520 20.080 ;
        RECT 108.220 19.740 108.900 36.370 ;
        RECT 109.600 19.740 110.280 36.370 ;
        RECT 108.220 18.040 110.280 19.740 ;
        RECT 110.980 31.640 111.660 36.370 ;
        RECT 112.360 31.640 113.040 36.370 ;
        RECT 110.980 28.920 113.040 31.640 ;
        RECT 113.740 28.920 114.420 36.370 ;
        RECT 110.980 26.540 114.420 28.920 ;
        RECT 115.120 29.260 115.800 36.370 ;
        RECT 116.500 31.980 117.180 36.370 ;
        RECT 117.880 31.980 118.560 36.370 ;
        RECT 116.500 29.260 118.560 31.980 ;
        RECT 115.120 26.540 118.560 29.260 ;
        RECT 110.980 23.480 118.560 26.540 ;
        RECT 119.260 26.200 119.940 36.370 ;
        RECT 120.640 28.580 121.320 36.370 ;
        RECT 122.020 28.580 122.700 36.370 ;
        RECT 120.640 26.200 122.700 28.580 ;
        RECT 119.260 23.480 122.700 26.200 ;
        RECT 110.980 20.420 122.700 23.480 ;
        RECT 123.400 23.820 124.080 36.370 ;
        RECT 123.400 20.420 124.560 23.820 ;
        RECT 110.980 18.040 124.560 20.420 ;
        RECT 87.980 17.360 124.560 18.040 ;
        RECT 0.560 14.940 124.560 17.360 ;
        RECT 0.560 12.220 121.320 14.940 ;
        RECT 0.560 9.840 46.340 12.220 ;
        RECT 0.560 6.780 33.920 9.840 ;
        RECT 0.560 4.090 2.640 6.780 ;
        RECT 3.340 4.090 8.620 6.780 ;
        RECT 9.320 4.090 15.060 6.780 ;
        RECT 15.760 4.090 21.040 6.780 ;
        RECT 21.740 4.090 27.480 6.780 ;
        RECT 28.180 4.090 33.920 6.780 ;
        RECT 34.620 6.780 46.340 9.840 ;
        RECT 34.620 4.090 39.900 6.780 ;
        RECT 40.600 4.090 46.340 6.780 ;
        RECT 47.040 4.090 52.320 12.220 ;
        RECT 53.020 4.090 58.760 12.220 ;
        RECT 59.460 9.840 83.600 12.220 ;
        RECT 59.460 6.780 77.620 9.840 ;
        RECT 59.460 4.090 65.200 6.780 ;
        RECT 65.900 6.440 77.620 6.780 ;
        RECT 65.900 4.090 71.180 6.440 ;
        RECT 71.880 4.090 77.620 6.440 ;
        RECT 78.320 4.090 83.600 9.840 ;
        RECT 84.300 4.090 90.040 12.220 ;
        RECT 90.740 4.090 96.480 12.220 ;
        RECT 97.180 4.090 102.460 12.220 ;
        RECT 103.160 11.880 121.320 12.220 ;
        RECT 103.160 7.490 114.880 11.880 ;
        RECT 103.160 4.090 108.900 7.490 ;
        RECT 109.600 4.090 114.880 7.490 ;
        RECT 115.580 4.090 121.320 11.880 ;
        RECT 122.020 4.090 124.560 14.940 ;
      LAYER met3 ;
        RECT 7.885 5.275 101.285 32.805 ;
  END
END S_term_RAM_IO
MACRO S_term_single
  CLASS BLOCK ;
  FOREIGN S_term_single ;
  ORIGIN 0.000 0.000 ;
  SIZE 223.275 BY 40.000 ;
  PIN Co
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.000 26.110 186.140 40.000 ;
    END
  END Co
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.680 0.000 5.820 6.160 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.000 0.000 117.140 6.500 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.040 0.000 128.180 6.500 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.540 0.000 139.680 6.500 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.580 0.000 150.720 6.500 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.620 0.000 161.760 6.500 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.660 0.000 172.800 6.500 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.160 0.000 184.300 6.500 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.200 0.000 195.340 6.500 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.240 0.000 206.380 6.500 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.280 0.000 217.420 6.500 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.720 0.000 16.860 6.160 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.760 0.000 27.900 6.500 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.800 0.000 38.940 6.500 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.300 0.000 50.440 6.500 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.340 0.000 61.480 6.500 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.380 0.000 72.520 6.500 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.420 0.000 83.560 6.500 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.920 0.000 95.060 6.500 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.960 0.000 106.100 6.500 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.840 29.540 187.980 40.000 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.780 32.260 205.920 40.000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.620 32.260 207.760 40.000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.000 29.540 209.140 40.000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.840 26.140 210.980 40.000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.680 29.200 212.820 40.000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.520 31.920 214.660 40.000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.360 23.760 216.500 40.000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.200 26.820 218.340 40.000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.040 28.860 220.180 40.000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.880 20.700 222.020 40.000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.680 32.260 189.820 40.000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.520 29.200 191.660 40.000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.360 26.820 193.500 40.000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.740 32.230 194.880 40.000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.580 26.480 196.720 40.000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.420 24.100 198.560 40.000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.260 32.230 200.400 40.000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.100 23.760 202.240 40.000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.940 20.360 204.080 40.000 ;
    END
  END FrameStrobe_O[9]
  PIN N1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.620 32.260 0.760 40.000 ;
    END
  END N1BEG[0]
  PIN N1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.000 29.540 2.140 40.000 ;
    END
  END N1BEG[1]
  PIN N1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.840 31.920 3.980 40.000 ;
    END
  END N1BEG[2]
  PIN N1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.680 31.240 5.820 40.000 ;
    END
  END N1BEG[3]
  PIN N2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.520 33.590 7.660 40.000 ;
    END
  END N2BEG[0]
  PIN N2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.360 26.820 9.500 40.000 ;
    END
  END N2BEG[1]
  PIN N2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.200 39.030 11.340 40.000 ;
    END
  END N2BEG[2]
  PIN N2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.040 32.260 13.180 40.000 ;
    END
  END N2BEG[3]
  PIN N2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.880 29.200 15.020 40.000 ;
    END
  END N2BEG[4]
  PIN N2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.260 31.920 16.400 40.000 ;
    END
  END N2BEG[5]
  PIN N2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.100 29.540 18.240 40.000 ;
    END
  END N2BEG[6]
  PIN N2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.940 32.060 20.080 40.000 ;
    END
  END N2BEG[7]
  PIN N2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.780 29.200 21.920 40.000 ;
    END
  END N2BEGb[0]
  PIN N2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.620 34.950 23.760 40.000 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.460 29.540 25.600 40.000 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.300 30.560 27.440 40.000 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.140 27.840 29.280 40.000 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.520 26.820 30.660 40.000 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.360 29.540 32.500 40.000 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.200 26.820 34.340 40.000 ;
    END
  END N2BEGb[7]
  PIN N4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.040 32.260 36.180 40.000 ;
    END
  END N4BEG[0]
  PIN N4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.980 32.260 54.120 40.000 ;
    END
  END N4BEG[10]
  PIN N4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.820 29.540 55.960 40.000 ;
    END
  END N4BEG[11]
  PIN N4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.660 39.030 57.800 40.000 ;
    END
  END N4BEG[12]
  PIN N4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.500 34.640 59.640 40.000 ;
    END
  END N4BEG[13]
  PIN N4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.880 26.820 61.020 40.000 ;
    END
  END N4BEG[14]
  PIN N4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.720 29.540 62.860 40.000 ;
    END
  END N4BEG[15]
  PIN N4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.880 26.820 38.020 40.000 ;
    END
  END N4BEG[1]
  PIN N4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.720 31.920 39.860 40.000 ;
    END
  END N4BEG[2]
  PIN N4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.560 33.590 41.700 40.000 ;
    END
  END N4BEG[3]
  PIN N4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.400 30.560 43.540 40.000 ;
    END
  END N4BEG[4]
  PIN N4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.240 28.860 45.380 40.000 ;
    END
  END N4BEG[5]
  PIN N4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.620 26.480 46.760 40.000 ;
    END
  END N4BEG[6]
  PIN N4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.460 29.540 48.600 40.000 ;
    END
  END N4BEG[7]
  PIN N4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.300 26.820 50.440 40.000 ;
    END
  END N4BEG[8]
  PIN N4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.140 24.100 52.280 40.000 ;
    END
  END N4BEG[9]
  PIN NN4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.560 32.260 64.700 40.000 ;
    END
  END NN4BEG[0]
  PIN NN4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.500 32.260 82.640 40.000 ;
    END
  END NN4BEG[10]
  PIN NN4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.340 34.950 84.480 40.000 ;
    END
  END NN4BEG[11]
  PIN NN4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.180 28.860 86.320 40.000 ;
    END
  END NN4BEG[12]
  PIN NN4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.020 29.540 88.160 40.000 ;
    END
  END NN4BEG[13]
  PIN NN4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.860 28.860 90.000 40.000 ;
    END
  END NN4BEG[14]
  PIN NN4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.240 33.590 91.380 40.000 ;
    END
  END NN4BEG[15]
  PIN NN4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.400 29.200 66.540 40.000 ;
    END
  END NN4BEG[1]
  PIN NN4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.240 31.920 68.380 40.000 ;
    END
  END NN4BEG[2]
  PIN NN4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.080 30.560 70.220 40.000 ;
    END
  END NN4BEG[3]
  PIN NN4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.920 26.820 72.060 40.000 ;
    END
  END NN4BEG[4]
  PIN NN4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.760 26.820 73.900 40.000 ;
    END
  END NN4BEG[5]
  PIN NN4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.140 32.060 75.280 40.000 ;
    END
  END NN4BEG[6]
  PIN NN4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.980 34.640 77.120 40.000 ;
    END
  END NN4BEG[7]
  PIN NN4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.820 26.820 78.960 40.000 ;
    END
  END NN4BEG[8]
  PIN NN4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.660 24.100 80.800 40.000 ;
    END
  END NN4BEG[9]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.080 31.580 93.220 40.000 ;
    END
  END S1END[0]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.920 28.860 95.060 40.000 ;
    END
  END S1END[1]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.760 30.900 96.900 40.000 ;
    END
  END S1END[2]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.600 39.030 98.740 40.000 ;
    END
  END S1END[3]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.440 25.800 100.580 40.000 ;
    END
  END S2END[0]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.280 32.910 102.420 40.000 ;
    END
  END S2END[1]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.120 23.080 104.260 40.000 ;
    END
  END S2END[2]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.500 32.910 105.640 40.000 ;
    END
  END S2END[3]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.340 22.740 107.480 40.000 ;
    END
  END S2END[4]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.180 20.700 109.320 40.000 ;
    END
  END S2END[5]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.020 30.360 111.160 40.000 ;
    END
  END S2END[6]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.860 39.030 113.000 40.000 ;
    END
  END S2END[7]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.700 39.030 114.840 40.000 ;
    END
  END S2MID[0]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.540 26.820 116.680 40.000 ;
    END
  END S2MID[1]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.380 23.420 118.520 40.000 ;
    END
  END S2MID[2]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.760 25.800 119.900 40.000 ;
    END
  END S2MID[3]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.600 23.760 121.740 40.000 ;
    END
  END S2MID[4]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.440 20.700 123.580 40.000 ;
    END
  END S2MID[5]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.280 23.760 125.420 40.000 ;
    END
  END S2MID[6]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.120 32.910 127.260 40.000 ;
    END
  END S2MID[7]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.960 23.420 129.100 40.000 ;
    END
  END S4END[0]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.900 39.030 147.040 40.000 ;
    END
  END S4END[10]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.740 32.910 148.880 40.000 ;
    END
  END S4END[11]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.120 26.480 150.260 40.000 ;
    END
  END S4END[12]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.960 28.860 152.100 40.000 ;
    END
  END S4END[13]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.800 25.800 153.940 40.000 ;
    END
  END S4END[14]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.640 28.860 155.780 40.000 ;
    END
  END S4END[15]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.800 32.910 130.940 40.000 ;
    END
  END S4END[1]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.640 23.420 132.780 40.000 ;
    END
  END S4END[2]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.480 32.910 134.620 40.000 ;
    END
  END S4END[3]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.860 39.030 136.000 40.000 ;
    END
  END S4END[4]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.700 23.420 137.840 40.000 ;
    END
  END S4END[5]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.540 30.190 139.680 40.000 ;
    END
  END S4END[6]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.380 22.740 141.520 40.000 ;
    END
  END S4END[7]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.220 30.190 143.360 40.000 ;
    END
  END S4END[8]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.060 23.420 145.200 40.000 ;
    END
  END S4END[9]
  PIN SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.480 27.640 157.620 40.000 ;
    END
  END SS4END[0]
  PIN SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.420 31.920 175.560 40.000 ;
    END
  END SS4END[10]
  PIN SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.260 28.860 177.400 40.000 ;
    END
  END SS4END[11]
  PIN SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.100 27.840 179.240 40.000 ;
    END
  END SS4END[12]
  PIN SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.480 35.630 180.620 40.000 ;
    END
  END SS4END[13]
  PIN SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.320 31.580 182.460 40.000 ;
    END
  END SS4END[14]
  PIN SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.160 28.320 184.300 40.000 ;
    END
  END SS4END[15]
  PIN SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.320 25.800 159.460 40.000 ;
    END
  END SS4END[1]
  PIN SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.160 23.080 161.300 40.000 ;
    END
  END SS4END[2]
  PIN SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.000 26.480 163.140 40.000 ;
    END
  END SS4END[3]
  PIN SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.380 23.080 164.520 40.000 ;
    END
  END SS4END[4]
  PIN SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.220 31.580 166.360 40.000 ;
    END
  END SS4END[5]
  PIN SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.060 31.920 168.200 40.000 ;
    END
  END SS4END[6]
  PIN SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.900 28.860 170.040 40.000 ;
    END
  END SS4END[7]
  PIN SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.740 26.140 171.880 40.000 ;
    END
  END SS4END[8]
  PIN SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.580 28.180 173.720 40.000 ;
    END
  END SS4END[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 40.090 5.200 41.690 32.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 110.835 5.200 112.435 32.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 181.580 5.200 183.180 32.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 75.465 5.200 77.065 32.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 146.210 5.200 147.810 32.880 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 217.580 39.695 ;
      LAYER met1 ;
        RECT 0.530 4.120 222.110 39.740 ;
      LAYER met2 ;
        RECT 1.040 31.980 1.720 39.850 ;
        RECT 0.560 29.260 1.720 31.980 ;
        RECT 2.420 31.640 3.560 39.850 ;
        RECT 4.260 31.640 5.400 39.850 ;
        RECT 2.420 30.960 5.400 31.640 ;
        RECT 6.100 33.310 7.240 39.850 ;
        RECT 7.940 33.310 9.080 39.850 ;
        RECT 6.100 30.960 9.080 33.310 ;
        RECT 2.420 29.260 9.080 30.960 ;
        RECT 0.560 26.540 9.080 29.260 ;
        RECT 9.780 38.750 10.920 39.850 ;
        RECT 11.620 38.750 12.760 39.850 ;
        RECT 9.780 31.980 12.760 38.750 ;
        RECT 13.460 31.980 14.600 39.850 ;
        RECT 9.780 28.920 14.600 31.980 ;
        RECT 15.300 31.640 15.980 39.850 ;
        RECT 16.680 31.640 17.820 39.850 ;
        RECT 15.300 29.260 17.820 31.640 ;
        RECT 18.520 31.780 19.660 39.850 ;
        RECT 20.360 31.780 21.500 39.850 ;
        RECT 18.520 29.260 21.500 31.780 ;
        RECT 15.300 28.920 21.500 29.260 ;
        RECT 22.200 34.670 23.340 39.850 ;
        RECT 24.040 34.670 25.180 39.850 ;
        RECT 22.200 29.260 25.180 34.670 ;
        RECT 25.880 30.280 27.020 39.850 ;
        RECT 27.720 30.280 28.860 39.850 ;
        RECT 25.880 29.260 28.860 30.280 ;
        RECT 22.200 28.920 28.860 29.260 ;
        RECT 9.780 27.560 28.860 28.920 ;
        RECT 29.560 27.560 30.240 39.850 ;
        RECT 9.780 26.540 30.240 27.560 ;
        RECT 30.940 29.260 32.080 39.850 ;
        RECT 32.780 29.260 33.920 39.850 ;
        RECT 30.940 26.540 33.920 29.260 ;
        RECT 34.620 31.980 35.760 39.850 ;
        RECT 36.460 31.980 37.600 39.850 ;
        RECT 34.620 26.540 37.600 31.980 ;
        RECT 38.300 31.640 39.440 39.850 ;
        RECT 40.140 33.310 41.280 39.850 ;
        RECT 41.980 33.310 43.120 39.850 ;
        RECT 40.140 31.640 43.120 33.310 ;
        RECT 38.300 30.280 43.120 31.640 ;
        RECT 43.820 30.280 44.960 39.850 ;
        RECT 38.300 28.580 44.960 30.280 ;
        RECT 45.660 28.580 46.340 39.850 ;
        RECT 38.300 26.540 46.340 28.580 ;
        RECT 0.560 26.200 46.340 26.540 ;
        RECT 47.040 29.260 48.180 39.850 ;
        RECT 48.880 29.260 50.020 39.850 ;
        RECT 47.040 26.540 50.020 29.260 ;
        RECT 50.720 26.540 51.860 39.850 ;
        RECT 47.040 26.200 51.860 26.540 ;
        RECT 0.560 23.820 51.860 26.200 ;
        RECT 52.560 31.980 53.700 39.850 ;
        RECT 54.400 31.980 55.540 39.850 ;
        RECT 52.560 29.260 55.540 31.980 ;
        RECT 56.240 38.750 57.380 39.850 ;
        RECT 58.080 38.750 59.220 39.850 ;
        RECT 56.240 34.360 59.220 38.750 ;
        RECT 59.920 34.360 60.600 39.850 ;
        RECT 56.240 29.260 60.600 34.360 ;
        RECT 52.560 26.540 60.600 29.260 ;
        RECT 61.300 29.260 62.440 39.850 ;
        RECT 63.140 31.980 64.280 39.850 ;
        RECT 64.980 31.980 66.120 39.850 ;
        RECT 63.140 29.260 66.120 31.980 ;
        RECT 61.300 28.920 66.120 29.260 ;
        RECT 66.820 31.640 67.960 39.850 ;
        RECT 68.660 31.640 69.800 39.850 ;
        RECT 66.820 30.280 69.800 31.640 ;
        RECT 70.500 30.280 71.640 39.850 ;
        RECT 66.820 28.920 71.640 30.280 ;
        RECT 61.300 26.540 71.640 28.920 ;
        RECT 72.340 26.540 73.480 39.850 ;
        RECT 74.180 31.780 74.860 39.850 ;
        RECT 75.560 34.360 76.700 39.850 ;
        RECT 77.400 34.360 78.540 39.850 ;
        RECT 75.560 31.780 78.540 34.360 ;
        RECT 74.180 26.540 78.540 31.780 ;
        RECT 79.240 26.540 80.380 39.850 ;
        RECT 52.560 23.820 80.380 26.540 ;
        RECT 81.080 31.980 82.220 39.850 ;
        RECT 82.920 34.670 84.060 39.850 ;
        RECT 84.760 34.670 85.900 39.850 ;
        RECT 82.920 31.980 85.900 34.670 ;
        RECT 81.080 28.580 85.900 31.980 ;
        RECT 86.600 29.260 87.740 39.850 ;
        RECT 88.440 29.260 89.580 39.850 ;
        RECT 86.600 28.580 89.580 29.260 ;
        RECT 90.280 33.310 90.960 39.850 ;
        RECT 91.660 33.310 92.800 39.850 ;
        RECT 90.280 31.300 92.800 33.310 ;
        RECT 93.500 31.300 94.640 39.850 ;
        RECT 90.280 28.580 94.640 31.300 ;
        RECT 95.340 30.620 96.480 39.850 ;
        RECT 97.180 38.750 98.320 39.850 ;
        RECT 99.020 38.750 100.160 39.850 ;
        RECT 97.180 30.620 100.160 38.750 ;
        RECT 95.340 28.580 100.160 30.620 ;
        RECT 81.080 25.520 100.160 28.580 ;
        RECT 100.860 32.630 102.000 39.850 ;
        RECT 102.700 32.630 103.840 39.850 ;
        RECT 100.860 25.520 103.840 32.630 ;
        RECT 81.080 23.820 103.840 25.520 ;
        RECT 0.560 22.800 103.840 23.820 ;
        RECT 104.540 32.630 105.220 39.850 ;
        RECT 105.920 32.630 107.060 39.850 ;
        RECT 104.540 22.800 107.060 32.630 ;
        RECT 0.560 22.460 107.060 22.800 ;
        RECT 107.760 22.460 108.900 39.850 ;
        RECT 0.560 20.420 108.900 22.460 ;
        RECT 109.600 30.080 110.740 39.850 ;
        RECT 111.440 38.750 112.580 39.850 ;
        RECT 113.280 38.750 114.420 39.850 ;
        RECT 115.120 38.750 116.260 39.850 ;
        RECT 111.440 30.080 116.260 38.750 ;
        RECT 109.600 26.540 116.260 30.080 ;
        RECT 116.960 26.540 118.100 39.850 ;
        RECT 109.600 23.140 118.100 26.540 ;
        RECT 118.800 25.520 119.480 39.850 ;
        RECT 120.180 25.520 121.320 39.850 ;
        RECT 118.800 23.480 121.320 25.520 ;
        RECT 122.020 23.480 123.160 39.850 ;
        RECT 118.800 23.140 123.160 23.480 ;
        RECT 109.600 20.420 123.160 23.140 ;
        RECT 123.860 23.480 125.000 39.850 ;
        RECT 125.700 32.630 126.840 39.850 ;
        RECT 127.540 32.630 128.680 39.850 ;
        RECT 125.700 23.480 128.680 32.630 ;
        RECT 123.860 23.140 128.680 23.480 ;
        RECT 129.380 32.630 130.520 39.850 ;
        RECT 131.220 32.630 132.360 39.850 ;
        RECT 129.380 23.140 132.360 32.630 ;
        RECT 133.060 32.630 134.200 39.850 ;
        RECT 134.900 38.750 135.580 39.850 ;
        RECT 136.280 38.750 137.420 39.850 ;
        RECT 134.900 32.630 137.420 38.750 ;
        RECT 133.060 23.140 137.420 32.630 ;
        RECT 138.120 29.910 139.260 39.850 ;
        RECT 139.960 29.910 141.100 39.850 ;
        RECT 138.120 23.140 141.100 29.910 ;
        RECT 123.860 22.460 141.100 23.140 ;
        RECT 141.800 29.910 142.940 39.850 ;
        RECT 143.640 29.910 144.780 39.850 ;
        RECT 141.800 23.140 144.780 29.910 ;
        RECT 145.480 38.750 146.620 39.850 ;
        RECT 147.320 38.750 148.460 39.850 ;
        RECT 145.480 32.630 148.460 38.750 ;
        RECT 149.160 32.630 149.840 39.850 ;
        RECT 145.480 26.200 149.840 32.630 ;
        RECT 150.540 28.580 151.680 39.850 ;
        RECT 152.380 28.580 153.520 39.850 ;
        RECT 150.540 26.200 153.520 28.580 ;
        RECT 145.480 25.520 153.520 26.200 ;
        RECT 154.220 28.580 155.360 39.850 ;
        RECT 156.060 28.580 157.200 39.850 ;
        RECT 154.220 27.360 157.200 28.580 ;
        RECT 157.900 27.360 159.040 39.850 ;
        RECT 154.220 25.520 159.040 27.360 ;
        RECT 159.740 25.520 160.880 39.850 ;
        RECT 145.480 23.140 160.880 25.520 ;
        RECT 141.800 22.800 160.880 23.140 ;
        RECT 161.580 26.200 162.720 39.850 ;
        RECT 163.420 26.200 164.100 39.850 ;
        RECT 161.580 22.800 164.100 26.200 ;
        RECT 164.800 31.300 165.940 39.850 ;
        RECT 166.640 31.640 167.780 39.850 ;
        RECT 168.480 31.640 169.620 39.850 ;
        RECT 166.640 31.300 169.620 31.640 ;
        RECT 164.800 28.580 169.620 31.300 ;
        RECT 170.320 28.580 171.460 39.850 ;
        RECT 164.800 25.860 171.460 28.580 ;
        RECT 172.160 27.900 173.300 39.850 ;
        RECT 174.000 31.640 175.140 39.850 ;
        RECT 175.840 31.640 176.980 39.850 ;
        RECT 174.000 28.580 176.980 31.640 ;
        RECT 177.680 28.580 178.820 39.850 ;
        RECT 174.000 27.900 178.820 28.580 ;
        RECT 172.160 27.560 178.820 27.900 ;
        RECT 179.520 35.350 180.200 39.850 ;
        RECT 180.900 35.350 182.040 39.850 ;
        RECT 179.520 31.300 182.040 35.350 ;
        RECT 182.740 31.300 183.880 39.850 ;
        RECT 179.520 28.040 183.880 31.300 ;
        RECT 184.580 28.040 185.720 39.850 ;
        RECT 179.520 27.560 185.720 28.040 ;
        RECT 172.160 25.860 185.720 27.560 ;
        RECT 164.800 25.830 185.720 25.860 ;
        RECT 186.420 29.260 187.560 39.850 ;
        RECT 188.260 31.980 189.400 39.850 ;
        RECT 190.100 31.980 191.240 39.850 ;
        RECT 188.260 29.260 191.240 31.980 ;
        RECT 186.420 28.920 191.240 29.260 ;
        RECT 191.940 28.920 193.080 39.850 ;
        RECT 186.420 26.540 193.080 28.920 ;
        RECT 193.780 31.950 194.460 39.850 ;
        RECT 195.160 31.950 196.300 39.850 ;
        RECT 193.780 26.540 196.300 31.950 ;
        RECT 186.420 26.200 196.300 26.540 ;
        RECT 197.000 26.200 198.140 39.850 ;
        RECT 186.420 25.830 198.140 26.200 ;
        RECT 164.800 23.820 198.140 25.830 ;
        RECT 198.840 31.950 199.980 39.850 ;
        RECT 200.680 31.950 201.820 39.850 ;
        RECT 198.840 23.820 201.820 31.950 ;
        RECT 164.800 23.480 201.820 23.820 ;
        RECT 202.520 23.480 203.660 39.850 ;
        RECT 164.800 22.800 203.660 23.480 ;
        RECT 141.800 22.460 203.660 22.800 ;
        RECT 123.860 20.420 203.660 22.460 ;
        RECT 0.560 20.080 203.660 20.420 ;
        RECT 204.360 31.980 205.500 39.850 ;
        RECT 206.200 31.980 207.340 39.850 ;
        RECT 208.040 31.980 208.720 39.850 ;
        RECT 204.360 29.260 208.720 31.980 ;
        RECT 209.420 29.260 210.560 39.850 ;
        RECT 204.360 25.860 210.560 29.260 ;
        RECT 211.260 28.920 212.400 39.850 ;
        RECT 213.100 31.640 214.240 39.850 ;
        RECT 214.940 31.640 216.080 39.850 ;
        RECT 213.100 28.920 216.080 31.640 ;
        RECT 211.260 25.860 216.080 28.920 ;
        RECT 204.360 23.480 216.080 25.860 ;
        RECT 216.780 26.540 217.920 39.850 ;
        RECT 218.620 28.580 219.760 39.850 ;
        RECT 220.460 28.580 221.600 39.850 ;
        RECT 218.620 26.540 221.600 28.580 ;
        RECT 216.780 23.480 221.600 26.540 ;
        RECT 204.360 20.420 221.600 23.480 ;
        RECT 204.360 20.080 222.080 20.420 ;
        RECT 0.560 6.780 222.080 20.080 ;
        RECT 0.560 6.440 27.480 6.780 ;
        RECT 0.560 4.090 5.400 6.440 ;
        RECT 6.100 4.090 16.440 6.440 ;
        RECT 17.140 4.090 27.480 6.440 ;
        RECT 28.180 4.090 38.520 6.780 ;
        RECT 39.220 4.090 50.020 6.780 ;
        RECT 50.720 4.090 61.060 6.780 ;
        RECT 61.760 4.090 72.100 6.780 ;
        RECT 72.800 4.090 83.140 6.780 ;
        RECT 83.840 4.090 94.640 6.780 ;
        RECT 95.340 4.090 105.680 6.780 ;
        RECT 106.380 4.090 116.720 6.780 ;
        RECT 117.420 4.090 127.760 6.780 ;
        RECT 128.460 4.090 139.260 6.780 ;
        RECT 139.960 4.090 150.300 6.780 ;
        RECT 151.000 4.090 161.340 6.780 ;
        RECT 162.040 4.090 172.380 6.780 ;
        RECT 173.080 4.090 183.880 6.780 ;
        RECT 184.580 4.090 194.920 6.780 ;
        RECT 195.620 4.090 205.960 6.780 ;
        RECT 206.660 4.090 217.000 6.780 ;
        RECT 217.700 4.090 222.080 6.780 ;
      LAYER met3 ;
        RECT 40.090 5.275 199.115 32.805 ;
  END
END S_term_single
MACRO S_term_single2
  CLASS BLOCK ;
  FOREIGN S_term_single2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 235.000 BY 40.000 ;
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.680 0.000 5.820 6.160 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.980 0.000 123.120 6.500 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.940 0.000 135.080 6.500 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.440 0.000 146.580 1.090 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.400 0.000 158.540 6.500 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.900 0.000 170.040 6.500 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.860 0.000 182.000 6.500 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.360 0.000 193.500 1.090 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.320 0.000 205.460 6.500 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.820 0.000 216.960 9.220 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.780 0.000 228.920 15.000 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.180 0.000 17.320 6.500 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.140 0.000 29.280 6.500 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.640 0.000 40.780 6.500 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.600 0.000 52.740 6.500 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.100 0.000 64.240 6.500 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.060 0.000 76.200 6.700 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.560 0.000 87.700 3.810 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.520 0.000 99.660 5.170 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.020 0.000 111.160 6.500 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.960 32.260 198.100 40.000 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.820 31.920 216.960 40.000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.660 31.920 218.800 40.000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.960 29.200 221.100 40.000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.800 26.480 222.940 40.000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.640 29.540 224.780 40.000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.480 32.260 226.620 40.000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.320 25.800 228.460 40.000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.160 28.860 230.300 40.000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.000 20.700 232.140 40.000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.840 23.760 233.980 40.000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.800 29.200 199.940 40.000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.640 31.920 201.780 40.000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.480 29.200 203.620 40.000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.780 26.480 205.920 40.000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.620 26.480 207.760 40.000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.460 23.760 209.600 40.000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.300 26.820 211.440 40.000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.140 23.760 213.280 40.000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.980 23.760 215.120 40.000 ;
    END
  END FrameStrobe_O[9]
  PIN N1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.080 31.920 1.220 40.000 ;
    END
  END N1BEG[0]
  PIN N1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.920 29.200 3.060 40.000 ;
    END
  END N1BEG[1]
  PIN N1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.760 32.260 4.900 40.000 ;
    END
  END N1BEG[2]
  PIN N1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.600 29.510 6.740 40.000 ;
    END
  END N1BEG[3]
  PIN N2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.440 31.920 8.580 40.000 ;
    END
  END N2BEG[0]
  PIN N2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.280 29.200 10.420 40.000 ;
    END
  END N2BEG[1]
  PIN N2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.120 39.030 12.260 40.000 ;
    END
  END N2BEG[2]
  PIN N2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.960 32.910 14.100 40.000 ;
    END
  END N2BEG[3]
  PIN N2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.800 29.200 15.940 40.000 ;
    END
  END N2BEG[4]
  PIN N2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.100 29.540 18.240 40.000 ;
    END
  END N2BEG[5]
  PIN N2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.940 32.230 20.080 40.000 ;
    END
  END N2BEG[6]
  PIN N2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.780 28.860 21.920 40.000 ;
    END
  END N2BEG[7]
  PIN N2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.620 31.240 23.760 40.000 ;
    END
  END N2BEGb[0]
  PIN N2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.460 29.200 25.600 40.000 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.300 33.590 27.440 40.000 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.140 29.540 29.280 40.000 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.980 34.950 31.120 40.000 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.280 29.200 33.420 40.000 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.120 26.480 35.260 40.000 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.960 31.240 37.100 40.000 ;
    END
  END N2BEGb[7]
  PIN N4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.800 26.480 38.940 40.000 ;
    END
  END N4BEG[0]
  PIN N4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.660 31.920 57.800 40.000 ;
    END
  END N4BEG[10]
  PIN N4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.500 31.920 59.640 40.000 ;
    END
  END N4BEG[11]
  PIN N4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.340 31.240 61.480 40.000 ;
    END
  END N4BEG[12]
  PIN N4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.180 29.200 63.320 40.000 ;
    END
  END N4BEG[13]
  PIN N4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.480 31.920 65.620 40.000 ;
    END
  END N4BEG[14]
  PIN N4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.320 29.200 67.460 40.000 ;
    END
  END N4BEG[15]
  PIN N4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.640 29.200 40.780 40.000 ;
    END
  END N4BEG[1]
  PIN N4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.480 32.260 42.620 40.000 ;
    END
  END N4BEG[2]
  PIN N4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.320 28.520 44.460 40.000 ;
    END
  END N4BEG[3]
  PIN N4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.160 31.240 46.300 40.000 ;
    END
  END N4BEG[4]
  PIN N4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.460 29.540 48.600 40.000 ;
    END
  END N4BEG[5]
  PIN N4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.300 26.480 50.440 40.000 ;
    END
  END N4BEG[6]
  PIN N4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.140 29.200 52.280 40.000 ;
    END
  END N4BEG[7]
  PIN N4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.980 29.540 54.120 40.000 ;
    END
  END N4BEG[8]
  PIN N4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.820 26.480 55.960 40.000 ;
    END
  END N4BEG[9]
  PIN NN4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.160 32.260 69.300 40.000 ;
    END
  END NN4BEG[0]
  PIN NN4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.020 31.920 88.160 40.000 ;
    END
  END NN4BEG[10]
  PIN NN4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.860 31.920 90.000 40.000 ;
    END
  END NN4BEG[11]
  PIN NN4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.700 29.200 91.840 40.000 ;
    END
  END NN4BEG[12]
  PIN NN4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.540 29.200 93.680 40.000 ;
    END
  END NN4BEG[13]
  PIN NN4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.840 29.540 95.980 40.000 ;
    END
  END NN4BEG[14]
  PIN NN4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.680 26.480 97.820 40.000 ;
    END
  END NN4BEG[15]
  PIN NN4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.000 29.200 71.140 40.000 ;
    END
  END NN4BEG[1]
  PIN NN4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.840 31.920 72.980 40.000 ;
    END
  END NN4BEG[2]
  PIN NN4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.680 29.200 74.820 40.000 ;
    END
  END NN4BEG[3]
  PIN NN4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.520 32.260 76.660 40.000 ;
    END
  END NN4BEG[4]
  PIN NN4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.360 32.060 78.500 40.000 ;
    END
  END NN4BEG[5]
  PIN NN4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.660 39.030 80.800 40.000 ;
    END
  END NN4BEG[6]
  PIN NN4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.500 28.830 82.640 40.000 ;
    END
  END NN4BEG[7]
  PIN NN4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.340 26.820 84.480 40.000 ;
    END
  END NN4BEG[8]
  PIN NN4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.180 26.480 86.320 40.000 ;
    END
  END NN4BEG[9]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.520 39.030 99.660 40.000 ;
    END
  END S1END[0]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.360 31.580 101.500 40.000 ;
    END
  END S1END[1]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.200 28.860 103.340 40.000 ;
    END
  END S1END[2]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.040 23.080 105.180 40.000 ;
    END
  END S1END[3]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.880 22.880 107.020 40.000 ;
    END
  END S2END[0]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.720 26.140 108.860 40.000 ;
    END
  END S2END[1]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.020 23.080 111.160 40.000 ;
    END
  END S2END[2]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.860 26.280 113.000 40.000 ;
    END
  END S2END[3]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.700 26.480 114.840 40.000 ;
    END
  END S2END[4]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.540 31.550 116.680 40.000 ;
    END
  END S2END[5]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.380 32.910 118.520 40.000 ;
    END
  END S2END[6]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.220 23.080 120.360 40.000 ;
    END
  END S2END[7]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.060 26.480 122.200 40.000 ;
    END
  END S2MID[0]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.900 23.080 124.040 40.000 ;
    END
  END S2MID[1]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.740 26.480 125.880 40.000 ;
    END
  END S2MID[2]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.040 23.080 128.180 40.000 ;
    END
  END S2MID[3]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.880 23.080 130.020 40.000 ;
    END
  END S2MID[4]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.720 32.910 131.860 40.000 ;
    END
  END S2MID[5]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.560 29.540 133.700 40.000 ;
    END
  END S2MID[6]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.400 26.480 135.540 40.000 ;
    END
  END S2MID[7]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.240 25.800 137.380 40.000 ;
    END
  END S4END[0]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.100 26.140 156.240 40.000 ;
    END
  END S4END[10]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.400 26.140 158.540 40.000 ;
    END
  END S4END[11]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.240 26.480 160.380 40.000 ;
    END
  END S4END[12]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.080 28.520 162.220 40.000 ;
    END
  END S4END[13]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.920 39.030 164.060 40.000 ;
    END
  END S4END[14]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.760 26.480 165.900 40.000 ;
    END
  END S4END[15]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.080 23.080 139.220 40.000 ;
    END
  END S4END[1]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.920 26.480 141.060 40.000 ;
    END
  END S4END[2]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.220 25.800 143.360 40.000 ;
    END
  END S4END[3]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.060 23.080 145.200 40.000 ;
    END
  END S4END[4]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.900 32.910 147.040 40.000 ;
    END
  END S4END[5]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.740 32.230 148.880 40.000 ;
    END
  END S4END[6]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.580 23.420 150.720 40.000 ;
    END
  END S4END[7]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.420 30.190 152.560 40.000 ;
    END
  END S4END[8]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.260 33.620 154.400 40.000 ;
    END
  END S4END[9]
  PIN SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.600 28.860 167.740 40.000 ;
    END
  END SS4END[0]
  PIN SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.460 31.920 186.600 40.000 ;
    END
  END SS4END[10]
  PIN SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.300 31.920 188.440 40.000 ;
    END
  END SS4END[11]
  PIN SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.600 28.520 190.740 40.000 ;
    END
  END SS4END[12]
  PIN SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.440 39.030 192.580 40.000 ;
    END
  END SS4END[13]
  PIN SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.280 31.920 194.420 40.000 ;
    END
  END SS4END[14]
  PIN SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.120 28.520 196.260 40.000 ;
    END
  END SS4END[15]
  PIN SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.440 26.480 169.580 40.000 ;
    END
  END SS4END[1]
  PIN SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.280 23.080 171.420 40.000 ;
    END
  END SS4END[2]
  PIN SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.580 26.820 173.720 40.000 ;
    END
  END SS4END[3]
  PIN SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.420 31.580 175.560 40.000 ;
    END
  END SS4END[4]
  PIN SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.260 28.860 177.400 40.000 ;
    END
  END SS4END[5]
  PIN SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.100 31.240 179.240 40.000 ;
    END
  END SS4END[6]
  PIN SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.940 28.860 181.080 40.000 ;
    END
  END SS4END[7]
  PIN SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.780 26.480 182.920 40.000 ;
    END
  END SS4END[8]
  PIN SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.620 23.080 184.760 40.000 ;
    END
  END SS4END[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 42.045 5.200 43.645 32.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 116.695 5.200 118.295 32.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 191.350 5.200 192.950 32.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 79.370 5.200 80.970 32.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 154.025 5.200 155.625 32.880 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 229.080 39.695 ;
      LAYER met1 ;
        RECT 34.430 40.000 88.160 40.020 ;
        RECT 0.990 4.120 234.070 40.000 ;
      LAYER met2 ;
        RECT 1.500 31.640 2.640 39.850 ;
        RECT 1.020 28.920 2.640 31.640 ;
        RECT 3.340 31.980 4.480 39.850 ;
        RECT 5.180 31.980 6.320 39.850 ;
        RECT 3.340 29.230 6.320 31.980 ;
        RECT 7.020 31.640 8.160 39.850 ;
        RECT 8.860 31.640 10.000 39.850 ;
        RECT 7.020 29.230 10.000 31.640 ;
        RECT 3.340 28.920 10.000 29.230 ;
        RECT 10.700 38.750 11.840 39.850 ;
        RECT 12.540 38.750 13.680 39.850 ;
        RECT 10.700 32.630 13.680 38.750 ;
        RECT 14.380 32.630 15.520 39.850 ;
        RECT 10.700 28.920 15.520 32.630 ;
        RECT 16.220 29.260 17.820 39.850 ;
        RECT 18.520 31.950 19.660 39.850 ;
        RECT 20.360 31.950 21.500 39.850 ;
        RECT 18.520 29.260 21.500 31.950 ;
        RECT 16.220 28.920 21.500 29.260 ;
        RECT 1.020 28.580 21.500 28.920 ;
        RECT 22.200 30.960 23.340 39.850 ;
        RECT 24.040 30.960 25.180 39.850 ;
        RECT 22.200 28.920 25.180 30.960 ;
        RECT 25.880 33.310 27.020 39.850 ;
        RECT 27.720 33.310 28.860 39.850 ;
        RECT 25.880 29.260 28.860 33.310 ;
        RECT 29.560 34.670 30.700 39.850 ;
        RECT 31.400 34.670 33.000 39.850 ;
        RECT 29.560 29.260 33.000 34.670 ;
        RECT 25.880 28.920 33.000 29.260 ;
        RECT 33.700 28.920 34.840 39.850 ;
        RECT 22.200 28.580 34.840 28.920 ;
        RECT 1.020 26.200 34.840 28.580 ;
        RECT 35.540 30.960 36.680 39.850 ;
        RECT 37.380 30.960 38.520 39.850 ;
        RECT 35.540 26.200 38.520 30.960 ;
        RECT 39.220 28.920 40.360 39.850 ;
        RECT 41.060 31.980 42.200 39.850 ;
        RECT 42.900 31.980 44.040 39.850 ;
        RECT 41.060 28.920 44.040 31.980 ;
        RECT 39.220 28.240 44.040 28.920 ;
        RECT 44.740 30.960 45.880 39.850 ;
        RECT 46.580 30.960 48.180 39.850 ;
        RECT 44.740 29.260 48.180 30.960 ;
        RECT 48.880 29.260 50.020 39.850 ;
        RECT 44.740 28.240 50.020 29.260 ;
        RECT 39.220 26.200 50.020 28.240 ;
        RECT 50.720 28.920 51.860 39.850 ;
        RECT 52.560 29.260 53.700 39.850 ;
        RECT 54.400 29.260 55.540 39.850 ;
        RECT 52.560 28.920 55.540 29.260 ;
        RECT 50.720 26.200 55.540 28.920 ;
        RECT 56.240 31.640 57.380 39.850 ;
        RECT 58.080 31.640 59.220 39.850 ;
        RECT 59.920 31.640 61.060 39.850 ;
        RECT 56.240 30.960 61.060 31.640 ;
        RECT 61.760 30.960 62.900 39.850 ;
        RECT 56.240 28.920 62.900 30.960 ;
        RECT 63.600 31.640 65.200 39.850 ;
        RECT 65.900 31.640 67.040 39.850 ;
        RECT 63.600 28.920 67.040 31.640 ;
        RECT 67.740 31.980 68.880 39.850 ;
        RECT 69.580 31.980 70.720 39.850 ;
        RECT 67.740 28.920 70.720 31.980 ;
        RECT 71.420 31.640 72.560 39.850 ;
        RECT 73.260 31.640 74.400 39.850 ;
        RECT 71.420 28.920 74.400 31.640 ;
        RECT 75.100 31.980 76.240 39.850 ;
        RECT 76.940 31.980 78.080 39.850 ;
        RECT 75.100 31.780 78.080 31.980 ;
        RECT 78.780 38.750 80.380 39.850 ;
        RECT 81.080 38.750 82.220 39.850 ;
        RECT 78.780 31.780 82.220 38.750 ;
        RECT 75.100 28.920 82.220 31.780 ;
        RECT 56.240 28.550 82.220 28.920 ;
        RECT 82.920 28.550 84.060 39.850 ;
        RECT 56.240 26.540 84.060 28.550 ;
        RECT 84.760 26.540 85.900 39.850 ;
        RECT 56.240 26.200 85.900 26.540 ;
        RECT 86.600 31.640 87.740 39.850 ;
        RECT 88.440 31.640 89.580 39.850 ;
        RECT 90.280 31.640 91.420 39.850 ;
        RECT 86.600 28.920 91.420 31.640 ;
        RECT 92.120 28.920 93.260 39.850 ;
        RECT 93.960 29.260 95.560 39.850 ;
        RECT 96.260 29.260 97.400 39.850 ;
        RECT 93.960 28.920 97.400 29.260 ;
        RECT 86.600 26.200 97.400 28.920 ;
        RECT 98.100 38.750 99.240 39.850 ;
        RECT 99.940 38.750 101.080 39.850 ;
        RECT 98.100 31.300 101.080 38.750 ;
        RECT 101.780 31.300 102.920 39.850 ;
        RECT 98.100 28.580 102.920 31.300 ;
        RECT 103.620 28.580 104.760 39.850 ;
        RECT 98.100 26.200 104.760 28.580 ;
        RECT 1.020 22.800 104.760 26.200 ;
        RECT 105.460 22.800 106.600 39.850 ;
        RECT 1.020 22.600 106.600 22.800 ;
        RECT 107.300 25.860 108.440 39.850 ;
        RECT 109.140 25.860 110.740 39.850 ;
        RECT 107.300 22.800 110.740 25.860 ;
        RECT 111.440 26.000 112.580 39.850 ;
        RECT 113.280 26.200 114.420 39.850 ;
        RECT 115.120 31.270 116.260 39.850 ;
        RECT 116.960 32.630 118.100 39.850 ;
        RECT 118.800 32.630 119.940 39.850 ;
        RECT 116.960 31.270 119.940 32.630 ;
        RECT 115.120 26.200 119.940 31.270 ;
        RECT 113.280 26.000 119.940 26.200 ;
        RECT 111.440 22.800 119.940 26.000 ;
        RECT 120.640 26.200 121.780 39.850 ;
        RECT 122.480 26.200 123.620 39.850 ;
        RECT 120.640 22.800 123.620 26.200 ;
        RECT 124.320 26.200 125.460 39.850 ;
        RECT 126.160 26.200 127.760 39.850 ;
        RECT 124.320 22.800 127.760 26.200 ;
        RECT 128.460 22.800 129.600 39.850 ;
        RECT 130.300 32.630 131.440 39.850 ;
        RECT 132.140 32.630 133.280 39.850 ;
        RECT 130.300 29.260 133.280 32.630 ;
        RECT 133.980 29.260 135.120 39.850 ;
        RECT 130.300 26.200 135.120 29.260 ;
        RECT 135.820 26.200 136.960 39.850 ;
        RECT 130.300 25.520 136.960 26.200 ;
        RECT 137.660 25.520 138.800 39.850 ;
        RECT 130.300 22.800 138.800 25.520 ;
        RECT 139.500 26.200 140.640 39.850 ;
        RECT 141.340 26.200 142.940 39.850 ;
        RECT 139.500 25.520 142.940 26.200 ;
        RECT 143.640 25.520 144.780 39.850 ;
        RECT 139.500 22.800 144.780 25.520 ;
        RECT 145.480 32.630 146.620 39.850 ;
        RECT 147.320 32.630 148.460 39.850 ;
        RECT 145.480 31.950 148.460 32.630 ;
        RECT 149.160 31.950 150.300 39.850 ;
        RECT 145.480 23.140 150.300 31.950 ;
        RECT 151.000 29.910 152.140 39.850 ;
        RECT 152.840 33.340 153.980 39.850 ;
        RECT 154.680 33.340 155.820 39.850 ;
        RECT 152.840 29.910 155.820 33.340 ;
        RECT 151.000 25.860 155.820 29.910 ;
        RECT 156.520 25.860 158.120 39.850 ;
        RECT 158.820 26.200 159.960 39.850 ;
        RECT 160.660 28.240 161.800 39.850 ;
        RECT 162.500 38.750 163.640 39.850 ;
        RECT 164.340 38.750 165.480 39.850 ;
        RECT 162.500 28.240 165.480 38.750 ;
        RECT 160.660 26.200 165.480 28.240 ;
        RECT 166.180 28.580 167.320 39.850 ;
        RECT 168.020 28.580 169.160 39.850 ;
        RECT 166.180 26.200 169.160 28.580 ;
        RECT 169.860 26.200 171.000 39.850 ;
        RECT 158.820 25.860 171.000 26.200 ;
        RECT 151.000 23.140 171.000 25.860 ;
        RECT 145.480 22.800 171.000 23.140 ;
        RECT 171.700 26.540 173.300 39.850 ;
        RECT 174.000 31.300 175.140 39.850 ;
        RECT 175.840 31.300 176.980 39.850 ;
        RECT 174.000 28.580 176.980 31.300 ;
        RECT 177.680 30.960 178.820 39.850 ;
        RECT 179.520 30.960 180.660 39.850 ;
        RECT 177.680 28.580 180.660 30.960 ;
        RECT 181.360 28.580 182.500 39.850 ;
        RECT 174.000 26.540 182.500 28.580 ;
        RECT 171.700 26.200 182.500 26.540 ;
        RECT 183.200 26.200 184.340 39.850 ;
        RECT 171.700 22.800 184.340 26.200 ;
        RECT 185.040 31.640 186.180 39.850 ;
        RECT 186.880 31.640 188.020 39.850 ;
        RECT 188.720 31.640 190.320 39.850 ;
        RECT 185.040 28.240 190.320 31.640 ;
        RECT 191.020 38.750 192.160 39.850 ;
        RECT 192.860 38.750 194.000 39.850 ;
        RECT 191.020 31.640 194.000 38.750 ;
        RECT 194.700 31.640 195.840 39.850 ;
        RECT 191.020 28.240 195.840 31.640 ;
        RECT 196.540 31.980 197.680 39.850 ;
        RECT 198.380 31.980 199.520 39.850 ;
        RECT 196.540 28.920 199.520 31.980 ;
        RECT 200.220 31.640 201.360 39.850 ;
        RECT 202.060 31.640 203.200 39.850 ;
        RECT 200.220 28.920 203.200 31.640 ;
        RECT 203.900 28.920 205.500 39.850 ;
        RECT 196.540 28.240 205.500 28.920 ;
        RECT 185.040 26.200 205.500 28.240 ;
        RECT 206.200 26.200 207.340 39.850 ;
        RECT 208.040 26.200 209.180 39.850 ;
        RECT 185.040 23.480 209.180 26.200 ;
        RECT 209.880 26.540 211.020 39.850 ;
        RECT 211.720 26.540 212.860 39.850 ;
        RECT 209.880 23.480 212.860 26.540 ;
        RECT 213.560 23.480 214.700 39.850 ;
        RECT 215.400 31.640 216.540 39.850 ;
        RECT 217.240 31.640 218.380 39.850 ;
        RECT 219.080 31.640 220.680 39.850 ;
        RECT 215.400 28.920 220.680 31.640 ;
        RECT 221.380 28.920 222.520 39.850 ;
        RECT 215.400 26.200 222.520 28.920 ;
        RECT 223.220 29.260 224.360 39.850 ;
        RECT 225.060 31.980 226.200 39.850 ;
        RECT 226.900 31.980 228.040 39.850 ;
        RECT 225.060 29.260 228.040 31.980 ;
        RECT 223.220 26.200 228.040 29.260 ;
        RECT 215.400 25.520 228.040 26.200 ;
        RECT 228.740 28.580 229.880 39.850 ;
        RECT 230.580 28.580 231.720 39.850 ;
        RECT 228.740 25.520 231.720 28.580 ;
        RECT 215.400 23.480 231.720 25.520 ;
        RECT 185.040 22.800 231.720 23.480 ;
        RECT 107.300 22.600 231.720 22.800 ;
        RECT 1.020 20.420 231.720 22.600 ;
        RECT 232.420 23.480 233.560 39.850 ;
        RECT 232.420 20.420 234.040 23.480 ;
        RECT 1.020 15.280 234.040 20.420 ;
        RECT 1.020 9.500 228.500 15.280 ;
        RECT 1.020 6.980 216.540 9.500 ;
        RECT 1.020 6.780 75.780 6.980 ;
        RECT 1.020 6.440 16.900 6.780 ;
        RECT 1.020 0.270 5.400 6.440 ;
        RECT 6.100 0.270 16.900 6.440 ;
        RECT 17.600 0.270 28.860 6.780 ;
        RECT 29.560 0.270 40.360 6.780 ;
        RECT 41.060 0.270 52.320 6.780 ;
        RECT 53.020 0.270 63.820 6.780 ;
        RECT 64.520 0.270 75.780 6.780 ;
        RECT 76.480 6.780 216.540 6.980 ;
        RECT 76.480 5.450 110.740 6.780 ;
        RECT 76.480 4.090 99.240 5.450 ;
        RECT 76.480 0.270 87.280 4.090 ;
        RECT 87.980 0.270 99.240 4.090 ;
        RECT 99.940 0.270 110.740 5.450 ;
        RECT 111.440 0.270 122.700 6.780 ;
        RECT 123.400 0.270 134.660 6.780 ;
        RECT 135.360 1.370 158.120 6.780 ;
        RECT 135.360 0.270 146.160 1.370 ;
        RECT 146.860 0.270 158.120 1.370 ;
        RECT 158.820 0.270 169.620 6.780 ;
        RECT 170.320 0.270 181.580 6.780 ;
        RECT 182.280 1.370 205.040 6.780 ;
        RECT 182.280 0.270 193.080 1.370 ;
        RECT 193.780 0.270 205.040 1.370 ;
        RECT 205.740 0.270 216.540 6.780 ;
        RECT 217.240 0.270 228.500 9.500 ;
        RECT 229.200 0.270 234.040 15.280 ;
      LAYER met3 ;
        RECT 40.085 5.275 199.575 38.585 ;
  END
END S_term_single2
MACRO W_IO
  CLASS BLOCK ;
  FOREIGN W_IO ;
  ORIGIN 0.000 0.000 ;
  SIZE 80.000 BY 223.115 ;
  PIN A_I_top
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.750 9.750 46.050 ;
    END
  END A_I_top
  PIN A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.550 6.990 35.850 ;
    END
  END A_O_top
  PIN A_T_top
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.990 10.210 41.290 ;
    END
  END A_T_top
  PIN A_config_C_bit0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.510 9.750 50.810 ;
    END
  END A_config_C_bit0
  PIN A_config_C_bit1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.270 10.210 55.570 ;
    END
  END A_config_C_bit1
  PIN A_config_C_bit2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.030 9.750 60.330 ;
    END
  END A_config_C_bit2
  PIN A_config_C_bit3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.790 13.890 65.090 ;
    END
  END A_config_C_bit3
  PIN B_I_top
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.750 9.750 12.050 ;
    END
  END B_I_top
  PIN B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.230 9.290 2.530 ;
    END
  END B_O_top
  PIN B_T_top
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.990 14.350 7.290 ;
    END
  END B_T_top
  PIN B_config_C_bit0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.510 9.750 16.810 ;
    END
  END B_config_C_bit0
  PIN B_config_C_bit1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.270 13.890 21.570 ;
    END
  END B_config_C_bit1
  PIN B_config_C_bit2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.030 9.750 26.330 ;
    END
  END B_config_C_bit2
  PIN B_config_C_bit3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.790 10.210 31.090 ;
    END
  END B_config_C_bit3
  PIN E1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.460 84.510 80.000 84.810 ;
    END
  END E1BEG[0]
  PIN E1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 57.870 85.870 80.000 86.170 ;
    END
  END E1BEG[1]
  PIN E1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 59.500 87.910 80.000 88.210 ;
    END
  END E1BEG[2]
  PIN E1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.750 89.270 80.000 89.570 ;
    END
  END E1BEG[3]
  PIN E2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 60.170 91.310 80.000 91.610 ;
    END
  END E2BEG[0]
  PIN E2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.950 92.670 80.000 92.970 ;
    END
  END E2BEG[1]
  PIN E2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 72.070 94.710 80.000 95.010 ;
    END
  END E2BEG[2]
  PIN E2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 68.910 96.070 80.000 96.370 ;
    END
  END E2BEG[3]
  PIN E2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 61.950 98.110 80.000 98.410 ;
    END
  END E2BEG[4]
  PIN E2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 78.570 100.150 80.000 100.450 ;
    END
  END E2BEG[5]
  PIN E2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 61.090 101.510 80.000 101.810 ;
    END
  END E2BEG[6]
  PIN E2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.810 103.550 80.000 103.850 ;
    END
  END E2BEG[7]
  PIN E2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 73.510 104.910 80.000 105.210 ;
    END
  END E2BEGb[0]
  PIN E2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 55.570 106.950 80.000 107.250 ;
    END
  END E2BEGb[1]
  PIN E2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 66.150 108.310 80.000 108.610 ;
    END
  END E2BEGb[2]
  PIN E2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 55.570 110.350 80.000 110.650 ;
    END
  END E2BEGb[3]
  PIN E2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 60.630 112.390 80.000 112.690 ;
    END
  END E2BEGb[4]
  PIN E2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 61.090 113.750 80.000 114.050 ;
    END
  END E2BEGb[5]
  PIN E2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 59.250 115.790 80.000 116.090 ;
    END
  END E2BEGb[6]
  PIN E2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.150 117.150 80.000 117.450 ;
    END
  END E2BEGb[7]
  PIN E6BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 60.630 147.070 80.000 147.370 ;
    END
  END E6BEG[0]
  PIN E6BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.290 164.070 80.000 164.370 ;
    END
  END E6BEG[10]
  PIN E6BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.350 166.110 80.000 166.410 ;
    END
  END E6BEG[11]
  PIN E6BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 67.990 148.430 80.000 148.730 ;
    END
  END E6BEG[1]
  PIN E6BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 58.330 150.470 80.000 150.770 ;
    END
  END E6BEG[2]
  PIN E6BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 55.570 151.830 80.000 152.130 ;
    END
  END E6BEG[3]
  PIN E6BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 58.330 153.870 80.000 154.170 ;
    END
  END E6BEG[4]
  PIN E6BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 61.950 155.910 80.000 156.210 ;
    END
  END E6BEG[5]
  PIN E6BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 58.330 157.270 80.000 157.570 ;
    END
  END E6BEG[6]
  PIN E6BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.490 159.310 80.000 159.610 ;
    END
  END E6BEG[7]
  PIN E6BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 68.910 160.670 80.000 160.970 ;
    END
  END E6BEG[8]
  PIN E6BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.810 162.710 80.000 163.010 ;
    END
  END E6BEG[9]
  PIN EE4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 57.410 119.190 80.000 119.490 ;
    END
  END EE4BEG[0]
  PIN EE4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 60.630 136.190 80.000 136.490 ;
    END
  END EE4BEG[10]
  PIN EE4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.150 138.230 80.000 138.530 ;
    END
  END EE4BEG[11]
  PIN EE4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 59.250 140.270 80.000 140.570 ;
    END
  END EE4BEG[12]
  PIN EE4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 60.630 141.630 80.000 141.930 ;
    END
  END EE4BEG[13]
  PIN EE4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.290 143.670 80.000 143.970 ;
    END
  END EE4BEG[14]
  PIN EE4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 61.950 145.030 80.000 145.330 ;
    END
  END EE4BEG[15]
  PIN EE4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 55.570 120.550 80.000 120.850 ;
    END
  END EE4BEG[1]
  PIN EE4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.150 122.590 80.000 122.890 ;
    END
  END EE4BEG[2]
  PIN EE4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.490 123.950 80.000 124.250 ;
    END
  END EE4BEG[3]
  PIN EE4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 61.950 125.990 80.000 126.290 ;
    END
  END EE4BEG[4]
  PIN EE4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.150 128.030 80.000 128.330 ;
    END
  END EE4BEG[5]
  PIN EE4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 55.570 129.390 80.000 129.690 ;
    END
  END EE4BEG[6]
  PIN EE4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.150 131.430 80.000 131.730 ;
    END
  END EE4BEG[7]
  PIN EE4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.150 132.790 80.000 133.090 ;
    END
  END EE4BEG[8]
  PIN EE4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.030 134.830 80.000 135.130 ;
    END
  END EE4BEG[9]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.550 6.990 69.850 ;
    END
  END FrameData[0]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.510 6.990 118.810 ;
    END
  END FrameData[10]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.270 6.990 123.570 ;
    END
  END FrameData[11]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.030 9.290 128.330 ;
    END
  END FrameData[12]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.790 9.290 133.090 ;
    END
  END FrameData[13]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.550 9.290 137.850 ;
    END
  END FrameData[14]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.310 9.290 142.610 ;
    END
  END FrameData[15]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.070 9.290 147.370 ;
    END
  END FrameData[16]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.510 6.990 152.810 ;
    END
  END FrameData[17]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.270 6.990 157.570 ;
    END
  END FrameData[18]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.030 6.990 162.330 ;
    END
  END FrameData[19]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.310 6.990 74.610 ;
    END
  END FrameData[1]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.790 6.990 167.090 ;
    END
  END FrameData[20]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.550 6.990 171.850 ;
    END
  END FrameData[21]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.310 9.290 176.610 ;
    END
  END FrameData[22]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 181.070 9.290 181.370 ;
    END
  END FrameData[23]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.830 6.990 186.130 ;
    END
  END FrameData[24]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.270 6.990 191.570 ;
    END
  END FrameData[25]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.030 9.290 196.330 ;
    END
  END FrameData[26]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.790 9.290 201.090 ;
    END
  END FrameData[27]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.550 9.290 205.850 ;
    END
  END FrameData[28]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.310 6.990 210.610 ;
    END
  END FrameData[29]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.750 6.990 80.050 ;
    END
  END FrameData[2]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.070 9.290 215.370 ;
    END
  END FrameData[30]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.830 8.830 220.130 ;
    END
  END FrameData[31]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.510 9.290 84.810 ;
    END
  END FrameData[3]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.270 9.290 89.570 ;
    END
  END FrameData[4]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.030 6.990 94.330 ;
    END
  END FrameData[5]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.790 9.290 99.090 ;
    END
  END FrameData[6]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.550 9.290 103.850 ;
    END
  END FrameData[7]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.310 9.290 108.610 ;
    END
  END FrameData[8]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.750 6.990 114.050 ;
    END
  END FrameData[9]
  PIN FrameData_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 67.990 168.150 80.000 168.450 ;
    END
  END FrameData_O[0]
  PIN FrameData_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.750 185.150 80.000 185.450 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.750 187.190 80.000 187.490 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 67.070 188.550 80.000 188.850 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.290 190.590 80.000 190.890 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.750 191.950 80.000 192.250 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 67.530 193.990 80.000 194.290 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 66.610 196.030 80.000 196.330 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.290 197.390 80.000 197.690 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 67.990 199.430 80.000 199.730 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 66.610 200.790 80.000 201.090 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 68.910 169.510 80.000 169.810 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.890 202.830 80.000 203.130 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 67.990 204.190 80.000 204.490 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 67.070 206.230 80.000 206.530 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.310 207.590 80.000 207.890 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 67.530 209.630 80.000 209.930 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 67.990 211.670 80.000 211.970 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.310 213.030 80.000 213.330 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 67.070 215.070 80.000 215.370 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 60.630 216.430 80.000 216.730 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 61.090 218.470 80.000 218.770 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.150 171.550 80.000 171.850 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 62.010 219.830 80.000 220.130 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.950 221.870 80.000 222.170 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 68.910 172.910 80.000 173.210 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 68.450 174.950 80.000 175.250 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 67.990 176.310 80.000 176.610 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 59.710 178.350 80.000 178.650 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 58.330 179.710 80.000 180.010 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 68.910 181.750 80.000 182.050 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 57.870 183.790 80.000 184.090 ;
    END
  END FrameData_O[9]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.000 0.000 2.140 9.560 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.020 0.000 42.160 1.090 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.700 0.000 45.840 6.840 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.840 0.000 49.980 2.420 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.980 0.000 54.120 7.520 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.660 0.000 57.800 3.440 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.800 0.000 61.940 1.090 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.940 0.000 66.080 11.260 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.620 0.000 69.760 5.170 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.760 0.000 73.900 9.900 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.900 0.000 78.040 15.680 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.680 0.000 5.820 6.160 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.820 0.000 9.960 6.500 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.960 0.000 14.100 9.560 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.640 0.000 17.780 6.530 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.780 0.000 21.920 9.560 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.920 0.000 26.060 17.380 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.600 0.000 29.740 20.440 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.740 0.000 33.880 14.660 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.880 0.000 38.020 16.700 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.000 217.220 2.140 223.115 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.720 216.880 39.860 223.115 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.860 217.220 44.000 223.115 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.540 213.790 47.680 223.115 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.220 221.950 51.360 223.115 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.360 211.440 55.500 223.115 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.040 209.060 59.180 223.115 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.720 221.950 62.860 223.115 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.400 210.760 66.540 223.115 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.540 201.920 70.680 223.115 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.220 210.080 74.360 223.115 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.680 213.820 5.820 223.115 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.360 217.190 9.500 223.115 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.040 216.880 13.180 223.115 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.180 221.950 17.320 223.115 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.860 217.220 21.000 223.115 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.540 216.880 24.680 223.115 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.680 221.950 28.820 223.115 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.360 221.950 32.500 223.115 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.040 213.820 36.180 223.115 ;
    END
  END FrameStrobe_O[9]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.900 200.560 78.040 223.115 ;
    END
  END UserCLK
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 27.705 5.200 29.305 217.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.690 5.200 52.290 217.840 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 16.215 5.200 17.815 217.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 39.200 5.200 40.800 217.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 62.185 5.200 63.785 217.840 ;
    END
  END VPWR
  PIN W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.030 0.870 80.000 1.170 ;
    END
  END W1END[0]
  PIN W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 55.570 2.230 80.000 2.530 ;
    END
  END W1END[1]
  PIN W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.950 4.270 80.000 4.570 ;
    END
  END W1END[2]
  PIN W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 57.410 5.630 80.000 5.930 ;
    END
  END W1END[3]
  PIN W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 68.910 21.270 80.000 21.570 ;
    END
  END W2END[0]
  PIN W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.890 23.310 80.000 23.610 ;
    END
  END W2END[1]
  PIN W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 76.670 24.670 80.000 24.970 ;
    END
  END W2END[2]
  PIN W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 60.170 26.710 80.000 27.010 ;
    END
  END W2END[3]
  PIN W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.030 28.750 80.000 29.050 ;
    END
  END W2END[4]
  PIN W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 76.670 30.110 80.000 30.410 ;
    END
  END W2END[5]
  PIN W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 55.570 32.150 80.000 32.450 ;
    END
  END W2END[6]
  PIN W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 59.250 33.510 80.000 33.810 ;
    END
  END W2END[7]
  PIN W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 68.910 7.670 80.000 7.970 ;
    END
  END W2MID[0]
  PIN W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 51.890 9.030 80.000 9.330 ;
    END
  END W2MID[1]
  PIN W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.490 11.070 80.000 11.370 ;
    END
  END W2MID[2]
  PIN W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 55.110 12.430 80.000 12.730 ;
    END
  END W2MID[3]
  PIN W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 68.910 14.470 80.000 14.770 ;
    END
  END W2MID[4]
  PIN W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.030 16.510 80.000 16.810 ;
    END
  END W2MID[5]
  PIN W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 68.450 17.870 80.000 18.170 ;
    END
  END W2MID[6]
  PIN W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 58.790 19.910 80.000 20.210 ;
    END
  END W2MID[7]
  PIN W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 62.010 63.430 80.000 63.730 ;
    END
  END W6END[0]
  PIN W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 59.710 80.430 80.000 80.730 ;
    END
  END W6END[10]
  PIN W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 55.570 82.470 80.000 82.770 ;
    END
  END W6END[11]
  PIN W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 66.610 64.790 80.000 65.090 ;
    END
  END W6END[1]
  PIN W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 57.870 66.830 80.000 67.130 ;
    END
  END W6END[2]
  PIN W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 66.150 68.190 80.000 68.490 ;
    END
  END W6END[3]
  PIN W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 58.330 70.230 80.000 70.530 ;
    END
  END W6END[4]
  PIN W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 57.410 72.270 80.000 72.570 ;
    END
  END W6END[5]
  PIN W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.460 73.630 80.000 73.930 ;
    END
  END W6END[6]
  PIN W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 54.650 75.670 80.000 75.970 ;
    END
  END W6END[7]
  PIN W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.950 77.030 80.000 77.330 ;
    END
  END W6END[8]
  PIN W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.460 79.070 80.000 79.370 ;
    END
  END W6END[9]
  PIN WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.150 35.550 80.000 35.850 ;
    END
  END WW4END[0]
  PIN WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 55.570 52.550 80.000 52.850 ;
    END
  END WW4END[10]
  PIN WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 58.040 54.590 80.000 54.890 ;
    END
  END WW4END[11]
  PIN WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 65.630 56.630 80.000 56.930 ;
    END
  END WW4END[12]
  PIN WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 67.070 57.990 80.000 58.290 ;
    END
  END WW4END[13]
  PIN WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 57.410 60.030 80.000 60.330 ;
    END
  END WW4END[14]
  PIN WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 61.090 61.390 80.000 61.690 ;
    END
  END WW4END[15]
  PIN WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 49.590 36.910 80.000 37.210 ;
    END
  END WW4END[1]
  PIN WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 55.570 38.950 80.000 39.250 ;
    END
  END WW4END[2]
  PIN WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.710 40.310 80.000 40.610 ;
    END
  END WW4END[3]
  PIN WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 66.610 42.350 80.000 42.650 ;
    END
  END WW4END[4]
  PIN WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 58.330 44.390 80.000 44.690 ;
    END
  END WW4END[5]
  PIN WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.150 45.750 80.000 46.050 ;
    END
  END WW4END[6]
  PIN WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 57.870 47.790 80.000 48.090 ;
    END
  END WW4END[7]
  PIN WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.030 49.150 80.000 49.450 ;
    END
  END WW4END[8]
  PIN WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 73.910 51.190 80.000 51.490 ;
    END
  END WW4END[9]
  OBS
      LAYER li1 ;
        RECT 5.520 1.445 79.895 217.685 ;
      LAYER met1 ;
        RECT 1.910 0.720 79.970 218.240 ;
      LAYER met2 ;
        RECT 2.420 216.940 5.400 222.770 ;
        RECT 1.940 213.540 5.400 216.940 ;
        RECT 6.100 216.910 9.080 222.770 ;
        RECT 9.780 216.910 12.760 222.770 ;
        RECT 6.100 216.600 12.760 216.910 ;
        RECT 13.460 221.670 16.900 222.770 ;
        RECT 17.600 221.670 20.580 222.770 ;
        RECT 13.460 216.940 20.580 221.670 ;
        RECT 21.280 216.940 24.260 222.770 ;
        RECT 13.460 216.600 24.260 216.940 ;
        RECT 24.960 221.670 28.400 222.770 ;
        RECT 29.100 221.670 32.080 222.770 ;
        RECT 32.780 221.670 35.760 222.770 ;
        RECT 24.960 216.600 35.760 221.670 ;
        RECT 6.100 213.540 35.760 216.600 ;
        RECT 36.460 216.600 39.440 222.770 ;
        RECT 40.140 216.940 43.580 222.770 ;
        RECT 44.280 216.940 47.260 222.770 ;
        RECT 40.140 216.600 47.260 216.940 ;
        RECT 36.460 213.540 47.260 216.600 ;
        RECT 1.940 213.510 47.260 213.540 ;
        RECT 47.960 221.670 50.940 222.770 ;
        RECT 51.640 221.670 55.080 222.770 ;
        RECT 47.960 213.510 55.080 221.670 ;
        RECT 1.940 211.160 55.080 213.510 ;
        RECT 55.780 211.160 58.760 222.770 ;
        RECT 1.940 208.780 58.760 211.160 ;
        RECT 59.460 221.670 62.440 222.770 ;
        RECT 63.140 221.670 66.120 222.770 ;
        RECT 59.460 210.480 66.120 221.670 ;
        RECT 66.820 210.480 70.260 222.770 ;
        RECT 59.460 208.780 70.260 210.480 ;
        RECT 1.940 201.640 70.260 208.780 ;
        RECT 70.960 209.800 73.940 222.770 ;
        RECT 74.640 209.800 77.620 222.770 ;
        RECT 70.960 201.640 77.620 209.800 ;
        RECT 1.940 200.280 77.620 201.640 ;
        RECT 78.320 200.280 79.940 222.770 ;
        RECT 1.940 20.720 79.940 200.280 ;
        RECT 1.940 17.660 29.320 20.720 ;
        RECT 1.940 9.840 25.640 17.660 ;
        RECT 2.420 6.780 13.680 9.840 ;
        RECT 2.420 6.440 9.540 6.780 ;
        RECT 2.420 0.270 5.400 6.440 ;
        RECT 6.100 0.270 9.540 6.440 ;
        RECT 10.240 0.270 13.680 6.780 ;
        RECT 14.380 6.810 21.500 9.840 ;
        RECT 14.380 0.270 17.360 6.810 ;
        RECT 18.060 0.270 21.500 6.810 ;
        RECT 22.200 0.270 25.640 9.840 ;
        RECT 26.340 0.270 29.320 17.660 ;
        RECT 30.020 16.980 79.940 20.720 ;
        RECT 30.020 14.940 37.600 16.980 ;
        RECT 30.020 0.270 33.460 14.940 ;
        RECT 34.160 0.270 37.600 14.940 ;
        RECT 38.300 15.960 79.940 16.980 ;
        RECT 38.300 11.540 77.620 15.960 ;
        RECT 38.300 7.800 65.660 11.540 ;
        RECT 38.300 7.120 53.700 7.800 ;
        RECT 38.300 1.370 45.420 7.120 ;
        RECT 38.300 0.270 41.740 1.370 ;
        RECT 42.440 0.270 45.420 1.370 ;
        RECT 46.120 2.700 53.700 7.120 ;
        RECT 46.120 0.270 49.560 2.700 ;
        RECT 50.260 0.270 53.700 2.700 ;
        RECT 54.400 3.720 65.660 7.800 ;
        RECT 54.400 0.270 57.380 3.720 ;
        RECT 58.080 1.370 65.660 3.720 ;
        RECT 58.080 0.270 61.520 1.370 ;
        RECT 62.220 0.270 65.660 1.370 ;
        RECT 66.360 10.180 77.620 11.540 ;
        RECT 66.360 5.450 73.480 10.180 ;
        RECT 66.360 0.270 69.340 5.450 ;
        RECT 70.040 0.270 73.480 5.450 ;
        RECT 74.180 0.270 77.620 10.180 ;
        RECT 78.320 0.270 79.940 15.960 ;
      LAYER met3 ;
        RECT 6.965 221.470 56.550 222.185 ;
        RECT 6.965 220.530 78.595 221.470 ;
        RECT 9.230 219.430 61.610 220.530 ;
        RECT 6.965 219.170 78.595 219.430 ;
        RECT 6.965 218.070 60.690 219.170 ;
        RECT 6.965 217.130 78.595 218.070 ;
        RECT 6.965 216.030 60.230 217.130 ;
        RECT 6.965 215.770 78.595 216.030 ;
        RECT 9.690 214.670 66.670 215.770 ;
        RECT 6.965 213.730 78.595 214.670 ;
        RECT 6.965 212.630 63.910 213.730 ;
        RECT 6.965 212.370 78.595 212.630 ;
        RECT 6.965 211.270 67.590 212.370 ;
        RECT 6.965 211.010 78.595 211.270 ;
        RECT 7.390 210.330 78.595 211.010 ;
        RECT 7.390 209.910 67.130 210.330 ;
        RECT 6.965 209.230 67.130 209.910 ;
        RECT 6.965 208.290 78.595 209.230 ;
        RECT 6.965 207.190 63.910 208.290 ;
        RECT 6.965 206.930 78.595 207.190 ;
        RECT 6.965 206.250 66.670 206.930 ;
        RECT 9.690 205.830 66.670 206.250 ;
        RECT 9.690 205.150 78.595 205.830 ;
        RECT 6.965 204.890 78.595 205.150 ;
        RECT 6.965 203.790 67.590 204.890 ;
        RECT 6.965 203.530 78.595 203.790 ;
        RECT 6.965 202.430 74.490 203.530 ;
        RECT 6.965 201.490 78.595 202.430 ;
        RECT 9.690 200.390 66.210 201.490 ;
        RECT 6.965 200.130 78.595 200.390 ;
        RECT 6.965 199.030 67.590 200.130 ;
        RECT 6.965 198.090 78.595 199.030 ;
        RECT 6.965 196.990 69.890 198.090 ;
        RECT 6.965 196.730 78.595 196.990 ;
        RECT 9.690 195.630 66.210 196.730 ;
        RECT 6.965 194.690 78.595 195.630 ;
        RECT 6.965 193.590 67.130 194.690 ;
        RECT 6.965 192.650 78.595 193.590 ;
        RECT 6.965 191.970 70.350 192.650 ;
        RECT 7.390 191.550 70.350 191.970 ;
        RECT 7.390 191.290 78.595 191.550 ;
        RECT 7.390 190.870 69.890 191.290 ;
        RECT 6.965 190.190 69.890 190.870 ;
        RECT 6.965 189.250 78.595 190.190 ;
        RECT 6.965 188.150 66.670 189.250 ;
        RECT 6.965 187.890 78.595 188.150 ;
        RECT 6.965 186.790 70.350 187.890 ;
        RECT 6.965 186.530 78.595 186.790 ;
        RECT 7.390 185.850 78.595 186.530 ;
        RECT 7.390 185.430 70.350 185.850 ;
        RECT 6.965 184.750 70.350 185.430 ;
        RECT 6.965 184.490 78.595 184.750 ;
        RECT 6.965 183.390 57.470 184.490 ;
        RECT 6.965 182.450 78.595 183.390 ;
        RECT 6.965 181.770 68.510 182.450 ;
        RECT 9.690 181.350 68.510 181.770 ;
        RECT 9.690 180.670 78.595 181.350 ;
        RECT 6.965 180.410 78.595 180.670 ;
        RECT 6.965 179.310 57.930 180.410 ;
        RECT 6.965 179.050 78.595 179.310 ;
        RECT 6.965 177.950 59.310 179.050 ;
        RECT 6.965 177.010 78.595 177.950 ;
        RECT 9.690 175.910 67.590 177.010 ;
        RECT 6.965 175.650 78.595 175.910 ;
        RECT 6.965 174.550 68.050 175.650 ;
        RECT 6.965 173.610 78.595 174.550 ;
        RECT 6.965 172.510 68.510 173.610 ;
        RECT 6.965 172.250 78.595 172.510 ;
        RECT 7.390 171.150 70.750 172.250 ;
        RECT 6.965 170.210 78.595 171.150 ;
        RECT 6.965 169.110 68.510 170.210 ;
        RECT 6.965 168.850 78.595 169.110 ;
        RECT 6.965 167.750 67.590 168.850 ;
        RECT 6.965 167.490 78.595 167.750 ;
        RECT 7.390 166.810 78.595 167.490 ;
        RECT 7.390 166.390 74.950 166.810 ;
        RECT 6.965 165.710 74.950 166.390 ;
        RECT 6.965 164.770 78.595 165.710 ;
        RECT 6.965 163.670 69.890 164.770 ;
        RECT 6.965 163.410 78.595 163.670 ;
        RECT 6.965 162.730 75.410 163.410 ;
        RECT 7.390 162.310 75.410 162.730 ;
        RECT 7.390 161.630 78.595 162.310 ;
        RECT 6.965 161.370 78.595 161.630 ;
        RECT 6.965 160.270 68.510 161.370 ;
        RECT 6.965 160.010 78.595 160.270 ;
        RECT 6.965 158.910 56.090 160.010 ;
        RECT 6.965 157.970 78.595 158.910 ;
        RECT 7.390 156.870 57.930 157.970 ;
        RECT 6.965 156.610 78.595 156.870 ;
        RECT 6.965 155.510 61.550 156.610 ;
        RECT 6.965 154.570 78.595 155.510 ;
        RECT 6.965 153.470 57.930 154.570 ;
        RECT 6.965 153.210 78.595 153.470 ;
        RECT 7.390 152.530 78.595 153.210 ;
        RECT 7.390 152.110 55.170 152.530 ;
        RECT 6.965 151.430 55.170 152.110 ;
        RECT 6.965 151.170 78.595 151.430 ;
        RECT 6.965 150.070 57.930 151.170 ;
        RECT 6.965 149.130 78.595 150.070 ;
        RECT 6.965 148.030 67.590 149.130 ;
        RECT 6.965 147.770 78.595 148.030 ;
        RECT 9.690 146.670 60.230 147.770 ;
        RECT 6.965 145.730 78.595 146.670 ;
        RECT 6.965 144.630 61.550 145.730 ;
        RECT 6.965 144.370 78.595 144.630 ;
        RECT 6.965 143.270 69.890 144.370 ;
        RECT 6.965 143.010 78.595 143.270 ;
        RECT 9.690 142.330 78.595 143.010 ;
        RECT 9.690 141.910 60.230 142.330 ;
        RECT 6.965 141.230 60.230 141.910 ;
        RECT 6.965 140.970 78.595 141.230 ;
        RECT 6.965 139.870 58.850 140.970 ;
        RECT 6.965 138.930 78.595 139.870 ;
        RECT 6.965 138.250 70.750 138.930 ;
        RECT 9.690 137.830 70.750 138.250 ;
        RECT 9.690 137.150 78.595 137.830 ;
        RECT 6.965 136.890 78.595 137.150 ;
        RECT 6.965 135.790 60.230 136.890 ;
        RECT 6.965 135.530 78.595 135.790 ;
        RECT 6.965 134.430 55.630 135.530 ;
        RECT 6.965 133.490 78.595 134.430 ;
        RECT 9.690 132.390 70.750 133.490 ;
        RECT 6.965 132.130 78.595 132.390 ;
        RECT 6.965 131.030 70.750 132.130 ;
        RECT 6.965 130.090 78.595 131.030 ;
        RECT 6.965 128.990 55.170 130.090 ;
        RECT 6.965 128.730 78.595 128.990 ;
        RECT 9.690 127.630 70.750 128.730 ;
        RECT 6.965 126.690 78.595 127.630 ;
        RECT 6.965 125.590 61.550 126.690 ;
        RECT 6.965 124.650 78.595 125.590 ;
        RECT 6.965 123.970 56.090 124.650 ;
        RECT 7.390 123.550 56.090 123.970 ;
        RECT 7.390 123.290 78.595 123.550 ;
        RECT 7.390 122.870 70.750 123.290 ;
        RECT 6.965 122.190 70.750 122.870 ;
        RECT 6.965 121.250 78.595 122.190 ;
        RECT 6.965 120.150 55.170 121.250 ;
        RECT 6.965 119.890 78.595 120.150 ;
        RECT 6.965 119.210 57.010 119.890 ;
        RECT 7.390 118.790 57.010 119.210 ;
        RECT 7.390 118.110 78.595 118.790 ;
        RECT 6.965 117.850 78.595 118.110 ;
        RECT 6.965 116.750 70.750 117.850 ;
        RECT 6.965 116.490 78.595 116.750 ;
        RECT 6.965 115.390 58.850 116.490 ;
        RECT 6.965 114.450 78.595 115.390 ;
        RECT 7.390 113.350 60.690 114.450 ;
        RECT 6.965 113.090 78.595 113.350 ;
        RECT 6.965 111.990 60.230 113.090 ;
        RECT 6.965 111.050 78.595 111.990 ;
        RECT 6.965 109.950 55.170 111.050 ;
        RECT 6.965 109.010 78.595 109.950 ;
        RECT 9.690 107.910 65.750 109.010 ;
        RECT 6.965 107.650 78.595 107.910 ;
        RECT 6.965 106.550 55.170 107.650 ;
        RECT 6.965 105.610 78.595 106.550 ;
        RECT 6.965 104.510 73.110 105.610 ;
        RECT 6.965 104.250 78.595 104.510 ;
        RECT 9.690 103.150 75.410 104.250 ;
        RECT 6.965 102.210 78.595 103.150 ;
        RECT 6.965 101.110 60.690 102.210 ;
        RECT 6.965 100.850 78.595 101.110 ;
        RECT 6.965 99.750 78.170 100.850 ;
        RECT 6.965 99.490 78.595 99.750 ;
        RECT 9.690 98.810 78.595 99.490 ;
        RECT 9.690 98.390 61.550 98.810 ;
        RECT 6.965 97.710 61.550 98.390 ;
        RECT 6.965 96.770 78.595 97.710 ;
        RECT 6.965 95.670 68.510 96.770 ;
        RECT 6.965 95.410 78.595 95.670 ;
        RECT 6.965 94.730 71.670 95.410 ;
        RECT 7.390 94.310 71.670 94.730 ;
        RECT 7.390 93.630 78.595 94.310 ;
        RECT 6.965 93.370 78.595 93.630 ;
        RECT 6.965 92.270 56.550 93.370 ;
        RECT 6.965 92.010 78.595 92.270 ;
        RECT 6.965 90.910 59.770 92.010 ;
        RECT 6.965 89.970 78.595 90.910 ;
        RECT 9.690 88.870 75.350 89.970 ;
        RECT 6.965 88.610 78.595 88.870 ;
        RECT 6.965 87.510 59.100 88.610 ;
        RECT 6.965 86.570 78.595 87.510 ;
        RECT 6.965 85.470 57.470 86.570 ;
        RECT 6.965 85.210 78.595 85.470 ;
        RECT 9.690 84.110 70.060 85.210 ;
        RECT 6.965 83.170 78.595 84.110 ;
        RECT 6.965 82.070 55.170 83.170 ;
        RECT 6.965 81.130 78.595 82.070 ;
        RECT 6.965 80.450 59.310 81.130 ;
        RECT 7.390 80.030 59.310 80.450 ;
        RECT 7.390 79.770 78.595 80.030 ;
        RECT 7.390 79.350 70.060 79.770 ;
        RECT 6.965 78.670 70.060 79.350 ;
        RECT 6.965 77.730 78.595 78.670 ;
        RECT 6.965 76.630 56.550 77.730 ;
        RECT 6.965 76.370 78.595 76.630 ;
        RECT 6.965 75.270 54.250 76.370 ;
        RECT 6.965 75.010 78.595 75.270 ;
        RECT 7.390 74.330 78.595 75.010 ;
        RECT 7.390 73.910 70.060 74.330 ;
        RECT 6.965 73.230 70.060 73.910 ;
        RECT 6.965 72.970 78.595 73.230 ;
        RECT 6.965 71.870 57.010 72.970 ;
        RECT 6.965 70.930 78.595 71.870 ;
        RECT 6.965 70.250 57.930 70.930 ;
        RECT 7.390 69.830 57.930 70.250 ;
        RECT 7.390 69.150 78.595 69.830 ;
        RECT 6.965 68.890 78.595 69.150 ;
        RECT 6.965 67.790 65.750 68.890 ;
        RECT 6.965 67.530 78.595 67.790 ;
        RECT 6.965 66.430 57.470 67.530 ;
        RECT 6.965 65.490 78.595 66.430 ;
        RECT 14.290 64.390 66.210 65.490 ;
        RECT 6.965 64.130 78.595 64.390 ;
        RECT 6.965 63.030 61.610 64.130 ;
        RECT 6.965 62.090 78.595 63.030 ;
        RECT 6.965 60.990 60.690 62.090 ;
        RECT 6.965 60.730 78.595 60.990 ;
        RECT 10.150 59.630 57.010 60.730 ;
        RECT 6.965 58.690 78.595 59.630 ;
        RECT 6.965 57.590 66.670 58.690 ;
        RECT 6.965 57.330 78.595 57.590 ;
        RECT 6.965 56.230 65.230 57.330 ;
        RECT 6.965 55.970 78.595 56.230 ;
        RECT 10.610 55.290 78.595 55.970 ;
        RECT 10.610 54.870 57.640 55.290 ;
        RECT 6.965 54.190 57.640 54.870 ;
        RECT 6.965 53.250 78.595 54.190 ;
        RECT 6.965 52.150 55.170 53.250 ;
        RECT 6.965 51.890 78.595 52.150 ;
        RECT 6.965 51.210 73.510 51.890 ;
        RECT 10.150 50.790 73.510 51.210 ;
        RECT 10.150 50.110 78.595 50.790 ;
        RECT 6.965 49.850 78.595 50.110 ;
        RECT 6.965 48.750 55.630 49.850 ;
        RECT 6.965 48.490 78.595 48.750 ;
        RECT 6.965 47.390 57.470 48.490 ;
        RECT 6.965 46.450 78.595 47.390 ;
        RECT 10.150 45.350 70.750 46.450 ;
        RECT 6.965 45.090 78.595 45.350 ;
        RECT 6.965 43.990 57.930 45.090 ;
        RECT 6.965 43.050 78.595 43.990 ;
        RECT 6.965 41.950 66.210 43.050 ;
        RECT 6.965 41.690 78.595 41.950 ;
        RECT 10.610 41.010 78.595 41.690 ;
        RECT 10.610 40.590 64.310 41.010 ;
        RECT 6.965 39.910 64.310 40.590 ;
        RECT 6.965 39.650 78.595 39.910 ;
        RECT 6.965 38.550 55.170 39.650 ;
        RECT 6.965 37.610 78.595 38.550 ;
        RECT 6.965 36.510 49.190 37.610 ;
        RECT 6.965 36.250 78.595 36.510 ;
        RECT 7.390 35.150 70.750 36.250 ;
        RECT 6.965 34.210 78.595 35.150 ;
        RECT 6.965 33.110 58.850 34.210 ;
        RECT 6.965 32.850 78.595 33.110 ;
        RECT 6.965 31.750 55.170 32.850 ;
        RECT 6.965 31.490 78.595 31.750 ;
        RECT 10.610 30.810 78.595 31.490 ;
        RECT 10.610 30.390 76.270 30.810 ;
        RECT 6.965 29.710 76.270 30.390 ;
        RECT 6.965 29.450 78.595 29.710 ;
        RECT 6.965 28.350 55.630 29.450 ;
        RECT 6.965 27.410 78.595 28.350 ;
        RECT 6.965 26.730 59.770 27.410 ;
        RECT 10.150 26.310 59.770 26.730 ;
        RECT 10.150 25.630 78.595 26.310 ;
        RECT 6.965 25.370 78.595 25.630 ;
        RECT 6.965 24.270 76.270 25.370 ;
        RECT 6.965 24.010 78.595 24.270 ;
        RECT 6.965 22.910 74.490 24.010 ;
        RECT 6.965 21.970 78.595 22.910 ;
        RECT 14.290 20.870 68.510 21.970 ;
        RECT 6.965 20.610 78.595 20.870 ;
        RECT 6.965 19.510 58.390 20.610 ;
        RECT 6.965 18.570 78.595 19.510 ;
        RECT 6.965 17.470 68.050 18.570 ;
        RECT 6.965 17.210 78.595 17.470 ;
        RECT 10.150 16.110 55.630 17.210 ;
        RECT 6.965 15.170 78.595 16.110 ;
        RECT 6.965 14.070 68.510 15.170 ;
        RECT 6.965 13.130 78.595 14.070 ;
        RECT 6.965 12.450 54.710 13.130 ;
        RECT 10.150 12.030 54.710 12.450 ;
        RECT 10.150 11.770 78.595 12.030 ;
        RECT 10.150 11.350 56.090 11.770 ;
        RECT 6.965 10.670 56.090 11.350 ;
        RECT 6.965 9.730 78.595 10.670 ;
        RECT 6.965 8.630 51.490 9.730 ;
        RECT 6.965 8.370 78.595 8.630 ;
        RECT 6.965 7.690 68.510 8.370 ;
        RECT 14.750 7.270 68.510 7.690 ;
        RECT 14.750 6.590 78.595 7.270 ;
        RECT 6.965 6.330 78.595 6.590 ;
        RECT 6.965 5.230 57.010 6.330 ;
        RECT 6.965 4.970 78.595 5.230 ;
        RECT 6.965 3.870 56.550 4.970 ;
        RECT 6.965 2.930 78.595 3.870 ;
        RECT 9.690 1.830 55.170 2.930 ;
        RECT 6.965 1.570 78.595 1.830 ;
        RECT 6.965 0.855 55.630 1.570 ;
      LAYER met4 ;
        RECT 18.215 5.200 27.305 217.840 ;
        RECT 29.705 5.200 38.800 217.840 ;
        RECT 41.200 5.200 50.290 217.840 ;
        RECT 52.690 5.200 61.785 217.840 ;
        RECT 64.185 5.200 69.625 217.840 ;
  END
END W_IO
MACRO sky130_sram_2kbyte_1rw1r_32x512_8
   CLASS BLOCK ;
   SIZE 683.1 BY 416.54 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  115.6 0.0 115.98 1.06 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  121.04 0.0 121.42 1.06 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  127.16 0.0 127.54 1.06 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  132.6 0.0 132.98 1.06 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  138.04 0.0 138.42 1.06 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  143.48 0.0 143.86 1.06 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  150.28 0.0 150.66 1.06 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  156.4 0.0 156.78 1.06 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  161.84 0.0 162.22 1.06 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  167.28 0.0 167.66 1.06 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  172.72 0.0 173.1 1.06 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  179.52 0.0 179.9 1.06 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  184.96 0.0 185.34 1.06 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  190.4 0.0 190.78 1.06 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  197.2 0.0 197.58 1.06 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  203.32 0.0 203.7 1.06 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  208.76 0.0 209.14 1.06 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  214.2 0.0 214.58 1.06 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  219.64 0.0 220.02 1.06 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  226.44 0.0 226.82 1.06 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  231.88 0.0 232.26 1.06 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  238.0 0.0 238.38 1.06 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  243.44 0.0 243.82 1.06 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  248.88 0.0 249.26 1.06 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  255.68 0.0 256.06 1.06 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  261.12 0.0 261.5 1.06 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  266.56 0.0 266.94 1.06 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  272.0 0.0 272.38 1.06 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  278.8 0.0 279.18 1.06 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  284.92 0.0 285.3 1.06 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  290.36 0.0 290.74 1.06 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  295.8 0.0 296.18 1.06 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  80.24 0.0 80.62 1.06 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  85.68 0.0 86.06 1.06 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 140.76 1.06 141.14 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 149.6 1.06 149.98 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 155.04 1.06 155.42 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 163.88 1.06 164.26 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 168.64 1.06 169.02 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 179.52 1.06 179.9 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 184.28 1.06 184.66 ;
      END
   END addr0[8]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  598.4 415.48 598.78 416.54 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  592.28 415.48 592.66 416.54 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  682.04 96.56 683.1 96.94 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  682.04 88.4 683.1 88.78 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  682.04 81.6 683.1 81.98 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  682.04 74.12 683.1 74.5 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  682.04 68.0 683.1 68.38 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  616.08 0.0 616.46 1.06 ;
      END
   END addr1[7]
   PIN addr1[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  616.76 0.0 617.14 1.06 ;
      END
   END addr1[8]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 40.12 1.06 40.5 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  682.04 395.76 683.1 396.14 ;
      END
   END csb1
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 49.64 1.06 50.02 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 41.48 1.06 41.86 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  654.16 415.48 654.54 416.54 ;
      END
   END clk1
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  91.12 0.0 91.5 1.06 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  97.92 0.0 98.3 1.06 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  102.68 0.0 103.06 1.06 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  108.8 0.0 109.18 1.06 ;
      END
   END wmask0[3]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  141.44 0.0 141.82 1.06 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  153.68 0.0 154.06 1.06 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  167.96 0.0 168.34 1.06 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  180.2 0.0 180.58 1.06 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  192.44 0.0 192.82 1.06 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  205.36 0.0 205.74 1.06 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  217.6 0.0 217.98 1.06 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  229.84 0.0 230.22 1.06 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  241.4 0.0 241.78 1.06 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  255.0 0.0 255.38 1.06 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  267.92 0.0 268.3 1.06 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  280.16 0.0 280.54 1.06 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  292.4 0.0 292.78 1.06 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  304.64 0.0 305.02 1.06 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  317.56 0.0 317.94 1.06 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  329.8 0.0 330.18 1.06 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  341.36 0.0 341.74 1.06 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  354.96 0.0 355.34 1.06 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  367.2 0.0 367.58 1.06 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  379.44 0.0 379.82 1.06 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  392.36 0.0 392.74 1.06 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  404.6 0.0 404.98 1.06 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  417.52 0.0 417.9 1.06 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  429.76 0.0 430.14 1.06 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  442.68 0.0 443.06 1.06 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  454.92 0.0 455.3 1.06 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  467.16 0.0 467.54 1.06 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  479.4 0.0 479.78 1.06 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  492.32 0.0 492.7 1.06 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  504.56 0.0 504.94 1.06 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  516.8 0.0 517.18 1.06 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  529.72 0.0 530.1 1.06 ;
      END
   END dout0[31]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  143.48 415.48 143.86 416.54 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  155.04 415.48 155.42 416.54 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  167.28 415.48 167.66 416.54 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  180.88 415.48 181.26 416.54 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  192.44 415.48 192.82 416.54 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  205.36 415.48 205.74 416.54 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  217.6 415.48 217.98 416.54 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  230.52 415.48 230.9 416.54 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  242.76 415.48 243.14 416.54 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  255.68 415.48 256.06 416.54 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  267.92 415.48 268.3 416.54 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  280.84 415.48 281.22 416.54 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  292.4 415.48 292.78 416.54 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  304.64 415.48 305.02 416.54 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  318.24 415.48 318.62 416.54 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  330.48 415.48 330.86 416.54 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  342.72 415.48 343.1 416.54 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  354.96 415.48 355.34 416.54 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  367.88 415.48 368.26 416.54 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  379.44 415.48 379.82 416.54 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  393.04 415.48 393.42 416.54 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  405.28 415.48 405.66 416.54 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  417.52 415.48 417.9 416.54 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  429.76 415.48 430.14 416.54 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  442.0 415.48 442.38 416.54 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  454.92 415.48 455.3 416.54 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  467.84 415.48 468.22 416.54 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  480.08 415.48 480.46 416.54 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  492.32 415.48 492.7 416.54 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  505.24 415.48 505.62 416.54 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  516.8 415.48 517.18 416.54 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  530.4 415.48 530.78 416.54 ;
      END
   END dout1[31]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  4.76 4.76 6.5 411.78 ;
         LAYER met4 ;
         RECT  676.6 4.76 678.34 411.78 ;
         LAYER met3 ;
         RECT  4.76 410.04 678.34 411.78 ;
         LAYER met3 ;
         RECT  4.76 4.76 678.34 6.5 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  680.0 1.36 681.74 415.18 ;
         LAYER met4 ;
         RECT  1.36 1.36 3.1 415.18 ;
         LAYER met3 ;
         RECT  1.36 1.36 681.74 3.1 ;
         LAYER met3 ;
         RECT  1.36 413.44 681.74 415.18 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 682.48 415.92 ;
   LAYER  met2 ;
      RECT  0.62 0.62 682.48 415.92 ;
   LAYER  met3 ;
      RECT  1.66 140.16 682.48 141.74 ;
      RECT  0.62 141.74 1.66 149.0 ;
      RECT  0.62 150.58 1.66 154.44 ;
      RECT  0.62 156.02 1.66 163.28 ;
      RECT  0.62 164.86 1.66 168.04 ;
      RECT  0.62 169.62 1.66 178.92 ;
      RECT  0.62 180.5 1.66 183.68 ;
      RECT  1.66 95.96 681.44 97.54 ;
      RECT  1.66 97.54 681.44 140.16 ;
      RECT  681.44 97.54 682.48 140.16 ;
      RECT  681.44 89.38 682.48 95.96 ;
      RECT  681.44 82.58 682.48 87.8 ;
      RECT  681.44 75.1 682.48 81.0 ;
      RECT  681.44 68.98 682.48 73.52 ;
      RECT  1.66 141.74 681.44 395.16 ;
      RECT  1.66 395.16 681.44 396.74 ;
      RECT  681.44 141.74 682.48 395.16 ;
      RECT  0.62 50.62 1.66 140.16 ;
      RECT  0.62 42.46 1.66 49.04 ;
      RECT  1.66 396.74 4.16 409.44 ;
      RECT  1.66 409.44 4.16 412.38 ;
      RECT  4.16 396.74 678.94 409.44 ;
      RECT  678.94 396.74 681.44 409.44 ;
      RECT  678.94 409.44 681.44 412.38 ;
      RECT  1.66 4.16 4.16 7.1 ;
      RECT  1.66 7.1 4.16 95.96 ;
      RECT  4.16 7.1 678.94 95.96 ;
      RECT  678.94 4.16 681.44 7.1 ;
      RECT  678.94 7.1 681.44 95.96 ;
      RECT  681.44 0.62 682.34 0.76 ;
      RECT  681.44 3.7 682.34 67.4 ;
      RECT  682.34 0.62 682.48 0.76 ;
      RECT  682.34 0.76 682.48 3.7 ;
      RECT  682.34 3.7 682.48 67.4 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 3.7 ;
      RECT  0.62 3.7 0.76 39.52 ;
      RECT  0.76 0.62 1.66 0.76 ;
      RECT  0.76 3.7 1.66 39.52 ;
      RECT  1.66 0.62 4.16 0.76 ;
      RECT  1.66 3.7 4.16 4.16 ;
      RECT  4.16 0.62 678.94 0.76 ;
      RECT  4.16 3.7 678.94 4.16 ;
      RECT  678.94 0.62 681.44 0.76 ;
      RECT  678.94 3.7 681.44 4.16 ;
      RECT  0.62 185.26 0.76 412.84 ;
      RECT  0.62 412.84 0.76 415.78 ;
      RECT  0.62 415.78 0.76 415.92 ;
      RECT  0.76 185.26 1.66 412.84 ;
      RECT  0.76 415.78 1.66 415.92 ;
      RECT  681.44 396.74 682.34 412.84 ;
      RECT  681.44 415.78 682.34 415.92 ;
      RECT  682.34 396.74 682.48 412.84 ;
      RECT  682.34 412.84 682.48 415.78 ;
      RECT  682.34 415.78 682.48 415.92 ;
      RECT  1.66 412.38 4.16 412.84 ;
      RECT  1.66 415.78 4.16 415.92 ;
      RECT  4.16 412.38 678.94 412.84 ;
      RECT  4.16 415.78 678.94 415.92 ;
      RECT  678.94 412.38 681.44 412.84 ;
      RECT  678.94 415.78 681.44 415.92 ;
   LAYER  met4 ;
      RECT  115.0 1.66 116.58 415.92 ;
      RECT  116.58 0.62 120.44 1.66 ;
      RECT  122.02 0.62 126.56 1.66 ;
      RECT  128.14 0.62 132.0 1.66 ;
      RECT  133.58 0.62 137.44 1.66 ;
      RECT  144.46 0.62 149.68 1.66 ;
      RECT  157.38 0.62 161.24 1.66 ;
      RECT  162.82 0.62 166.68 1.66 ;
      RECT  173.7 0.62 178.92 1.66 ;
      RECT  185.94 0.62 189.8 1.66 ;
      RECT  198.18 0.62 202.72 1.66 ;
      RECT  209.74 0.62 213.6 1.66 ;
      RECT  220.62 0.62 225.84 1.66 ;
      RECT  232.86 0.62 237.4 1.66 ;
      RECT  244.42 0.62 248.28 1.66 ;
      RECT  256.66 0.62 260.52 1.66 ;
      RECT  262.1 0.62 265.96 1.66 ;
      RECT  272.98 0.62 278.2 1.66 ;
      RECT  285.9 0.62 289.76 1.66 ;
      RECT  81.22 0.62 85.08 1.66 ;
      RECT  116.58 1.66 597.8 414.88 ;
      RECT  597.8 1.66 599.38 414.88 ;
      RECT  593.26 414.88 597.8 415.92 ;
      RECT  599.38 414.88 653.56 415.92 ;
      RECT  86.66 0.62 90.52 1.66 ;
      RECT  92.1 0.62 97.32 1.66 ;
      RECT  98.9 0.62 102.08 1.66 ;
      RECT  103.66 0.62 108.2 1.66 ;
      RECT  109.78 0.62 115.0 1.66 ;
      RECT  139.02 0.62 140.84 1.66 ;
      RECT  142.42 0.62 142.88 1.66 ;
      RECT  151.26 0.62 153.08 1.66 ;
      RECT  154.66 0.62 155.8 1.66 ;
      RECT  168.94 0.62 172.12 1.66 ;
      RECT  181.18 0.62 184.36 1.66 ;
      RECT  191.38 0.62 191.84 1.66 ;
      RECT  193.42 0.62 196.6 1.66 ;
      RECT  204.3 0.62 204.76 1.66 ;
      RECT  206.34 0.62 208.16 1.66 ;
      RECT  215.18 0.62 217.0 1.66 ;
      RECT  218.58 0.62 219.04 1.66 ;
      RECT  227.42 0.62 229.24 1.66 ;
      RECT  230.82 0.62 231.28 1.66 ;
      RECT  238.98 0.62 240.8 1.66 ;
      RECT  242.38 0.62 242.84 1.66 ;
      RECT  249.86 0.62 254.4 1.66 ;
      RECT  268.9 0.62 271.4 1.66 ;
      RECT  281.14 0.62 284.32 1.66 ;
      RECT  291.34 0.62 291.8 1.66 ;
      RECT  293.38 0.62 295.2 1.66 ;
      RECT  296.78 0.62 304.04 1.66 ;
      RECT  305.62 0.62 316.96 1.66 ;
      RECT  318.54 0.62 329.2 1.66 ;
      RECT  330.78 0.62 340.76 1.66 ;
      RECT  342.34 0.62 354.36 1.66 ;
      RECT  355.94 0.62 366.6 1.66 ;
      RECT  368.18 0.62 378.84 1.66 ;
      RECT  380.42 0.62 391.76 1.66 ;
      RECT  393.34 0.62 404.0 1.66 ;
      RECT  405.58 0.62 416.92 1.66 ;
      RECT  418.5 0.62 429.16 1.66 ;
      RECT  430.74 0.62 442.08 1.66 ;
      RECT  443.66 0.62 454.32 1.66 ;
      RECT  455.9 0.62 466.56 1.66 ;
      RECT  468.14 0.62 478.8 1.66 ;
      RECT  480.38 0.62 491.72 1.66 ;
      RECT  493.3 0.62 503.96 1.66 ;
      RECT  505.54 0.62 516.2 1.66 ;
      RECT  517.78 0.62 529.12 1.66 ;
      RECT  530.7 0.62 615.48 1.66 ;
      RECT  116.58 414.88 142.88 415.92 ;
      RECT  144.46 414.88 154.44 415.92 ;
      RECT  156.02 414.88 166.68 415.92 ;
      RECT  168.26 414.88 180.28 415.92 ;
      RECT  181.86 414.88 191.84 415.92 ;
      RECT  193.42 414.88 204.76 415.92 ;
      RECT  206.34 414.88 217.0 415.92 ;
      RECT  218.58 414.88 229.92 415.92 ;
      RECT  231.5 414.88 242.16 415.92 ;
      RECT  243.74 414.88 255.08 415.92 ;
      RECT  256.66 414.88 267.32 415.92 ;
      RECT  268.9 414.88 280.24 415.92 ;
      RECT  281.82 414.88 291.8 415.92 ;
      RECT  293.38 414.88 304.04 415.92 ;
      RECT  305.62 414.88 317.64 415.92 ;
      RECT  319.22 414.88 329.88 415.92 ;
      RECT  331.46 414.88 342.12 415.92 ;
      RECT  343.7 414.88 354.36 415.92 ;
      RECT  355.94 414.88 367.28 415.92 ;
      RECT  368.86 414.88 378.84 415.92 ;
      RECT  380.42 414.88 392.44 415.92 ;
      RECT  394.02 414.88 404.68 415.92 ;
      RECT  406.26 414.88 416.92 415.92 ;
      RECT  418.5 414.88 429.16 415.92 ;
      RECT  430.74 414.88 441.4 415.92 ;
      RECT  442.98 414.88 454.32 415.92 ;
      RECT  455.9 414.88 467.24 415.92 ;
      RECT  468.82 414.88 479.48 415.92 ;
      RECT  481.06 414.88 491.72 415.92 ;
      RECT  493.3 414.88 504.64 415.92 ;
      RECT  506.22 414.88 516.2 415.92 ;
      RECT  517.78 414.88 529.8 415.92 ;
      RECT  531.38 414.88 591.68 415.92 ;
      RECT  4.16 1.66 7.1 4.16 ;
      RECT  4.16 412.38 7.1 415.92 ;
      RECT  7.1 1.66 115.0 4.16 ;
      RECT  7.1 4.16 115.0 412.38 ;
      RECT  7.1 412.38 115.0 415.92 ;
      RECT  599.38 1.66 676.0 4.16 ;
      RECT  599.38 4.16 676.0 412.38 ;
      RECT  599.38 412.38 676.0 414.88 ;
      RECT  676.0 1.66 678.94 4.16 ;
      RECT  676.0 412.38 678.94 414.88 ;
      RECT  617.74 0.62 679.4 0.76 ;
      RECT  617.74 0.76 679.4 1.66 ;
      RECT  679.4 0.62 682.34 0.76 ;
      RECT  682.34 0.62 682.48 0.76 ;
      RECT  682.34 0.76 682.48 1.66 ;
      RECT  655.14 414.88 679.4 415.78 ;
      RECT  655.14 415.78 679.4 415.92 ;
      RECT  679.4 415.78 682.34 415.92 ;
      RECT  682.34 414.88 682.48 415.78 ;
      RECT  682.34 415.78 682.48 415.92 ;
      RECT  678.94 1.66 679.4 4.16 ;
      RECT  682.34 1.66 682.48 4.16 ;
      RECT  678.94 4.16 679.4 412.38 ;
      RECT  682.34 4.16 682.48 412.38 ;
      RECT  678.94 412.38 679.4 414.88 ;
      RECT  682.34 412.38 682.48 414.88 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 1.66 ;
      RECT  0.76 0.62 3.7 0.76 ;
      RECT  3.7 0.62 79.64 0.76 ;
      RECT  3.7 0.76 79.64 1.66 ;
      RECT  0.62 1.66 0.76 4.16 ;
      RECT  3.7 1.66 4.16 4.16 ;
      RECT  0.62 4.16 0.76 412.38 ;
      RECT  3.7 4.16 4.16 412.38 ;
      RECT  0.62 412.38 0.76 415.78 ;
      RECT  0.62 415.78 0.76 415.92 ;
      RECT  0.76 415.78 3.7 415.92 ;
      RECT  3.7 412.38 4.16 415.78 ;
      RECT  3.7 415.78 4.16 415.92 ;
   END
END    sky130_sram_2kbyte_1rw1r_32x512_8
MACRO LUT4AB
  CLASS BLOCK ;
  FOREIGN LUT4AB ;
  ORIGIN 0.000 0.000 ;
  SIZE 223.275 BY 223.115 ;
  PIN Ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.460 0.000 186.600 7.000 ;
    END
  END Ci
  PIN Co
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.000 217.220 186.140 223.115 ;
    END
  END Co
  PIN E1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 204.610 84.510 223.275 84.810 ;
    END
  END E1BEG[0]
  PIN E1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 219.790 85.870 223.275 86.170 ;
    END
  END E1BEG[1]
  PIN E1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.620 87.910 223.275 88.210 ;
    END
  END E1BEG[2]
  PIN E1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 219.790 89.270 223.275 89.570 ;
    END
  END E1BEG[3]
  PIN E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.510 6.990 84.810 ;
    END
  END E1END[0]
  PIN E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.870 7.450 86.170 ;
    END
  END E1END[1]
  PIN E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.910 6.530 88.210 ;
    END
  END E1END[2]
  PIN E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.270 20.330 89.570 ;
    END
  END E1END[3]
  PIN E2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 219.790 91.310 223.275 91.610 ;
    END
  END E2BEG[0]
  PIN E2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.850 92.670 223.275 92.970 ;
    END
  END E2BEG[1]
  PIN E2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 219.790 94.710 223.275 95.010 ;
    END
  END E2BEG[2]
  PIN E2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 200.470 96.070 223.275 96.370 ;
    END
  END E2BEG[3]
  PIN E2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 200.930 98.110 223.275 98.410 ;
    END
  END E2BEG[4]
  PIN E2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 100.150 223.275 100.450 ;
    END
  END E2BEG[5]
  PIN E2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 101.510 223.275 101.810 ;
    END
  END E2BEG[6]
  PIN E2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 219.790 103.550 223.275 103.850 ;
    END
  END E2BEG[7]
  PIN E2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 219.790 104.910 223.275 105.210 ;
    END
  END E2BEGb[0]
  PIN E2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 219.790 106.950 223.275 107.250 ;
    END
  END E2BEGb[1]
  PIN E2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.390 108.310 223.275 108.610 ;
    END
  END E2BEGb[2]
  PIN E2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 219.790 110.350 223.275 110.650 ;
    END
  END E2BEGb[3]
  PIN E2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 204.610 112.390 223.275 112.690 ;
    END
  END E2BEGb[4]
  PIN E2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 205.530 113.750 223.275 114.050 ;
    END
  END E2BEGb[5]
  PIN E2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 219.790 115.790 223.275 116.090 ;
    END
  END E2BEGb[6]
  PIN E2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 203.230 117.150 223.275 117.450 ;
    END
  END E2BEGb[7]
  PIN E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.910 20.330 105.210 ;
    END
  END E2END[0]
  PIN E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.950 19.870 107.250 ;
    END
  END E2END[1]
  PIN E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.310 9.290 108.610 ;
    END
  END E2END[2]
  PIN E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.350 5.610 110.650 ;
    END
  END E2END[3]
  PIN E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.390 18.950 112.690 ;
    END
  END E2END[4]
  PIN E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.750 27.690 114.050 ;
    END
  END E2END[5]
  PIN E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.790 17.570 116.090 ;
    END
  END E2END[6]
  PIN E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.150 6.990 117.450 ;
    END
  END E2END[7]
  PIN E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.310 20.790 91.610 ;
    END
  END E2MID[0]
  PIN E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.670 11.590 92.970 ;
    END
  END E2MID[1]
  PIN E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.710 17.860 95.010 ;
    END
  END E2MID[2]
  PIN E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.070 16.650 96.370 ;
    END
  END E2MID[3]
  PIN E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.110 20.330 98.410 ;
    END
  END E2MID[4]
  PIN E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.150 6.530 100.450 ;
    END
  END E2MID[5]
  PIN E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.510 15.270 101.810 ;
    END
  END E2MID[6]
  PIN E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.550 18.030 103.850 ;
    END
  END E2MID[7]
  PIN E6BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 147.070 223.275 147.370 ;
    END
  END E6BEG[0]
  PIN E6BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 164.070 223.275 164.370 ;
    END
  END E6BEG[10]
  PIN E6BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 166.110 223.275 166.410 ;
    END
  END E6BEG[11]
  PIN E6BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 148.430 223.275 148.730 ;
    END
  END E6BEG[1]
  PIN E6BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 150.470 223.275 150.770 ;
    END
  END E6BEG[2]
  PIN E6BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 151.830 223.275 152.130 ;
    END
  END E6BEG[3]
  PIN E6BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 153.870 223.275 154.170 ;
    END
  END E6BEG[4]
  PIN E6BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.410 155.910 223.275 156.210 ;
    END
  END E6BEG[5]
  PIN E6BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.410 157.270 223.275 157.570 ;
    END
  END E6BEG[6]
  PIN E6BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 159.310 223.275 159.610 ;
    END
  END E6BEG[7]
  PIN E6BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.410 160.670 223.275 160.970 ;
    END
  END E6BEG[8]
  PIN E6BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.590 162.710 223.275 163.010 ;
    END
  END E6BEG[9]
  PIN E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.070 7.450 147.370 ;
    END
  END E6END[0]
  PIN E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.070 9.750 164.370 ;
    END
  END E6END[10]
  PIN E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.110 19.410 166.410 ;
    END
  END E6END[11]
  PIN E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.430 7.450 148.730 ;
    END
  END E6END[1]
  PIN E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 150.470 20.790 150.770 ;
    END
  END E6END[2]
  PIN E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.830 16.940 152.130 ;
    END
  END E6END[3]
  PIN E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.870 14.350 154.170 ;
    END
  END E6END[4]
  PIN E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.910 18.030 156.210 ;
    END
  END E6END[5]
  PIN E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.270 18.780 157.570 ;
    END
  END E6END[6]
  PIN E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.310 20.330 159.610 ;
    END
  END E6END[7]
  PIN E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.670 19.410 160.970 ;
    END
  END E6END[8]
  PIN E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.710 13.430 163.010 ;
    END
  END E6END[9]
  PIN EE4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 208.290 119.190 223.275 119.490 ;
    END
  END EE4BEG[0]
  PIN EE4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 200.930 136.190 223.275 136.490 ;
    END
  END EE4BEG[10]
  PIN EE4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.590 138.230 223.275 138.530 ;
    END
  END EE4BEG[11]
  PIN EE4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 200.930 140.270 223.275 140.570 ;
    END
  END EE4BEG[12]
  PIN EE4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 200.470 141.630 223.275 141.930 ;
    END
  END EE4BEG[13]
  PIN EE4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 200.470 143.670 223.275 143.970 ;
    END
  END EE4BEG[14]
  PIN EE4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.850 145.030 223.275 145.330 ;
    END
  END EE4BEG[15]
  PIN EE4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.850 120.550 223.275 120.850 ;
    END
  END EE4BEG[1]
  PIN EE4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 193.110 122.590 223.275 122.890 ;
    END
  END EE4BEG[2]
  PIN EE4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.850 123.950 223.275 124.250 ;
    END
  END EE4BEG[3]
  PIN EE4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 199.090 125.990 223.275 126.290 ;
    END
  END EE4BEG[4]
  PIN EE4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.390 128.030 223.275 128.330 ;
    END
  END EE4BEG[5]
  PIN EE4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.750 129.390 223.275 129.690 ;
    END
  END EE4BEG[6]
  PIN EE4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 200.470 131.430 223.275 131.730 ;
    END
  END EE4BEG[7]
  PIN EE4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 202.310 132.790 223.275 133.090 ;
    END
  END EE4BEG[8]
  PIN EE4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 202.770 134.830 223.275 135.130 ;
    END
  END EE4BEG[9]
  PIN EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.190 7.450 119.490 ;
    END
  END EE4END[0]
  PIN EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.190 35.510 136.490 ;
    END
  END EE4END[10]
  PIN EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.230 18.700 138.530 ;
    END
  END EE4END[11]
  PIN EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.270 8.370 140.570 ;
    END
  END EE4END[12]
  PIN EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.630 7.050 141.930 ;
    END
  END EE4END[13]
  PIN EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.670 20.330 143.970 ;
    END
  END EE4END[14]
  PIN EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.030 21.710 145.330 ;
    END
  END EE4END[15]
  PIN EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.550 13.890 120.850 ;
    END
  END EE4END[1]
  PIN EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.590 16.650 122.890 ;
    END
  END EE4END[2]
  PIN EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.950 9.290 124.250 ;
    END
  END EE4END[3]
  PIN EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.990 34.130 126.290 ;
    END
  END EE4END[4]
  PIN EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.030 19.870 128.330 ;
    END
  END EE4END[5]
  PIN EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.390 13.430 129.690 ;
    END
  END EE4END[6]
  PIN EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.430 20.790 131.730 ;
    END
  END EE4END[7]
  PIN EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.790 18.700 133.090 ;
    END
  END EE4END[8]
  PIN EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.830 14.810 135.130 ;
    END
  END EE4END[9]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.150 6.990 168.450 ;
    END
  END FrameData[0]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.150 6.990 185.450 ;
    END
  END FrameData[10]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.190 6.990 187.490 ;
    END
  END FrameData[11]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 188.550 6.530 188.850 ;
    END
  END FrameData[12]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.590 6.990 190.890 ;
    END
  END FrameData[13]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.950 6.530 192.250 ;
    END
  END FrameData[14]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.990 7.450 194.290 ;
    END
  END FrameData[15]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.030 6.990 196.330 ;
    END
  END FrameData[16]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.390 6.530 197.690 ;
    END
  END FrameData[17]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.430 7.910 199.730 ;
    END
  END FrameData[18]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.790 18.950 201.090 ;
    END
  END FrameData[19]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 169.510 6.530 169.810 ;
    END
  END FrameData[1]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.830 7.450 203.130 ;
    END
  END FrameData[20]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.190 16.190 204.490 ;
    END
  END FrameData[21]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.230 6.530 206.530 ;
    END
  END FrameData[22]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.590 18.950 207.890 ;
    END
  END FrameData[23]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.630 6.990 209.930 ;
    END
  END FrameData[24]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 211.670 18.950 211.970 ;
    END
  END FrameData[25]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.030 16.190 213.330 ;
    END
  END FrameData[26]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.070 18.950 215.370 ;
    END
  END FrameData[27]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.430 14.810 216.730 ;
    END
  END FrameData[28]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 218.470 19.410 218.770 ;
    END
  END FrameData[29]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.550 6.990 171.850 ;
    END
  END FrameData[2]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.830 20.330 220.130 ;
    END
  END FrameData[30]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.870 20.330 222.170 ;
    END
  END FrameData[31]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.910 7.450 173.210 ;
    END
  END FrameData[3]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.950 6.530 175.250 ;
    END
  END FrameData[4]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.310 12.970 176.610 ;
    END
  END FrameData[5]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.350 16.190 178.650 ;
    END
  END FrameData[6]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.710 20.330 180.010 ;
    END
  END FrameData[7]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 181.750 19.870 182.050 ;
    END
  END FrameData[8]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.790 19.870 184.090 ;
    END
  END FrameData[9]
  PIN FrameData_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 168.150 223.275 168.450 ;
    END
  END FrameData_O[0]
  PIN FrameData_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 185.150 223.275 185.450 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 187.190 223.275 187.490 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.630 188.550 223.275 188.850 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 190.590 223.275 190.890 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.730 191.950 223.275 192.250 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 193.990 223.275 194.290 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 196.030 223.275 196.330 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 197.390 223.275 197.690 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 199.430 223.275 199.730 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 200.790 223.275 201.090 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 169.510 223.275 169.810 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.730 202.830 223.275 203.130 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.210 204.190 223.275 204.490 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 206.230 223.275 206.530 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.590 207.590 223.275 207.890 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.270 209.630 223.275 209.930 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 211.670 223.275 211.970 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.590 213.030 223.275 213.330 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.210 215.070 223.275 215.370 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 205.990 216.430 223.275 216.730 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 218.470 223.275 218.770 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.810 171.550 223.275 171.850 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.450 219.830 223.275 220.130 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 203.230 221.870 223.275 222.170 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 221.630 172.910 223.275 173.210 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 220.250 174.950 223.275 175.250 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.590 176.310 223.275 176.610 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.910 178.350 223.275 178.650 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 211.510 179.710 223.275 180.010 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.670 181.750 223.275 182.050 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.590 183.790 223.275 184.090 ;
    END
  END FrameData_O[9]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.300 0.000 188.440 6.500 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.780 0.000 205.920 11.940 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.620 0.000 207.760 9.560 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.460 0.000 209.600 17.040 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.300 0.000 211.440 15.000 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.680 0.000 212.820 8.570 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.520 0.000 214.660 6.160 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.360 0.000 216.500 22.820 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.200 0.000 218.340 16.700 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.040 0.000 220.180 3.780 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.880 0.000 222.020 6.500 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.680 0.000 189.820 11.940 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.520 0.000 191.660 15.000 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.360 0.000 193.500 5.850 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.200 0.000 195.340 20.440 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.040 0.000 197.180 22.820 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.880 0.000 199.020 9.220 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.260 0.000 200.400 25.880 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.100 0.000 202.240 13.980 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.940 0.000 204.080 13.870 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.840 216.880 187.980 223.115 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.780 217.190 205.920 223.115 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.620 208.720 207.760 223.115 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.000 215.830 209.140 223.115 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.840 217.220 210.980 223.115 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.680 211.780 212.820 223.115 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.520 209.060 214.660 223.115 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.360 213.820 216.500 223.115 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.200 203.280 218.340 223.115 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.040 202.940 220.180 223.115 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.880 219.940 222.020 223.115 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.680 213.820 189.820 223.115 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.520 211.780 191.660 223.115 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.360 209.060 193.500 223.115 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.740 213.140 194.880 223.115 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.580 206.340 196.720 223.115 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.420 206.340 198.560 223.115 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.260 203.620 200.400 223.115 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.100 200.220 202.240 223.115 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.940 211.750 204.080 223.115 ;
    END
  END FrameStrobe_O[9]
  PIN N1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.620 206.340 0.760 223.115 ;
    END
  END N1BEG[0]
  PIN N1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.000 204.980 2.140 223.115 ;
    END
  END N1BEG[1]
  PIN N1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.840 199.880 3.980 223.115 ;
    END
  END N1BEG[2]
  PIN N1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.680 206.000 5.820 223.115 ;
    END
  END N1BEG[3]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.620 0.000 0.760 11.600 ;
    END
  END N1END[0]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.000 0.000 2.140 17.380 ;
    END
  END N1END[1]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.840 0.000 3.980 6.500 ;
    END
  END N1END[2]
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.680 0.000 5.820 11.940 ;
    END
  END N1END[3]
  PIN N2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.520 215.520 7.660 223.115 ;
    END
  END N2BEG[0]
  PIN N2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.360 200.900 9.500 223.115 ;
    END
  END N2BEG[1]
  PIN N2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.200 204.640 11.340 223.115 ;
    END
  END N2BEG[2]
  PIN N2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.040 213.790 13.180 223.115 ;
    END
  END N2BEG[3]
  PIN N2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.880 218.920 15.020 223.115 ;
    END
  END N2BEG[4]
  PIN N2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.260 217.870 16.400 223.115 ;
    END
  END N2BEG[5]
  PIN N2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.100 213.820 18.240 223.115 ;
    END
  END N2BEG[6]
  PIN N2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.940 219.940 20.080 223.115 ;
    END
  END N2BEG[7]
  PIN N2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.780 221.950 21.920 223.115 ;
    END
  END N2BEGb[0]
  PIN N2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.620 216.510 23.760 223.115 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.460 221.950 25.600 223.115 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.300 219.600 27.440 223.115 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.140 216.340 29.280 223.115 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.520 217.870 30.660 223.115 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.360 203.620 32.500 223.115 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.200 218.580 34.340 223.115 ;
    END
  END N2BEGb[7]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.780 0.000 21.920 6.500 ;
    END
  END N2END[0]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.620 0.000 23.760 5.820 ;
    END
  END N2END[1]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.000 0.000 25.140 7.210 ;
    END
  END N2END[2]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.840 0.000 26.980 9.220 ;
    END
  END N2END[3]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.680 0.000 28.820 4.800 ;
    END
  END N2END[4]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.520 0.000 30.660 5.820 ;
    END
  END N2END[5]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.360 0.000 32.500 11.600 ;
    END
  END N2END[6]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.200 0.000 34.340 9.560 ;
    END
  END N2END[7]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.520 0.000 7.660 13.870 ;
    END
  END N2MID[0]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.360 0.000 9.500 20.440 ;
    END
  END N2MID[1]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.200 0.000 11.340 4.490 ;
    END
  END N2MID[2]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.580 0.000 12.720 15.340 ;
    END
  END N2MID[3]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.420 0.000 14.560 17.380 ;
    END
  END N2MID[4]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.260 0.000 16.400 6.500 ;
    END
  END N2MID[5]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.100 0.000 18.240 1.060 ;
    END
  END N2MID[6]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.940 0.000 20.080 7.520 ;
    END
  END N2MID[7]
  PIN N4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.040 202.910 36.180 223.115 ;
    END
  END N4BEG[0]
  PIN N4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.980 218.550 54.120 223.115 ;
    END
  END N4BEG[10]
  PIN N4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.820 219.600 55.960 223.115 ;
    END
  END N4BEG[11]
  PIN N4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.660 211.780 57.800 223.115 ;
    END
  END N4BEG[12]
  PIN N4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.500 213.820 59.640 223.115 ;
    END
  END N4BEG[13]
  PIN N4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.880 211.780 61.020 223.115 ;
    END
  END N4BEG[14]
  PIN N4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.720 216.680 62.860 223.115 ;
    END
  END N4BEG[15]
  PIN N4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.880 221.300 38.020 223.115 ;
    END
  END N4BEG[1]
  PIN N4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.720 221.950 39.860 223.115 ;
    END
  END N4BEG[2]
  PIN N4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.560 220.280 41.700 223.115 ;
    END
  END N4BEG[3]
  PIN N4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.400 221.950 43.540 223.115 ;
    END
  END N4BEG[4]
  PIN N4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.240 217.190 45.380 223.115 ;
    END
  END N4BEG[5]
  PIN N4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.620 220.280 46.760 223.115 ;
    END
  END N4BEG[6]
  PIN N4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.460 205.160 48.600 223.115 ;
    END
  END N4BEG[7]
  PIN N4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.300 215.860 50.440 223.115 ;
    END
  END N4BEG[8]
  PIN N4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.140 217.190 52.280 223.115 ;
    END
  END N4BEG[9]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.580 0.000 35.720 6.500 ;
    END
  END N4END[0]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.520 0.000 53.660 15.000 ;
    END
  END N4END[10]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.360 0.000 55.500 20.780 ;
    END
  END N4END[11]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.200 0.000 57.340 13.870 ;
    END
  END N4END[12]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.040 0.000 59.180 3.130 ;
    END
  END N4END[13]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.420 0.000 60.560 1.090 ;
    END
  END N4END[14]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.260 0.000 62.400 4.120 ;
    END
  END N4END[15]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.420 0.000 37.560 17.380 ;
    END
  END N4END[1]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.260 0.000 39.400 9.220 ;
    END
  END N4END[2]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.100 0.000 41.240 6.500 ;
    END
  END N4END[3]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.940 0.000 43.080 17.040 ;
    END
  END N4END[4]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.780 0.000 44.920 9.040 ;
    END
  END N4END[5]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.620 0.000 46.760 13.980 ;
    END
  END N4END[6]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.000 0.000 48.140 1.090 ;
    END
  END N4END[7]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.840 0.000 49.980 1.090 ;
    END
  END N4END[8]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.680 0.000 51.820 29.440 ;
    END
  END N4END[9]
  PIN NN4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.560 216.510 64.700 223.115 ;
    END
  END NN4BEG[0]
  PIN NN4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.500 217.220 82.640 223.115 ;
    END
  END NN4BEG[10]
  PIN NN4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.340 214.500 84.480 223.115 ;
    END
  END NN4BEG[11]
  PIN NN4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.180 213.820 86.320 223.115 ;
    END
  END NN4BEG[12]
  PIN NN4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.020 211.440 88.160 223.115 ;
    END
  END NN4BEG[13]
  PIN NN4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.860 209.060 90.000 223.115 ;
    END
  END NN4BEG[14]
  PIN NN4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.240 214.160 91.380 223.115 ;
    END
  END NN4BEG[15]
  PIN NN4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.400 213.820 66.540 223.115 ;
    END
  END NN4BEG[1]
  PIN NN4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.240 210.080 68.380 223.115 ;
    END
  END NN4BEG[2]
  PIN NN4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.080 221.950 70.220 223.115 ;
    END
  END NN4BEG[3]
  PIN NN4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.920 209.060 72.060 223.115 ;
    END
  END NN4BEG[4]
  PIN NN4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.760 207.360 73.900 223.115 ;
    END
  END NN4BEG[5]
  PIN NN4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.140 212.800 75.280 223.115 ;
    END
  END NN4BEG[6]
  PIN NN4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.980 206.340 77.120 223.115 ;
    END
  END NN4BEG[7]
  PIN NN4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.820 221.950 78.960 223.115 ;
    END
  END NN4BEG[8]
  PIN NN4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.660 211.440 80.800 223.115 ;
    END
  END NN4BEG[9]
  PIN NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.100 0.000 64.240 6.160 ;
    END
  END NN4END[0]
  PIN NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.040 0.000 82.180 6.020 ;
    END
  END NN4END[10]
  PIN NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.420 0.000 83.560 36.760 ;
    END
  END NN4END[11]
  PIN NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.260 0.000 85.400 5.850 ;
    END
  END NN4END[12]
  PIN NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.100 0.000 87.240 4.960 ;
    END
  END NN4END[13]
  PIN NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.940 0.000 89.080 13.870 ;
    END
  END NN4END[14]
  PIN NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.780 0.000 90.920 44.580 ;
    END
  END NN4END[15]
  PIN NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.940 0.000 66.080 6.160 ;
    END
  END NN4END[1]
  PIN NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.780 0.000 67.920 11.600 ;
    END
  END NN4END[2]
  PIN NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.620 0.000 69.760 15.340 ;
    END
  END NN4END[3]
  PIN NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.000 0.000 71.140 39.140 ;
    END
  END NN4END[4]
  PIN NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.840 0.000 72.980 19.920 ;
    END
  END NN4END[5]
  PIN NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.680 0.000 74.820 12.650 ;
    END
  END NN4END[6]
  PIN NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.520 0.000 76.660 47.640 ;
    END
  END NN4END[7]
  PIN NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.360 0.000 78.500 50.020 ;
    END
  END NN4END[8]
  PIN NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.200 0.000 80.340 7.180 ;
    END
  END NN4END[9]
  PIN S1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.620 0.000 92.760 6.160 ;
    END
  END S1BEG[0]
  PIN S1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.460 0.000 94.600 8.540 ;
    END
  END S1BEG[1]
  PIN S1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.840 0.000 95.980 4.490 ;
    END
  END S1BEG[2]
  PIN S1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.680 0.000 97.820 4.460 ;
    END
  END S1BEG[3]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.080 219.230 93.220 223.115 ;
    END
  END S1END[0]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.920 216.540 95.060 223.115 ;
    END
  END S1END[1]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.760 213.480 96.900 223.115 ;
    END
  END S1END[2]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.600 221.950 98.740 223.115 ;
    END
  END S1END[3]
  PIN S2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.780 0.000 113.920 3.130 ;
    END
  END S2BEG[0]
  PIN S2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.620 0.000 115.760 6.160 ;
    END
  END S2BEG[1]
  PIN S2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.460 0.000 117.600 3.130 ;
    END
  END S2BEG[2]
  PIN S2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.840 0.000 118.980 11.260 ;
    END
  END S2BEG[3]
  PIN S2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.680 0.000 120.820 2.760 ;
    END
  END S2BEG[4]
  PIN S2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.520 0.000 122.660 2.420 ;
    END
  END S2BEG[5]
  PIN S2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.360 0.000 124.500 4.490 ;
    END
  END S2BEG[6]
  PIN S2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.200 0.000 126.340 3.780 ;
    END
  END S2BEG[7]
  PIN S2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.520 0.000 99.660 4.490 ;
    END
  END S2BEGb[0]
  PIN S2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.360 0.000 101.500 17.040 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.200 0.000 103.340 19.420 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.040 0.000 105.180 14.180 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.420 0.000 106.560 1.090 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.260 0.000 108.400 7.210 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.100 0.000 110.240 17.040 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.940 0.000 112.080 18.400 ;
    END
  END S2BEGb[7]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.440 211.100 100.580 223.115 ;
    END
  END S2END[0]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.280 219.230 102.420 223.115 ;
    END
  END S2END[1]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.120 213.140 104.260 223.115 ;
    END
  END S2END[2]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.500 217.220 105.640 223.115 ;
    END
  END S2END[3]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.340 211.100 107.480 223.115 ;
    END
  END S2END[4]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.180 221.950 109.320 223.115 ;
    END
  END S2END[5]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.020 221.950 111.160 223.115 ;
    END
  END S2END[6]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.860 213.140 113.000 223.115 ;
    END
  END S2END[7]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.700 211.440 114.840 223.115 ;
    END
  END S2MID[0]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.540 208.040 116.680 223.115 ;
    END
  END S2MID[1]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.380 208.380 118.520 223.115 ;
    END
  END S2MID[2]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.760 216.880 119.900 223.115 ;
    END
  END S2MID[3]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.600 217.220 121.740 223.115 ;
    END
  END S2MID[4]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.440 213.480 123.580 223.115 ;
    END
  END S2MID[5]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.280 213.110 125.420 223.115 ;
    END
  END S2MID[6]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.120 203.620 127.260 223.115 ;
    END
  END S2MID[7]
  PIN S4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.040 0.000 128.180 2.080 ;
    END
  END S4BEG[0]
  PIN S4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.520 0.000 145.660 8.540 ;
    END
  END S4BEG[10]
  PIN S4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.360 0.000 147.500 11.260 ;
    END
  END S4BEG[11]
  PIN S4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.200 0.000 149.340 1.090 ;
    END
  END S4BEG[12]
  PIN S4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.040 0.000 151.180 11.940 ;
    END
  END S4BEG[13]
  PIN S4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.880 0.000 153.020 5.820 ;
    END
  END S4BEG[14]
  PIN S4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.260 0.000 154.400 8.540 ;
    END
  END S4BEG[15]
  PIN S4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.420 0.000 129.560 7.210 ;
    END
  END S4BEG[1]
  PIN S4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.260 0.000 131.400 16.700 ;
    END
  END S4BEG[2]
  PIN S4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.100 0.000 133.240 25.200 ;
    END
  END S4BEG[3]
  PIN S4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.940 0.000 135.080 17.040 ;
    END
  END S4BEG[4]
  PIN S4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.780 0.000 136.920 18.060 ;
    END
  END S4BEG[5]
  PIN S4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.620 0.000 138.760 1.400 ;
    END
  END S4BEG[6]
  PIN S4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.460 0.000 140.600 16.700 ;
    END
  END S4BEG[7]
  PIN S4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.840 0.000 141.980 19.420 ;
    END
  END S4BEG[8]
  PIN S4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.680 0.000 143.820 8.360 ;
    END
  END S4BEG[9]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.960 205.660 129.100 223.115 ;
    END
  END S4END[0]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.900 194.920 147.040 223.115 ;
    END
  END S4END[10]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.740 211.280 148.880 223.115 ;
    END
  END S4END[11]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.120 213.140 150.260 223.115 ;
    END
  END S4END[12]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.960 214.470 152.100 223.115 ;
    END
  END S4END[13]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.800 204.440 153.940 223.115 ;
    END
  END S4END[14]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.640 214.470 155.780 223.115 ;
    END
  END S4END[15]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.800 221.950 130.940 223.115 ;
    END
  END S4END[1]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.640 206.340 132.780 223.115 ;
    END
  END S4END[2]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.480 221.300 134.620 223.115 ;
    END
  END S4END[3]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.860 221.950 136.000 223.115 ;
    END
  END S4END[4]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.700 200.560 137.840 223.115 ;
    END
  END S4END[5]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.540 201.920 139.680 223.115 ;
    END
  END S4END[6]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.380 214.470 141.520 223.115 ;
    END
  END S4END[7]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.220 218.580 143.360 223.115 ;
    END
  END S4END[8]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.060 220.960 145.200 223.115 ;
    END
  END S4END[9]
  PIN SS4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.100 0.000 156.240 14.320 ;
    END
  END SS4BEG[0]
  PIN SS4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.040 0.000 174.180 12.620 ;
    END
  END SS4BEG[10]
  PIN SS4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.880 0.000 176.020 3.130 ;
    END
  END SS4BEG[11]
  PIN SS4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.260 0.000 177.400 7.210 ;
    END
  END SS4BEG[12]
  PIN SS4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.100 0.000 179.240 12.960 ;
    END
  END SS4BEG[13]
  PIN SS4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.940 0.000 181.080 16.700 ;
    END
  END SS4BEG[14]
  PIN SS4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.780 0.000 182.920 7.210 ;
    END
  END SS4BEG[15]
  PIN SS4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.940 0.000 158.080 1.090 ;
    END
  END SS4BEG[1]
  PIN SS4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.780 0.000 159.920 0.920 ;
    END
  END SS4BEG[2]
  PIN SS4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.620 0.000 161.760 8.360 ;
    END
  END SS4BEG[3]
  PIN SS4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.460 0.000 163.600 9.720 ;
    END
  END SS4BEG[4]
  PIN SS4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.840 0.000 164.980 10.400 ;
    END
  END SS4BEG[5]
  PIN SS4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.680 0.000 166.820 7.210 ;
    END
  END SS4BEG[6]
  PIN SS4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.520 0.000 168.660 16.520 ;
    END
  END SS4BEG[7]
  PIN SS4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.360 0.000 170.500 0.920 ;
    END
  END SS4BEG[8]
  PIN SS4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.200 0.000 172.340 13.800 ;
    END
  END SS4BEG[9]
  PIN SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.480 216.540 157.620 223.115 ;
    END
  END SS4END[0]
  PIN SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.420 215.860 175.560 223.115 ;
    END
  END SS4END[10]
  PIN SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.260 217.400 177.400 223.115 ;
    END
  END SS4END[11]
  PIN SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.100 218.580 179.240 223.115 ;
    END
  END SS4END[12]
  PIN SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.480 209.920 180.620 223.115 ;
    END
  END SS4END[13]
  PIN SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.320 205.660 182.460 223.115 ;
    END
  END SS4END[14]
  PIN SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.160 139.880 184.300 223.115 ;
    END
  END SS4END[15]
  PIN SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.320 213.140 159.460 223.115 ;
    END
  END SS4END[1]
  PIN SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.160 216.540 161.300 223.115 ;
    END
  END SS4END[2]
  PIN SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.000 207.670 163.140 223.115 ;
    END
  END SS4END[3]
  PIN SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.380 212.800 164.520 223.115 ;
    END
  END SS4END[4]
  PIN SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.220 214.470 166.360 223.115 ;
    END
  END SS4END[5]
  PIN SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.060 214.470 168.200 223.115 ;
    END
  END SS4END[6]
  PIN SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.900 221.950 170.040 223.115 ;
    END
  END SS4END[7]
  PIN SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.740 214.470 171.880 223.115 ;
    END
  END SS4END[8]
  PIN SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.580 214.300 173.720 223.115 ;
    END
  END SS4END[9]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.620 0.000 184.760 10.400 ;
    END
  END UserCLK
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 5.200 99.440 217.840 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 5.200 22.640 217.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 5.200 176.240 217.840 ;
    END
  END VPWR
  PIN W1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.870 15.270 1.170 ;
    END
  END W1BEG[0]
  PIN W1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.230 9.750 2.530 ;
    END
  END W1BEG[1]
  PIN W1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.270 18.950 4.570 ;
    END
  END W1BEG[2]
  PIN W1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.630 13.890 5.930 ;
    END
  END W1BEG[3]
  PIN W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 202.770 0.870 223.275 1.170 ;
    END
  END W1END[0]
  PIN W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 200.930 2.230 223.275 2.530 ;
    END
  END W1END[1]
  PIN W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 200.010 4.270 223.275 4.570 ;
    END
  END W1END[2]
  PIN W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 200.930 5.630 223.275 5.930 ;
    END
  END W1END[3]
  PIN W2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.670 15.730 7.970 ;
    END
  END W2BEG[0]
  PIN W2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.030 16.190 9.330 ;
    END
  END W2BEG[1]
  PIN W2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.070 18.490 11.370 ;
    END
  END W2BEG[2]
  PIN W2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.430 19.410 12.730 ;
    END
  END W2BEG[3]
  PIN W2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.470 20.330 14.770 ;
    END
  END W2BEG[4]
  PIN W2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.510 14.810 16.810 ;
    END
  END W2BEG[5]
  PIN W2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.870 10.210 18.170 ;
    END
  END W2BEG[6]
  PIN W2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.910 18.950 20.210 ;
    END
  END W2BEG[7]
  PIN W2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.270 6.990 21.570 ;
    END
  END W2BEGb[0]
  PIN W2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.310 19.410 23.610 ;
    END
  END W2BEGb[1]
  PIN W2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.670 7.450 24.970 ;
    END
  END W2BEGb[2]
  PIN W2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.710 19.700 27.010 ;
    END
  END W2BEGb[3]
  PIN W2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.750 14.350 29.050 ;
    END
  END W2BEGb[4]
  PIN W2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.110 1.470 30.410 ;
    END
  END W2BEGb[5]
  PIN W2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.150 20.330 32.450 ;
    END
  END W2BEGb[6]
  PIN W2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.510 9.750 33.810 ;
    END
  END W2BEGb[7]
  PIN W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 212.890 21.270 223.275 21.570 ;
    END
  END W2END[0]
  PIN W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 212.430 23.310 223.275 23.610 ;
    END
  END W2END[1]
  PIN W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 200.930 24.670 223.275 24.970 ;
    END
  END W2END[2]
  PIN W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.850 26.710 223.275 27.010 ;
    END
  END W2END[3]
  PIN W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.450 28.750 223.275 29.050 ;
    END
  END W2END[4]
  PIN W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.910 30.110 223.275 30.410 ;
    END
  END W2END[5]
  PIN W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 212.890 32.150 223.275 32.450 ;
    END
  END W2END[6]
  PIN W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 205.990 33.510 223.275 33.810 ;
    END
  END W2END[7]
  PIN W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 200.930 7.670 223.275 7.970 ;
    END
  END W2MID[0]
  PIN W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 212.890 9.030 223.275 9.330 ;
    END
  END W2MID[1]
  PIN W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 205.070 11.070 223.275 11.370 ;
    END
  END W2MID[2]
  PIN W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 205.530 12.430 223.275 12.730 ;
    END
  END W2MID[3]
  PIN W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.390 14.470 223.275 14.770 ;
    END
  END W2MID[4]
  PIN W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 200.930 16.510 223.275 16.810 ;
    END
  END W2MID[5]
  PIN W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 200.010 17.870 223.275 18.170 ;
    END
  END W2MID[6]
  PIN W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.850 19.910 223.275 20.210 ;
    END
  END W2MID[7]
  PIN W6BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.430 10.210 63.730 ;
    END
  END W6BEG[0]
  PIN W6BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.430 9.750 80.730 ;
    END
  END W6BEG[10]
  PIN W6BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.470 14.350 82.770 ;
    END
  END W6BEG[11]
  PIN W6BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.790 9.750 65.090 ;
    END
  END W6BEG[1]
  PIN W6BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.830 13.890 67.130 ;
    END
  END W6BEG[2]
  PIN W6BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.190 16.650 68.490 ;
    END
  END W6BEG[3]
  PIN W6BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.230 18.950 70.530 ;
    END
  END W6BEG[4]
  PIN W6BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.270 25.390 72.570 ;
    END
  END W6BEG[5]
  PIN W6BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.630 17.110 73.930 ;
    END
  END W6BEG[6]
  PIN W6BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.670 18.490 75.970 ;
    END
  END W6BEG[7]
  PIN W6BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.030 7.050 77.330 ;
    END
  END W6BEG[8]
  PIN W6BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.070 20.330 79.370 ;
    END
  END W6BEG[9]
  PIN W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 211.970 63.430 223.275 63.730 ;
    END
  END W6END[0]
  PIN W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 197.250 80.430 223.275 80.730 ;
    END
  END W6END[10]
  PIN W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 200.930 82.470 223.275 82.770 ;
    END
  END W6END[11]
  PIN W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 202.770 64.790 223.275 65.090 ;
    END
  END W6END[1]
  PIN W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.850 66.830 223.275 67.130 ;
    END
  END W6END[2]
  PIN W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 200.470 68.190 223.275 68.490 ;
    END
  END W6END[3]
  PIN W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 168.270 70.230 223.275 70.530 ;
    END
  END W6END[4]
  PIN W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.670 72.270 223.275 72.570 ;
    END
  END W6END[5]
  PIN W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.670 73.630 223.275 73.930 ;
    END
  END W6END[6]
  PIN W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 200.470 75.670 223.275 75.970 ;
    END
  END W6END[7]
  PIN W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.390 77.030 223.275 77.330 ;
    END
  END W6END[8]
  PIN W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 203.690 79.070 223.275 79.370 ;
    END
  END W6END[9]
  PIN WW4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.550 16.650 35.850 ;
    END
  END WW4BEG[0]
  PIN WW4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.550 6.990 52.850 ;
    END
  END WW4BEG[10]
  PIN WW4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.590 19.870 54.890 ;
    END
  END WW4BEG[11]
  PIN WW4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.630 13.890 56.930 ;
    END
  END WW4BEG[12]
  PIN WW4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.990 20.330 58.290 ;
    END
  END WW4BEG[13]
  PIN WW4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.030 23.090 60.330 ;
    END
  END WW4BEG[14]
  PIN WW4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.390 23.090 61.690 ;
    END
  END WW4BEG[15]
  PIN WW4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.910 24.010 37.210 ;
    END
  END WW4BEG[1]
  PIN WW4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.950 17.110 39.250 ;
    END
  END WW4BEG[2]
  PIN WW4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.310 20.330 40.610 ;
    END
  END WW4BEG[3]
  PIN WW4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.350 20.330 42.650 ;
    END
  END WW4BEG[4]
  PIN WW4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.390 18.490 44.690 ;
    END
  END WW4BEG[5]
  PIN WW4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.750 20.330 46.050 ;
    END
  END WW4BEG[6]
  PIN WW4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.790 20.330 48.090 ;
    END
  END WW4BEG[7]
  PIN WW4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.150 18.950 49.450 ;
    END
  END WW4BEG[8]
  PIN WW4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.190 20.330 51.490 ;
    END
  END WW4BEG[9]
  PIN WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 211.510 35.550 223.275 35.850 ;
    END
  END WW4END[0]
  PIN WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 200.470 52.550 223.275 52.850 ;
    END
  END WW4END[10]
  PIN WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 200.470 54.590 223.275 54.890 ;
    END
  END WW4END[11]
  PIN WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 202.310 56.630 223.275 56.930 ;
    END
  END WW4END[12]
  PIN WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.750 57.990 223.275 58.290 ;
    END
  END WW4END[13]
  PIN WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 219.790 60.030 223.275 60.330 ;
    END
  END WW4END[14]
  PIN WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 194.030 61.390 223.275 61.690 ;
    END
  END WW4END[15]
  PIN WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.070 36.910 223.275 37.210 ;
    END
  END WW4END[1]
  PIN WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.390 38.950 223.275 39.250 ;
    END
  END WW4END[2]
  PIN WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.850 40.310 223.275 40.610 ;
    END
  END WW4END[3]
  PIN WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 190.140 42.350 223.275 42.650 ;
    END
  END WW4END[4]
  PIN WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 203.690 44.390 223.275 44.690 ;
    END
  END WW4END[5]
  PIN WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 200.470 45.750 223.275 46.050 ;
    END
  END WW4END[6]
  PIN WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 199.950 47.790 223.275 48.090 ;
    END
  END WW4END[7]
  PIN WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 210.590 49.150 223.275 49.450 ;
    END
  END WW4END[8]
  PIN WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 200.470 51.190 223.275 51.490 ;
    END
  END WW4END[9]
  OBS
      LAYER li1 ;
        RECT 5.520 0.765 222.955 220.235 ;
      LAYER met1 ;
        RECT 0.530 0.720 223.030 222.320 ;
      LAYER met2 ;
        RECT 1.040 206.060 1.720 222.770 ;
        RECT 0.560 204.700 1.720 206.060 ;
        RECT 2.420 204.700 3.560 222.770 ;
        RECT 0.560 199.600 3.560 204.700 ;
        RECT 4.260 205.720 5.400 222.770 ;
        RECT 6.100 215.240 7.240 222.770 ;
        RECT 7.940 215.240 9.080 222.770 ;
        RECT 6.100 205.720 9.080 215.240 ;
        RECT 4.260 200.620 9.080 205.720 ;
        RECT 9.780 204.360 10.920 222.770 ;
        RECT 11.620 213.510 12.760 222.770 ;
        RECT 13.460 218.640 14.600 222.770 ;
        RECT 15.300 218.640 15.980 222.770 ;
        RECT 13.460 217.590 15.980 218.640 ;
        RECT 16.680 217.590 17.820 222.770 ;
        RECT 13.460 213.540 17.820 217.590 ;
        RECT 18.520 219.660 19.660 222.770 ;
        RECT 20.360 221.670 21.500 222.770 ;
        RECT 22.200 221.670 23.340 222.770 ;
        RECT 20.360 219.660 23.340 221.670 ;
        RECT 18.520 216.230 23.340 219.660 ;
        RECT 24.040 221.670 25.180 222.770 ;
        RECT 25.880 221.670 27.020 222.770 ;
        RECT 24.040 219.320 27.020 221.670 ;
        RECT 27.720 219.320 28.860 222.770 ;
        RECT 24.040 216.230 28.860 219.320 ;
        RECT 18.520 216.060 28.860 216.230 ;
        RECT 29.560 217.590 30.240 222.770 ;
        RECT 30.940 217.590 32.080 222.770 ;
        RECT 29.560 216.060 32.080 217.590 ;
        RECT 18.520 213.540 32.080 216.060 ;
        RECT 13.460 213.510 32.080 213.540 ;
        RECT 11.620 204.360 32.080 213.510 ;
        RECT 9.780 203.340 32.080 204.360 ;
        RECT 32.780 218.300 33.920 222.770 ;
        RECT 34.620 218.300 35.760 222.770 ;
        RECT 32.780 203.340 35.760 218.300 ;
        RECT 9.780 202.630 35.760 203.340 ;
        RECT 36.460 221.020 37.600 222.770 ;
        RECT 38.300 221.670 39.440 222.770 ;
        RECT 40.140 221.670 41.280 222.770 ;
        RECT 38.300 221.020 41.280 221.670 ;
        RECT 36.460 220.000 41.280 221.020 ;
        RECT 41.980 221.670 43.120 222.770 ;
        RECT 43.820 221.670 44.960 222.770 ;
        RECT 41.980 220.000 44.960 221.670 ;
        RECT 36.460 216.910 44.960 220.000 ;
        RECT 45.660 220.000 46.340 222.770 ;
        RECT 47.040 220.000 48.180 222.770 ;
        RECT 45.660 216.910 48.180 220.000 ;
        RECT 36.460 204.880 48.180 216.910 ;
        RECT 48.880 215.580 50.020 222.770 ;
        RECT 50.720 216.910 51.860 222.770 ;
        RECT 52.560 218.270 53.700 222.770 ;
        RECT 54.400 219.320 55.540 222.770 ;
        RECT 56.240 219.320 57.380 222.770 ;
        RECT 54.400 218.270 57.380 219.320 ;
        RECT 52.560 216.910 57.380 218.270 ;
        RECT 50.720 215.580 57.380 216.910 ;
        RECT 48.880 211.500 57.380 215.580 ;
        RECT 58.080 213.540 59.220 222.770 ;
        RECT 59.920 213.540 60.600 222.770 ;
        RECT 58.080 211.500 60.600 213.540 ;
        RECT 61.300 216.400 62.440 222.770 ;
        RECT 63.140 216.400 64.280 222.770 ;
        RECT 61.300 216.230 64.280 216.400 ;
        RECT 64.980 216.230 66.120 222.770 ;
        RECT 61.300 213.540 66.120 216.230 ;
        RECT 66.820 213.540 67.960 222.770 ;
        RECT 61.300 211.500 67.960 213.540 ;
        RECT 48.880 209.800 67.960 211.500 ;
        RECT 68.660 221.670 69.800 222.770 ;
        RECT 70.500 221.670 71.640 222.770 ;
        RECT 68.660 209.800 71.640 221.670 ;
        RECT 48.880 208.780 71.640 209.800 ;
        RECT 72.340 208.780 73.480 222.770 ;
        RECT 48.880 207.080 73.480 208.780 ;
        RECT 74.180 212.520 74.860 222.770 ;
        RECT 75.560 212.520 76.700 222.770 ;
        RECT 74.180 207.080 76.700 212.520 ;
        RECT 48.880 206.060 76.700 207.080 ;
        RECT 77.400 221.670 78.540 222.770 ;
        RECT 79.240 221.670 80.380 222.770 ;
        RECT 77.400 211.160 80.380 221.670 ;
        RECT 81.080 216.940 82.220 222.770 ;
        RECT 82.920 216.940 84.060 222.770 ;
        RECT 81.080 214.220 84.060 216.940 ;
        RECT 84.760 214.220 85.900 222.770 ;
        RECT 81.080 213.540 85.900 214.220 ;
        RECT 86.600 213.540 87.740 222.770 ;
        RECT 81.080 211.160 87.740 213.540 ;
        RECT 88.440 211.160 89.580 222.770 ;
        RECT 77.400 208.780 89.580 211.160 ;
        RECT 90.280 213.880 90.960 222.770 ;
        RECT 91.660 218.950 92.800 222.770 ;
        RECT 93.500 218.950 94.640 222.770 ;
        RECT 91.660 216.260 94.640 218.950 ;
        RECT 95.340 216.260 96.480 222.770 ;
        RECT 91.660 213.880 96.480 216.260 ;
        RECT 90.280 213.200 96.480 213.880 ;
        RECT 97.180 221.670 98.320 222.770 ;
        RECT 99.020 221.670 100.160 222.770 ;
        RECT 97.180 213.200 100.160 221.670 ;
        RECT 90.280 210.820 100.160 213.200 ;
        RECT 100.860 218.950 102.000 222.770 ;
        RECT 102.700 218.950 103.840 222.770 ;
        RECT 100.860 212.860 103.840 218.950 ;
        RECT 104.540 216.940 105.220 222.770 ;
        RECT 105.920 216.940 107.060 222.770 ;
        RECT 104.540 212.860 107.060 216.940 ;
        RECT 100.860 210.820 107.060 212.860 ;
        RECT 107.760 221.670 108.900 222.770 ;
        RECT 109.600 221.670 110.740 222.770 ;
        RECT 111.440 221.670 112.580 222.770 ;
        RECT 107.760 212.860 112.580 221.670 ;
        RECT 113.280 212.860 114.420 222.770 ;
        RECT 107.760 211.160 114.420 212.860 ;
        RECT 115.120 211.160 116.260 222.770 ;
        RECT 107.760 210.820 116.260 211.160 ;
        RECT 90.280 208.780 116.260 210.820 ;
        RECT 77.400 207.760 116.260 208.780 ;
        RECT 116.960 208.100 118.100 222.770 ;
        RECT 118.800 216.600 119.480 222.770 ;
        RECT 120.180 216.940 121.320 222.770 ;
        RECT 122.020 216.940 123.160 222.770 ;
        RECT 120.180 216.600 123.160 216.940 ;
        RECT 118.800 213.200 123.160 216.600 ;
        RECT 123.860 213.200 125.000 222.770 ;
        RECT 118.800 212.830 125.000 213.200 ;
        RECT 125.700 212.830 126.840 222.770 ;
        RECT 118.800 208.100 126.840 212.830 ;
        RECT 116.960 207.760 126.840 208.100 ;
        RECT 77.400 206.060 126.840 207.760 ;
        RECT 48.880 204.880 126.840 206.060 ;
        RECT 36.460 203.340 126.840 204.880 ;
        RECT 127.540 205.380 128.680 222.770 ;
        RECT 129.380 221.670 130.520 222.770 ;
        RECT 131.220 221.670 132.360 222.770 ;
        RECT 129.380 206.060 132.360 221.670 ;
        RECT 133.060 221.020 134.200 222.770 ;
        RECT 134.900 221.670 135.580 222.770 ;
        RECT 136.280 221.670 137.420 222.770 ;
        RECT 134.900 221.020 137.420 221.670 ;
        RECT 133.060 206.060 137.420 221.020 ;
        RECT 129.380 205.380 137.420 206.060 ;
        RECT 127.540 203.340 137.420 205.380 ;
        RECT 36.460 202.630 137.420 203.340 ;
        RECT 9.780 200.620 137.420 202.630 ;
        RECT 4.260 200.280 137.420 200.620 ;
        RECT 138.120 201.640 139.260 222.770 ;
        RECT 139.960 214.190 141.100 222.770 ;
        RECT 141.800 218.300 142.940 222.770 ;
        RECT 143.640 220.680 144.780 222.770 ;
        RECT 145.480 220.680 146.620 222.770 ;
        RECT 143.640 218.300 146.620 220.680 ;
        RECT 141.800 214.190 146.620 218.300 ;
        RECT 139.960 201.640 146.620 214.190 ;
        RECT 138.120 200.280 146.620 201.640 ;
        RECT 4.260 199.600 146.620 200.280 ;
        RECT 0.560 194.640 146.620 199.600 ;
        RECT 147.320 211.000 148.460 222.770 ;
        RECT 149.160 212.860 149.840 222.770 ;
        RECT 150.540 214.190 151.680 222.770 ;
        RECT 152.380 214.190 153.520 222.770 ;
        RECT 150.540 212.860 153.520 214.190 ;
        RECT 149.160 211.000 153.520 212.860 ;
        RECT 147.320 204.160 153.520 211.000 ;
        RECT 154.220 214.190 155.360 222.770 ;
        RECT 156.060 216.260 157.200 222.770 ;
        RECT 157.900 216.260 159.040 222.770 ;
        RECT 156.060 214.190 159.040 216.260 ;
        RECT 154.220 212.860 159.040 214.190 ;
        RECT 159.740 216.260 160.880 222.770 ;
        RECT 161.580 216.260 162.720 222.770 ;
        RECT 159.740 212.860 162.720 216.260 ;
        RECT 154.220 207.390 162.720 212.860 ;
        RECT 163.420 212.520 164.100 222.770 ;
        RECT 164.800 214.190 165.940 222.770 ;
        RECT 166.640 214.190 167.780 222.770 ;
        RECT 168.480 221.670 169.620 222.770 ;
        RECT 170.320 221.670 171.460 222.770 ;
        RECT 168.480 214.190 171.460 221.670 ;
        RECT 172.160 214.190 173.300 222.770 ;
        RECT 164.800 214.020 173.300 214.190 ;
        RECT 174.000 215.580 175.140 222.770 ;
        RECT 175.840 217.120 176.980 222.770 ;
        RECT 177.680 218.300 178.820 222.770 ;
        RECT 179.520 218.300 180.200 222.770 ;
        RECT 177.680 217.120 180.200 218.300 ;
        RECT 175.840 215.580 180.200 217.120 ;
        RECT 174.000 214.020 180.200 215.580 ;
        RECT 164.800 212.520 180.200 214.020 ;
        RECT 163.420 209.640 180.200 212.520 ;
        RECT 180.900 209.640 182.040 222.770 ;
        RECT 163.420 207.390 182.040 209.640 ;
        RECT 154.220 205.380 182.040 207.390 ;
        RECT 182.740 205.380 183.880 222.770 ;
        RECT 154.220 204.160 183.880 205.380 ;
        RECT 147.320 194.640 183.880 204.160 ;
        RECT 0.560 139.600 183.880 194.640 ;
        RECT 184.580 216.940 185.720 222.770 ;
        RECT 186.420 216.940 187.560 222.770 ;
        RECT 184.580 216.600 187.560 216.940 ;
        RECT 188.260 216.600 189.400 222.770 ;
        RECT 184.580 213.540 189.400 216.600 ;
        RECT 190.100 213.540 191.240 222.770 ;
        RECT 184.580 211.500 191.240 213.540 ;
        RECT 191.940 211.500 193.080 222.770 ;
        RECT 184.580 208.780 193.080 211.500 ;
        RECT 193.780 212.860 194.460 222.770 ;
        RECT 195.160 212.860 196.300 222.770 ;
        RECT 193.780 208.780 196.300 212.860 ;
        RECT 184.580 206.060 196.300 208.780 ;
        RECT 197.000 206.060 198.140 222.770 ;
        RECT 198.840 206.060 199.980 222.770 ;
        RECT 184.580 203.340 199.980 206.060 ;
        RECT 200.680 203.340 201.820 222.770 ;
        RECT 184.580 199.940 201.820 203.340 ;
        RECT 202.520 211.470 203.660 222.770 ;
        RECT 204.360 216.910 205.500 222.770 ;
        RECT 206.200 216.910 207.340 222.770 ;
        RECT 204.360 211.470 207.340 216.910 ;
        RECT 202.520 208.440 207.340 211.470 ;
        RECT 208.040 215.550 208.720 222.770 ;
        RECT 209.420 216.940 210.560 222.770 ;
        RECT 211.260 216.940 212.400 222.770 ;
        RECT 209.420 215.550 212.400 216.940 ;
        RECT 208.040 211.500 212.400 215.550 ;
        RECT 213.100 211.500 214.240 222.770 ;
        RECT 208.040 208.780 214.240 211.500 ;
        RECT 214.940 213.540 216.080 222.770 ;
        RECT 216.780 213.540 217.920 222.770 ;
        RECT 214.940 208.780 217.920 213.540 ;
        RECT 208.040 208.440 217.920 208.780 ;
        RECT 202.520 203.000 217.920 208.440 ;
        RECT 218.620 203.000 219.760 222.770 ;
        RECT 202.520 202.660 219.760 203.000 ;
        RECT 220.460 219.660 221.600 222.770 ;
        RECT 222.300 219.660 223.000 222.770 ;
        RECT 220.460 202.660 223.000 219.660 ;
        RECT 202.520 199.940 223.000 202.660 ;
        RECT 184.580 139.600 223.000 199.940 ;
        RECT 0.560 50.300 223.000 139.600 ;
        RECT 0.560 47.920 78.080 50.300 ;
        RECT 0.560 39.420 76.240 47.920 ;
        RECT 0.560 29.720 70.720 39.420 ;
        RECT 0.560 20.720 51.400 29.720 ;
        RECT 0.560 17.660 9.080 20.720 ;
        RECT 0.560 11.880 1.720 17.660 ;
        RECT 1.040 0.155 1.720 11.880 ;
        RECT 2.420 14.150 9.080 17.660 ;
        RECT 2.420 12.220 7.240 14.150 ;
        RECT 2.420 6.780 5.400 12.220 ;
        RECT 2.420 0.155 3.560 6.780 ;
        RECT 4.260 0.155 5.400 6.780 ;
        RECT 6.100 0.155 7.240 12.220 ;
        RECT 7.940 0.155 9.080 14.150 ;
        RECT 9.780 17.660 51.400 20.720 ;
        RECT 9.780 15.620 14.140 17.660 ;
        RECT 9.780 4.770 12.300 15.620 ;
        RECT 9.780 0.155 10.920 4.770 ;
        RECT 11.620 0.155 12.300 4.770 ;
        RECT 13.000 0.155 14.140 15.620 ;
        RECT 14.840 11.880 37.140 17.660 ;
        RECT 14.840 9.500 32.080 11.880 ;
        RECT 14.840 7.800 26.560 9.500 ;
        RECT 14.840 6.780 19.660 7.800 ;
        RECT 14.840 0.155 15.980 6.780 ;
        RECT 16.680 1.340 19.660 6.780 ;
        RECT 16.680 0.155 17.820 1.340 ;
        RECT 18.520 0.155 19.660 1.340 ;
        RECT 20.360 7.490 26.560 7.800 ;
        RECT 20.360 6.780 24.720 7.490 ;
        RECT 20.360 0.155 21.500 6.780 ;
        RECT 22.200 6.100 24.720 6.780 ;
        RECT 22.200 0.155 23.340 6.100 ;
        RECT 24.040 0.155 24.720 6.100 ;
        RECT 25.420 0.155 26.560 7.490 ;
        RECT 27.260 6.100 32.080 9.500 ;
        RECT 27.260 5.080 30.240 6.100 ;
        RECT 27.260 0.155 28.400 5.080 ;
        RECT 29.100 0.155 30.240 5.080 ;
        RECT 30.940 0.155 32.080 6.100 ;
        RECT 32.780 9.840 37.140 11.880 ;
        RECT 32.780 0.155 33.920 9.840 ;
        RECT 34.620 6.780 37.140 9.840 ;
        RECT 34.620 0.155 35.300 6.780 ;
        RECT 36.000 0.155 37.140 6.780 ;
        RECT 37.840 17.320 51.400 17.660 ;
        RECT 37.840 9.500 42.660 17.320 ;
        RECT 37.840 0.155 38.980 9.500 ;
        RECT 39.680 6.780 42.660 9.500 ;
        RECT 39.680 0.155 40.820 6.780 ;
        RECT 41.520 0.155 42.660 6.780 ;
        RECT 43.360 14.260 51.400 17.320 ;
        RECT 43.360 9.320 46.340 14.260 ;
        RECT 43.360 0.155 44.500 9.320 ;
        RECT 45.200 0.155 46.340 9.320 ;
        RECT 47.040 1.370 51.400 14.260 ;
        RECT 47.040 0.155 47.720 1.370 ;
        RECT 48.420 0.155 49.560 1.370 ;
        RECT 50.260 0.155 51.400 1.370 ;
        RECT 52.100 21.060 70.720 29.720 ;
        RECT 52.100 15.280 55.080 21.060 ;
        RECT 52.100 0.155 53.240 15.280 ;
        RECT 53.940 0.155 55.080 15.280 ;
        RECT 55.780 15.620 70.720 21.060 ;
        RECT 55.780 14.150 69.340 15.620 ;
        RECT 55.780 0.155 56.920 14.150 ;
        RECT 57.620 11.880 69.340 14.150 ;
        RECT 57.620 6.440 67.500 11.880 ;
        RECT 57.620 4.400 63.820 6.440 ;
        RECT 57.620 3.410 61.980 4.400 ;
        RECT 57.620 0.155 58.760 3.410 ;
        RECT 59.460 1.370 61.980 3.410 ;
        RECT 59.460 0.155 60.140 1.370 ;
        RECT 60.840 0.155 61.980 1.370 ;
        RECT 62.680 0.155 63.820 4.400 ;
        RECT 64.520 0.155 65.660 6.440 ;
        RECT 66.360 0.155 67.500 6.440 ;
        RECT 68.200 0.155 69.340 11.880 ;
        RECT 70.040 0.155 70.720 15.620 ;
        RECT 71.420 20.200 76.240 39.420 ;
        RECT 71.420 0.155 72.560 20.200 ;
        RECT 73.260 12.930 76.240 20.200 ;
        RECT 73.260 0.155 74.400 12.930 ;
        RECT 75.100 0.155 76.240 12.930 ;
        RECT 76.940 0.155 78.080 47.920 ;
        RECT 78.780 44.860 223.000 50.300 ;
        RECT 78.780 37.040 90.500 44.860 ;
        RECT 78.780 7.460 83.140 37.040 ;
        RECT 78.780 0.155 79.920 7.460 ;
        RECT 80.620 6.300 83.140 7.460 ;
        RECT 80.620 0.155 81.760 6.300 ;
        RECT 82.460 0.155 83.140 6.300 ;
        RECT 83.840 14.150 90.500 37.040 ;
        RECT 83.840 6.130 88.660 14.150 ;
        RECT 83.840 0.155 84.980 6.130 ;
        RECT 85.680 5.240 88.660 6.130 ;
        RECT 85.680 0.155 86.820 5.240 ;
        RECT 87.520 0.155 88.660 5.240 ;
        RECT 89.360 0.155 90.500 14.150 ;
        RECT 91.200 26.160 223.000 44.860 ;
        RECT 91.200 25.480 199.980 26.160 ;
        RECT 91.200 19.700 132.820 25.480 ;
        RECT 91.200 17.320 102.920 19.700 ;
        RECT 91.200 8.820 101.080 17.320 ;
        RECT 91.200 6.440 94.180 8.820 ;
        RECT 91.200 0.155 92.340 6.440 ;
        RECT 93.040 0.155 94.180 6.440 ;
        RECT 94.880 4.770 101.080 8.820 ;
        RECT 94.880 0.155 95.560 4.770 ;
        RECT 96.260 4.740 99.240 4.770 ;
        RECT 96.260 0.155 97.400 4.740 ;
        RECT 98.100 0.155 99.240 4.740 ;
        RECT 99.940 0.155 101.080 4.770 ;
        RECT 101.780 0.155 102.920 17.320 ;
        RECT 103.620 18.680 132.820 19.700 ;
        RECT 103.620 17.320 111.660 18.680 ;
        RECT 103.620 14.460 109.820 17.320 ;
        RECT 103.620 0.155 104.760 14.460 ;
        RECT 105.460 7.490 109.820 14.460 ;
        RECT 105.460 1.370 107.980 7.490 ;
        RECT 105.460 0.155 106.140 1.370 ;
        RECT 106.840 0.155 107.980 1.370 ;
        RECT 108.680 0.155 109.820 7.490 ;
        RECT 110.520 0.155 111.660 17.320 ;
        RECT 112.360 16.980 132.820 18.680 ;
        RECT 112.360 11.540 130.980 16.980 ;
        RECT 112.360 6.440 118.560 11.540 ;
        RECT 112.360 3.410 115.340 6.440 ;
        RECT 112.360 0.155 113.500 3.410 ;
        RECT 114.200 0.155 115.340 3.410 ;
        RECT 116.040 3.410 118.560 6.440 ;
        RECT 116.040 0.155 117.180 3.410 ;
        RECT 117.880 0.155 118.560 3.410 ;
        RECT 119.260 7.490 130.980 11.540 ;
        RECT 119.260 4.770 129.140 7.490 ;
        RECT 119.260 3.040 124.080 4.770 ;
        RECT 119.260 0.155 120.400 3.040 ;
        RECT 121.100 2.700 124.080 3.040 ;
        RECT 121.100 0.155 122.240 2.700 ;
        RECT 122.940 0.155 124.080 2.700 ;
        RECT 124.780 4.060 129.140 4.770 ;
        RECT 124.780 0.155 125.920 4.060 ;
        RECT 126.620 2.360 129.140 4.060 ;
        RECT 126.620 0.155 127.760 2.360 ;
        RECT 128.460 0.155 129.140 2.360 ;
        RECT 129.840 0.155 130.980 7.490 ;
        RECT 131.680 0.155 132.820 16.980 ;
        RECT 133.520 23.100 199.980 25.480 ;
        RECT 133.520 20.720 196.760 23.100 ;
        RECT 133.520 19.700 194.920 20.720 ;
        RECT 133.520 18.340 141.560 19.700 ;
        RECT 133.520 17.320 136.500 18.340 ;
        RECT 133.520 0.155 134.660 17.320 ;
        RECT 135.360 0.155 136.500 17.320 ;
        RECT 137.200 16.980 141.560 18.340 ;
        RECT 137.200 1.680 140.180 16.980 ;
        RECT 137.200 0.155 138.340 1.680 ;
        RECT 139.040 0.155 140.180 1.680 ;
        RECT 140.880 0.155 141.560 16.980 ;
        RECT 142.260 16.980 194.920 19.700 ;
        RECT 142.260 16.800 180.660 16.980 ;
        RECT 142.260 14.600 168.240 16.800 ;
        RECT 142.260 12.220 155.820 14.600 ;
        RECT 142.260 11.540 150.760 12.220 ;
        RECT 142.260 8.820 147.080 11.540 ;
        RECT 142.260 8.640 145.240 8.820 ;
        RECT 142.260 0.155 143.400 8.640 ;
        RECT 144.100 0.155 145.240 8.640 ;
        RECT 145.940 0.155 147.080 8.820 ;
        RECT 147.780 1.370 150.760 11.540 ;
        RECT 147.780 0.155 148.920 1.370 ;
        RECT 149.620 0.155 150.760 1.370 ;
        RECT 151.460 8.820 155.820 12.220 ;
        RECT 151.460 6.100 153.980 8.820 ;
        RECT 151.460 0.155 152.600 6.100 ;
        RECT 153.300 0.155 153.980 6.100 ;
        RECT 154.680 0.155 155.820 8.820 ;
        RECT 156.520 10.680 168.240 14.600 ;
        RECT 156.520 10.000 164.560 10.680 ;
        RECT 156.520 8.640 163.180 10.000 ;
        RECT 156.520 1.370 161.340 8.640 ;
        RECT 156.520 0.155 157.660 1.370 ;
        RECT 158.360 1.200 161.340 1.370 ;
        RECT 158.360 0.155 159.500 1.200 ;
        RECT 160.200 0.155 161.340 1.200 ;
        RECT 162.040 0.155 163.180 8.640 ;
        RECT 163.880 0.155 164.560 10.000 ;
        RECT 165.260 7.490 168.240 10.680 ;
        RECT 165.260 0.155 166.400 7.490 ;
        RECT 167.100 0.155 168.240 7.490 ;
        RECT 168.940 14.080 180.660 16.800 ;
        RECT 168.940 1.200 171.920 14.080 ;
        RECT 168.940 0.155 170.080 1.200 ;
        RECT 170.780 0.155 171.920 1.200 ;
        RECT 172.620 13.240 180.660 14.080 ;
        RECT 172.620 12.900 178.820 13.240 ;
        RECT 172.620 0.155 173.760 12.900 ;
        RECT 174.460 7.490 178.820 12.900 ;
        RECT 174.460 3.410 176.980 7.490 ;
        RECT 174.460 0.155 175.600 3.410 ;
        RECT 176.300 0.155 176.980 3.410 ;
        RECT 177.680 0.155 178.820 7.490 ;
        RECT 179.520 0.155 180.660 13.240 ;
        RECT 181.360 15.280 194.920 16.980 ;
        RECT 181.360 12.220 191.240 15.280 ;
        RECT 181.360 10.680 189.400 12.220 ;
        RECT 181.360 7.490 184.340 10.680 ;
        RECT 181.360 0.155 182.500 7.490 ;
        RECT 183.200 0.155 184.340 7.490 ;
        RECT 185.040 7.280 189.400 10.680 ;
        RECT 185.040 0.155 186.180 7.280 ;
        RECT 186.880 6.780 189.400 7.280 ;
        RECT 186.880 0.155 188.020 6.780 ;
        RECT 188.720 0.155 189.400 6.780 ;
        RECT 190.100 0.155 191.240 12.220 ;
        RECT 191.940 6.130 194.920 15.280 ;
        RECT 191.940 0.155 193.080 6.130 ;
        RECT 193.780 0.155 194.920 6.130 ;
        RECT 195.620 0.155 196.760 20.720 ;
        RECT 197.460 9.500 199.980 23.100 ;
        RECT 197.460 0.155 198.600 9.500 ;
        RECT 199.300 0.155 199.980 9.500 ;
        RECT 200.680 23.100 223.000 26.160 ;
        RECT 200.680 17.320 216.080 23.100 ;
        RECT 200.680 14.260 209.180 17.320 ;
        RECT 200.680 0.155 201.820 14.260 ;
        RECT 202.520 14.150 209.180 14.260 ;
        RECT 202.520 0.155 203.660 14.150 ;
        RECT 204.360 12.220 209.180 14.150 ;
        RECT 204.360 0.155 205.500 12.220 ;
        RECT 206.200 9.840 209.180 12.220 ;
        RECT 206.200 0.155 207.340 9.840 ;
        RECT 208.040 0.155 209.180 9.840 ;
        RECT 209.880 15.280 216.080 17.320 ;
        RECT 209.880 0.155 211.020 15.280 ;
        RECT 211.720 8.850 216.080 15.280 ;
        RECT 211.720 0.155 212.400 8.850 ;
        RECT 213.100 6.440 216.080 8.850 ;
        RECT 213.100 0.155 214.240 6.440 ;
        RECT 214.940 0.155 216.080 6.440 ;
        RECT 216.780 16.980 223.000 23.100 ;
        RECT 216.780 0.155 217.920 16.980 ;
        RECT 218.620 6.780 223.000 16.980 ;
        RECT 218.620 4.060 221.600 6.780 ;
        RECT 218.620 0.155 219.760 4.060 ;
        RECT 220.460 0.155 221.600 4.060 ;
        RECT 222.300 0.155 223.000 6.780 ;
      LAYER met3 ;
        RECT 20.730 221.470 202.830 222.185 ;
        RECT 1.445 220.530 222.115 221.470 ;
        RECT 20.730 219.430 206.050 220.530 ;
        RECT 1.445 219.170 222.115 219.430 ;
        RECT 19.810 218.070 209.270 219.170 ;
        RECT 1.445 217.130 222.115 218.070 ;
        RECT 15.210 216.030 205.590 217.130 ;
        RECT 1.445 215.770 222.115 216.030 ;
        RECT 19.350 214.670 208.810 215.770 ;
        RECT 1.445 213.730 222.115 214.670 ;
        RECT 16.590 212.630 210.190 213.730 ;
        RECT 1.445 212.370 222.115 212.630 ;
        RECT 19.350 211.270 213.410 212.370 ;
        RECT 1.445 210.330 222.115 211.270 ;
        RECT 7.390 209.230 213.870 210.330 ;
        RECT 1.445 208.290 222.115 209.230 ;
        RECT 19.350 207.190 210.190 208.290 ;
        RECT 1.445 206.930 222.115 207.190 ;
        RECT 6.930 205.830 213.410 206.930 ;
        RECT 1.445 204.890 222.115 205.830 ;
        RECT 16.590 203.790 208.810 204.890 ;
        RECT 1.445 203.530 222.115 203.790 ;
        RECT 7.850 202.430 214.330 203.530 ;
        RECT 1.445 201.490 222.115 202.430 ;
        RECT 19.350 200.390 213.870 201.490 ;
        RECT 1.445 200.130 222.115 200.390 ;
        RECT 8.310 199.030 209.270 200.130 ;
        RECT 1.445 198.090 222.115 199.030 ;
        RECT 6.930 196.990 213.410 198.090 ;
        RECT 1.445 196.730 222.115 196.990 ;
        RECT 7.390 195.630 213.870 196.730 ;
        RECT 1.445 194.690 222.115 195.630 ;
        RECT 7.850 193.590 209.270 194.690 ;
        RECT 1.445 192.650 222.115 193.590 ;
        RECT 6.930 191.550 214.330 192.650 ;
        RECT 1.445 191.290 222.115 191.550 ;
        RECT 7.390 190.190 213.410 191.290 ;
        RECT 1.445 189.250 222.115 190.190 ;
        RECT 6.930 188.150 221.230 189.250 ;
        RECT 1.445 187.890 222.115 188.150 ;
        RECT 7.390 186.790 213.870 187.890 ;
        RECT 1.445 185.850 222.115 186.790 ;
        RECT 7.390 184.750 213.410 185.850 ;
        RECT 1.445 184.490 222.115 184.750 ;
        RECT 20.270 183.390 210.190 184.490 ;
        RECT 1.445 182.450 222.115 183.390 ;
        RECT 20.270 181.350 209.270 182.450 ;
        RECT 1.445 180.410 222.115 181.350 ;
        RECT 20.730 179.310 211.110 180.410 ;
        RECT 1.445 179.050 222.115 179.310 ;
        RECT 16.590 177.950 206.510 179.050 ;
        RECT 1.445 177.010 222.115 177.950 ;
        RECT 13.370 175.910 210.190 177.010 ;
        RECT 1.445 175.650 222.115 175.910 ;
        RECT 6.930 174.550 219.850 175.650 ;
        RECT 1.445 173.610 222.115 174.550 ;
        RECT 7.850 172.510 221.230 173.610 ;
        RECT 1.445 172.250 222.115 172.510 ;
        RECT 7.390 171.150 213.410 172.250 ;
        RECT 1.445 170.210 222.115 171.150 ;
        RECT 6.930 169.110 209.270 170.210 ;
        RECT 1.445 168.850 222.115 169.110 ;
        RECT 7.390 167.750 213.870 168.850 ;
        RECT 1.445 166.810 222.115 167.750 ;
        RECT 19.810 165.710 213.870 166.810 ;
        RECT 1.445 164.770 222.115 165.710 ;
        RECT 10.150 163.670 213.870 164.770 ;
        RECT 1.445 163.410 222.115 163.670 ;
        RECT 13.830 162.310 210.190 163.410 ;
        RECT 1.445 161.370 222.115 162.310 ;
        RECT 19.810 160.270 218.010 161.370 ;
        RECT 1.445 160.010 222.115 160.270 ;
        RECT 20.730 158.910 209.270 160.010 ;
        RECT 1.445 157.970 222.115 158.910 ;
        RECT 19.180 156.870 218.010 157.970 ;
        RECT 1.445 156.610 222.115 156.870 ;
        RECT 18.430 155.510 218.010 156.610 ;
        RECT 1.445 154.570 222.115 155.510 ;
        RECT 14.750 153.470 213.410 154.570 ;
        RECT 1.445 152.530 222.115 153.470 ;
        RECT 17.340 151.430 213.870 152.530 ;
        RECT 1.445 151.170 222.115 151.430 ;
        RECT 21.190 150.070 213.410 151.170 ;
        RECT 1.445 149.130 222.115 150.070 ;
        RECT 7.850 148.030 213.870 149.130 ;
        RECT 1.445 147.770 222.115 148.030 ;
        RECT 7.850 146.670 213.870 147.770 ;
        RECT 1.445 145.730 222.115 146.670 ;
        RECT 22.110 144.630 201.450 145.730 ;
        RECT 1.445 144.370 222.115 144.630 ;
        RECT 20.730 143.270 200.070 144.370 ;
        RECT 1.445 142.330 222.115 143.270 ;
        RECT 7.450 141.230 200.070 142.330 ;
        RECT 1.445 140.970 222.115 141.230 ;
        RECT 8.770 139.870 200.530 140.970 ;
        RECT 1.445 138.930 222.115 139.870 ;
        RECT 19.100 137.830 210.190 138.930 ;
        RECT 1.445 136.890 222.115 137.830 ;
        RECT 35.910 135.790 200.530 136.890 ;
        RECT 1.445 135.530 222.115 135.790 ;
        RECT 15.210 134.430 202.370 135.530 ;
        RECT 1.445 133.490 222.115 134.430 ;
        RECT 19.100 132.390 201.910 133.490 ;
        RECT 1.445 132.130 222.115 132.390 ;
        RECT 21.190 131.030 200.070 132.130 ;
        RECT 1.445 130.090 222.115 131.030 ;
        RECT 13.830 128.990 213.350 130.090 ;
        RECT 1.445 128.730 222.115 128.990 ;
        RECT 20.270 127.630 200.990 128.730 ;
        RECT 1.445 126.690 222.115 127.630 ;
        RECT 34.530 125.590 198.690 126.690 ;
        RECT 1.445 124.650 222.115 125.590 ;
        RECT 9.690 123.550 206.450 124.650 ;
        RECT 1.445 123.290 222.115 123.550 ;
        RECT 17.050 122.190 192.710 123.290 ;
        RECT 1.445 121.250 222.115 122.190 ;
        RECT 14.290 120.150 201.450 121.250 ;
        RECT 1.445 119.890 222.115 120.150 ;
        RECT 7.850 118.790 207.890 119.890 ;
        RECT 1.445 117.850 222.115 118.790 ;
        RECT 7.390 116.750 202.830 117.850 ;
        RECT 1.445 116.490 222.115 116.750 ;
        RECT 17.970 115.390 219.390 116.490 ;
        RECT 1.445 114.450 222.115 115.390 ;
        RECT 28.090 113.350 205.130 114.450 ;
        RECT 1.445 113.090 222.115 113.350 ;
        RECT 19.350 111.990 204.210 113.090 ;
        RECT 1.445 111.050 222.115 111.990 ;
        RECT 6.010 109.950 219.390 111.050 ;
        RECT 1.445 109.010 222.115 109.950 ;
        RECT 9.690 107.910 200.990 109.010 ;
        RECT 1.445 107.650 222.115 107.910 ;
        RECT 20.270 106.550 219.390 107.650 ;
        RECT 1.445 105.610 222.115 106.550 ;
        RECT 20.730 104.510 219.390 105.610 ;
        RECT 1.445 104.250 222.115 104.510 ;
        RECT 18.430 103.150 219.390 104.250 ;
        RECT 1.445 102.210 222.115 103.150 ;
        RECT 15.670 101.110 209.270 102.210 ;
        RECT 1.445 100.850 222.115 101.110 ;
        RECT 6.930 99.750 213.410 100.850 ;
        RECT 1.445 98.810 222.115 99.750 ;
        RECT 20.730 97.710 200.530 98.810 ;
        RECT 1.445 96.770 222.115 97.710 ;
        RECT 17.050 95.670 200.070 96.770 ;
        RECT 1.445 95.410 222.115 95.670 ;
        RECT 18.260 94.310 219.390 95.410 ;
        RECT 1.445 93.370 222.115 94.310 ;
        RECT 11.990 92.270 201.450 93.370 ;
        RECT 1.445 92.010 222.115 92.270 ;
        RECT 21.190 90.910 219.390 92.010 ;
        RECT 1.445 89.970 222.115 90.910 ;
        RECT 20.730 88.870 219.390 89.970 ;
        RECT 1.445 88.610 222.115 88.870 ;
        RECT 6.930 87.510 206.220 88.610 ;
        RECT 1.445 86.570 222.115 87.510 ;
        RECT 7.850 85.470 219.390 86.570 ;
        RECT 1.445 85.210 222.115 85.470 ;
        RECT 7.390 84.110 204.210 85.210 ;
        RECT 1.445 83.170 222.115 84.110 ;
        RECT 14.750 82.070 200.530 83.170 ;
        RECT 1.445 81.130 222.115 82.070 ;
        RECT 10.150 80.030 196.850 81.130 ;
        RECT 1.445 79.770 222.115 80.030 ;
        RECT 20.730 78.670 203.290 79.770 ;
        RECT 1.445 77.730 222.115 78.670 ;
        RECT 7.450 76.630 200.990 77.730 ;
        RECT 1.445 76.370 222.115 76.630 ;
        RECT 18.890 75.270 200.070 76.370 ;
        RECT 1.445 74.330 222.115 75.270 ;
        RECT 17.510 73.230 214.270 74.330 ;
        RECT 1.445 72.970 222.115 73.230 ;
        RECT 25.790 71.870 214.270 72.970 ;
        RECT 1.445 70.930 222.115 71.870 ;
        RECT 19.350 69.830 167.870 70.930 ;
        RECT 1.445 68.890 222.115 69.830 ;
        RECT 17.050 67.790 200.070 68.890 ;
        RECT 1.445 67.530 222.115 67.790 ;
        RECT 14.290 66.430 206.450 67.530 ;
        RECT 1.445 65.490 222.115 66.430 ;
        RECT 10.150 64.390 202.370 65.490 ;
        RECT 1.445 64.130 222.115 64.390 ;
        RECT 10.610 63.030 211.570 64.130 ;
        RECT 1.445 62.090 222.115 63.030 ;
        RECT 23.490 60.990 193.630 62.090 ;
        RECT 1.445 60.730 222.115 60.990 ;
        RECT 23.490 59.630 219.390 60.730 ;
        RECT 1.445 58.690 222.115 59.630 ;
        RECT 20.730 57.590 213.350 58.690 ;
        RECT 1.445 57.330 222.115 57.590 ;
        RECT 14.290 56.230 201.910 57.330 ;
        RECT 1.445 55.290 222.115 56.230 ;
        RECT 20.270 54.190 200.070 55.290 ;
        RECT 1.445 53.250 222.115 54.190 ;
        RECT 7.390 52.150 200.070 53.250 ;
        RECT 1.445 51.890 222.115 52.150 ;
        RECT 20.730 50.790 200.070 51.890 ;
        RECT 1.445 49.850 222.115 50.790 ;
        RECT 19.350 48.750 210.190 49.850 ;
        RECT 1.445 48.490 222.115 48.750 ;
        RECT 20.730 47.390 199.550 48.490 ;
        RECT 1.445 46.450 222.115 47.390 ;
        RECT 20.730 45.350 200.070 46.450 ;
        RECT 1.445 45.090 222.115 45.350 ;
        RECT 18.890 43.990 203.290 45.090 ;
        RECT 1.445 43.050 222.115 43.990 ;
        RECT 20.730 41.950 189.740 43.050 ;
        RECT 1.445 41.010 222.115 41.950 ;
        RECT 20.730 39.910 201.450 41.010 ;
        RECT 1.445 39.650 222.115 39.910 ;
        RECT 17.510 38.550 200.990 39.650 ;
        RECT 1.445 37.610 222.115 38.550 ;
        RECT 24.410 36.510 209.670 37.610 ;
        RECT 1.445 36.250 222.115 36.510 ;
        RECT 17.050 35.150 211.110 36.250 ;
        RECT 1.445 34.210 222.115 35.150 ;
        RECT 10.150 33.110 205.590 34.210 ;
        RECT 1.445 32.850 222.115 33.110 ;
        RECT 20.730 31.750 212.490 32.850 ;
        RECT 1.445 30.810 222.115 31.750 ;
        RECT 1.870 29.710 206.510 30.810 ;
        RECT 1.445 29.450 222.115 29.710 ;
        RECT 14.750 28.350 206.050 29.450 ;
        RECT 1.445 27.410 222.115 28.350 ;
        RECT 20.100 26.310 201.450 27.410 ;
        RECT 1.445 25.370 222.115 26.310 ;
        RECT 7.850 24.270 200.530 25.370 ;
        RECT 1.445 24.010 222.115 24.270 ;
        RECT 19.810 22.910 212.030 24.010 ;
        RECT 1.445 21.970 222.115 22.910 ;
        RECT 7.390 20.870 212.490 21.970 ;
        RECT 1.445 20.610 222.115 20.870 ;
        RECT 19.350 19.510 201.450 20.610 ;
        RECT 1.445 18.570 222.115 19.510 ;
        RECT 10.610 17.470 199.610 18.570 ;
        RECT 1.445 17.210 222.115 17.470 ;
        RECT 15.210 16.110 200.530 17.210 ;
        RECT 1.445 15.170 222.115 16.110 ;
        RECT 20.730 14.070 200.990 15.170 ;
        RECT 1.445 13.130 222.115 14.070 ;
        RECT 19.810 12.030 205.130 13.130 ;
        RECT 1.445 11.770 222.115 12.030 ;
        RECT 18.890 10.670 204.670 11.770 ;
        RECT 1.445 9.730 222.115 10.670 ;
        RECT 16.590 8.630 212.490 9.730 ;
        RECT 1.445 8.370 222.115 8.630 ;
        RECT 16.130 7.270 200.530 8.370 ;
        RECT 1.445 6.330 222.115 7.270 ;
        RECT 14.290 5.230 200.530 6.330 ;
        RECT 1.445 4.970 222.115 5.230 ;
        RECT 19.350 3.870 199.610 4.970 ;
        RECT 1.445 2.930 222.115 3.870 ;
        RECT 10.150 1.830 200.530 2.930 ;
        RECT 1.445 1.570 222.115 1.830 ;
        RECT 15.670 0.470 202.370 1.570 ;
        RECT 1.445 0.175 222.115 0.470 ;
      LAYER met4 ;
        RECT 13.175 4.800 20.640 217.425 ;
        RECT 23.040 4.800 97.440 217.425 ;
        RECT 99.840 4.800 174.240 217.425 ;
        RECT 176.640 4.800 208.545 217.425 ;
        RECT 13.175 1.535 208.545 4.800 ;
  END
END LUT4AB
END LIBRARY