module counter (out);
   output out;
   DFFPOSX1 \x0/d0 (.Q(out));
endmodule

