# macro with bus bit (intentionally reverse order of liberty)

VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MACRO bus4
 SIZE 50 BY 20 ;
 PIN in[0] DIRECTION INPUT ; END in[0]
 PIN in[1] DIRECTION INPUT ; END in[1]
 PIN in[2] DIRECTION INPUT ; END in[2]
 PIN in[3] DIRECTION INPUT ; END in[3]
 PIN out[0] DIRECTION OUTPUT ; END out[0]
 PIN out[1] DIRECTION OUTPUT ; END out[1]
 PIN out[2] DIRECTION OUTPUT ; END out[2]
 PIN out[3] DIRECTION OUTPUT ; END out[3]
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END bus4

END LIBRARY

