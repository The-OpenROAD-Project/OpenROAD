sky130_fd_sc_hs_merged.lef