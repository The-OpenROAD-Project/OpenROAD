# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_io__overlay_gpiov2
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 80 BY 200 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 1.270000 56.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 53.125000 80.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 1.270000 51.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 48.365000 80.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN PAD
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 31.870000 127.605000 53.410000 149.150000 ;
    END
  END PAD
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT  0.000000  8.885000  1.270000  9.105000 ;
        RECT  0.000000  9.105000 80.000000 13.315000 ;
        RECT  0.000000 13.315000  1.270000 13.535000 ;
        RECT 78.730000  8.885000 80.000000  9.105000 ;
        RECT 78.730000 13.315000 80.000000 13.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 8.985000 80.000000 13.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT  0.000000 2.035000  1.270000 2.255000 ;
        RECT  0.000000 2.255000 80.000000 7.265000 ;
        RECT  0.000000 7.265000  1.270000 7.485000 ;
        RECT 78.730000 2.035000 80.000000 2.255000 ;
        RECT 78.730000 7.265000 80.000000 7.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 2.135000 80.000000 7.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 14.935000  0.965000 15.155000 ;
        RECT 0.000000 15.155000 78.970000 18.165000 ;
        RECT 0.000000 18.165000  0.965000 18.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 79.035000 14.935000 80.000000 18.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 15.035000 80.000000 18.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT  0.000000 19.785000  1.270000 20.005000 ;
        RECT  0.000000 20.005000 80.000000 24.215000 ;
        RECT  0.000000 24.215000  1.270000 24.435000 ;
        RECT 78.730000 19.785000 80.000000 20.005000 ;
        RECT 78.730000 24.215000 80.000000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT  0.000000 70.035000  1.270000 70.155000 ;
        RECT  0.000000 70.155000 80.000000 94.865000 ;
        RECT  0.000000 94.865000  1.270000 95.000000 ;
        RECT 78.730000 70.035000 80.000000 70.155000 ;
        RECT 78.730000 94.865000 80.000000 95.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 19.885000 80.000000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 70.035000 80.000000 94.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT  0.000000 64.085000  1.270000 64.305000 ;
        RECT  0.000000 64.305000 80.000000 68.315000 ;
        RECT  0.000000 68.315000  1.270000 68.535000 ;
        RECT 78.730000 64.085000 80.000000 64.305000 ;
        RECT 78.730000 68.315000 80.000000 68.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 64.185000 80.000000 68.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT  0.000000 36.735000  1.270000 36.955000 ;
        RECT  0.000000 36.955000 80.000000 39.965000 ;
        RECT  0.000000 39.965000  1.270000 40.185000 ;
        RECT 78.730000 36.735000 80.000000 36.955000 ;
        RECT 78.730000 39.965000 80.000000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 47.735000 1.270000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 51.645000 80.000000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 56.405000 1.270000 56.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 47.735000 80.000000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 56.405000 80.000000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 36.835000 80.000000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 47.735000 80.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT  0.000000 41.585000  1.270000 41.805000 ;
        RECT  0.000000 41.805000 80.000000 46.015000 ;
        RECT  0.000000 46.015000  1.270000 46.235000 ;
        RECT 78.730000 41.585000 80.000000 41.805000 ;
        RECT 78.730000 46.015000 80.000000 46.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 41.685000 80.000000 46.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT  0.000000 175.785000  1.270000 175.910000 ;
        RECT  0.000000 175.910000 80.000000 199.880000 ;
        RECT  0.000000 199.880000  1.270000 200.000000 ;
        RECT 78.730000 175.785000 80.000000 175.910000 ;
        RECT 78.730000 199.880000 80.000000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT  0.000000 25.835000  1.270000 26.055000 ;
        RECT  0.000000 26.055000 80.000000 30.265000 ;
        RECT  0.000000 30.265000  1.270000 30.485000 ;
        RECT 78.730000 25.835000 80.000000 26.055000 ;
        RECT 78.730000 30.265000 80.000000 30.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 175.785000 80.000000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 25.935000 80.000000 30.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT  0.000000 58.235000  1.270000 58.455000 ;
        RECT  0.000000 58.455000 80.000000 62.465000 ;
        RECT  0.000000 62.465000  1.270000 62.685000 ;
        RECT 78.730000 58.235000 80.000000 58.455000 ;
        RECT 78.730000 62.465000 80.000000 62.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 58.335000 80.000000 62.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT  0.000000 31.885000  1.270000 32.105000 ;
        RECT  0.000000 32.105000 80.000000 35.115000 ;
        RECT  0.000000 35.115000  1.270000 35.335000 ;
        RECT 78.730000 31.885000 80.000000 32.105000 ;
        RECT 78.730000 35.115000 80.000000 35.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 31.985000 80.000000 35.235000 ;
    END
  END VSWITCH
  OBS
    LAYER via4 ;
      RECT  0.995000  20.195000  1.795000  20.995000 ;
      RECT  0.995000  23.225000  1.795000  24.025000 ;
      RECT  0.995000  26.245000  1.795000  27.045000 ;
      RECT  0.995000  29.275000  1.795000  30.075000 ;
      RECT  1.000000   2.450000  1.800000   3.250000 ;
      RECT  1.000000   4.360000  1.800000   5.160000 ;
      RECT  1.000000   6.270000  1.800000   7.070000 ;
      RECT  1.000000  15.345000  1.800000  16.145000 ;
      RECT  1.000000  17.175000  1.800000  17.975000 ;
      RECT  1.000000  32.295000  1.800000  33.095000 ;
      RECT  1.000000  34.125000  1.800000  34.925000 ;
      RECT  1.000000  37.145000  1.800000  37.945000 ;
      RECT  1.000000  38.975000  1.800000  39.775000 ;
      RECT  1.000000  41.995000  1.800000  42.795000 ;
      RECT  1.000000  45.025000  1.800000  45.825000 ;
      RECT  1.000000  51.835000  1.800000  52.635000 ;
      RECT  1.000000  58.645000  1.800000  59.445000 ;
      RECT  1.000000  61.475000  1.800000  62.275000 ;
      RECT  1.000000  64.495000  1.800000  65.295000 ;
      RECT  1.000000  67.325000  1.800000  68.125000 ;
      RECT  1.000000  70.350000  1.800000  71.150000 ;
      RECT  1.000000  72.030000  1.800000  72.830000 ;
      RECT  1.000000  73.710000  1.800000  74.510000 ;
      RECT  1.000000  75.390000  1.800000  76.190000 ;
      RECT  1.000000  77.070000  1.800000  77.870000 ;
      RECT  1.000000  78.750000  1.800000  79.550000 ;
      RECT  1.000000  80.430000  1.800000  81.230000 ;
      RECT  1.000000  82.110000  1.800000  82.910000 ;
      RECT  1.000000  83.790000  1.800000  84.590000 ;
      RECT  1.000000  85.470000  1.800000  86.270000 ;
      RECT  1.000000  87.150000  1.800000  87.950000 ;
      RECT  1.000000  88.830000  1.800000  89.630000 ;
      RECT  1.000000  90.510000  1.800000  91.310000 ;
      RECT  1.000000  92.190000  1.800000  92.990000 ;
      RECT  1.000000  93.870000  1.800000  94.670000 ;
      RECT  1.000000 176.155000  1.800000 176.955000 ;
      RECT  1.000000 177.775000  1.800000 178.575000 ;
      RECT  1.000000 179.395000  1.800000 180.195000 ;
      RECT  1.000000 181.015000  1.800000 181.815000 ;
      RECT  1.000000 182.635000  1.800000 183.435000 ;
      RECT  1.000000 184.255000  1.800000 185.055000 ;
      RECT  1.000000 185.875000  1.800000 186.675000 ;
      RECT  1.000000 187.495000  1.800000 188.295000 ;
      RECT  1.000000 189.115000  1.800000 189.915000 ;
      RECT  1.000000 190.735000  1.800000 191.535000 ;
      RECT  1.000000 192.355000  1.800000 193.155000 ;
      RECT  1.000000 193.975000  1.800000 194.775000 ;
      RECT  1.000000 195.595000  1.800000 196.395000 ;
      RECT  1.000000 197.215000  1.800000 198.015000 ;
      RECT  1.000000 198.835000  1.800000 199.635000 ;
      RECT  1.005000   9.295000  1.805000  10.095000 ;
      RECT  1.005000  12.325000  1.805000  13.125000 ;
      RECT  2.600000  20.195000  3.400000  20.995000 ;
      RECT  2.600000  23.225000  3.400000  24.025000 ;
      RECT  2.600000  26.245000  3.400000  27.045000 ;
      RECT  2.600000  29.275000  3.400000  30.075000 ;
      RECT  2.605000   2.450000  3.405000   3.250000 ;
      RECT  2.605000   4.360000  3.405000   5.160000 ;
      RECT  2.605000   6.270000  3.405000   7.070000 ;
      RECT  2.605000  15.345000  3.405000  16.145000 ;
      RECT  2.605000  17.175000  3.405000  17.975000 ;
      RECT  2.605000  32.295000  3.405000  33.095000 ;
      RECT  2.605000  34.125000  3.405000  34.925000 ;
      RECT  2.605000  37.145000  3.405000  37.945000 ;
      RECT  2.605000  38.975000  3.405000  39.775000 ;
      RECT  2.605000  41.995000  3.405000  42.795000 ;
      RECT  2.605000  45.025000  3.405000  45.825000 ;
      RECT  2.605000  51.835000  3.405000  52.635000 ;
      RECT  2.605000  58.645000  3.405000  59.445000 ;
      RECT  2.605000  61.475000  3.405000  62.275000 ;
      RECT  2.605000  64.495000  3.405000  65.295000 ;
      RECT  2.605000  67.325000  3.405000  68.125000 ;
      RECT  2.605000  70.350000  3.405000  71.150000 ;
      RECT  2.605000  72.030000  3.405000  72.830000 ;
      RECT  2.605000  73.710000  3.405000  74.510000 ;
      RECT  2.605000  75.390000  3.405000  76.190000 ;
      RECT  2.605000  77.070000  3.405000  77.870000 ;
      RECT  2.605000  78.750000  3.405000  79.550000 ;
      RECT  2.605000  80.430000  3.405000  81.230000 ;
      RECT  2.605000  82.110000  3.405000  82.910000 ;
      RECT  2.605000  83.790000  3.405000  84.590000 ;
      RECT  2.605000  85.470000  3.405000  86.270000 ;
      RECT  2.605000  87.150000  3.405000  87.950000 ;
      RECT  2.605000  88.830000  3.405000  89.630000 ;
      RECT  2.605000  90.510000  3.405000  91.310000 ;
      RECT  2.605000  92.190000  3.405000  92.990000 ;
      RECT  2.605000  93.870000  3.405000  94.670000 ;
      RECT  2.605000 176.155000  3.405000 176.955000 ;
      RECT  2.605000 177.775000  3.405000 178.575000 ;
      RECT  2.605000 179.395000  3.405000 180.195000 ;
      RECT  2.605000 181.015000  3.405000 181.815000 ;
      RECT  2.605000 182.635000  3.405000 183.435000 ;
      RECT  2.605000 184.255000  3.405000 185.055000 ;
      RECT  2.605000 185.875000  3.405000 186.675000 ;
      RECT  2.605000 187.495000  3.405000 188.295000 ;
      RECT  2.605000 189.115000  3.405000 189.915000 ;
      RECT  2.605000 190.735000  3.405000 191.535000 ;
      RECT  2.605000 192.355000  3.405000 193.155000 ;
      RECT  2.605000 193.975000  3.405000 194.775000 ;
      RECT  2.605000 195.595000  3.405000 196.395000 ;
      RECT  2.605000 197.215000  3.405000 198.015000 ;
      RECT  2.605000 198.835000  3.405000 199.635000 ;
      RECT  2.610000   9.295000  3.410000  10.095000 ;
      RECT  2.610000  12.325000  3.410000  13.125000 ;
      RECT  4.205000  20.195000  5.005000  20.995000 ;
      RECT  4.205000  23.225000  5.005000  24.025000 ;
      RECT  4.205000  26.245000  5.005000  27.045000 ;
      RECT  4.205000  29.275000  5.005000  30.075000 ;
      RECT  4.210000   2.450000  5.010000   3.250000 ;
      RECT  4.210000   4.360000  5.010000   5.160000 ;
      RECT  4.210000   6.270000  5.010000   7.070000 ;
      RECT  4.210000  15.345000  5.010000  16.145000 ;
      RECT  4.210000  17.175000  5.010000  17.975000 ;
      RECT  4.210000  32.295000  5.010000  33.095000 ;
      RECT  4.210000  34.125000  5.010000  34.925000 ;
      RECT  4.210000  37.145000  5.010000  37.945000 ;
      RECT  4.210000  38.975000  5.010000  39.775000 ;
      RECT  4.210000  41.995000  5.010000  42.795000 ;
      RECT  4.210000  45.025000  5.010000  45.825000 ;
      RECT  4.210000  51.835000  5.010000  52.635000 ;
      RECT  4.210000  58.645000  5.010000  59.445000 ;
      RECT  4.210000  61.475000  5.010000  62.275000 ;
      RECT  4.210000  64.495000  5.010000  65.295000 ;
      RECT  4.210000  67.325000  5.010000  68.125000 ;
      RECT  4.210000  70.350000  5.010000  71.150000 ;
      RECT  4.210000  72.030000  5.010000  72.830000 ;
      RECT  4.210000  73.710000  5.010000  74.510000 ;
      RECT  4.210000  75.390000  5.010000  76.190000 ;
      RECT  4.210000  77.070000  5.010000  77.870000 ;
      RECT  4.210000  78.750000  5.010000  79.550000 ;
      RECT  4.210000  80.430000  5.010000  81.230000 ;
      RECT  4.210000  82.110000  5.010000  82.910000 ;
      RECT  4.210000  83.790000  5.010000  84.590000 ;
      RECT  4.210000  85.470000  5.010000  86.270000 ;
      RECT  4.210000  87.150000  5.010000  87.950000 ;
      RECT  4.210000  88.830000  5.010000  89.630000 ;
      RECT  4.210000  90.510000  5.010000  91.310000 ;
      RECT  4.210000  92.190000  5.010000  92.990000 ;
      RECT  4.210000  93.870000  5.010000  94.670000 ;
      RECT  4.210000 176.155000  5.010000 176.955000 ;
      RECT  4.210000 177.775000  5.010000 178.575000 ;
      RECT  4.210000 179.395000  5.010000 180.195000 ;
      RECT  4.210000 181.015000  5.010000 181.815000 ;
      RECT  4.210000 182.635000  5.010000 183.435000 ;
      RECT  4.210000 184.255000  5.010000 185.055000 ;
      RECT  4.210000 185.875000  5.010000 186.675000 ;
      RECT  4.210000 187.495000  5.010000 188.295000 ;
      RECT  4.210000 189.115000  5.010000 189.915000 ;
      RECT  4.210000 190.735000  5.010000 191.535000 ;
      RECT  4.210000 192.355000  5.010000 193.155000 ;
      RECT  4.210000 193.975000  5.010000 194.775000 ;
      RECT  4.210000 195.595000  5.010000 196.395000 ;
      RECT  4.210000 197.215000  5.010000 198.015000 ;
      RECT  4.210000 198.835000  5.010000 199.635000 ;
      RECT  4.215000   9.295000  5.015000  10.095000 ;
      RECT  4.215000  12.325000  5.015000  13.125000 ;
      RECT  5.810000  20.195000  6.610000  20.995000 ;
      RECT  5.810000  23.225000  6.610000  24.025000 ;
      RECT  5.810000  26.245000  6.610000  27.045000 ;
      RECT  5.810000  29.275000  6.610000  30.075000 ;
      RECT  5.815000   2.450000  6.615000   3.250000 ;
      RECT  5.815000   4.360000  6.615000   5.160000 ;
      RECT  5.815000   6.270000  6.615000   7.070000 ;
      RECT  5.815000  15.345000  6.615000  16.145000 ;
      RECT  5.815000  17.175000  6.615000  17.975000 ;
      RECT  5.815000  32.295000  6.615000  33.095000 ;
      RECT  5.815000  34.125000  6.615000  34.925000 ;
      RECT  5.815000  37.145000  6.615000  37.945000 ;
      RECT  5.815000  38.975000  6.615000  39.775000 ;
      RECT  5.815000  41.995000  6.615000  42.795000 ;
      RECT  5.815000  45.025000  6.615000  45.825000 ;
      RECT  5.815000  51.835000  6.615000  52.635000 ;
      RECT  5.815000  58.645000  6.615000  59.445000 ;
      RECT  5.815000  61.475000  6.615000  62.275000 ;
      RECT  5.815000  64.495000  6.615000  65.295000 ;
      RECT  5.815000  67.325000  6.615000  68.125000 ;
      RECT  5.815000  70.350000  6.615000  71.150000 ;
      RECT  5.815000  72.030000  6.615000  72.830000 ;
      RECT  5.815000  73.710000  6.615000  74.510000 ;
      RECT  5.815000  75.390000  6.615000  76.190000 ;
      RECT  5.815000  77.070000  6.615000  77.870000 ;
      RECT  5.815000  78.750000  6.615000  79.550000 ;
      RECT  5.815000  80.430000  6.615000  81.230000 ;
      RECT  5.815000  82.110000  6.615000  82.910000 ;
      RECT  5.815000  83.790000  6.615000  84.590000 ;
      RECT  5.815000  85.470000  6.615000  86.270000 ;
      RECT  5.815000  87.150000  6.615000  87.950000 ;
      RECT  5.815000  88.830000  6.615000  89.630000 ;
      RECT  5.815000  90.510000  6.615000  91.310000 ;
      RECT  5.815000  92.190000  6.615000  92.990000 ;
      RECT  5.815000  93.870000  6.615000  94.670000 ;
      RECT  5.815000 176.155000  6.615000 176.955000 ;
      RECT  5.815000 177.775000  6.615000 178.575000 ;
      RECT  5.815000 179.395000  6.615000 180.195000 ;
      RECT  5.815000 181.015000  6.615000 181.815000 ;
      RECT  5.815000 182.635000  6.615000 183.435000 ;
      RECT  5.815000 184.255000  6.615000 185.055000 ;
      RECT  5.815000 185.875000  6.615000 186.675000 ;
      RECT  5.815000 187.495000  6.615000 188.295000 ;
      RECT  5.815000 189.115000  6.615000 189.915000 ;
      RECT  5.815000 190.735000  6.615000 191.535000 ;
      RECT  5.815000 192.355000  6.615000 193.155000 ;
      RECT  5.815000 193.975000  6.615000 194.775000 ;
      RECT  5.815000 195.595000  6.615000 196.395000 ;
      RECT  5.815000 197.215000  6.615000 198.015000 ;
      RECT  5.815000 198.835000  6.615000 199.635000 ;
      RECT  5.820000   9.295000  6.620000  10.095000 ;
      RECT  5.820000  12.325000  6.620000  13.125000 ;
      RECT  7.415000  20.195000  8.215000  20.995000 ;
      RECT  7.415000  23.225000  8.215000  24.025000 ;
      RECT  7.415000  26.245000  8.215000  27.045000 ;
      RECT  7.415000  29.275000  8.215000  30.075000 ;
      RECT  7.420000   2.450000  8.220000   3.250000 ;
      RECT  7.420000   4.360000  8.220000   5.160000 ;
      RECT  7.420000   6.270000  8.220000   7.070000 ;
      RECT  7.420000  15.345000  8.220000  16.145000 ;
      RECT  7.420000  17.175000  8.220000  17.975000 ;
      RECT  7.420000  32.295000  8.220000  33.095000 ;
      RECT  7.420000  34.125000  8.220000  34.925000 ;
      RECT  7.420000  37.145000  8.220000  37.945000 ;
      RECT  7.420000  38.975000  8.220000  39.775000 ;
      RECT  7.420000  41.995000  8.220000  42.795000 ;
      RECT  7.420000  45.025000  8.220000  45.825000 ;
      RECT  7.420000  51.835000  8.220000  52.635000 ;
      RECT  7.420000  58.645000  8.220000  59.445000 ;
      RECT  7.420000  61.475000  8.220000  62.275000 ;
      RECT  7.420000  64.495000  8.220000  65.295000 ;
      RECT  7.420000  67.325000  8.220000  68.125000 ;
      RECT  7.420000  70.350000  8.220000  71.150000 ;
      RECT  7.420000  72.030000  8.220000  72.830000 ;
      RECT  7.420000  73.710000  8.220000  74.510000 ;
      RECT  7.420000  75.390000  8.220000  76.190000 ;
      RECT  7.420000  77.070000  8.220000  77.870000 ;
      RECT  7.420000  78.750000  8.220000  79.550000 ;
      RECT  7.420000  80.430000  8.220000  81.230000 ;
      RECT  7.420000  82.110000  8.220000  82.910000 ;
      RECT  7.420000  83.790000  8.220000  84.590000 ;
      RECT  7.420000  85.470000  8.220000  86.270000 ;
      RECT  7.420000  87.150000  8.220000  87.950000 ;
      RECT  7.420000  88.830000  8.220000  89.630000 ;
      RECT  7.420000  90.510000  8.220000  91.310000 ;
      RECT  7.420000  92.190000  8.220000  92.990000 ;
      RECT  7.420000  93.870000  8.220000  94.670000 ;
      RECT  7.420000 176.155000  8.220000 176.955000 ;
      RECT  7.420000 177.775000  8.220000 178.575000 ;
      RECT  7.420000 179.395000  8.220000 180.195000 ;
      RECT  7.420000 181.015000  8.220000 181.815000 ;
      RECT  7.420000 182.635000  8.220000 183.435000 ;
      RECT  7.420000 184.255000  8.220000 185.055000 ;
      RECT  7.420000 185.875000  8.220000 186.675000 ;
      RECT  7.420000 187.495000  8.220000 188.295000 ;
      RECT  7.420000 189.115000  8.220000 189.915000 ;
      RECT  7.420000 190.735000  8.220000 191.535000 ;
      RECT  7.420000 192.355000  8.220000 193.155000 ;
      RECT  7.420000 193.975000  8.220000 194.775000 ;
      RECT  7.420000 195.595000  8.220000 196.395000 ;
      RECT  7.420000 197.215000  8.220000 198.015000 ;
      RECT  7.420000 198.835000  8.220000 199.635000 ;
      RECT  7.425000   9.295000  8.225000  10.095000 ;
      RECT  7.425000  12.325000  8.225000  13.125000 ;
      RECT  9.020000  20.195000  9.820000  20.995000 ;
      RECT  9.020000  23.225000  9.820000  24.025000 ;
      RECT  9.020000  26.245000  9.820000  27.045000 ;
      RECT  9.020000  29.275000  9.820000  30.075000 ;
      RECT  9.025000   2.450000  9.825000   3.250000 ;
      RECT  9.025000   4.360000  9.825000   5.160000 ;
      RECT  9.025000   6.270000  9.825000   7.070000 ;
      RECT  9.025000  15.345000  9.825000  16.145000 ;
      RECT  9.025000  17.175000  9.825000  17.975000 ;
      RECT  9.025000  32.295000  9.825000  33.095000 ;
      RECT  9.025000  34.125000  9.825000  34.925000 ;
      RECT  9.025000  37.145000  9.825000  37.945000 ;
      RECT  9.025000  38.975000  9.825000  39.775000 ;
      RECT  9.025000  41.995000  9.825000  42.795000 ;
      RECT  9.025000  45.025000  9.825000  45.825000 ;
      RECT  9.025000  51.835000  9.825000  52.635000 ;
      RECT  9.025000  58.645000  9.825000  59.445000 ;
      RECT  9.025000  61.475000  9.825000  62.275000 ;
      RECT  9.025000  64.495000  9.825000  65.295000 ;
      RECT  9.025000  67.325000  9.825000  68.125000 ;
      RECT  9.025000  70.350000  9.825000  71.150000 ;
      RECT  9.025000  72.030000  9.825000  72.830000 ;
      RECT  9.025000  73.710000  9.825000  74.510000 ;
      RECT  9.025000  75.390000  9.825000  76.190000 ;
      RECT  9.025000  77.070000  9.825000  77.870000 ;
      RECT  9.025000  78.750000  9.825000  79.550000 ;
      RECT  9.025000  80.430000  9.825000  81.230000 ;
      RECT  9.025000  82.110000  9.825000  82.910000 ;
      RECT  9.025000  83.790000  9.825000  84.590000 ;
      RECT  9.025000  85.470000  9.825000  86.270000 ;
      RECT  9.025000  87.150000  9.825000  87.950000 ;
      RECT  9.025000  88.830000  9.825000  89.630000 ;
      RECT  9.025000  90.510000  9.825000  91.310000 ;
      RECT  9.025000  92.190000  9.825000  92.990000 ;
      RECT  9.025000  93.870000  9.825000  94.670000 ;
      RECT  9.025000 176.155000  9.825000 176.955000 ;
      RECT  9.025000 177.775000  9.825000 178.575000 ;
      RECT  9.025000 179.395000  9.825000 180.195000 ;
      RECT  9.025000 181.015000  9.825000 181.815000 ;
      RECT  9.025000 182.635000  9.825000 183.435000 ;
      RECT  9.025000 184.255000  9.825000 185.055000 ;
      RECT  9.025000 185.875000  9.825000 186.675000 ;
      RECT  9.025000 187.495000  9.825000 188.295000 ;
      RECT  9.025000 189.115000  9.825000 189.915000 ;
      RECT  9.025000 190.735000  9.825000 191.535000 ;
      RECT  9.025000 192.355000  9.825000 193.155000 ;
      RECT  9.025000 193.975000  9.825000 194.775000 ;
      RECT  9.025000 195.595000  9.825000 196.395000 ;
      RECT  9.025000 197.215000  9.825000 198.015000 ;
      RECT  9.025000 198.835000  9.825000 199.635000 ;
      RECT  9.030000   9.295000  9.830000  10.095000 ;
      RECT  9.030000  12.325000  9.830000  13.125000 ;
      RECT 10.625000  20.195000 11.425000  20.995000 ;
      RECT 10.625000  23.225000 11.425000  24.025000 ;
      RECT 10.625000  26.245000 11.425000  27.045000 ;
      RECT 10.625000  29.275000 11.425000  30.075000 ;
      RECT 10.630000   2.450000 11.430000   3.250000 ;
      RECT 10.630000   4.360000 11.430000   5.160000 ;
      RECT 10.630000   6.270000 11.430000   7.070000 ;
      RECT 10.630000  15.345000 11.430000  16.145000 ;
      RECT 10.630000  17.175000 11.430000  17.975000 ;
      RECT 10.630000  32.295000 11.430000  33.095000 ;
      RECT 10.630000  34.125000 11.430000  34.925000 ;
      RECT 10.630000  37.145000 11.430000  37.945000 ;
      RECT 10.630000  38.975000 11.430000  39.775000 ;
      RECT 10.630000  41.995000 11.430000  42.795000 ;
      RECT 10.630000  45.025000 11.430000  45.825000 ;
      RECT 10.630000  51.835000 11.430000  52.635000 ;
      RECT 10.630000  58.645000 11.430000  59.445000 ;
      RECT 10.630000  61.475000 11.430000  62.275000 ;
      RECT 10.630000  64.495000 11.430000  65.295000 ;
      RECT 10.630000  67.325000 11.430000  68.125000 ;
      RECT 10.630000  70.350000 11.430000  71.150000 ;
      RECT 10.630000  72.030000 11.430000  72.830000 ;
      RECT 10.630000  73.710000 11.430000  74.510000 ;
      RECT 10.630000  75.390000 11.430000  76.190000 ;
      RECT 10.630000  77.070000 11.430000  77.870000 ;
      RECT 10.630000  78.750000 11.430000  79.550000 ;
      RECT 10.630000  80.430000 11.430000  81.230000 ;
      RECT 10.630000  82.110000 11.430000  82.910000 ;
      RECT 10.630000  83.790000 11.430000  84.590000 ;
      RECT 10.630000  85.470000 11.430000  86.270000 ;
      RECT 10.630000  87.150000 11.430000  87.950000 ;
      RECT 10.630000  88.830000 11.430000  89.630000 ;
      RECT 10.630000  90.510000 11.430000  91.310000 ;
      RECT 10.630000  92.190000 11.430000  92.990000 ;
      RECT 10.630000  93.870000 11.430000  94.670000 ;
      RECT 10.630000 176.155000 11.430000 176.955000 ;
      RECT 10.630000 177.775000 11.430000 178.575000 ;
      RECT 10.630000 179.395000 11.430000 180.195000 ;
      RECT 10.630000 181.015000 11.430000 181.815000 ;
      RECT 10.630000 182.635000 11.430000 183.435000 ;
      RECT 10.630000 184.255000 11.430000 185.055000 ;
      RECT 10.630000 185.875000 11.430000 186.675000 ;
      RECT 10.630000 187.495000 11.430000 188.295000 ;
      RECT 10.630000 189.115000 11.430000 189.915000 ;
      RECT 10.630000 190.735000 11.430000 191.535000 ;
      RECT 10.630000 192.355000 11.430000 193.155000 ;
      RECT 10.630000 193.975000 11.430000 194.775000 ;
      RECT 10.630000 195.595000 11.430000 196.395000 ;
      RECT 10.630000 197.215000 11.430000 198.015000 ;
      RECT 10.630000 198.835000 11.430000 199.635000 ;
      RECT 10.635000   9.295000 11.435000  10.095000 ;
      RECT 10.635000  12.325000 11.435000  13.125000 ;
      RECT 12.230000  20.195000 13.030000  20.995000 ;
      RECT 12.230000  23.225000 13.030000  24.025000 ;
      RECT 12.230000  26.245000 13.030000  27.045000 ;
      RECT 12.230000  29.275000 13.030000  30.075000 ;
      RECT 12.235000   2.450000 13.035000   3.250000 ;
      RECT 12.235000   4.360000 13.035000   5.160000 ;
      RECT 12.235000   6.270000 13.035000   7.070000 ;
      RECT 12.235000  15.345000 13.035000  16.145000 ;
      RECT 12.235000  17.175000 13.035000  17.975000 ;
      RECT 12.235000  32.295000 13.035000  33.095000 ;
      RECT 12.235000  34.125000 13.035000  34.925000 ;
      RECT 12.235000  37.145000 13.035000  37.945000 ;
      RECT 12.235000  38.975000 13.035000  39.775000 ;
      RECT 12.235000  41.995000 13.035000  42.795000 ;
      RECT 12.235000  45.025000 13.035000  45.825000 ;
      RECT 12.235000  51.835000 13.035000  52.635000 ;
      RECT 12.235000  58.645000 13.035000  59.445000 ;
      RECT 12.235000  61.475000 13.035000  62.275000 ;
      RECT 12.235000  64.495000 13.035000  65.295000 ;
      RECT 12.235000  67.325000 13.035000  68.125000 ;
      RECT 12.235000  70.350000 13.035000  71.150000 ;
      RECT 12.235000  72.030000 13.035000  72.830000 ;
      RECT 12.235000  73.710000 13.035000  74.510000 ;
      RECT 12.235000  75.390000 13.035000  76.190000 ;
      RECT 12.235000  77.070000 13.035000  77.870000 ;
      RECT 12.235000  78.750000 13.035000  79.550000 ;
      RECT 12.235000  80.430000 13.035000  81.230000 ;
      RECT 12.235000  82.110000 13.035000  82.910000 ;
      RECT 12.235000  83.790000 13.035000  84.590000 ;
      RECT 12.235000  85.470000 13.035000  86.270000 ;
      RECT 12.235000  87.150000 13.035000  87.950000 ;
      RECT 12.235000  88.830000 13.035000  89.630000 ;
      RECT 12.235000  90.510000 13.035000  91.310000 ;
      RECT 12.235000  92.190000 13.035000  92.990000 ;
      RECT 12.235000  93.870000 13.035000  94.670000 ;
      RECT 12.235000 176.155000 13.035000 176.955000 ;
      RECT 12.235000 177.775000 13.035000 178.575000 ;
      RECT 12.235000 179.395000 13.035000 180.195000 ;
      RECT 12.235000 181.015000 13.035000 181.815000 ;
      RECT 12.235000 182.635000 13.035000 183.435000 ;
      RECT 12.235000 184.255000 13.035000 185.055000 ;
      RECT 12.235000 185.875000 13.035000 186.675000 ;
      RECT 12.235000 187.495000 13.035000 188.295000 ;
      RECT 12.235000 189.115000 13.035000 189.915000 ;
      RECT 12.235000 190.735000 13.035000 191.535000 ;
      RECT 12.235000 192.355000 13.035000 193.155000 ;
      RECT 12.235000 193.975000 13.035000 194.775000 ;
      RECT 12.235000 195.595000 13.035000 196.395000 ;
      RECT 12.235000 197.215000 13.035000 198.015000 ;
      RECT 12.235000 198.835000 13.035000 199.635000 ;
      RECT 12.240000   9.295000 13.040000  10.095000 ;
      RECT 12.240000  12.325000 13.040000  13.125000 ;
      RECT 13.835000  20.195000 14.635000  20.995000 ;
      RECT 13.835000  23.225000 14.635000  24.025000 ;
      RECT 13.835000  26.245000 14.635000  27.045000 ;
      RECT 13.835000  29.275000 14.635000  30.075000 ;
      RECT 13.840000   2.450000 14.640000   3.250000 ;
      RECT 13.840000   4.360000 14.640000   5.160000 ;
      RECT 13.840000   6.270000 14.640000   7.070000 ;
      RECT 13.840000  15.345000 14.640000  16.145000 ;
      RECT 13.840000  17.175000 14.640000  17.975000 ;
      RECT 13.840000  32.295000 14.640000  33.095000 ;
      RECT 13.840000  34.125000 14.640000  34.925000 ;
      RECT 13.840000  37.145000 14.640000  37.945000 ;
      RECT 13.840000  38.975000 14.640000  39.775000 ;
      RECT 13.840000  41.995000 14.640000  42.795000 ;
      RECT 13.840000  45.025000 14.640000  45.825000 ;
      RECT 13.840000  51.835000 14.640000  52.635000 ;
      RECT 13.840000  58.645000 14.640000  59.445000 ;
      RECT 13.840000  61.475000 14.640000  62.275000 ;
      RECT 13.840000  64.495000 14.640000  65.295000 ;
      RECT 13.840000  67.325000 14.640000  68.125000 ;
      RECT 13.840000  70.350000 14.640000  71.150000 ;
      RECT 13.840000  72.030000 14.640000  72.830000 ;
      RECT 13.840000  73.710000 14.640000  74.510000 ;
      RECT 13.840000  75.390000 14.640000  76.190000 ;
      RECT 13.840000  77.070000 14.640000  77.870000 ;
      RECT 13.840000  78.750000 14.640000  79.550000 ;
      RECT 13.840000  80.430000 14.640000  81.230000 ;
      RECT 13.840000  82.110000 14.640000  82.910000 ;
      RECT 13.840000  83.790000 14.640000  84.590000 ;
      RECT 13.840000  85.470000 14.640000  86.270000 ;
      RECT 13.840000  87.150000 14.640000  87.950000 ;
      RECT 13.840000  88.830000 14.640000  89.630000 ;
      RECT 13.840000  90.510000 14.640000  91.310000 ;
      RECT 13.840000  92.190000 14.640000  92.990000 ;
      RECT 13.840000  93.870000 14.640000  94.670000 ;
      RECT 13.840000 176.155000 14.640000 176.955000 ;
      RECT 13.840000 177.775000 14.640000 178.575000 ;
      RECT 13.840000 179.395000 14.640000 180.195000 ;
      RECT 13.840000 181.015000 14.640000 181.815000 ;
      RECT 13.840000 182.635000 14.640000 183.435000 ;
      RECT 13.840000 184.255000 14.640000 185.055000 ;
      RECT 13.840000 185.875000 14.640000 186.675000 ;
      RECT 13.840000 187.495000 14.640000 188.295000 ;
      RECT 13.840000 189.115000 14.640000 189.915000 ;
      RECT 13.840000 190.735000 14.640000 191.535000 ;
      RECT 13.840000 192.355000 14.640000 193.155000 ;
      RECT 13.840000 193.975000 14.640000 194.775000 ;
      RECT 13.840000 195.595000 14.640000 196.395000 ;
      RECT 13.840000 197.215000 14.640000 198.015000 ;
      RECT 13.840000 198.835000 14.640000 199.635000 ;
      RECT 13.845000   9.295000 14.645000  10.095000 ;
      RECT 13.845000  12.325000 14.645000  13.125000 ;
      RECT 15.440000  20.195000 16.240000  20.995000 ;
      RECT 15.440000  23.225000 16.240000  24.025000 ;
      RECT 15.440000  26.245000 16.240000  27.045000 ;
      RECT 15.440000  29.275000 16.240000  30.075000 ;
      RECT 15.445000   2.450000 16.245000   3.250000 ;
      RECT 15.445000   4.360000 16.245000   5.160000 ;
      RECT 15.445000   6.270000 16.245000   7.070000 ;
      RECT 15.445000  15.345000 16.245000  16.145000 ;
      RECT 15.445000  17.175000 16.245000  17.975000 ;
      RECT 15.445000  32.295000 16.245000  33.095000 ;
      RECT 15.445000  34.125000 16.245000  34.925000 ;
      RECT 15.445000  37.145000 16.245000  37.945000 ;
      RECT 15.445000  38.975000 16.245000  39.775000 ;
      RECT 15.445000  41.995000 16.245000  42.795000 ;
      RECT 15.445000  45.025000 16.245000  45.825000 ;
      RECT 15.445000  51.835000 16.245000  52.635000 ;
      RECT 15.445000  58.645000 16.245000  59.445000 ;
      RECT 15.445000  61.475000 16.245000  62.275000 ;
      RECT 15.445000  64.495000 16.245000  65.295000 ;
      RECT 15.445000  67.325000 16.245000  68.125000 ;
      RECT 15.445000  70.350000 16.245000  71.150000 ;
      RECT 15.445000  72.030000 16.245000  72.830000 ;
      RECT 15.445000  73.710000 16.245000  74.510000 ;
      RECT 15.445000  75.390000 16.245000  76.190000 ;
      RECT 15.445000  77.070000 16.245000  77.870000 ;
      RECT 15.445000  78.750000 16.245000  79.550000 ;
      RECT 15.445000  80.430000 16.245000  81.230000 ;
      RECT 15.445000  82.110000 16.245000  82.910000 ;
      RECT 15.445000  83.790000 16.245000  84.590000 ;
      RECT 15.445000  85.470000 16.245000  86.270000 ;
      RECT 15.445000  87.150000 16.245000  87.950000 ;
      RECT 15.445000  88.830000 16.245000  89.630000 ;
      RECT 15.445000  90.510000 16.245000  91.310000 ;
      RECT 15.445000  92.190000 16.245000  92.990000 ;
      RECT 15.445000  93.870000 16.245000  94.670000 ;
      RECT 15.445000 176.155000 16.245000 176.955000 ;
      RECT 15.445000 177.775000 16.245000 178.575000 ;
      RECT 15.445000 179.395000 16.245000 180.195000 ;
      RECT 15.445000 181.015000 16.245000 181.815000 ;
      RECT 15.445000 182.635000 16.245000 183.435000 ;
      RECT 15.445000 184.255000 16.245000 185.055000 ;
      RECT 15.445000 185.875000 16.245000 186.675000 ;
      RECT 15.445000 187.495000 16.245000 188.295000 ;
      RECT 15.445000 189.115000 16.245000 189.915000 ;
      RECT 15.445000 190.735000 16.245000 191.535000 ;
      RECT 15.445000 192.355000 16.245000 193.155000 ;
      RECT 15.445000 193.975000 16.245000 194.775000 ;
      RECT 15.445000 195.595000 16.245000 196.395000 ;
      RECT 15.445000 197.215000 16.245000 198.015000 ;
      RECT 15.445000 198.835000 16.245000 199.635000 ;
      RECT 15.450000   9.295000 16.250000  10.095000 ;
      RECT 15.450000  12.325000 16.250000  13.125000 ;
      RECT 17.045000  20.195000 17.845000  20.995000 ;
      RECT 17.045000  23.225000 17.845000  24.025000 ;
      RECT 17.045000  26.245000 17.845000  27.045000 ;
      RECT 17.045000  29.275000 17.845000  30.075000 ;
      RECT 17.050000   2.450000 17.850000   3.250000 ;
      RECT 17.050000   4.360000 17.850000   5.160000 ;
      RECT 17.050000   6.270000 17.850000   7.070000 ;
      RECT 17.050000  15.345000 17.850000  16.145000 ;
      RECT 17.050000  17.175000 17.850000  17.975000 ;
      RECT 17.050000  32.295000 17.850000  33.095000 ;
      RECT 17.050000  34.125000 17.850000  34.925000 ;
      RECT 17.050000  37.145000 17.850000  37.945000 ;
      RECT 17.050000  38.975000 17.850000  39.775000 ;
      RECT 17.050000  41.995000 17.850000  42.795000 ;
      RECT 17.050000  45.025000 17.850000  45.825000 ;
      RECT 17.050000  51.835000 17.850000  52.635000 ;
      RECT 17.050000  58.645000 17.850000  59.445000 ;
      RECT 17.050000  61.475000 17.850000  62.275000 ;
      RECT 17.050000  64.495000 17.850000  65.295000 ;
      RECT 17.050000  67.325000 17.850000  68.125000 ;
      RECT 17.050000  70.350000 17.850000  71.150000 ;
      RECT 17.050000  72.030000 17.850000  72.830000 ;
      RECT 17.050000  73.710000 17.850000  74.510000 ;
      RECT 17.050000  75.390000 17.850000  76.190000 ;
      RECT 17.050000  77.070000 17.850000  77.870000 ;
      RECT 17.050000  78.750000 17.850000  79.550000 ;
      RECT 17.050000  80.430000 17.850000  81.230000 ;
      RECT 17.050000  82.110000 17.850000  82.910000 ;
      RECT 17.050000  83.790000 17.850000  84.590000 ;
      RECT 17.050000  85.470000 17.850000  86.270000 ;
      RECT 17.050000  87.150000 17.850000  87.950000 ;
      RECT 17.050000  88.830000 17.850000  89.630000 ;
      RECT 17.050000  90.510000 17.850000  91.310000 ;
      RECT 17.050000  92.190000 17.850000  92.990000 ;
      RECT 17.050000  93.870000 17.850000  94.670000 ;
      RECT 17.050000 176.155000 17.850000 176.955000 ;
      RECT 17.050000 177.775000 17.850000 178.575000 ;
      RECT 17.050000 179.395000 17.850000 180.195000 ;
      RECT 17.050000 181.015000 17.850000 181.815000 ;
      RECT 17.050000 182.635000 17.850000 183.435000 ;
      RECT 17.050000 184.255000 17.850000 185.055000 ;
      RECT 17.050000 185.875000 17.850000 186.675000 ;
      RECT 17.050000 187.495000 17.850000 188.295000 ;
      RECT 17.050000 189.115000 17.850000 189.915000 ;
      RECT 17.050000 190.735000 17.850000 191.535000 ;
      RECT 17.050000 192.355000 17.850000 193.155000 ;
      RECT 17.050000 193.975000 17.850000 194.775000 ;
      RECT 17.050000 195.595000 17.850000 196.395000 ;
      RECT 17.050000 197.215000 17.850000 198.015000 ;
      RECT 17.050000 198.835000 17.850000 199.635000 ;
      RECT 17.055000   9.295000 17.855000  10.095000 ;
      RECT 17.055000  12.325000 17.855000  13.125000 ;
      RECT 18.650000  20.195000 19.450000  20.995000 ;
      RECT 18.650000  23.225000 19.450000  24.025000 ;
      RECT 18.650000  26.245000 19.450000  27.045000 ;
      RECT 18.650000  29.275000 19.450000  30.075000 ;
      RECT 18.655000   2.450000 19.455000   3.250000 ;
      RECT 18.655000   4.360000 19.455000   5.160000 ;
      RECT 18.655000   6.270000 19.455000   7.070000 ;
      RECT 18.655000  15.345000 19.455000  16.145000 ;
      RECT 18.655000  17.175000 19.455000  17.975000 ;
      RECT 18.655000  32.295000 19.455000  33.095000 ;
      RECT 18.655000  34.125000 19.455000  34.925000 ;
      RECT 18.655000  37.145000 19.455000  37.945000 ;
      RECT 18.655000  38.975000 19.455000  39.775000 ;
      RECT 18.655000  41.995000 19.455000  42.795000 ;
      RECT 18.655000  45.025000 19.455000  45.825000 ;
      RECT 18.655000  51.835000 19.455000  52.635000 ;
      RECT 18.655000  58.645000 19.455000  59.445000 ;
      RECT 18.655000  61.475000 19.455000  62.275000 ;
      RECT 18.655000  64.495000 19.455000  65.295000 ;
      RECT 18.655000  67.325000 19.455000  68.125000 ;
      RECT 18.655000  70.350000 19.455000  71.150000 ;
      RECT 18.655000  72.030000 19.455000  72.830000 ;
      RECT 18.655000  73.710000 19.455000  74.510000 ;
      RECT 18.655000  75.390000 19.455000  76.190000 ;
      RECT 18.655000  77.070000 19.455000  77.870000 ;
      RECT 18.655000  78.750000 19.455000  79.550000 ;
      RECT 18.655000  80.430000 19.455000  81.230000 ;
      RECT 18.655000  82.110000 19.455000  82.910000 ;
      RECT 18.655000  83.790000 19.455000  84.590000 ;
      RECT 18.655000  85.470000 19.455000  86.270000 ;
      RECT 18.655000  87.150000 19.455000  87.950000 ;
      RECT 18.655000  88.830000 19.455000  89.630000 ;
      RECT 18.655000  90.510000 19.455000  91.310000 ;
      RECT 18.655000  92.190000 19.455000  92.990000 ;
      RECT 18.655000  93.870000 19.455000  94.670000 ;
      RECT 18.655000 176.155000 19.455000 176.955000 ;
      RECT 18.655000 177.775000 19.455000 178.575000 ;
      RECT 18.655000 179.395000 19.455000 180.195000 ;
      RECT 18.655000 181.015000 19.455000 181.815000 ;
      RECT 18.655000 182.635000 19.455000 183.435000 ;
      RECT 18.655000 184.255000 19.455000 185.055000 ;
      RECT 18.655000 185.875000 19.455000 186.675000 ;
      RECT 18.655000 187.495000 19.455000 188.295000 ;
      RECT 18.655000 189.115000 19.455000 189.915000 ;
      RECT 18.655000 190.735000 19.455000 191.535000 ;
      RECT 18.655000 192.355000 19.455000 193.155000 ;
      RECT 18.655000 193.975000 19.455000 194.775000 ;
      RECT 18.655000 195.595000 19.455000 196.395000 ;
      RECT 18.655000 197.215000 19.455000 198.015000 ;
      RECT 18.655000 198.835000 19.455000 199.635000 ;
      RECT 18.660000   9.295000 19.460000  10.095000 ;
      RECT 18.660000  12.325000 19.460000  13.125000 ;
      RECT 20.255000  20.195000 21.055000  20.995000 ;
      RECT 20.255000  23.225000 21.055000  24.025000 ;
      RECT 20.255000  26.245000 21.055000  27.045000 ;
      RECT 20.255000  29.275000 21.055000  30.075000 ;
      RECT 20.260000   2.450000 21.060000   3.250000 ;
      RECT 20.260000   4.360000 21.060000   5.160000 ;
      RECT 20.260000   6.270000 21.060000   7.070000 ;
      RECT 20.260000  15.345000 21.060000  16.145000 ;
      RECT 20.260000  17.175000 21.060000  17.975000 ;
      RECT 20.260000  32.295000 21.060000  33.095000 ;
      RECT 20.260000  34.125000 21.060000  34.925000 ;
      RECT 20.260000  37.145000 21.060000  37.945000 ;
      RECT 20.260000  38.975000 21.060000  39.775000 ;
      RECT 20.260000  41.995000 21.060000  42.795000 ;
      RECT 20.260000  45.025000 21.060000  45.825000 ;
      RECT 20.260000  51.835000 21.060000  52.635000 ;
      RECT 20.260000  58.645000 21.060000  59.445000 ;
      RECT 20.260000  61.475000 21.060000  62.275000 ;
      RECT 20.260000  64.495000 21.060000  65.295000 ;
      RECT 20.260000  67.325000 21.060000  68.125000 ;
      RECT 20.260000  70.350000 21.060000  71.150000 ;
      RECT 20.260000  72.030000 21.060000  72.830000 ;
      RECT 20.260000  73.710000 21.060000  74.510000 ;
      RECT 20.260000  75.390000 21.060000  76.190000 ;
      RECT 20.260000  77.070000 21.060000  77.870000 ;
      RECT 20.260000  78.750000 21.060000  79.550000 ;
      RECT 20.260000  80.430000 21.060000  81.230000 ;
      RECT 20.260000  82.110000 21.060000  82.910000 ;
      RECT 20.260000  83.790000 21.060000  84.590000 ;
      RECT 20.260000  85.470000 21.060000  86.270000 ;
      RECT 20.260000  87.150000 21.060000  87.950000 ;
      RECT 20.260000  88.830000 21.060000  89.630000 ;
      RECT 20.260000  90.510000 21.060000  91.310000 ;
      RECT 20.260000  92.190000 21.060000  92.990000 ;
      RECT 20.260000  93.870000 21.060000  94.670000 ;
      RECT 20.260000 176.155000 21.060000 176.955000 ;
      RECT 20.260000 177.775000 21.060000 178.575000 ;
      RECT 20.260000 179.395000 21.060000 180.195000 ;
      RECT 20.260000 181.015000 21.060000 181.815000 ;
      RECT 20.260000 182.635000 21.060000 183.435000 ;
      RECT 20.260000 184.255000 21.060000 185.055000 ;
      RECT 20.260000 185.875000 21.060000 186.675000 ;
      RECT 20.260000 187.495000 21.060000 188.295000 ;
      RECT 20.260000 189.115000 21.060000 189.915000 ;
      RECT 20.260000 190.735000 21.060000 191.535000 ;
      RECT 20.260000 192.355000 21.060000 193.155000 ;
      RECT 20.260000 193.975000 21.060000 194.775000 ;
      RECT 20.260000 195.595000 21.060000 196.395000 ;
      RECT 20.260000 197.215000 21.060000 198.015000 ;
      RECT 20.260000 198.835000 21.060000 199.635000 ;
      RECT 20.265000   9.295000 21.065000  10.095000 ;
      RECT 20.265000  12.325000 21.065000  13.125000 ;
      RECT 21.860000  20.195000 22.660000  20.995000 ;
      RECT 21.860000  23.225000 22.660000  24.025000 ;
      RECT 21.860000  26.245000 22.660000  27.045000 ;
      RECT 21.860000  29.275000 22.660000  30.075000 ;
      RECT 21.865000   2.450000 22.665000   3.250000 ;
      RECT 21.865000   4.360000 22.665000   5.160000 ;
      RECT 21.865000   6.270000 22.665000   7.070000 ;
      RECT 21.865000  15.345000 22.665000  16.145000 ;
      RECT 21.865000  17.175000 22.665000  17.975000 ;
      RECT 21.865000  32.295000 22.665000  33.095000 ;
      RECT 21.865000  34.125000 22.665000  34.925000 ;
      RECT 21.865000  37.145000 22.665000  37.945000 ;
      RECT 21.865000  38.975000 22.665000  39.775000 ;
      RECT 21.865000  41.995000 22.665000  42.795000 ;
      RECT 21.865000  45.025000 22.665000  45.825000 ;
      RECT 21.865000  51.835000 22.665000  52.635000 ;
      RECT 21.865000  58.645000 22.665000  59.445000 ;
      RECT 21.865000  61.475000 22.665000  62.275000 ;
      RECT 21.865000  64.495000 22.665000  65.295000 ;
      RECT 21.865000  67.325000 22.665000  68.125000 ;
      RECT 21.865000  70.350000 22.665000  71.150000 ;
      RECT 21.865000  72.030000 22.665000  72.830000 ;
      RECT 21.865000  73.710000 22.665000  74.510000 ;
      RECT 21.865000  75.390000 22.665000  76.190000 ;
      RECT 21.865000  77.070000 22.665000  77.870000 ;
      RECT 21.865000  78.750000 22.665000  79.550000 ;
      RECT 21.865000  80.430000 22.665000  81.230000 ;
      RECT 21.865000  82.110000 22.665000  82.910000 ;
      RECT 21.865000  83.790000 22.665000  84.590000 ;
      RECT 21.865000  85.470000 22.665000  86.270000 ;
      RECT 21.865000  87.150000 22.665000  87.950000 ;
      RECT 21.865000  88.830000 22.665000  89.630000 ;
      RECT 21.865000  90.510000 22.665000  91.310000 ;
      RECT 21.865000  92.190000 22.665000  92.990000 ;
      RECT 21.865000  93.870000 22.665000  94.670000 ;
      RECT 21.865000 176.155000 22.665000 176.955000 ;
      RECT 21.865000 177.775000 22.665000 178.575000 ;
      RECT 21.865000 179.395000 22.665000 180.195000 ;
      RECT 21.865000 181.015000 22.665000 181.815000 ;
      RECT 21.865000 182.635000 22.665000 183.435000 ;
      RECT 21.865000 184.255000 22.665000 185.055000 ;
      RECT 21.865000 185.875000 22.665000 186.675000 ;
      RECT 21.865000 187.495000 22.665000 188.295000 ;
      RECT 21.865000 189.115000 22.665000 189.915000 ;
      RECT 21.865000 190.735000 22.665000 191.535000 ;
      RECT 21.865000 192.355000 22.665000 193.155000 ;
      RECT 21.865000 193.975000 22.665000 194.775000 ;
      RECT 21.865000 195.595000 22.665000 196.395000 ;
      RECT 21.865000 197.215000 22.665000 198.015000 ;
      RECT 21.865000 198.835000 22.665000 199.635000 ;
      RECT 21.870000   9.295000 22.670000  10.095000 ;
      RECT 21.870000  12.325000 22.670000  13.125000 ;
      RECT 23.465000  20.195000 24.265000  20.995000 ;
      RECT 23.465000  23.225000 24.265000  24.025000 ;
      RECT 23.465000  26.245000 24.265000  27.045000 ;
      RECT 23.465000  29.275000 24.265000  30.075000 ;
      RECT 23.470000   2.450000 24.270000   3.250000 ;
      RECT 23.470000   4.360000 24.270000   5.160000 ;
      RECT 23.470000   6.270000 24.270000   7.070000 ;
      RECT 23.470000  15.345000 24.270000  16.145000 ;
      RECT 23.470000  17.175000 24.270000  17.975000 ;
      RECT 23.470000  32.295000 24.270000  33.095000 ;
      RECT 23.470000  34.125000 24.270000  34.925000 ;
      RECT 23.470000  37.145000 24.270000  37.945000 ;
      RECT 23.470000  38.975000 24.270000  39.775000 ;
      RECT 23.470000  41.995000 24.270000  42.795000 ;
      RECT 23.470000  45.025000 24.270000  45.825000 ;
      RECT 23.470000  51.835000 24.270000  52.635000 ;
      RECT 23.470000  58.645000 24.270000  59.445000 ;
      RECT 23.470000  61.475000 24.270000  62.275000 ;
      RECT 23.470000  64.495000 24.270000  65.295000 ;
      RECT 23.470000  67.325000 24.270000  68.125000 ;
      RECT 23.470000  70.350000 24.270000  71.150000 ;
      RECT 23.470000  72.030000 24.270000  72.830000 ;
      RECT 23.470000  73.710000 24.270000  74.510000 ;
      RECT 23.470000  75.390000 24.270000  76.190000 ;
      RECT 23.470000  77.070000 24.270000  77.870000 ;
      RECT 23.470000  78.750000 24.270000  79.550000 ;
      RECT 23.470000  80.430000 24.270000  81.230000 ;
      RECT 23.470000  82.110000 24.270000  82.910000 ;
      RECT 23.470000  83.790000 24.270000  84.590000 ;
      RECT 23.470000  85.470000 24.270000  86.270000 ;
      RECT 23.470000  87.150000 24.270000  87.950000 ;
      RECT 23.470000  88.830000 24.270000  89.630000 ;
      RECT 23.470000  90.510000 24.270000  91.310000 ;
      RECT 23.470000  92.190000 24.270000  92.990000 ;
      RECT 23.470000  93.870000 24.270000  94.670000 ;
      RECT 23.470000 176.155000 24.270000 176.955000 ;
      RECT 23.470000 177.775000 24.270000 178.575000 ;
      RECT 23.470000 179.395000 24.270000 180.195000 ;
      RECT 23.470000 181.015000 24.270000 181.815000 ;
      RECT 23.470000 182.635000 24.270000 183.435000 ;
      RECT 23.470000 184.255000 24.270000 185.055000 ;
      RECT 23.470000 185.875000 24.270000 186.675000 ;
      RECT 23.470000 187.495000 24.270000 188.295000 ;
      RECT 23.470000 189.115000 24.270000 189.915000 ;
      RECT 23.470000 190.735000 24.270000 191.535000 ;
      RECT 23.470000 192.355000 24.270000 193.155000 ;
      RECT 23.470000 193.975000 24.270000 194.775000 ;
      RECT 23.470000 195.595000 24.270000 196.395000 ;
      RECT 23.470000 197.215000 24.270000 198.015000 ;
      RECT 23.470000 198.835000 24.270000 199.635000 ;
      RECT 23.475000   9.295000 24.275000  10.095000 ;
      RECT 23.475000  12.325000 24.275000  13.125000 ;
      RECT 25.070000  20.195000 25.870000  20.995000 ;
      RECT 25.070000  23.225000 25.870000  24.025000 ;
      RECT 25.070000  26.245000 25.870000  27.045000 ;
      RECT 25.070000  29.275000 25.870000  30.075000 ;
      RECT 25.075000   2.450000 25.875000   3.250000 ;
      RECT 25.075000   4.360000 25.875000   5.160000 ;
      RECT 25.075000   6.270000 25.875000   7.070000 ;
      RECT 25.075000  15.345000 25.875000  16.145000 ;
      RECT 25.075000  17.175000 25.875000  17.975000 ;
      RECT 25.075000  32.295000 25.875000  33.095000 ;
      RECT 25.075000  34.125000 25.875000  34.925000 ;
      RECT 25.075000  37.145000 25.875000  37.945000 ;
      RECT 25.075000  38.975000 25.875000  39.775000 ;
      RECT 25.075000  41.995000 25.875000  42.795000 ;
      RECT 25.075000  45.025000 25.875000  45.825000 ;
      RECT 25.075000  51.835000 25.875000  52.635000 ;
      RECT 25.075000  58.645000 25.875000  59.445000 ;
      RECT 25.075000  61.475000 25.875000  62.275000 ;
      RECT 25.075000  64.495000 25.875000  65.295000 ;
      RECT 25.075000  67.325000 25.875000  68.125000 ;
      RECT 25.075000  70.350000 25.875000  71.150000 ;
      RECT 25.075000  72.030000 25.875000  72.830000 ;
      RECT 25.075000  73.710000 25.875000  74.510000 ;
      RECT 25.075000  75.390000 25.875000  76.190000 ;
      RECT 25.075000  77.070000 25.875000  77.870000 ;
      RECT 25.075000  78.750000 25.875000  79.550000 ;
      RECT 25.075000  80.430000 25.875000  81.230000 ;
      RECT 25.075000  82.110000 25.875000  82.910000 ;
      RECT 25.075000  83.790000 25.875000  84.590000 ;
      RECT 25.075000  85.470000 25.875000  86.270000 ;
      RECT 25.075000  87.150000 25.875000  87.950000 ;
      RECT 25.075000  88.830000 25.875000  89.630000 ;
      RECT 25.075000  90.510000 25.875000  91.310000 ;
      RECT 25.075000  92.190000 25.875000  92.990000 ;
      RECT 25.075000  93.870000 25.875000  94.670000 ;
      RECT 25.075000 176.155000 25.875000 176.955000 ;
      RECT 25.075000 177.775000 25.875000 178.575000 ;
      RECT 25.075000 179.395000 25.875000 180.195000 ;
      RECT 25.075000 181.015000 25.875000 181.815000 ;
      RECT 25.075000 182.635000 25.875000 183.435000 ;
      RECT 25.075000 184.255000 25.875000 185.055000 ;
      RECT 25.075000 185.875000 25.875000 186.675000 ;
      RECT 25.075000 187.495000 25.875000 188.295000 ;
      RECT 25.075000 189.115000 25.875000 189.915000 ;
      RECT 25.075000 190.735000 25.875000 191.535000 ;
      RECT 25.075000 192.355000 25.875000 193.155000 ;
      RECT 25.075000 193.975000 25.875000 194.775000 ;
      RECT 25.075000 195.595000 25.875000 196.395000 ;
      RECT 25.075000 197.215000 25.875000 198.015000 ;
      RECT 25.075000 198.835000 25.875000 199.635000 ;
      RECT 25.080000   9.295000 25.880000  10.095000 ;
      RECT 25.080000  12.325000 25.880000  13.125000 ;
      RECT 26.675000  20.195000 27.475000  20.995000 ;
      RECT 26.675000  23.225000 27.475000  24.025000 ;
      RECT 26.675000  26.245000 27.475000  27.045000 ;
      RECT 26.675000  29.275000 27.475000  30.075000 ;
      RECT 26.680000   2.450000 27.480000   3.250000 ;
      RECT 26.680000   4.360000 27.480000   5.160000 ;
      RECT 26.680000   6.270000 27.480000   7.070000 ;
      RECT 26.680000  15.345000 27.480000  16.145000 ;
      RECT 26.680000  17.175000 27.480000  17.975000 ;
      RECT 26.680000  32.295000 27.480000  33.095000 ;
      RECT 26.680000  34.125000 27.480000  34.925000 ;
      RECT 26.680000  37.145000 27.480000  37.945000 ;
      RECT 26.680000  38.975000 27.480000  39.775000 ;
      RECT 26.680000  41.995000 27.480000  42.795000 ;
      RECT 26.680000  45.025000 27.480000  45.825000 ;
      RECT 26.680000  51.835000 27.480000  52.635000 ;
      RECT 26.680000  58.645000 27.480000  59.445000 ;
      RECT 26.680000  61.475000 27.480000  62.275000 ;
      RECT 26.680000  64.495000 27.480000  65.295000 ;
      RECT 26.680000  67.325000 27.480000  68.125000 ;
      RECT 26.680000  70.350000 27.480000  71.150000 ;
      RECT 26.680000  72.030000 27.480000  72.830000 ;
      RECT 26.680000  73.710000 27.480000  74.510000 ;
      RECT 26.680000  75.390000 27.480000  76.190000 ;
      RECT 26.680000  77.070000 27.480000  77.870000 ;
      RECT 26.680000  78.750000 27.480000  79.550000 ;
      RECT 26.680000  80.430000 27.480000  81.230000 ;
      RECT 26.680000  82.110000 27.480000  82.910000 ;
      RECT 26.680000  83.790000 27.480000  84.590000 ;
      RECT 26.680000  85.470000 27.480000  86.270000 ;
      RECT 26.680000  87.150000 27.480000  87.950000 ;
      RECT 26.680000  88.830000 27.480000  89.630000 ;
      RECT 26.680000  90.510000 27.480000  91.310000 ;
      RECT 26.680000  92.190000 27.480000  92.990000 ;
      RECT 26.680000  93.870000 27.480000  94.670000 ;
      RECT 26.680000 176.155000 27.480000 176.955000 ;
      RECT 26.680000 177.775000 27.480000 178.575000 ;
      RECT 26.680000 179.395000 27.480000 180.195000 ;
      RECT 26.680000 181.015000 27.480000 181.815000 ;
      RECT 26.680000 182.635000 27.480000 183.435000 ;
      RECT 26.680000 184.255000 27.480000 185.055000 ;
      RECT 26.680000 185.875000 27.480000 186.675000 ;
      RECT 26.680000 187.495000 27.480000 188.295000 ;
      RECT 26.680000 189.115000 27.480000 189.915000 ;
      RECT 26.680000 190.735000 27.480000 191.535000 ;
      RECT 26.680000 192.355000 27.480000 193.155000 ;
      RECT 26.680000 193.975000 27.480000 194.775000 ;
      RECT 26.680000 195.595000 27.480000 196.395000 ;
      RECT 26.680000 197.215000 27.480000 198.015000 ;
      RECT 26.680000 198.835000 27.480000 199.635000 ;
      RECT 26.685000   9.295000 27.485000  10.095000 ;
      RECT 26.685000  12.325000 27.485000  13.125000 ;
      RECT 28.280000  20.195000 29.080000  20.995000 ;
      RECT 28.280000  23.225000 29.080000  24.025000 ;
      RECT 28.280000  26.245000 29.080000  27.045000 ;
      RECT 28.280000  29.275000 29.080000  30.075000 ;
      RECT 28.285000   2.450000 29.085000   3.250000 ;
      RECT 28.285000   4.360000 29.085000   5.160000 ;
      RECT 28.285000   6.270000 29.085000   7.070000 ;
      RECT 28.285000  15.345000 29.085000  16.145000 ;
      RECT 28.285000  17.175000 29.085000  17.975000 ;
      RECT 28.285000  32.295000 29.085000  33.095000 ;
      RECT 28.285000  34.125000 29.085000  34.925000 ;
      RECT 28.285000  37.145000 29.085000  37.945000 ;
      RECT 28.285000  38.975000 29.085000  39.775000 ;
      RECT 28.285000  41.995000 29.085000  42.795000 ;
      RECT 28.285000  45.025000 29.085000  45.825000 ;
      RECT 28.285000  51.835000 29.085000  52.635000 ;
      RECT 28.285000  58.645000 29.085000  59.445000 ;
      RECT 28.285000  61.475000 29.085000  62.275000 ;
      RECT 28.285000  64.495000 29.085000  65.295000 ;
      RECT 28.285000  67.325000 29.085000  68.125000 ;
      RECT 28.285000  70.350000 29.085000  71.150000 ;
      RECT 28.285000  72.030000 29.085000  72.830000 ;
      RECT 28.285000  73.710000 29.085000  74.510000 ;
      RECT 28.285000  75.390000 29.085000  76.190000 ;
      RECT 28.285000  77.070000 29.085000  77.870000 ;
      RECT 28.285000  78.750000 29.085000  79.550000 ;
      RECT 28.285000  80.430000 29.085000  81.230000 ;
      RECT 28.285000  82.110000 29.085000  82.910000 ;
      RECT 28.285000  83.790000 29.085000  84.590000 ;
      RECT 28.285000  85.470000 29.085000  86.270000 ;
      RECT 28.285000  87.150000 29.085000  87.950000 ;
      RECT 28.285000  88.830000 29.085000  89.630000 ;
      RECT 28.285000  90.510000 29.085000  91.310000 ;
      RECT 28.285000  92.190000 29.085000  92.990000 ;
      RECT 28.285000  93.870000 29.085000  94.670000 ;
      RECT 28.285000 176.155000 29.085000 176.955000 ;
      RECT 28.285000 177.775000 29.085000 178.575000 ;
      RECT 28.285000 179.395000 29.085000 180.195000 ;
      RECT 28.285000 181.015000 29.085000 181.815000 ;
      RECT 28.285000 182.635000 29.085000 183.435000 ;
      RECT 28.285000 184.255000 29.085000 185.055000 ;
      RECT 28.285000 185.875000 29.085000 186.675000 ;
      RECT 28.285000 187.495000 29.085000 188.295000 ;
      RECT 28.285000 189.115000 29.085000 189.915000 ;
      RECT 28.285000 190.735000 29.085000 191.535000 ;
      RECT 28.285000 192.355000 29.085000 193.155000 ;
      RECT 28.285000 193.975000 29.085000 194.775000 ;
      RECT 28.285000 195.595000 29.085000 196.395000 ;
      RECT 28.285000 197.215000 29.085000 198.015000 ;
      RECT 28.285000 198.835000 29.085000 199.635000 ;
      RECT 28.290000   9.295000 29.090000  10.095000 ;
      RECT 28.290000  12.325000 29.090000  13.125000 ;
      RECT 29.885000  20.195000 30.685000  20.995000 ;
      RECT 29.885000  23.225000 30.685000  24.025000 ;
      RECT 29.885000  26.245000 30.685000  27.045000 ;
      RECT 29.885000  29.275000 30.685000  30.075000 ;
      RECT 29.890000   2.450000 30.690000   3.250000 ;
      RECT 29.890000   4.360000 30.690000   5.160000 ;
      RECT 29.890000   6.270000 30.690000   7.070000 ;
      RECT 29.890000  15.345000 30.690000  16.145000 ;
      RECT 29.890000  17.175000 30.690000  17.975000 ;
      RECT 29.890000  32.295000 30.690000  33.095000 ;
      RECT 29.890000  34.125000 30.690000  34.925000 ;
      RECT 29.890000  37.145000 30.690000  37.945000 ;
      RECT 29.890000  38.975000 30.690000  39.775000 ;
      RECT 29.890000  41.995000 30.690000  42.795000 ;
      RECT 29.890000  45.025000 30.690000  45.825000 ;
      RECT 29.890000  51.835000 30.690000  52.635000 ;
      RECT 29.890000  58.645000 30.690000  59.445000 ;
      RECT 29.890000  61.475000 30.690000  62.275000 ;
      RECT 29.890000  64.495000 30.690000  65.295000 ;
      RECT 29.890000  67.325000 30.690000  68.125000 ;
      RECT 29.890000  70.350000 30.690000  71.150000 ;
      RECT 29.890000  72.030000 30.690000  72.830000 ;
      RECT 29.890000  73.710000 30.690000  74.510000 ;
      RECT 29.890000  75.390000 30.690000  76.190000 ;
      RECT 29.890000  77.070000 30.690000  77.870000 ;
      RECT 29.890000  78.750000 30.690000  79.550000 ;
      RECT 29.890000  80.430000 30.690000  81.230000 ;
      RECT 29.890000  82.110000 30.690000  82.910000 ;
      RECT 29.890000  83.790000 30.690000  84.590000 ;
      RECT 29.890000  85.470000 30.690000  86.270000 ;
      RECT 29.890000  87.150000 30.690000  87.950000 ;
      RECT 29.890000  88.830000 30.690000  89.630000 ;
      RECT 29.890000  90.510000 30.690000  91.310000 ;
      RECT 29.890000  92.190000 30.690000  92.990000 ;
      RECT 29.890000  93.870000 30.690000  94.670000 ;
      RECT 29.890000 176.155000 30.690000 176.955000 ;
      RECT 29.890000 177.775000 30.690000 178.575000 ;
      RECT 29.890000 179.395000 30.690000 180.195000 ;
      RECT 29.890000 181.015000 30.690000 181.815000 ;
      RECT 29.890000 182.635000 30.690000 183.435000 ;
      RECT 29.890000 184.255000 30.690000 185.055000 ;
      RECT 29.890000 185.875000 30.690000 186.675000 ;
      RECT 29.890000 187.495000 30.690000 188.295000 ;
      RECT 29.890000 189.115000 30.690000 189.915000 ;
      RECT 29.890000 190.735000 30.690000 191.535000 ;
      RECT 29.890000 192.355000 30.690000 193.155000 ;
      RECT 29.890000 193.975000 30.690000 194.775000 ;
      RECT 29.890000 195.595000 30.690000 196.395000 ;
      RECT 29.890000 197.215000 30.690000 198.015000 ;
      RECT 29.890000 198.835000 30.690000 199.635000 ;
      RECT 29.895000   9.295000 30.695000  10.095000 ;
      RECT 29.895000  12.325000 30.695000  13.125000 ;
      RECT 31.490000  20.195000 32.290000  20.995000 ;
      RECT 31.490000  23.225000 32.290000  24.025000 ;
      RECT 31.490000  26.245000 32.290000  27.045000 ;
      RECT 31.490000  29.275000 32.290000  30.075000 ;
      RECT 31.495000   2.450000 32.295000   3.250000 ;
      RECT 31.495000   4.360000 32.295000   5.160000 ;
      RECT 31.495000   6.270000 32.295000   7.070000 ;
      RECT 31.495000  15.345000 32.295000  16.145000 ;
      RECT 31.495000  17.175000 32.295000  17.975000 ;
      RECT 31.495000  32.295000 32.295000  33.095000 ;
      RECT 31.495000  34.125000 32.295000  34.925000 ;
      RECT 31.495000  37.145000 32.295000  37.945000 ;
      RECT 31.495000  38.975000 32.295000  39.775000 ;
      RECT 31.495000  41.995000 32.295000  42.795000 ;
      RECT 31.495000  45.025000 32.295000  45.825000 ;
      RECT 31.495000  51.835000 32.295000  52.635000 ;
      RECT 31.495000  58.645000 32.295000  59.445000 ;
      RECT 31.495000  61.475000 32.295000  62.275000 ;
      RECT 31.495000  64.495000 32.295000  65.295000 ;
      RECT 31.495000  67.325000 32.295000  68.125000 ;
      RECT 31.495000  70.350000 32.295000  71.150000 ;
      RECT 31.495000  72.030000 32.295000  72.830000 ;
      RECT 31.495000  73.710000 32.295000  74.510000 ;
      RECT 31.495000  75.390000 32.295000  76.190000 ;
      RECT 31.495000  77.070000 32.295000  77.870000 ;
      RECT 31.495000  78.750000 32.295000  79.550000 ;
      RECT 31.495000  80.430000 32.295000  81.230000 ;
      RECT 31.495000  82.110000 32.295000  82.910000 ;
      RECT 31.495000  83.790000 32.295000  84.590000 ;
      RECT 31.495000  85.470000 32.295000  86.270000 ;
      RECT 31.495000  87.150000 32.295000  87.950000 ;
      RECT 31.495000  88.830000 32.295000  89.630000 ;
      RECT 31.495000  90.510000 32.295000  91.310000 ;
      RECT 31.495000  92.190000 32.295000  92.990000 ;
      RECT 31.495000  93.870000 32.295000  94.670000 ;
      RECT 31.495000 176.155000 32.295000 176.955000 ;
      RECT 31.495000 177.775000 32.295000 178.575000 ;
      RECT 31.495000 179.395000 32.295000 180.195000 ;
      RECT 31.495000 181.015000 32.295000 181.815000 ;
      RECT 31.495000 182.635000 32.295000 183.435000 ;
      RECT 31.495000 184.255000 32.295000 185.055000 ;
      RECT 31.495000 185.875000 32.295000 186.675000 ;
      RECT 31.495000 187.495000 32.295000 188.295000 ;
      RECT 31.495000 189.115000 32.295000 189.915000 ;
      RECT 31.495000 190.735000 32.295000 191.535000 ;
      RECT 31.495000 192.355000 32.295000 193.155000 ;
      RECT 31.495000 193.975000 32.295000 194.775000 ;
      RECT 31.495000 195.595000 32.295000 196.395000 ;
      RECT 31.495000 197.215000 32.295000 198.015000 ;
      RECT 31.495000 198.835000 32.295000 199.635000 ;
      RECT 31.500000   9.295000 32.300000  10.095000 ;
      RECT 31.500000  12.325000 32.300000  13.125000 ;
      RECT 33.095000  20.195000 33.895000  20.995000 ;
      RECT 33.095000  23.225000 33.895000  24.025000 ;
      RECT 33.095000  26.245000 33.895000  27.045000 ;
      RECT 33.095000  29.275000 33.895000  30.075000 ;
      RECT 33.100000   2.450000 33.900000   3.250000 ;
      RECT 33.100000   4.360000 33.900000   5.160000 ;
      RECT 33.100000   6.270000 33.900000   7.070000 ;
      RECT 33.100000  15.345000 33.900000  16.145000 ;
      RECT 33.100000  17.175000 33.900000  17.975000 ;
      RECT 33.100000  32.295000 33.900000  33.095000 ;
      RECT 33.100000  34.125000 33.900000  34.925000 ;
      RECT 33.100000  37.145000 33.900000  37.945000 ;
      RECT 33.100000  38.975000 33.900000  39.775000 ;
      RECT 33.100000  41.995000 33.900000  42.795000 ;
      RECT 33.100000  45.025000 33.900000  45.825000 ;
      RECT 33.100000  51.835000 33.900000  52.635000 ;
      RECT 33.100000  58.645000 33.900000  59.445000 ;
      RECT 33.100000  61.475000 33.900000  62.275000 ;
      RECT 33.100000  64.495000 33.900000  65.295000 ;
      RECT 33.100000  67.325000 33.900000  68.125000 ;
      RECT 33.100000  70.350000 33.900000  71.150000 ;
      RECT 33.100000  72.030000 33.900000  72.830000 ;
      RECT 33.100000  73.710000 33.900000  74.510000 ;
      RECT 33.100000  75.390000 33.900000  76.190000 ;
      RECT 33.100000  77.070000 33.900000  77.870000 ;
      RECT 33.100000  78.750000 33.900000  79.550000 ;
      RECT 33.100000  80.430000 33.900000  81.230000 ;
      RECT 33.100000  82.110000 33.900000  82.910000 ;
      RECT 33.100000  83.790000 33.900000  84.590000 ;
      RECT 33.100000  85.470000 33.900000  86.270000 ;
      RECT 33.100000  87.150000 33.900000  87.950000 ;
      RECT 33.100000  88.830000 33.900000  89.630000 ;
      RECT 33.100000  90.510000 33.900000  91.310000 ;
      RECT 33.100000  92.190000 33.900000  92.990000 ;
      RECT 33.100000  93.870000 33.900000  94.670000 ;
      RECT 33.100000 176.155000 33.900000 176.955000 ;
      RECT 33.100000 177.775000 33.900000 178.575000 ;
      RECT 33.100000 179.395000 33.900000 180.195000 ;
      RECT 33.100000 181.015000 33.900000 181.815000 ;
      RECT 33.100000 182.635000 33.900000 183.435000 ;
      RECT 33.100000 184.255000 33.900000 185.055000 ;
      RECT 33.100000 185.875000 33.900000 186.675000 ;
      RECT 33.100000 187.495000 33.900000 188.295000 ;
      RECT 33.100000 189.115000 33.900000 189.915000 ;
      RECT 33.100000 190.735000 33.900000 191.535000 ;
      RECT 33.100000 192.355000 33.900000 193.155000 ;
      RECT 33.100000 193.975000 33.900000 194.775000 ;
      RECT 33.100000 195.595000 33.900000 196.395000 ;
      RECT 33.100000 197.215000 33.900000 198.015000 ;
      RECT 33.100000 198.835000 33.900000 199.635000 ;
      RECT 33.105000   9.295000 33.905000  10.095000 ;
      RECT 33.105000  12.325000 33.905000  13.125000 ;
      RECT 34.700000  20.195000 35.500000  20.995000 ;
      RECT 34.700000  23.225000 35.500000  24.025000 ;
      RECT 34.700000  26.245000 35.500000  27.045000 ;
      RECT 34.700000  29.275000 35.500000  30.075000 ;
      RECT 34.705000   2.450000 35.505000   3.250000 ;
      RECT 34.705000   4.360000 35.505000   5.160000 ;
      RECT 34.705000   6.270000 35.505000   7.070000 ;
      RECT 34.705000  15.345000 35.505000  16.145000 ;
      RECT 34.705000  17.175000 35.505000  17.975000 ;
      RECT 34.705000  32.295000 35.505000  33.095000 ;
      RECT 34.705000  34.125000 35.505000  34.925000 ;
      RECT 34.705000  37.145000 35.505000  37.945000 ;
      RECT 34.705000  38.975000 35.505000  39.775000 ;
      RECT 34.705000  41.995000 35.505000  42.795000 ;
      RECT 34.705000  45.025000 35.505000  45.825000 ;
      RECT 34.705000  51.835000 35.505000  52.635000 ;
      RECT 34.705000  58.645000 35.505000  59.445000 ;
      RECT 34.705000  61.475000 35.505000  62.275000 ;
      RECT 34.705000  64.495000 35.505000  65.295000 ;
      RECT 34.705000  67.325000 35.505000  68.125000 ;
      RECT 34.705000  70.350000 35.505000  71.150000 ;
      RECT 34.705000  72.030000 35.505000  72.830000 ;
      RECT 34.705000  73.710000 35.505000  74.510000 ;
      RECT 34.705000  75.390000 35.505000  76.190000 ;
      RECT 34.705000  77.070000 35.505000  77.870000 ;
      RECT 34.705000  78.750000 35.505000  79.550000 ;
      RECT 34.705000  80.430000 35.505000  81.230000 ;
      RECT 34.705000  82.110000 35.505000  82.910000 ;
      RECT 34.705000  83.790000 35.505000  84.590000 ;
      RECT 34.705000  85.470000 35.505000  86.270000 ;
      RECT 34.705000  87.150000 35.505000  87.950000 ;
      RECT 34.705000  88.830000 35.505000  89.630000 ;
      RECT 34.705000  90.510000 35.505000  91.310000 ;
      RECT 34.705000  92.190000 35.505000  92.990000 ;
      RECT 34.705000  93.870000 35.505000  94.670000 ;
      RECT 34.705000 176.155000 35.505000 176.955000 ;
      RECT 34.705000 177.775000 35.505000 178.575000 ;
      RECT 34.705000 179.395000 35.505000 180.195000 ;
      RECT 34.705000 181.015000 35.505000 181.815000 ;
      RECT 34.705000 182.635000 35.505000 183.435000 ;
      RECT 34.705000 184.255000 35.505000 185.055000 ;
      RECT 34.705000 185.875000 35.505000 186.675000 ;
      RECT 34.705000 187.495000 35.505000 188.295000 ;
      RECT 34.705000 189.115000 35.505000 189.915000 ;
      RECT 34.705000 190.735000 35.505000 191.535000 ;
      RECT 34.705000 192.355000 35.505000 193.155000 ;
      RECT 34.705000 193.975000 35.505000 194.775000 ;
      RECT 34.705000 195.595000 35.505000 196.395000 ;
      RECT 34.705000 197.215000 35.505000 198.015000 ;
      RECT 34.705000 198.835000 35.505000 199.635000 ;
      RECT 34.710000   9.295000 35.510000  10.095000 ;
      RECT 34.710000  12.325000 35.510000  13.125000 ;
      RECT 36.305000  20.195000 37.105000  20.995000 ;
      RECT 36.305000  23.225000 37.105000  24.025000 ;
      RECT 36.305000  26.245000 37.105000  27.045000 ;
      RECT 36.305000  29.275000 37.105000  30.075000 ;
      RECT 36.310000   2.450000 37.110000   3.250000 ;
      RECT 36.310000   4.360000 37.110000   5.160000 ;
      RECT 36.310000   6.270000 37.110000   7.070000 ;
      RECT 36.310000  15.345000 37.110000  16.145000 ;
      RECT 36.310000  17.175000 37.110000  17.975000 ;
      RECT 36.310000  32.295000 37.110000  33.095000 ;
      RECT 36.310000  34.125000 37.110000  34.925000 ;
      RECT 36.310000  37.145000 37.110000  37.945000 ;
      RECT 36.310000  38.975000 37.110000  39.775000 ;
      RECT 36.310000  41.995000 37.110000  42.795000 ;
      RECT 36.310000  45.025000 37.110000  45.825000 ;
      RECT 36.310000  51.835000 37.110000  52.635000 ;
      RECT 36.310000  58.645000 37.110000  59.445000 ;
      RECT 36.310000  61.475000 37.110000  62.275000 ;
      RECT 36.310000  64.495000 37.110000  65.295000 ;
      RECT 36.310000  67.325000 37.110000  68.125000 ;
      RECT 36.310000  70.350000 37.110000  71.150000 ;
      RECT 36.310000  72.030000 37.110000  72.830000 ;
      RECT 36.310000  73.710000 37.110000  74.510000 ;
      RECT 36.310000  75.390000 37.110000  76.190000 ;
      RECT 36.310000  77.070000 37.110000  77.870000 ;
      RECT 36.310000  78.750000 37.110000  79.550000 ;
      RECT 36.310000  80.430000 37.110000  81.230000 ;
      RECT 36.310000  82.110000 37.110000  82.910000 ;
      RECT 36.310000  83.790000 37.110000  84.590000 ;
      RECT 36.310000  85.470000 37.110000  86.270000 ;
      RECT 36.310000  87.150000 37.110000  87.950000 ;
      RECT 36.310000  88.830000 37.110000  89.630000 ;
      RECT 36.310000  90.510000 37.110000  91.310000 ;
      RECT 36.310000  92.190000 37.110000  92.990000 ;
      RECT 36.310000  93.870000 37.110000  94.670000 ;
      RECT 36.310000 176.155000 37.110000 176.955000 ;
      RECT 36.310000 177.775000 37.110000 178.575000 ;
      RECT 36.310000 179.395000 37.110000 180.195000 ;
      RECT 36.310000 181.015000 37.110000 181.815000 ;
      RECT 36.310000 182.635000 37.110000 183.435000 ;
      RECT 36.310000 184.255000 37.110000 185.055000 ;
      RECT 36.310000 185.875000 37.110000 186.675000 ;
      RECT 36.310000 187.495000 37.110000 188.295000 ;
      RECT 36.310000 189.115000 37.110000 189.915000 ;
      RECT 36.310000 190.735000 37.110000 191.535000 ;
      RECT 36.310000 192.355000 37.110000 193.155000 ;
      RECT 36.310000 193.975000 37.110000 194.775000 ;
      RECT 36.310000 195.595000 37.110000 196.395000 ;
      RECT 36.310000 197.215000 37.110000 198.015000 ;
      RECT 36.310000 198.835000 37.110000 199.635000 ;
      RECT 36.315000   9.295000 37.115000  10.095000 ;
      RECT 36.315000  12.325000 37.115000  13.125000 ;
      RECT 37.910000  20.195000 38.710000  20.995000 ;
      RECT 37.910000  23.225000 38.710000  24.025000 ;
      RECT 37.910000  26.245000 38.710000  27.045000 ;
      RECT 37.910000  29.275000 38.710000  30.075000 ;
      RECT 37.915000   2.450000 38.715000   3.250000 ;
      RECT 37.915000   4.360000 38.715000   5.160000 ;
      RECT 37.915000   6.270000 38.715000   7.070000 ;
      RECT 37.915000  15.345000 38.715000  16.145000 ;
      RECT 37.915000  17.175000 38.715000  17.975000 ;
      RECT 37.915000  32.295000 38.715000  33.095000 ;
      RECT 37.915000  34.125000 38.715000  34.925000 ;
      RECT 37.915000  37.145000 38.715000  37.945000 ;
      RECT 37.915000  38.975000 38.715000  39.775000 ;
      RECT 37.915000  41.995000 38.715000  42.795000 ;
      RECT 37.915000  45.025000 38.715000  45.825000 ;
      RECT 37.915000  51.835000 38.715000  52.635000 ;
      RECT 37.915000  58.645000 38.715000  59.445000 ;
      RECT 37.915000  61.475000 38.715000  62.275000 ;
      RECT 37.915000  64.495000 38.715000  65.295000 ;
      RECT 37.915000  67.325000 38.715000  68.125000 ;
      RECT 37.915000  70.350000 38.715000  71.150000 ;
      RECT 37.915000  72.030000 38.715000  72.830000 ;
      RECT 37.915000  73.710000 38.715000  74.510000 ;
      RECT 37.915000  75.390000 38.715000  76.190000 ;
      RECT 37.915000  77.070000 38.715000  77.870000 ;
      RECT 37.915000  78.750000 38.715000  79.550000 ;
      RECT 37.915000  80.430000 38.715000  81.230000 ;
      RECT 37.915000  82.110000 38.715000  82.910000 ;
      RECT 37.915000  83.790000 38.715000  84.590000 ;
      RECT 37.915000  85.470000 38.715000  86.270000 ;
      RECT 37.915000  87.150000 38.715000  87.950000 ;
      RECT 37.915000  88.830000 38.715000  89.630000 ;
      RECT 37.915000  90.510000 38.715000  91.310000 ;
      RECT 37.915000  92.190000 38.715000  92.990000 ;
      RECT 37.915000  93.870000 38.715000  94.670000 ;
      RECT 37.915000 176.155000 38.715000 176.955000 ;
      RECT 37.915000 177.775000 38.715000 178.575000 ;
      RECT 37.915000 179.395000 38.715000 180.195000 ;
      RECT 37.915000 181.015000 38.715000 181.815000 ;
      RECT 37.915000 182.635000 38.715000 183.435000 ;
      RECT 37.915000 184.255000 38.715000 185.055000 ;
      RECT 37.915000 185.875000 38.715000 186.675000 ;
      RECT 37.915000 187.495000 38.715000 188.295000 ;
      RECT 37.915000 189.115000 38.715000 189.915000 ;
      RECT 37.915000 190.735000 38.715000 191.535000 ;
      RECT 37.915000 192.355000 38.715000 193.155000 ;
      RECT 37.915000 193.975000 38.715000 194.775000 ;
      RECT 37.915000 195.595000 38.715000 196.395000 ;
      RECT 37.915000 197.215000 38.715000 198.015000 ;
      RECT 37.915000 198.835000 38.715000 199.635000 ;
      RECT 37.920000   9.295000 38.720000  10.095000 ;
      RECT 37.920000  12.325000 38.720000  13.125000 ;
      RECT 39.515000  20.195000 40.315000  20.995000 ;
      RECT 39.515000  23.225000 40.315000  24.025000 ;
      RECT 39.515000  26.245000 40.315000  27.045000 ;
      RECT 39.515000  29.275000 40.315000  30.075000 ;
      RECT 39.520000   2.450000 40.320000   3.250000 ;
      RECT 39.520000   4.360000 40.320000   5.160000 ;
      RECT 39.520000   6.270000 40.320000   7.070000 ;
      RECT 39.520000  15.345000 40.320000  16.145000 ;
      RECT 39.520000  17.175000 40.320000  17.975000 ;
      RECT 39.520000  32.295000 40.320000  33.095000 ;
      RECT 39.520000  34.125000 40.320000  34.925000 ;
      RECT 39.520000  37.145000 40.320000  37.945000 ;
      RECT 39.520000  38.975000 40.320000  39.775000 ;
      RECT 39.520000  41.995000 40.320000  42.795000 ;
      RECT 39.520000  45.025000 40.320000  45.825000 ;
      RECT 39.520000  51.835000 40.320000  52.635000 ;
      RECT 39.520000  58.645000 40.320000  59.445000 ;
      RECT 39.520000  61.475000 40.320000  62.275000 ;
      RECT 39.520000  64.495000 40.320000  65.295000 ;
      RECT 39.520000  67.325000 40.320000  68.125000 ;
      RECT 39.520000  70.350000 40.320000  71.150000 ;
      RECT 39.520000  72.030000 40.320000  72.830000 ;
      RECT 39.520000  73.710000 40.320000  74.510000 ;
      RECT 39.520000  75.390000 40.320000  76.190000 ;
      RECT 39.520000  77.070000 40.320000  77.870000 ;
      RECT 39.520000  78.750000 40.320000  79.550000 ;
      RECT 39.520000  80.430000 40.320000  81.230000 ;
      RECT 39.520000  82.110000 40.320000  82.910000 ;
      RECT 39.520000  83.790000 40.320000  84.590000 ;
      RECT 39.520000  85.470000 40.320000  86.270000 ;
      RECT 39.520000  87.150000 40.320000  87.950000 ;
      RECT 39.520000  88.830000 40.320000  89.630000 ;
      RECT 39.520000  90.510000 40.320000  91.310000 ;
      RECT 39.520000  92.190000 40.320000  92.990000 ;
      RECT 39.520000  93.870000 40.320000  94.670000 ;
      RECT 39.520000 176.155000 40.320000 176.955000 ;
      RECT 39.520000 177.775000 40.320000 178.575000 ;
      RECT 39.520000 179.395000 40.320000 180.195000 ;
      RECT 39.520000 181.015000 40.320000 181.815000 ;
      RECT 39.520000 182.635000 40.320000 183.435000 ;
      RECT 39.520000 184.255000 40.320000 185.055000 ;
      RECT 39.520000 185.875000 40.320000 186.675000 ;
      RECT 39.520000 187.495000 40.320000 188.295000 ;
      RECT 39.520000 189.115000 40.320000 189.915000 ;
      RECT 39.520000 190.735000 40.320000 191.535000 ;
      RECT 39.520000 192.355000 40.320000 193.155000 ;
      RECT 39.520000 193.975000 40.320000 194.775000 ;
      RECT 39.520000 195.595000 40.320000 196.395000 ;
      RECT 39.520000 197.215000 40.320000 198.015000 ;
      RECT 39.520000 198.835000 40.320000 199.635000 ;
      RECT 39.525000   9.295000 40.325000  10.095000 ;
      RECT 39.525000  12.325000 40.325000  13.125000 ;
      RECT 41.120000  20.195000 41.920000  20.995000 ;
      RECT 41.120000  23.225000 41.920000  24.025000 ;
      RECT 41.120000  26.245000 41.920000  27.045000 ;
      RECT 41.120000  29.275000 41.920000  30.075000 ;
      RECT 41.125000   2.450000 41.925000   3.250000 ;
      RECT 41.125000   4.360000 41.925000   5.160000 ;
      RECT 41.125000   6.270000 41.925000   7.070000 ;
      RECT 41.125000  15.345000 41.925000  16.145000 ;
      RECT 41.125000  17.175000 41.925000  17.975000 ;
      RECT 41.125000  32.295000 41.925000  33.095000 ;
      RECT 41.125000  34.125000 41.925000  34.925000 ;
      RECT 41.125000  37.145000 41.925000  37.945000 ;
      RECT 41.125000  38.975000 41.925000  39.775000 ;
      RECT 41.125000  41.995000 41.925000  42.795000 ;
      RECT 41.125000  45.025000 41.925000  45.825000 ;
      RECT 41.125000  51.835000 41.925000  52.635000 ;
      RECT 41.125000  58.645000 41.925000  59.445000 ;
      RECT 41.125000  61.475000 41.925000  62.275000 ;
      RECT 41.125000  64.495000 41.925000  65.295000 ;
      RECT 41.125000  67.325000 41.925000  68.125000 ;
      RECT 41.125000  70.350000 41.925000  71.150000 ;
      RECT 41.125000  72.030000 41.925000  72.830000 ;
      RECT 41.125000  73.710000 41.925000  74.510000 ;
      RECT 41.125000  75.390000 41.925000  76.190000 ;
      RECT 41.125000  77.070000 41.925000  77.870000 ;
      RECT 41.125000  78.750000 41.925000  79.550000 ;
      RECT 41.125000  80.430000 41.925000  81.230000 ;
      RECT 41.125000  82.110000 41.925000  82.910000 ;
      RECT 41.125000  83.790000 41.925000  84.590000 ;
      RECT 41.125000  85.470000 41.925000  86.270000 ;
      RECT 41.125000  87.150000 41.925000  87.950000 ;
      RECT 41.125000  88.830000 41.925000  89.630000 ;
      RECT 41.125000  90.510000 41.925000  91.310000 ;
      RECT 41.125000  92.190000 41.925000  92.990000 ;
      RECT 41.125000  93.870000 41.925000  94.670000 ;
      RECT 41.125000 176.155000 41.925000 176.955000 ;
      RECT 41.125000 177.775000 41.925000 178.575000 ;
      RECT 41.125000 179.395000 41.925000 180.195000 ;
      RECT 41.125000 181.015000 41.925000 181.815000 ;
      RECT 41.125000 182.635000 41.925000 183.435000 ;
      RECT 41.125000 184.255000 41.925000 185.055000 ;
      RECT 41.125000 185.875000 41.925000 186.675000 ;
      RECT 41.125000 187.495000 41.925000 188.295000 ;
      RECT 41.125000 189.115000 41.925000 189.915000 ;
      RECT 41.125000 190.735000 41.925000 191.535000 ;
      RECT 41.125000 192.355000 41.925000 193.155000 ;
      RECT 41.125000 193.975000 41.925000 194.775000 ;
      RECT 41.125000 195.595000 41.925000 196.395000 ;
      RECT 41.125000 197.215000 41.925000 198.015000 ;
      RECT 41.125000 198.835000 41.925000 199.635000 ;
      RECT 41.130000   9.295000 41.930000  10.095000 ;
      RECT 41.130000  12.325000 41.930000  13.125000 ;
      RECT 42.725000  20.195000 43.525000  20.995000 ;
      RECT 42.725000  23.225000 43.525000  24.025000 ;
      RECT 42.725000  26.245000 43.525000  27.045000 ;
      RECT 42.725000  29.275000 43.525000  30.075000 ;
      RECT 42.730000   2.450000 43.530000   3.250000 ;
      RECT 42.730000   4.360000 43.530000   5.160000 ;
      RECT 42.730000   6.270000 43.530000   7.070000 ;
      RECT 42.730000  15.345000 43.530000  16.145000 ;
      RECT 42.730000  17.175000 43.530000  17.975000 ;
      RECT 42.730000  32.295000 43.530000  33.095000 ;
      RECT 42.730000  34.125000 43.530000  34.925000 ;
      RECT 42.730000  37.145000 43.530000  37.945000 ;
      RECT 42.730000  38.975000 43.530000  39.775000 ;
      RECT 42.730000  41.995000 43.530000  42.795000 ;
      RECT 42.730000  45.025000 43.530000  45.825000 ;
      RECT 42.730000  51.835000 43.530000  52.635000 ;
      RECT 42.730000  58.645000 43.530000  59.445000 ;
      RECT 42.730000  61.475000 43.530000  62.275000 ;
      RECT 42.730000  64.495000 43.530000  65.295000 ;
      RECT 42.730000  67.325000 43.530000  68.125000 ;
      RECT 42.730000  70.350000 43.530000  71.150000 ;
      RECT 42.730000  72.030000 43.530000  72.830000 ;
      RECT 42.730000  73.710000 43.530000  74.510000 ;
      RECT 42.730000  75.390000 43.530000  76.190000 ;
      RECT 42.730000  77.070000 43.530000  77.870000 ;
      RECT 42.730000  78.750000 43.530000  79.550000 ;
      RECT 42.730000  80.430000 43.530000  81.230000 ;
      RECT 42.730000  82.110000 43.530000  82.910000 ;
      RECT 42.730000  83.790000 43.530000  84.590000 ;
      RECT 42.730000  85.470000 43.530000  86.270000 ;
      RECT 42.730000  87.150000 43.530000  87.950000 ;
      RECT 42.730000  88.830000 43.530000  89.630000 ;
      RECT 42.730000  90.510000 43.530000  91.310000 ;
      RECT 42.730000  92.190000 43.530000  92.990000 ;
      RECT 42.730000  93.870000 43.530000  94.670000 ;
      RECT 42.730000 176.155000 43.530000 176.955000 ;
      RECT 42.730000 177.775000 43.530000 178.575000 ;
      RECT 42.730000 179.395000 43.530000 180.195000 ;
      RECT 42.730000 181.015000 43.530000 181.815000 ;
      RECT 42.730000 182.635000 43.530000 183.435000 ;
      RECT 42.730000 184.255000 43.530000 185.055000 ;
      RECT 42.730000 185.875000 43.530000 186.675000 ;
      RECT 42.730000 187.495000 43.530000 188.295000 ;
      RECT 42.730000 189.115000 43.530000 189.915000 ;
      RECT 42.730000 190.735000 43.530000 191.535000 ;
      RECT 42.730000 192.355000 43.530000 193.155000 ;
      RECT 42.730000 193.975000 43.530000 194.775000 ;
      RECT 42.730000 195.595000 43.530000 196.395000 ;
      RECT 42.730000 197.215000 43.530000 198.015000 ;
      RECT 42.730000 198.835000 43.530000 199.635000 ;
      RECT 42.735000   9.295000 43.535000  10.095000 ;
      RECT 42.735000  12.325000 43.535000  13.125000 ;
      RECT 44.330000  20.195000 45.130000  20.995000 ;
      RECT 44.330000  23.225000 45.130000  24.025000 ;
      RECT 44.330000  26.245000 45.130000  27.045000 ;
      RECT 44.330000  29.275000 45.130000  30.075000 ;
      RECT 44.335000   2.450000 45.135000   3.250000 ;
      RECT 44.335000   4.360000 45.135000   5.160000 ;
      RECT 44.335000   6.270000 45.135000   7.070000 ;
      RECT 44.335000  15.345000 45.135000  16.145000 ;
      RECT 44.335000  17.175000 45.135000  17.975000 ;
      RECT 44.335000  32.295000 45.135000  33.095000 ;
      RECT 44.335000  34.125000 45.135000  34.925000 ;
      RECT 44.335000  37.145000 45.135000  37.945000 ;
      RECT 44.335000  38.975000 45.135000  39.775000 ;
      RECT 44.335000  41.995000 45.135000  42.795000 ;
      RECT 44.335000  45.025000 45.135000  45.825000 ;
      RECT 44.335000  51.835000 45.135000  52.635000 ;
      RECT 44.335000  58.645000 45.135000  59.445000 ;
      RECT 44.335000  61.475000 45.135000  62.275000 ;
      RECT 44.335000  64.495000 45.135000  65.295000 ;
      RECT 44.335000  67.325000 45.135000  68.125000 ;
      RECT 44.335000  70.350000 45.135000  71.150000 ;
      RECT 44.335000  72.030000 45.135000  72.830000 ;
      RECT 44.335000  73.710000 45.135000  74.510000 ;
      RECT 44.335000  75.390000 45.135000  76.190000 ;
      RECT 44.335000  77.070000 45.135000  77.870000 ;
      RECT 44.335000  78.750000 45.135000  79.550000 ;
      RECT 44.335000  80.430000 45.135000  81.230000 ;
      RECT 44.335000  82.110000 45.135000  82.910000 ;
      RECT 44.335000  83.790000 45.135000  84.590000 ;
      RECT 44.335000  85.470000 45.135000  86.270000 ;
      RECT 44.335000  87.150000 45.135000  87.950000 ;
      RECT 44.335000  88.830000 45.135000  89.630000 ;
      RECT 44.335000  90.510000 45.135000  91.310000 ;
      RECT 44.335000  92.190000 45.135000  92.990000 ;
      RECT 44.335000  93.870000 45.135000  94.670000 ;
      RECT 44.335000 176.155000 45.135000 176.955000 ;
      RECT 44.335000 177.775000 45.135000 178.575000 ;
      RECT 44.335000 179.395000 45.135000 180.195000 ;
      RECT 44.335000 181.015000 45.135000 181.815000 ;
      RECT 44.335000 182.635000 45.135000 183.435000 ;
      RECT 44.335000 184.255000 45.135000 185.055000 ;
      RECT 44.335000 185.875000 45.135000 186.675000 ;
      RECT 44.335000 187.495000 45.135000 188.295000 ;
      RECT 44.335000 189.115000 45.135000 189.915000 ;
      RECT 44.335000 190.735000 45.135000 191.535000 ;
      RECT 44.335000 192.355000 45.135000 193.155000 ;
      RECT 44.335000 193.975000 45.135000 194.775000 ;
      RECT 44.335000 195.595000 45.135000 196.395000 ;
      RECT 44.335000 197.215000 45.135000 198.015000 ;
      RECT 44.335000 198.835000 45.135000 199.635000 ;
      RECT 44.340000   9.295000 45.140000  10.095000 ;
      RECT 44.340000  12.325000 45.140000  13.125000 ;
      RECT 45.935000  20.195000 46.735000  20.995000 ;
      RECT 45.935000  23.225000 46.735000  24.025000 ;
      RECT 45.935000  26.245000 46.735000  27.045000 ;
      RECT 45.935000  29.275000 46.735000  30.075000 ;
      RECT 45.940000   2.450000 46.740000   3.250000 ;
      RECT 45.940000   4.360000 46.740000   5.160000 ;
      RECT 45.940000   6.270000 46.740000   7.070000 ;
      RECT 45.940000  15.345000 46.740000  16.145000 ;
      RECT 45.940000  17.175000 46.740000  17.975000 ;
      RECT 45.940000  32.295000 46.740000  33.095000 ;
      RECT 45.940000  34.125000 46.740000  34.925000 ;
      RECT 45.940000  37.145000 46.740000  37.945000 ;
      RECT 45.940000  38.975000 46.740000  39.775000 ;
      RECT 45.940000  41.995000 46.740000  42.795000 ;
      RECT 45.940000  45.025000 46.740000  45.825000 ;
      RECT 45.940000  51.835000 46.740000  52.635000 ;
      RECT 45.940000  58.645000 46.740000  59.445000 ;
      RECT 45.940000  61.475000 46.740000  62.275000 ;
      RECT 45.940000  64.495000 46.740000  65.295000 ;
      RECT 45.940000  67.325000 46.740000  68.125000 ;
      RECT 45.940000  70.350000 46.740000  71.150000 ;
      RECT 45.940000  72.030000 46.740000  72.830000 ;
      RECT 45.940000  73.710000 46.740000  74.510000 ;
      RECT 45.940000  75.390000 46.740000  76.190000 ;
      RECT 45.940000  77.070000 46.740000  77.870000 ;
      RECT 45.940000  78.750000 46.740000  79.550000 ;
      RECT 45.940000  80.430000 46.740000  81.230000 ;
      RECT 45.940000  82.110000 46.740000  82.910000 ;
      RECT 45.940000  83.790000 46.740000  84.590000 ;
      RECT 45.940000  85.470000 46.740000  86.270000 ;
      RECT 45.940000  87.150000 46.740000  87.950000 ;
      RECT 45.940000  88.830000 46.740000  89.630000 ;
      RECT 45.940000  90.510000 46.740000  91.310000 ;
      RECT 45.940000  92.190000 46.740000  92.990000 ;
      RECT 45.940000  93.870000 46.740000  94.670000 ;
      RECT 45.940000 176.155000 46.740000 176.955000 ;
      RECT 45.940000 177.775000 46.740000 178.575000 ;
      RECT 45.940000 179.395000 46.740000 180.195000 ;
      RECT 45.940000 181.015000 46.740000 181.815000 ;
      RECT 45.940000 182.635000 46.740000 183.435000 ;
      RECT 45.940000 184.255000 46.740000 185.055000 ;
      RECT 45.940000 185.875000 46.740000 186.675000 ;
      RECT 45.940000 187.495000 46.740000 188.295000 ;
      RECT 45.940000 189.115000 46.740000 189.915000 ;
      RECT 45.940000 190.735000 46.740000 191.535000 ;
      RECT 45.940000 192.355000 46.740000 193.155000 ;
      RECT 45.940000 193.975000 46.740000 194.775000 ;
      RECT 45.940000 195.595000 46.740000 196.395000 ;
      RECT 45.940000 197.215000 46.740000 198.015000 ;
      RECT 45.940000 198.835000 46.740000 199.635000 ;
      RECT 45.945000   9.295000 46.745000  10.095000 ;
      RECT 45.945000  12.325000 46.745000  13.125000 ;
      RECT 47.540000  20.195000 48.340000  20.995000 ;
      RECT 47.540000  23.225000 48.340000  24.025000 ;
      RECT 47.540000  26.245000 48.340000  27.045000 ;
      RECT 47.540000  29.275000 48.340000  30.075000 ;
      RECT 47.545000   2.450000 48.345000   3.250000 ;
      RECT 47.545000   4.360000 48.345000   5.160000 ;
      RECT 47.545000   6.270000 48.345000   7.070000 ;
      RECT 47.545000  15.345000 48.345000  16.145000 ;
      RECT 47.545000  17.175000 48.345000  17.975000 ;
      RECT 47.545000  32.295000 48.345000  33.095000 ;
      RECT 47.545000  34.125000 48.345000  34.925000 ;
      RECT 47.545000  37.145000 48.345000  37.945000 ;
      RECT 47.545000  38.975000 48.345000  39.775000 ;
      RECT 47.545000  41.995000 48.345000  42.795000 ;
      RECT 47.545000  45.025000 48.345000  45.825000 ;
      RECT 47.545000  51.835000 48.345000  52.635000 ;
      RECT 47.545000  58.645000 48.345000  59.445000 ;
      RECT 47.545000  61.475000 48.345000  62.275000 ;
      RECT 47.545000  64.495000 48.345000  65.295000 ;
      RECT 47.545000  67.325000 48.345000  68.125000 ;
      RECT 47.545000  70.350000 48.345000  71.150000 ;
      RECT 47.545000  72.030000 48.345000  72.830000 ;
      RECT 47.545000  73.710000 48.345000  74.510000 ;
      RECT 47.545000  75.390000 48.345000  76.190000 ;
      RECT 47.545000  77.070000 48.345000  77.870000 ;
      RECT 47.545000  78.750000 48.345000  79.550000 ;
      RECT 47.545000  80.430000 48.345000  81.230000 ;
      RECT 47.545000  82.110000 48.345000  82.910000 ;
      RECT 47.545000  83.790000 48.345000  84.590000 ;
      RECT 47.545000  85.470000 48.345000  86.270000 ;
      RECT 47.545000  87.150000 48.345000  87.950000 ;
      RECT 47.545000  88.830000 48.345000  89.630000 ;
      RECT 47.545000  90.510000 48.345000  91.310000 ;
      RECT 47.545000  92.190000 48.345000  92.990000 ;
      RECT 47.545000  93.870000 48.345000  94.670000 ;
      RECT 47.545000 176.155000 48.345000 176.955000 ;
      RECT 47.545000 177.775000 48.345000 178.575000 ;
      RECT 47.545000 179.395000 48.345000 180.195000 ;
      RECT 47.545000 181.015000 48.345000 181.815000 ;
      RECT 47.545000 182.635000 48.345000 183.435000 ;
      RECT 47.545000 184.255000 48.345000 185.055000 ;
      RECT 47.545000 185.875000 48.345000 186.675000 ;
      RECT 47.545000 187.495000 48.345000 188.295000 ;
      RECT 47.545000 189.115000 48.345000 189.915000 ;
      RECT 47.545000 190.735000 48.345000 191.535000 ;
      RECT 47.545000 192.355000 48.345000 193.155000 ;
      RECT 47.545000 193.975000 48.345000 194.775000 ;
      RECT 47.545000 195.595000 48.345000 196.395000 ;
      RECT 47.545000 197.215000 48.345000 198.015000 ;
      RECT 47.545000 198.835000 48.345000 199.635000 ;
      RECT 47.550000   9.295000 48.350000  10.095000 ;
      RECT 47.550000  12.325000 48.350000  13.125000 ;
      RECT 49.145000  20.195000 49.945000  20.995000 ;
      RECT 49.145000  23.225000 49.945000  24.025000 ;
      RECT 49.145000  26.245000 49.945000  27.045000 ;
      RECT 49.145000  29.275000 49.945000  30.075000 ;
      RECT 49.150000   2.450000 49.950000   3.250000 ;
      RECT 49.150000   4.360000 49.950000   5.160000 ;
      RECT 49.150000   6.270000 49.950000   7.070000 ;
      RECT 49.150000  15.345000 49.950000  16.145000 ;
      RECT 49.150000  17.175000 49.950000  17.975000 ;
      RECT 49.150000  32.295000 49.950000  33.095000 ;
      RECT 49.150000  34.125000 49.950000  34.925000 ;
      RECT 49.150000  37.145000 49.950000  37.945000 ;
      RECT 49.150000  38.975000 49.950000  39.775000 ;
      RECT 49.150000  41.995000 49.950000  42.795000 ;
      RECT 49.150000  45.025000 49.950000  45.825000 ;
      RECT 49.150000  51.835000 49.950000  52.635000 ;
      RECT 49.150000  58.645000 49.950000  59.445000 ;
      RECT 49.150000  61.475000 49.950000  62.275000 ;
      RECT 49.150000  64.495000 49.950000  65.295000 ;
      RECT 49.150000  67.325000 49.950000  68.125000 ;
      RECT 49.150000  70.350000 49.950000  71.150000 ;
      RECT 49.150000  72.030000 49.950000  72.830000 ;
      RECT 49.150000  73.710000 49.950000  74.510000 ;
      RECT 49.150000  75.390000 49.950000  76.190000 ;
      RECT 49.150000  77.070000 49.950000  77.870000 ;
      RECT 49.150000  78.750000 49.950000  79.550000 ;
      RECT 49.150000  80.430000 49.950000  81.230000 ;
      RECT 49.150000  82.110000 49.950000  82.910000 ;
      RECT 49.150000  83.790000 49.950000  84.590000 ;
      RECT 49.150000  85.470000 49.950000  86.270000 ;
      RECT 49.150000  87.150000 49.950000  87.950000 ;
      RECT 49.150000  88.830000 49.950000  89.630000 ;
      RECT 49.150000  90.510000 49.950000  91.310000 ;
      RECT 49.150000  92.190000 49.950000  92.990000 ;
      RECT 49.150000  93.870000 49.950000  94.670000 ;
      RECT 49.150000 176.155000 49.950000 176.955000 ;
      RECT 49.150000 177.775000 49.950000 178.575000 ;
      RECT 49.150000 179.395000 49.950000 180.195000 ;
      RECT 49.150000 181.015000 49.950000 181.815000 ;
      RECT 49.150000 182.635000 49.950000 183.435000 ;
      RECT 49.150000 184.255000 49.950000 185.055000 ;
      RECT 49.150000 185.875000 49.950000 186.675000 ;
      RECT 49.150000 187.495000 49.950000 188.295000 ;
      RECT 49.150000 189.115000 49.950000 189.915000 ;
      RECT 49.150000 190.735000 49.950000 191.535000 ;
      RECT 49.150000 192.355000 49.950000 193.155000 ;
      RECT 49.150000 193.975000 49.950000 194.775000 ;
      RECT 49.150000 195.595000 49.950000 196.395000 ;
      RECT 49.150000 197.215000 49.950000 198.015000 ;
      RECT 49.150000 198.835000 49.950000 199.635000 ;
      RECT 49.155000   9.295000 49.955000  10.095000 ;
      RECT 49.155000  12.325000 49.955000  13.125000 ;
      RECT 50.750000  20.195000 51.550000  20.995000 ;
      RECT 50.750000  23.225000 51.550000  24.025000 ;
      RECT 50.750000  26.245000 51.550000  27.045000 ;
      RECT 50.750000  29.275000 51.550000  30.075000 ;
      RECT 50.755000   2.450000 51.555000   3.250000 ;
      RECT 50.755000   4.360000 51.555000   5.160000 ;
      RECT 50.755000   6.270000 51.555000   7.070000 ;
      RECT 50.755000  15.345000 51.555000  16.145000 ;
      RECT 50.755000  17.175000 51.555000  17.975000 ;
      RECT 50.755000  32.295000 51.555000  33.095000 ;
      RECT 50.755000  34.125000 51.555000  34.925000 ;
      RECT 50.755000  37.145000 51.555000  37.945000 ;
      RECT 50.755000  38.975000 51.555000  39.775000 ;
      RECT 50.755000  41.995000 51.555000  42.795000 ;
      RECT 50.755000  45.025000 51.555000  45.825000 ;
      RECT 50.755000  51.835000 51.555000  52.635000 ;
      RECT 50.755000  58.645000 51.555000  59.445000 ;
      RECT 50.755000  61.475000 51.555000  62.275000 ;
      RECT 50.755000  64.495000 51.555000  65.295000 ;
      RECT 50.755000  67.325000 51.555000  68.125000 ;
      RECT 50.755000  70.350000 51.555000  71.150000 ;
      RECT 50.755000  72.030000 51.555000  72.830000 ;
      RECT 50.755000  73.710000 51.555000  74.510000 ;
      RECT 50.755000  75.390000 51.555000  76.190000 ;
      RECT 50.755000  77.070000 51.555000  77.870000 ;
      RECT 50.755000  78.750000 51.555000  79.550000 ;
      RECT 50.755000  80.430000 51.555000  81.230000 ;
      RECT 50.755000  82.110000 51.555000  82.910000 ;
      RECT 50.755000  83.790000 51.555000  84.590000 ;
      RECT 50.755000  85.470000 51.555000  86.270000 ;
      RECT 50.755000  87.150000 51.555000  87.950000 ;
      RECT 50.755000  88.830000 51.555000  89.630000 ;
      RECT 50.755000  90.510000 51.555000  91.310000 ;
      RECT 50.755000  92.190000 51.555000  92.990000 ;
      RECT 50.755000  93.870000 51.555000  94.670000 ;
      RECT 50.755000 176.155000 51.555000 176.955000 ;
      RECT 50.755000 177.775000 51.555000 178.575000 ;
      RECT 50.755000 179.395000 51.555000 180.195000 ;
      RECT 50.755000 181.015000 51.555000 181.815000 ;
      RECT 50.755000 182.635000 51.555000 183.435000 ;
      RECT 50.755000 184.255000 51.555000 185.055000 ;
      RECT 50.755000 185.875000 51.555000 186.675000 ;
      RECT 50.755000 187.495000 51.555000 188.295000 ;
      RECT 50.755000 189.115000 51.555000 189.915000 ;
      RECT 50.755000 190.735000 51.555000 191.535000 ;
      RECT 50.755000 192.355000 51.555000 193.155000 ;
      RECT 50.755000 193.975000 51.555000 194.775000 ;
      RECT 50.755000 195.595000 51.555000 196.395000 ;
      RECT 50.755000 197.215000 51.555000 198.015000 ;
      RECT 50.755000 198.835000 51.555000 199.635000 ;
      RECT 50.760000   9.295000 51.560000  10.095000 ;
      RECT 50.760000  12.325000 51.560000  13.125000 ;
      RECT 52.355000  20.195000 53.155000  20.995000 ;
      RECT 52.355000  23.225000 53.155000  24.025000 ;
      RECT 52.355000  26.245000 53.155000  27.045000 ;
      RECT 52.355000  29.275000 53.155000  30.075000 ;
      RECT 52.360000   2.450000 53.160000   3.250000 ;
      RECT 52.360000   4.360000 53.160000   5.160000 ;
      RECT 52.360000   6.270000 53.160000   7.070000 ;
      RECT 52.360000  15.345000 53.160000  16.145000 ;
      RECT 52.360000  17.175000 53.160000  17.975000 ;
      RECT 52.360000  32.295000 53.160000  33.095000 ;
      RECT 52.360000  34.125000 53.160000  34.925000 ;
      RECT 52.360000  37.145000 53.160000  37.945000 ;
      RECT 52.360000  38.975000 53.160000  39.775000 ;
      RECT 52.360000  41.995000 53.160000  42.795000 ;
      RECT 52.360000  45.025000 53.160000  45.825000 ;
      RECT 52.360000  51.835000 53.160000  52.635000 ;
      RECT 52.360000  58.645000 53.160000  59.445000 ;
      RECT 52.360000  61.475000 53.160000  62.275000 ;
      RECT 52.360000  64.495000 53.160000  65.295000 ;
      RECT 52.360000  67.325000 53.160000  68.125000 ;
      RECT 52.360000  70.350000 53.160000  71.150000 ;
      RECT 52.360000  72.030000 53.160000  72.830000 ;
      RECT 52.360000  73.710000 53.160000  74.510000 ;
      RECT 52.360000  75.390000 53.160000  76.190000 ;
      RECT 52.360000  77.070000 53.160000  77.870000 ;
      RECT 52.360000  78.750000 53.160000  79.550000 ;
      RECT 52.360000  80.430000 53.160000  81.230000 ;
      RECT 52.360000  82.110000 53.160000  82.910000 ;
      RECT 52.360000  83.790000 53.160000  84.590000 ;
      RECT 52.360000  85.470000 53.160000  86.270000 ;
      RECT 52.360000  87.150000 53.160000  87.950000 ;
      RECT 52.360000  88.830000 53.160000  89.630000 ;
      RECT 52.360000  90.510000 53.160000  91.310000 ;
      RECT 52.360000  92.190000 53.160000  92.990000 ;
      RECT 52.360000  93.870000 53.160000  94.670000 ;
      RECT 52.360000 176.155000 53.160000 176.955000 ;
      RECT 52.360000 177.775000 53.160000 178.575000 ;
      RECT 52.360000 179.395000 53.160000 180.195000 ;
      RECT 52.360000 181.015000 53.160000 181.815000 ;
      RECT 52.360000 182.635000 53.160000 183.435000 ;
      RECT 52.360000 184.255000 53.160000 185.055000 ;
      RECT 52.360000 185.875000 53.160000 186.675000 ;
      RECT 52.360000 187.495000 53.160000 188.295000 ;
      RECT 52.360000 189.115000 53.160000 189.915000 ;
      RECT 52.360000 190.735000 53.160000 191.535000 ;
      RECT 52.360000 192.355000 53.160000 193.155000 ;
      RECT 52.360000 193.975000 53.160000 194.775000 ;
      RECT 52.360000 195.595000 53.160000 196.395000 ;
      RECT 52.360000 197.215000 53.160000 198.015000 ;
      RECT 52.360000 198.835000 53.160000 199.635000 ;
      RECT 52.365000   9.295000 53.165000  10.095000 ;
      RECT 52.365000  12.325000 53.165000  13.125000 ;
      RECT 53.960000  20.195000 54.760000  20.995000 ;
      RECT 53.960000  23.225000 54.760000  24.025000 ;
      RECT 53.960000  26.245000 54.760000  27.045000 ;
      RECT 53.960000  29.275000 54.760000  30.075000 ;
      RECT 53.965000   2.450000 54.765000   3.250000 ;
      RECT 53.965000   4.360000 54.765000   5.160000 ;
      RECT 53.965000   6.270000 54.765000   7.070000 ;
      RECT 53.965000  15.345000 54.765000  16.145000 ;
      RECT 53.965000  17.175000 54.765000  17.975000 ;
      RECT 53.965000  32.295000 54.765000  33.095000 ;
      RECT 53.965000  34.125000 54.765000  34.925000 ;
      RECT 53.965000  37.145000 54.765000  37.945000 ;
      RECT 53.965000  38.975000 54.765000  39.775000 ;
      RECT 53.965000  41.995000 54.765000  42.795000 ;
      RECT 53.965000  45.025000 54.765000  45.825000 ;
      RECT 53.965000  51.835000 54.765000  52.635000 ;
      RECT 53.965000  58.645000 54.765000  59.445000 ;
      RECT 53.965000  61.475000 54.765000  62.275000 ;
      RECT 53.965000  64.495000 54.765000  65.295000 ;
      RECT 53.965000  67.325000 54.765000  68.125000 ;
      RECT 53.965000  70.350000 54.765000  71.150000 ;
      RECT 53.965000  72.030000 54.765000  72.830000 ;
      RECT 53.965000  73.710000 54.765000  74.510000 ;
      RECT 53.965000  75.390000 54.765000  76.190000 ;
      RECT 53.965000  77.070000 54.765000  77.870000 ;
      RECT 53.965000  78.750000 54.765000  79.550000 ;
      RECT 53.965000  80.430000 54.765000  81.230000 ;
      RECT 53.965000  82.110000 54.765000  82.910000 ;
      RECT 53.965000  83.790000 54.765000  84.590000 ;
      RECT 53.965000  85.470000 54.765000  86.270000 ;
      RECT 53.965000  87.150000 54.765000  87.950000 ;
      RECT 53.965000  88.830000 54.765000  89.630000 ;
      RECT 53.965000  90.510000 54.765000  91.310000 ;
      RECT 53.965000  92.190000 54.765000  92.990000 ;
      RECT 53.965000  93.870000 54.765000  94.670000 ;
      RECT 53.965000 176.155000 54.765000 176.955000 ;
      RECT 53.965000 177.775000 54.765000 178.575000 ;
      RECT 53.965000 179.395000 54.765000 180.195000 ;
      RECT 53.965000 181.015000 54.765000 181.815000 ;
      RECT 53.965000 182.635000 54.765000 183.435000 ;
      RECT 53.965000 184.255000 54.765000 185.055000 ;
      RECT 53.965000 185.875000 54.765000 186.675000 ;
      RECT 53.965000 187.495000 54.765000 188.295000 ;
      RECT 53.965000 189.115000 54.765000 189.915000 ;
      RECT 53.965000 190.735000 54.765000 191.535000 ;
      RECT 53.965000 192.355000 54.765000 193.155000 ;
      RECT 53.965000 193.975000 54.765000 194.775000 ;
      RECT 53.965000 195.595000 54.765000 196.395000 ;
      RECT 53.965000 197.215000 54.765000 198.015000 ;
      RECT 53.965000 198.835000 54.765000 199.635000 ;
      RECT 53.970000   9.295000 54.770000  10.095000 ;
      RECT 53.970000  12.325000 54.770000  13.125000 ;
      RECT 55.565000  20.195000 56.365000  20.995000 ;
      RECT 55.565000  23.225000 56.365000  24.025000 ;
      RECT 55.565000  26.245000 56.365000  27.045000 ;
      RECT 55.565000  29.275000 56.365000  30.075000 ;
      RECT 55.570000   2.450000 56.370000   3.250000 ;
      RECT 55.570000   4.360000 56.370000   5.160000 ;
      RECT 55.570000   6.270000 56.370000   7.070000 ;
      RECT 55.570000  15.345000 56.370000  16.145000 ;
      RECT 55.570000  17.175000 56.370000  17.975000 ;
      RECT 55.570000  32.295000 56.370000  33.095000 ;
      RECT 55.570000  34.125000 56.370000  34.925000 ;
      RECT 55.570000  37.145000 56.370000  37.945000 ;
      RECT 55.570000  38.975000 56.370000  39.775000 ;
      RECT 55.570000  41.995000 56.370000  42.795000 ;
      RECT 55.570000  45.025000 56.370000  45.825000 ;
      RECT 55.570000  51.835000 56.370000  52.635000 ;
      RECT 55.570000  58.645000 56.370000  59.445000 ;
      RECT 55.570000  61.475000 56.370000  62.275000 ;
      RECT 55.570000  64.495000 56.370000  65.295000 ;
      RECT 55.570000  67.325000 56.370000  68.125000 ;
      RECT 55.570000  70.350000 56.370000  71.150000 ;
      RECT 55.570000  72.030000 56.370000  72.830000 ;
      RECT 55.570000  73.710000 56.370000  74.510000 ;
      RECT 55.570000  75.390000 56.370000  76.190000 ;
      RECT 55.570000  77.070000 56.370000  77.870000 ;
      RECT 55.570000  78.750000 56.370000  79.550000 ;
      RECT 55.570000  80.430000 56.370000  81.230000 ;
      RECT 55.570000  82.110000 56.370000  82.910000 ;
      RECT 55.570000  83.790000 56.370000  84.590000 ;
      RECT 55.570000  85.470000 56.370000  86.270000 ;
      RECT 55.570000  87.150000 56.370000  87.950000 ;
      RECT 55.570000  88.830000 56.370000  89.630000 ;
      RECT 55.570000  90.510000 56.370000  91.310000 ;
      RECT 55.570000  92.190000 56.370000  92.990000 ;
      RECT 55.570000  93.870000 56.370000  94.670000 ;
      RECT 55.570000 176.155000 56.370000 176.955000 ;
      RECT 55.570000 177.775000 56.370000 178.575000 ;
      RECT 55.570000 179.395000 56.370000 180.195000 ;
      RECT 55.570000 181.015000 56.370000 181.815000 ;
      RECT 55.570000 182.635000 56.370000 183.435000 ;
      RECT 55.570000 184.255000 56.370000 185.055000 ;
      RECT 55.570000 185.875000 56.370000 186.675000 ;
      RECT 55.570000 187.495000 56.370000 188.295000 ;
      RECT 55.570000 189.115000 56.370000 189.915000 ;
      RECT 55.570000 190.735000 56.370000 191.535000 ;
      RECT 55.570000 192.355000 56.370000 193.155000 ;
      RECT 55.570000 193.975000 56.370000 194.775000 ;
      RECT 55.570000 195.595000 56.370000 196.395000 ;
      RECT 55.570000 197.215000 56.370000 198.015000 ;
      RECT 55.570000 198.835000 56.370000 199.635000 ;
      RECT 55.575000   9.295000 56.375000  10.095000 ;
      RECT 55.575000  12.325000 56.375000  13.125000 ;
      RECT 57.170000  20.195000 57.970000  20.995000 ;
      RECT 57.170000  23.225000 57.970000  24.025000 ;
      RECT 57.170000  26.245000 57.970000  27.045000 ;
      RECT 57.170000  29.275000 57.970000  30.075000 ;
      RECT 57.175000   2.450000 57.975000   3.250000 ;
      RECT 57.175000   4.360000 57.975000   5.160000 ;
      RECT 57.175000   6.270000 57.975000   7.070000 ;
      RECT 57.175000   9.295000 57.975000  10.095000 ;
      RECT 57.175000  12.325000 57.975000  13.125000 ;
      RECT 57.175000  15.345000 57.975000  16.145000 ;
      RECT 57.175000  17.175000 57.975000  17.975000 ;
      RECT 57.175000  32.295000 57.975000  33.095000 ;
      RECT 57.175000  34.125000 57.975000  34.925000 ;
      RECT 57.175000  37.145000 57.975000  37.945000 ;
      RECT 57.175000  38.975000 57.975000  39.775000 ;
      RECT 57.175000  41.995000 57.975000  42.795000 ;
      RECT 57.175000  45.025000 57.975000  45.825000 ;
      RECT 57.175000  51.835000 57.975000  52.635000 ;
      RECT 57.175000  58.645000 57.975000  59.445000 ;
      RECT 57.175000  61.475000 57.975000  62.275000 ;
      RECT 57.175000  64.495000 57.975000  65.295000 ;
      RECT 57.175000  67.325000 57.975000  68.125000 ;
      RECT 57.175000  70.350000 57.975000  71.150000 ;
      RECT 57.175000  72.030000 57.975000  72.830000 ;
      RECT 57.175000  73.710000 57.975000  74.510000 ;
      RECT 57.175000  75.390000 57.975000  76.190000 ;
      RECT 57.175000  77.070000 57.975000  77.870000 ;
      RECT 57.175000  78.750000 57.975000  79.550000 ;
      RECT 57.175000  80.430000 57.975000  81.230000 ;
      RECT 57.175000  82.110000 57.975000  82.910000 ;
      RECT 57.175000  83.790000 57.975000  84.590000 ;
      RECT 57.175000  85.470000 57.975000  86.270000 ;
      RECT 57.175000  87.150000 57.975000  87.950000 ;
      RECT 57.175000  88.830000 57.975000  89.630000 ;
      RECT 57.175000  90.510000 57.975000  91.310000 ;
      RECT 57.175000  92.190000 57.975000  92.990000 ;
      RECT 57.175000  93.870000 57.975000  94.670000 ;
      RECT 57.175000 176.155000 57.975000 176.955000 ;
      RECT 57.175000 177.775000 57.975000 178.575000 ;
      RECT 57.175000 179.395000 57.975000 180.195000 ;
      RECT 57.175000 181.015000 57.975000 181.815000 ;
      RECT 57.175000 182.635000 57.975000 183.435000 ;
      RECT 57.175000 184.255000 57.975000 185.055000 ;
      RECT 57.175000 185.875000 57.975000 186.675000 ;
      RECT 57.175000 187.495000 57.975000 188.295000 ;
      RECT 57.175000 189.115000 57.975000 189.915000 ;
      RECT 57.175000 190.735000 57.975000 191.535000 ;
      RECT 57.175000 192.355000 57.975000 193.155000 ;
      RECT 57.175000 193.975000 57.975000 194.775000 ;
      RECT 57.175000 195.595000 57.975000 196.395000 ;
      RECT 57.175000 197.215000 57.975000 198.015000 ;
      RECT 57.175000 198.835000 57.975000 199.635000 ;
      RECT 58.775000   9.295000 59.575000  10.095000 ;
      RECT 58.775000  12.325000 59.575000  13.125000 ;
      RECT 58.775000  20.195000 59.575000  20.995000 ;
      RECT 58.775000  23.225000 59.575000  24.025000 ;
      RECT 58.775000  26.245000 59.575000  27.045000 ;
      RECT 58.775000  29.275000 59.575000  30.075000 ;
      RECT 58.775000  41.995000 59.575000  42.795000 ;
      RECT 58.775000  45.025000 59.575000  45.825000 ;
      RECT 58.780000   2.450000 59.580000   3.250000 ;
      RECT 58.780000   4.360000 59.580000   5.160000 ;
      RECT 58.780000   6.270000 59.580000   7.070000 ;
      RECT 58.780000  15.345000 59.580000  16.145000 ;
      RECT 58.780000  17.175000 59.580000  17.975000 ;
      RECT 58.780000  32.295000 59.580000  33.095000 ;
      RECT 58.780000  34.125000 59.580000  34.925000 ;
      RECT 58.780000  37.145000 59.580000  37.945000 ;
      RECT 58.780000  38.975000 59.580000  39.775000 ;
      RECT 58.780000  51.835000 59.580000  52.635000 ;
      RECT 58.780000  58.645000 59.580000  59.445000 ;
      RECT 58.780000  61.475000 59.580000  62.275000 ;
      RECT 58.780000  64.495000 59.580000  65.295000 ;
      RECT 58.780000  67.325000 59.580000  68.125000 ;
      RECT 58.780000  70.350000 59.580000  71.150000 ;
      RECT 58.780000  72.030000 59.580000  72.830000 ;
      RECT 58.780000  73.710000 59.580000  74.510000 ;
      RECT 58.780000  75.390000 59.580000  76.190000 ;
      RECT 58.780000  77.070000 59.580000  77.870000 ;
      RECT 58.780000  78.750000 59.580000  79.550000 ;
      RECT 58.780000  80.430000 59.580000  81.230000 ;
      RECT 58.780000  82.110000 59.580000  82.910000 ;
      RECT 58.780000  83.790000 59.580000  84.590000 ;
      RECT 58.780000  85.470000 59.580000  86.270000 ;
      RECT 58.780000  87.150000 59.580000  87.950000 ;
      RECT 58.780000  88.830000 59.580000  89.630000 ;
      RECT 58.780000  90.510000 59.580000  91.310000 ;
      RECT 58.780000  92.190000 59.580000  92.990000 ;
      RECT 58.780000  93.870000 59.580000  94.670000 ;
      RECT 58.780000 176.155000 59.580000 176.955000 ;
      RECT 58.780000 177.775000 59.580000 178.575000 ;
      RECT 58.780000 179.395000 59.580000 180.195000 ;
      RECT 58.780000 181.015000 59.580000 181.815000 ;
      RECT 58.780000 182.635000 59.580000 183.435000 ;
      RECT 58.780000 184.255000 59.580000 185.055000 ;
      RECT 58.780000 185.875000 59.580000 186.675000 ;
      RECT 58.780000 187.495000 59.580000 188.295000 ;
      RECT 58.780000 189.115000 59.580000 189.915000 ;
      RECT 58.780000 190.735000 59.580000 191.535000 ;
      RECT 58.780000 192.355000 59.580000 193.155000 ;
      RECT 58.780000 193.975000 59.580000 194.775000 ;
      RECT 58.780000 195.595000 59.580000 196.395000 ;
      RECT 58.780000 197.215000 59.580000 198.015000 ;
      RECT 58.780000 198.835000 59.580000 199.635000 ;
      RECT 60.375000   9.295000 61.175000  10.095000 ;
      RECT 60.375000  12.325000 61.175000  13.125000 ;
      RECT 60.375000  20.195000 61.175000  20.995000 ;
      RECT 60.375000  23.225000 61.175000  24.025000 ;
      RECT 60.375000  41.995000 61.175000  42.795000 ;
      RECT 60.375000  45.025000 61.175000  45.825000 ;
      RECT 60.380000   2.450000 61.180000   3.250000 ;
      RECT 60.380000   4.360000 61.180000   5.160000 ;
      RECT 60.380000   6.270000 61.180000   7.070000 ;
      RECT 60.380000  15.345000 61.180000  16.145000 ;
      RECT 60.380000  17.175000 61.180000  17.975000 ;
      RECT 60.380000  26.245000 61.180000  27.045000 ;
      RECT 60.380000  29.275000 61.180000  30.075000 ;
      RECT 60.380000  32.295000 61.180000  33.095000 ;
      RECT 60.380000  34.125000 61.180000  34.925000 ;
      RECT 60.380000  51.835000 61.180000  52.635000 ;
      RECT 60.380000  64.495000 61.180000  65.295000 ;
      RECT 60.380000  67.325000 61.180000  68.125000 ;
      RECT 60.380000  70.350000 61.180000  71.150000 ;
      RECT 60.380000  72.030000 61.180000  72.830000 ;
      RECT 60.380000  73.710000 61.180000  74.510000 ;
      RECT 60.380000  75.390000 61.180000  76.190000 ;
      RECT 60.380000  77.070000 61.180000  77.870000 ;
      RECT 60.380000  78.750000 61.180000  79.550000 ;
      RECT 60.380000  80.430000 61.180000  81.230000 ;
      RECT 60.380000  82.110000 61.180000  82.910000 ;
      RECT 60.380000  83.790000 61.180000  84.590000 ;
      RECT 60.380000  85.470000 61.180000  86.270000 ;
      RECT 60.380000  87.150000 61.180000  87.950000 ;
      RECT 60.380000  88.830000 61.180000  89.630000 ;
      RECT 60.380000  90.510000 61.180000  91.310000 ;
      RECT 60.380000  92.190000 61.180000  92.990000 ;
      RECT 60.380000  93.870000 61.180000  94.670000 ;
      RECT 60.380000 176.155000 61.180000 176.955000 ;
      RECT 60.380000 177.775000 61.180000 178.575000 ;
      RECT 60.380000 179.395000 61.180000 180.195000 ;
      RECT 60.380000 181.015000 61.180000 181.815000 ;
      RECT 60.380000 182.635000 61.180000 183.435000 ;
      RECT 60.380000 184.255000 61.180000 185.055000 ;
      RECT 60.380000 185.875000 61.180000 186.675000 ;
      RECT 60.380000 187.495000 61.180000 188.295000 ;
      RECT 60.380000 189.115000 61.180000 189.915000 ;
      RECT 60.380000 190.735000 61.180000 191.535000 ;
      RECT 60.380000 192.355000 61.180000 193.155000 ;
      RECT 60.380000 193.975000 61.180000 194.775000 ;
      RECT 60.380000 195.595000 61.180000 196.395000 ;
      RECT 60.380000 197.215000 61.180000 198.015000 ;
      RECT 60.380000 198.835000 61.180000 199.635000 ;
      RECT 60.385000  37.145000 61.185000  37.945000 ;
      RECT 60.385000  38.975000 61.185000  39.775000 ;
      RECT 60.385000  58.645000 61.185000  59.445000 ;
      RECT 60.385000  61.475000 61.185000  62.275000 ;
      RECT 61.975000   9.295000 62.775000  10.095000 ;
      RECT 61.975000  12.325000 62.775000  13.125000 ;
      RECT 61.975000  20.195000 62.775000  20.995000 ;
      RECT 61.975000  23.225000 62.775000  24.025000 ;
      RECT 61.975000  41.995000 62.775000  42.795000 ;
      RECT 61.975000  45.025000 62.775000  45.825000 ;
      RECT 61.980000   2.450000 62.780000   3.250000 ;
      RECT 61.980000   4.360000 62.780000   5.160000 ;
      RECT 61.980000   6.270000 62.780000   7.070000 ;
      RECT 61.980000  15.345000 62.780000  16.145000 ;
      RECT 61.980000  17.175000 62.780000  17.975000 ;
      RECT 61.980000  26.245000 62.780000  27.045000 ;
      RECT 61.980000  29.275000 62.780000  30.075000 ;
      RECT 61.980000  32.295000 62.780000  33.095000 ;
      RECT 61.980000  34.125000 62.780000  34.925000 ;
      RECT 61.980000  51.835000 62.780000  52.635000 ;
      RECT 61.980000  64.495000 62.780000  65.295000 ;
      RECT 61.980000  67.325000 62.780000  68.125000 ;
      RECT 61.980000  70.350000 62.780000  71.150000 ;
      RECT 61.980000  72.030000 62.780000  72.830000 ;
      RECT 61.980000  73.710000 62.780000  74.510000 ;
      RECT 61.980000  75.390000 62.780000  76.190000 ;
      RECT 61.980000  77.070000 62.780000  77.870000 ;
      RECT 61.980000  78.750000 62.780000  79.550000 ;
      RECT 61.980000  80.430000 62.780000  81.230000 ;
      RECT 61.980000  82.110000 62.780000  82.910000 ;
      RECT 61.980000  83.790000 62.780000  84.590000 ;
      RECT 61.980000  85.470000 62.780000  86.270000 ;
      RECT 61.980000  87.150000 62.780000  87.950000 ;
      RECT 61.980000  88.830000 62.780000  89.630000 ;
      RECT 61.980000  90.510000 62.780000  91.310000 ;
      RECT 61.980000  92.190000 62.780000  92.990000 ;
      RECT 61.980000  93.870000 62.780000  94.670000 ;
      RECT 61.980000 176.155000 62.780000 176.955000 ;
      RECT 61.980000 177.775000 62.780000 178.575000 ;
      RECT 61.980000 179.395000 62.780000 180.195000 ;
      RECT 61.980000 181.015000 62.780000 181.815000 ;
      RECT 61.980000 182.635000 62.780000 183.435000 ;
      RECT 61.980000 184.255000 62.780000 185.055000 ;
      RECT 61.980000 185.875000 62.780000 186.675000 ;
      RECT 61.980000 187.495000 62.780000 188.295000 ;
      RECT 61.980000 189.115000 62.780000 189.915000 ;
      RECT 61.980000 190.735000 62.780000 191.535000 ;
      RECT 61.980000 192.355000 62.780000 193.155000 ;
      RECT 61.980000 193.975000 62.780000 194.775000 ;
      RECT 61.980000 195.595000 62.780000 196.395000 ;
      RECT 61.980000 197.215000 62.780000 198.015000 ;
      RECT 61.980000 198.835000 62.780000 199.635000 ;
      RECT 61.985000  37.145000 62.785000  37.945000 ;
      RECT 61.985000  38.975000 62.785000  39.775000 ;
      RECT 61.985000  58.645000 62.785000  59.445000 ;
      RECT 61.985000  61.475000 62.785000  62.275000 ;
      RECT 63.575000   9.295000 64.375000  10.095000 ;
      RECT 63.575000  12.325000 64.375000  13.125000 ;
      RECT 63.575000  20.195000 64.375000  20.995000 ;
      RECT 63.575000  23.225000 64.375000  24.025000 ;
      RECT 63.575000  41.995000 64.375000  42.795000 ;
      RECT 63.575000  45.025000 64.375000  45.825000 ;
      RECT 63.580000   2.450000 64.380000   3.250000 ;
      RECT 63.580000   4.360000 64.380000   5.160000 ;
      RECT 63.580000   6.270000 64.380000   7.070000 ;
      RECT 63.580000  15.345000 64.380000  16.145000 ;
      RECT 63.580000  17.175000 64.380000  17.975000 ;
      RECT 63.580000  26.245000 64.380000  27.045000 ;
      RECT 63.580000  29.275000 64.380000  30.075000 ;
      RECT 63.580000  32.295000 64.380000  33.095000 ;
      RECT 63.580000  34.125000 64.380000  34.925000 ;
      RECT 63.580000  51.835000 64.380000  52.635000 ;
      RECT 63.580000  64.495000 64.380000  65.295000 ;
      RECT 63.580000  67.325000 64.380000  68.125000 ;
      RECT 63.580000  70.350000 64.380000  71.150000 ;
      RECT 63.580000  72.030000 64.380000  72.830000 ;
      RECT 63.580000  73.710000 64.380000  74.510000 ;
      RECT 63.580000  75.390000 64.380000  76.190000 ;
      RECT 63.580000  77.070000 64.380000  77.870000 ;
      RECT 63.580000  78.750000 64.380000  79.550000 ;
      RECT 63.580000  80.430000 64.380000  81.230000 ;
      RECT 63.580000  82.110000 64.380000  82.910000 ;
      RECT 63.580000  83.790000 64.380000  84.590000 ;
      RECT 63.580000  85.470000 64.380000  86.270000 ;
      RECT 63.580000  87.150000 64.380000  87.950000 ;
      RECT 63.580000  88.830000 64.380000  89.630000 ;
      RECT 63.580000  90.510000 64.380000  91.310000 ;
      RECT 63.580000  92.190000 64.380000  92.990000 ;
      RECT 63.580000  93.870000 64.380000  94.670000 ;
      RECT 63.580000 176.155000 64.380000 176.955000 ;
      RECT 63.580000 177.775000 64.380000 178.575000 ;
      RECT 63.580000 179.395000 64.380000 180.195000 ;
      RECT 63.580000 181.015000 64.380000 181.815000 ;
      RECT 63.580000 182.635000 64.380000 183.435000 ;
      RECT 63.580000 184.255000 64.380000 185.055000 ;
      RECT 63.580000 185.875000 64.380000 186.675000 ;
      RECT 63.580000 187.495000 64.380000 188.295000 ;
      RECT 63.580000 189.115000 64.380000 189.915000 ;
      RECT 63.580000 190.735000 64.380000 191.535000 ;
      RECT 63.580000 192.355000 64.380000 193.155000 ;
      RECT 63.580000 193.975000 64.380000 194.775000 ;
      RECT 63.580000 195.595000 64.380000 196.395000 ;
      RECT 63.580000 197.215000 64.380000 198.015000 ;
      RECT 63.580000 198.835000 64.380000 199.635000 ;
      RECT 63.585000  37.145000 64.385000  37.945000 ;
      RECT 63.585000  38.975000 64.385000  39.775000 ;
      RECT 63.585000  58.645000 64.385000  59.445000 ;
      RECT 63.585000  61.475000 64.385000  62.275000 ;
      RECT 65.175000   9.295000 65.975000  10.095000 ;
      RECT 65.175000  12.325000 65.975000  13.125000 ;
      RECT 65.175000  20.195000 65.975000  20.995000 ;
      RECT 65.175000  23.225000 65.975000  24.025000 ;
      RECT 65.175000  41.995000 65.975000  42.795000 ;
      RECT 65.175000  45.025000 65.975000  45.825000 ;
      RECT 65.180000   2.450000 65.980000   3.250000 ;
      RECT 65.180000   4.360000 65.980000   5.160000 ;
      RECT 65.180000   6.270000 65.980000   7.070000 ;
      RECT 65.180000  15.345000 65.980000  16.145000 ;
      RECT 65.180000  17.175000 65.980000  17.975000 ;
      RECT 65.180000  26.245000 65.980000  27.045000 ;
      RECT 65.180000  29.275000 65.980000  30.075000 ;
      RECT 65.180000  32.295000 65.980000  33.095000 ;
      RECT 65.180000  34.125000 65.980000  34.925000 ;
      RECT 65.180000  51.835000 65.980000  52.635000 ;
      RECT 65.180000  64.495000 65.980000  65.295000 ;
      RECT 65.180000  67.325000 65.980000  68.125000 ;
      RECT 65.180000  70.350000 65.980000  71.150000 ;
      RECT 65.180000  72.030000 65.980000  72.830000 ;
      RECT 65.180000  73.710000 65.980000  74.510000 ;
      RECT 65.180000  75.390000 65.980000  76.190000 ;
      RECT 65.180000  77.070000 65.980000  77.870000 ;
      RECT 65.180000  78.750000 65.980000  79.550000 ;
      RECT 65.180000  80.430000 65.980000  81.230000 ;
      RECT 65.180000  82.110000 65.980000  82.910000 ;
      RECT 65.180000  83.790000 65.980000  84.590000 ;
      RECT 65.180000  85.470000 65.980000  86.270000 ;
      RECT 65.180000  87.150000 65.980000  87.950000 ;
      RECT 65.180000  88.830000 65.980000  89.630000 ;
      RECT 65.180000  90.510000 65.980000  91.310000 ;
      RECT 65.180000  92.190000 65.980000  92.990000 ;
      RECT 65.180000  93.870000 65.980000  94.670000 ;
      RECT 65.180000 176.155000 65.980000 176.955000 ;
      RECT 65.180000 177.775000 65.980000 178.575000 ;
      RECT 65.180000 179.395000 65.980000 180.195000 ;
      RECT 65.180000 181.015000 65.980000 181.815000 ;
      RECT 65.180000 182.635000 65.980000 183.435000 ;
      RECT 65.180000 184.255000 65.980000 185.055000 ;
      RECT 65.180000 185.875000 65.980000 186.675000 ;
      RECT 65.180000 187.495000 65.980000 188.295000 ;
      RECT 65.180000 189.115000 65.980000 189.915000 ;
      RECT 65.180000 190.735000 65.980000 191.535000 ;
      RECT 65.180000 192.355000 65.980000 193.155000 ;
      RECT 65.180000 193.975000 65.980000 194.775000 ;
      RECT 65.180000 195.595000 65.980000 196.395000 ;
      RECT 65.180000 197.215000 65.980000 198.015000 ;
      RECT 65.180000 198.835000 65.980000 199.635000 ;
      RECT 65.185000  37.145000 65.985000  37.945000 ;
      RECT 65.185000  38.975000 65.985000  39.775000 ;
      RECT 65.185000  58.645000 65.985000  59.445000 ;
      RECT 65.185000  61.475000 65.985000  62.275000 ;
      RECT 66.775000   9.295000 67.575000  10.095000 ;
      RECT 66.775000  12.325000 67.575000  13.125000 ;
      RECT 66.775000  20.195000 67.575000  20.995000 ;
      RECT 66.775000  23.225000 67.575000  24.025000 ;
      RECT 66.775000  41.995000 67.575000  42.795000 ;
      RECT 66.775000  45.025000 67.575000  45.825000 ;
      RECT 66.780000   2.450000 67.580000   3.250000 ;
      RECT 66.780000   4.360000 67.580000   5.160000 ;
      RECT 66.780000   6.270000 67.580000   7.070000 ;
      RECT 66.780000  15.345000 67.580000  16.145000 ;
      RECT 66.780000  17.175000 67.580000  17.975000 ;
      RECT 66.780000  26.245000 67.580000  27.045000 ;
      RECT 66.780000  29.275000 67.580000  30.075000 ;
      RECT 66.780000  32.295000 67.580000  33.095000 ;
      RECT 66.780000  34.125000 67.580000  34.925000 ;
      RECT 66.780000  51.835000 67.580000  52.635000 ;
      RECT 66.780000  64.495000 67.580000  65.295000 ;
      RECT 66.780000  67.325000 67.580000  68.125000 ;
      RECT 66.780000  70.350000 67.580000  71.150000 ;
      RECT 66.780000  72.030000 67.580000  72.830000 ;
      RECT 66.780000  73.710000 67.580000  74.510000 ;
      RECT 66.780000  75.390000 67.580000  76.190000 ;
      RECT 66.780000  77.070000 67.580000  77.870000 ;
      RECT 66.780000  78.750000 67.580000  79.550000 ;
      RECT 66.780000  80.430000 67.580000  81.230000 ;
      RECT 66.780000  82.110000 67.580000  82.910000 ;
      RECT 66.780000  83.790000 67.580000  84.590000 ;
      RECT 66.780000  85.470000 67.580000  86.270000 ;
      RECT 66.780000  87.150000 67.580000  87.950000 ;
      RECT 66.780000  88.830000 67.580000  89.630000 ;
      RECT 66.780000  90.510000 67.580000  91.310000 ;
      RECT 66.780000  92.190000 67.580000  92.990000 ;
      RECT 66.780000  93.870000 67.580000  94.670000 ;
      RECT 66.780000 176.155000 67.580000 176.955000 ;
      RECT 66.780000 177.775000 67.580000 178.575000 ;
      RECT 66.780000 179.395000 67.580000 180.195000 ;
      RECT 66.780000 181.015000 67.580000 181.815000 ;
      RECT 66.780000 182.635000 67.580000 183.435000 ;
      RECT 66.780000 184.255000 67.580000 185.055000 ;
      RECT 66.780000 185.875000 67.580000 186.675000 ;
      RECT 66.780000 187.495000 67.580000 188.295000 ;
      RECT 66.780000 189.115000 67.580000 189.915000 ;
      RECT 66.780000 190.735000 67.580000 191.535000 ;
      RECT 66.780000 192.355000 67.580000 193.155000 ;
      RECT 66.780000 193.975000 67.580000 194.775000 ;
      RECT 66.780000 195.595000 67.580000 196.395000 ;
      RECT 66.780000 197.215000 67.580000 198.015000 ;
      RECT 66.780000 198.835000 67.580000 199.635000 ;
      RECT 66.785000  37.145000 67.585000  37.945000 ;
      RECT 66.785000  38.975000 67.585000  39.775000 ;
      RECT 66.785000  58.645000 67.585000  59.445000 ;
      RECT 66.785000  61.475000 67.585000  62.275000 ;
      RECT 68.375000   9.295000 69.175000  10.095000 ;
      RECT 68.375000  12.325000 69.175000  13.125000 ;
      RECT 68.375000  20.195000 69.175000  20.995000 ;
      RECT 68.375000  23.225000 69.175000  24.025000 ;
      RECT 68.375000  41.995000 69.175000  42.795000 ;
      RECT 68.375000  45.025000 69.175000  45.825000 ;
      RECT 68.380000   2.450000 69.180000   3.250000 ;
      RECT 68.380000   4.360000 69.180000   5.160000 ;
      RECT 68.380000   6.270000 69.180000   7.070000 ;
      RECT 68.380000  15.345000 69.180000  16.145000 ;
      RECT 68.380000  17.175000 69.180000  17.975000 ;
      RECT 68.380000  26.245000 69.180000  27.045000 ;
      RECT 68.380000  29.275000 69.180000  30.075000 ;
      RECT 68.380000  32.295000 69.180000  33.095000 ;
      RECT 68.380000  34.125000 69.180000  34.925000 ;
      RECT 68.380000  51.835000 69.180000  52.635000 ;
      RECT 68.380000  64.495000 69.180000  65.295000 ;
      RECT 68.380000  67.325000 69.180000  68.125000 ;
      RECT 68.380000  70.350000 69.180000  71.150000 ;
      RECT 68.380000  72.030000 69.180000  72.830000 ;
      RECT 68.380000  73.710000 69.180000  74.510000 ;
      RECT 68.380000  75.390000 69.180000  76.190000 ;
      RECT 68.380000  77.070000 69.180000  77.870000 ;
      RECT 68.380000  78.750000 69.180000  79.550000 ;
      RECT 68.380000  80.430000 69.180000  81.230000 ;
      RECT 68.380000  82.110000 69.180000  82.910000 ;
      RECT 68.380000  83.790000 69.180000  84.590000 ;
      RECT 68.380000  85.470000 69.180000  86.270000 ;
      RECT 68.380000  87.150000 69.180000  87.950000 ;
      RECT 68.380000  88.830000 69.180000  89.630000 ;
      RECT 68.380000  90.510000 69.180000  91.310000 ;
      RECT 68.380000  92.190000 69.180000  92.990000 ;
      RECT 68.380000  93.870000 69.180000  94.670000 ;
      RECT 68.380000 176.155000 69.180000 176.955000 ;
      RECT 68.380000 177.775000 69.180000 178.575000 ;
      RECT 68.380000 179.395000 69.180000 180.195000 ;
      RECT 68.380000 181.015000 69.180000 181.815000 ;
      RECT 68.380000 182.635000 69.180000 183.435000 ;
      RECT 68.380000 184.255000 69.180000 185.055000 ;
      RECT 68.380000 185.875000 69.180000 186.675000 ;
      RECT 68.380000 187.495000 69.180000 188.295000 ;
      RECT 68.380000 189.115000 69.180000 189.915000 ;
      RECT 68.380000 190.735000 69.180000 191.535000 ;
      RECT 68.380000 192.355000 69.180000 193.155000 ;
      RECT 68.380000 193.975000 69.180000 194.775000 ;
      RECT 68.380000 195.595000 69.180000 196.395000 ;
      RECT 68.380000 197.215000 69.180000 198.015000 ;
      RECT 68.380000 198.835000 69.180000 199.635000 ;
      RECT 68.385000  37.145000 69.185000  37.945000 ;
      RECT 68.385000  38.975000 69.185000  39.775000 ;
      RECT 68.385000  58.645000 69.185000  59.445000 ;
      RECT 68.385000  61.475000 69.185000  62.275000 ;
      RECT 69.975000   9.295000 70.775000  10.095000 ;
      RECT 69.975000  12.325000 70.775000  13.125000 ;
      RECT 69.975000  20.195000 70.775000  20.995000 ;
      RECT 69.975000  23.225000 70.775000  24.025000 ;
      RECT 69.975000  41.995000 70.775000  42.795000 ;
      RECT 69.975000  45.025000 70.775000  45.825000 ;
      RECT 69.980000   2.450000 70.780000   3.250000 ;
      RECT 69.980000   4.360000 70.780000   5.160000 ;
      RECT 69.980000   6.270000 70.780000   7.070000 ;
      RECT 69.980000  15.345000 70.780000  16.145000 ;
      RECT 69.980000  17.175000 70.780000  17.975000 ;
      RECT 69.980000  26.245000 70.780000  27.045000 ;
      RECT 69.980000  29.275000 70.780000  30.075000 ;
      RECT 69.980000  32.295000 70.780000  33.095000 ;
      RECT 69.980000  34.125000 70.780000  34.925000 ;
      RECT 69.980000  51.835000 70.780000  52.635000 ;
      RECT 69.980000  64.495000 70.780000  65.295000 ;
      RECT 69.980000  67.325000 70.780000  68.125000 ;
      RECT 69.980000  70.350000 70.780000  71.150000 ;
      RECT 69.980000  72.030000 70.780000  72.830000 ;
      RECT 69.980000  73.710000 70.780000  74.510000 ;
      RECT 69.980000  75.390000 70.780000  76.190000 ;
      RECT 69.980000  77.070000 70.780000  77.870000 ;
      RECT 69.980000  78.750000 70.780000  79.550000 ;
      RECT 69.980000  80.430000 70.780000  81.230000 ;
      RECT 69.980000  82.110000 70.780000  82.910000 ;
      RECT 69.980000  83.790000 70.780000  84.590000 ;
      RECT 69.980000  85.470000 70.780000  86.270000 ;
      RECT 69.980000  87.150000 70.780000  87.950000 ;
      RECT 69.980000  88.830000 70.780000  89.630000 ;
      RECT 69.980000  90.510000 70.780000  91.310000 ;
      RECT 69.980000  92.190000 70.780000  92.990000 ;
      RECT 69.980000  93.870000 70.780000  94.670000 ;
      RECT 69.980000 176.155000 70.780000 176.955000 ;
      RECT 69.980000 177.775000 70.780000 178.575000 ;
      RECT 69.980000 179.395000 70.780000 180.195000 ;
      RECT 69.980000 181.015000 70.780000 181.815000 ;
      RECT 69.980000 182.635000 70.780000 183.435000 ;
      RECT 69.980000 184.255000 70.780000 185.055000 ;
      RECT 69.980000 185.875000 70.780000 186.675000 ;
      RECT 69.980000 187.495000 70.780000 188.295000 ;
      RECT 69.980000 189.115000 70.780000 189.915000 ;
      RECT 69.980000 190.735000 70.780000 191.535000 ;
      RECT 69.980000 192.355000 70.780000 193.155000 ;
      RECT 69.980000 193.975000 70.780000 194.775000 ;
      RECT 69.980000 195.595000 70.780000 196.395000 ;
      RECT 69.980000 197.215000 70.780000 198.015000 ;
      RECT 69.980000 198.835000 70.780000 199.635000 ;
      RECT 69.985000  37.145000 70.785000  37.945000 ;
      RECT 69.985000  38.975000 70.785000  39.775000 ;
      RECT 69.985000  58.645000 70.785000  59.445000 ;
      RECT 69.985000  61.475000 70.785000  62.275000 ;
      RECT 71.575000   9.295000 72.375000  10.095000 ;
      RECT 71.575000  12.325000 72.375000  13.125000 ;
      RECT 71.575000  20.195000 72.375000  20.995000 ;
      RECT 71.575000  23.225000 72.375000  24.025000 ;
      RECT 71.575000  41.995000 72.375000  42.795000 ;
      RECT 71.575000  45.025000 72.375000  45.825000 ;
      RECT 71.580000   2.450000 72.380000   3.250000 ;
      RECT 71.580000   4.360000 72.380000   5.160000 ;
      RECT 71.580000   6.270000 72.380000   7.070000 ;
      RECT 71.580000  15.345000 72.380000  16.145000 ;
      RECT 71.580000  17.175000 72.380000  17.975000 ;
      RECT 71.580000  26.245000 72.380000  27.045000 ;
      RECT 71.580000  29.275000 72.380000  30.075000 ;
      RECT 71.580000  32.295000 72.380000  33.095000 ;
      RECT 71.580000  34.125000 72.380000  34.925000 ;
      RECT 71.580000  51.835000 72.380000  52.635000 ;
      RECT 71.580000  64.495000 72.380000  65.295000 ;
      RECT 71.580000  67.325000 72.380000  68.125000 ;
      RECT 71.580000  70.350000 72.380000  71.150000 ;
      RECT 71.580000  72.030000 72.380000  72.830000 ;
      RECT 71.580000  73.710000 72.380000  74.510000 ;
      RECT 71.580000  75.390000 72.380000  76.190000 ;
      RECT 71.580000  77.070000 72.380000  77.870000 ;
      RECT 71.580000  78.750000 72.380000  79.550000 ;
      RECT 71.580000  80.430000 72.380000  81.230000 ;
      RECT 71.580000  82.110000 72.380000  82.910000 ;
      RECT 71.580000  83.790000 72.380000  84.590000 ;
      RECT 71.580000  85.470000 72.380000  86.270000 ;
      RECT 71.580000  87.150000 72.380000  87.950000 ;
      RECT 71.580000  88.830000 72.380000  89.630000 ;
      RECT 71.580000  90.510000 72.380000  91.310000 ;
      RECT 71.580000  92.190000 72.380000  92.990000 ;
      RECT 71.580000  93.870000 72.380000  94.670000 ;
      RECT 71.580000 176.155000 72.380000 176.955000 ;
      RECT 71.580000 177.775000 72.380000 178.575000 ;
      RECT 71.580000 179.395000 72.380000 180.195000 ;
      RECT 71.580000 181.015000 72.380000 181.815000 ;
      RECT 71.580000 182.635000 72.380000 183.435000 ;
      RECT 71.580000 184.255000 72.380000 185.055000 ;
      RECT 71.580000 185.875000 72.380000 186.675000 ;
      RECT 71.580000 187.495000 72.380000 188.295000 ;
      RECT 71.580000 189.115000 72.380000 189.915000 ;
      RECT 71.580000 190.735000 72.380000 191.535000 ;
      RECT 71.580000 192.355000 72.380000 193.155000 ;
      RECT 71.580000 193.975000 72.380000 194.775000 ;
      RECT 71.580000 195.595000 72.380000 196.395000 ;
      RECT 71.580000 197.215000 72.380000 198.015000 ;
      RECT 71.580000 198.835000 72.380000 199.635000 ;
      RECT 71.585000  37.145000 72.385000  37.945000 ;
      RECT 71.585000  38.975000 72.385000  39.775000 ;
      RECT 71.585000  58.645000 72.385000  59.445000 ;
      RECT 71.585000  61.475000 72.385000  62.275000 ;
      RECT 73.175000   9.295000 73.975000  10.095000 ;
      RECT 73.175000  12.325000 73.975000  13.125000 ;
      RECT 73.175000  20.195000 73.975000  20.995000 ;
      RECT 73.175000  23.225000 73.975000  24.025000 ;
      RECT 73.175000  41.995000 73.975000  42.795000 ;
      RECT 73.175000  45.025000 73.975000  45.825000 ;
      RECT 73.180000   2.450000 73.980000   3.250000 ;
      RECT 73.180000   4.360000 73.980000   5.160000 ;
      RECT 73.180000   6.270000 73.980000   7.070000 ;
      RECT 73.180000  15.345000 73.980000  16.145000 ;
      RECT 73.180000  17.175000 73.980000  17.975000 ;
      RECT 73.180000  26.245000 73.980000  27.045000 ;
      RECT 73.180000  29.275000 73.980000  30.075000 ;
      RECT 73.180000  32.295000 73.980000  33.095000 ;
      RECT 73.180000  34.125000 73.980000  34.925000 ;
      RECT 73.180000  51.835000 73.980000  52.635000 ;
      RECT 73.180000  64.495000 73.980000  65.295000 ;
      RECT 73.180000  67.325000 73.980000  68.125000 ;
      RECT 73.180000  70.350000 73.980000  71.150000 ;
      RECT 73.180000  72.030000 73.980000  72.830000 ;
      RECT 73.180000  73.710000 73.980000  74.510000 ;
      RECT 73.180000  75.390000 73.980000  76.190000 ;
      RECT 73.180000  77.070000 73.980000  77.870000 ;
      RECT 73.180000  78.750000 73.980000  79.550000 ;
      RECT 73.180000  80.430000 73.980000  81.230000 ;
      RECT 73.180000  82.110000 73.980000  82.910000 ;
      RECT 73.180000  83.790000 73.980000  84.590000 ;
      RECT 73.180000  85.470000 73.980000  86.270000 ;
      RECT 73.180000  87.150000 73.980000  87.950000 ;
      RECT 73.180000  88.830000 73.980000  89.630000 ;
      RECT 73.180000  90.510000 73.980000  91.310000 ;
      RECT 73.180000  92.190000 73.980000  92.990000 ;
      RECT 73.180000  93.870000 73.980000  94.670000 ;
      RECT 73.180000 176.155000 73.980000 176.955000 ;
      RECT 73.180000 177.775000 73.980000 178.575000 ;
      RECT 73.180000 179.395000 73.980000 180.195000 ;
      RECT 73.180000 181.015000 73.980000 181.815000 ;
      RECT 73.180000 182.635000 73.980000 183.435000 ;
      RECT 73.180000 184.255000 73.980000 185.055000 ;
      RECT 73.180000 185.875000 73.980000 186.675000 ;
      RECT 73.180000 187.495000 73.980000 188.295000 ;
      RECT 73.180000 189.115000 73.980000 189.915000 ;
      RECT 73.180000 190.735000 73.980000 191.535000 ;
      RECT 73.180000 192.355000 73.980000 193.155000 ;
      RECT 73.180000 193.975000 73.980000 194.775000 ;
      RECT 73.180000 195.595000 73.980000 196.395000 ;
      RECT 73.180000 197.215000 73.980000 198.015000 ;
      RECT 73.180000 198.835000 73.980000 199.635000 ;
      RECT 73.185000  37.145000 73.985000  37.945000 ;
      RECT 73.185000  38.975000 73.985000  39.775000 ;
      RECT 73.185000  58.645000 73.985000  59.445000 ;
      RECT 73.185000  61.475000 73.985000  62.275000 ;
      RECT 74.775000   9.295000 75.575000  10.095000 ;
      RECT 74.775000  12.325000 75.575000  13.125000 ;
      RECT 74.775000  20.195000 75.575000  20.995000 ;
      RECT 74.775000  23.225000 75.575000  24.025000 ;
      RECT 74.775000  41.995000 75.575000  42.795000 ;
      RECT 74.775000  45.025000 75.575000  45.825000 ;
      RECT 74.780000   2.450000 75.580000   3.250000 ;
      RECT 74.780000   4.360000 75.580000   5.160000 ;
      RECT 74.780000   6.270000 75.580000   7.070000 ;
      RECT 74.780000  15.345000 75.580000  16.145000 ;
      RECT 74.780000  17.175000 75.580000  17.975000 ;
      RECT 74.780000  26.245000 75.580000  27.045000 ;
      RECT 74.780000  29.275000 75.580000  30.075000 ;
      RECT 74.780000  32.295000 75.580000  33.095000 ;
      RECT 74.780000  34.125000 75.580000  34.925000 ;
      RECT 74.780000  51.835000 75.580000  52.635000 ;
      RECT 74.780000  64.495000 75.580000  65.295000 ;
      RECT 74.780000  67.325000 75.580000  68.125000 ;
      RECT 74.780000  70.350000 75.580000  71.150000 ;
      RECT 74.780000  72.030000 75.580000  72.830000 ;
      RECT 74.780000  73.710000 75.580000  74.510000 ;
      RECT 74.780000  75.390000 75.580000  76.190000 ;
      RECT 74.780000  77.070000 75.580000  77.870000 ;
      RECT 74.780000  78.750000 75.580000  79.550000 ;
      RECT 74.780000  80.430000 75.580000  81.230000 ;
      RECT 74.780000  82.110000 75.580000  82.910000 ;
      RECT 74.780000  83.790000 75.580000  84.590000 ;
      RECT 74.780000  85.470000 75.580000  86.270000 ;
      RECT 74.780000  87.150000 75.580000  87.950000 ;
      RECT 74.780000  88.830000 75.580000  89.630000 ;
      RECT 74.780000  90.510000 75.580000  91.310000 ;
      RECT 74.780000  92.190000 75.580000  92.990000 ;
      RECT 74.780000  93.870000 75.580000  94.670000 ;
      RECT 74.780000 176.155000 75.580000 176.955000 ;
      RECT 74.780000 177.775000 75.580000 178.575000 ;
      RECT 74.780000 179.395000 75.580000 180.195000 ;
      RECT 74.780000 181.015000 75.580000 181.815000 ;
      RECT 74.780000 182.635000 75.580000 183.435000 ;
      RECT 74.780000 184.255000 75.580000 185.055000 ;
      RECT 74.780000 185.875000 75.580000 186.675000 ;
      RECT 74.780000 187.495000 75.580000 188.295000 ;
      RECT 74.780000 189.115000 75.580000 189.915000 ;
      RECT 74.780000 190.735000 75.580000 191.535000 ;
      RECT 74.780000 192.355000 75.580000 193.155000 ;
      RECT 74.780000 193.975000 75.580000 194.775000 ;
      RECT 74.780000 195.595000 75.580000 196.395000 ;
      RECT 74.780000 197.215000 75.580000 198.015000 ;
      RECT 74.780000 198.835000 75.580000 199.635000 ;
      RECT 74.785000  37.145000 75.585000  37.945000 ;
      RECT 74.785000  38.975000 75.585000  39.775000 ;
      RECT 74.785000  58.645000 75.585000  59.445000 ;
      RECT 74.785000  61.475000 75.585000  62.275000 ;
      RECT 76.375000   9.295000 77.175000  10.095000 ;
      RECT 76.375000  12.325000 77.175000  13.125000 ;
      RECT 76.375000  20.195000 77.175000  20.995000 ;
      RECT 76.375000  23.225000 77.175000  24.025000 ;
      RECT 76.375000  41.995000 77.175000  42.795000 ;
      RECT 76.375000  45.025000 77.175000  45.825000 ;
      RECT 76.380000   2.450000 77.180000   3.250000 ;
      RECT 76.380000   4.360000 77.180000   5.160000 ;
      RECT 76.380000   6.270000 77.180000   7.070000 ;
      RECT 76.380000  15.345000 77.180000  16.145000 ;
      RECT 76.380000  17.175000 77.180000  17.975000 ;
      RECT 76.380000  26.245000 77.180000  27.045000 ;
      RECT 76.380000  29.275000 77.180000  30.075000 ;
      RECT 76.380000  32.295000 77.180000  33.095000 ;
      RECT 76.380000  34.125000 77.180000  34.925000 ;
      RECT 76.380000  51.835000 77.180000  52.635000 ;
      RECT 76.380000  64.495000 77.180000  65.295000 ;
      RECT 76.380000  67.325000 77.180000  68.125000 ;
      RECT 76.380000  70.350000 77.180000  71.150000 ;
      RECT 76.380000  72.030000 77.180000  72.830000 ;
      RECT 76.380000  73.710000 77.180000  74.510000 ;
      RECT 76.380000  75.390000 77.180000  76.190000 ;
      RECT 76.380000  77.070000 77.180000  77.870000 ;
      RECT 76.380000  78.750000 77.180000  79.550000 ;
      RECT 76.380000  80.430000 77.180000  81.230000 ;
      RECT 76.380000  82.110000 77.180000  82.910000 ;
      RECT 76.380000  83.790000 77.180000  84.590000 ;
      RECT 76.380000  85.470000 77.180000  86.270000 ;
      RECT 76.380000  87.150000 77.180000  87.950000 ;
      RECT 76.380000  88.830000 77.180000  89.630000 ;
      RECT 76.380000  90.510000 77.180000  91.310000 ;
      RECT 76.380000  92.190000 77.180000  92.990000 ;
      RECT 76.380000  93.870000 77.180000  94.670000 ;
      RECT 76.380000 176.155000 77.180000 176.955000 ;
      RECT 76.380000 177.775000 77.180000 178.575000 ;
      RECT 76.380000 179.395000 77.180000 180.195000 ;
      RECT 76.380000 181.015000 77.180000 181.815000 ;
      RECT 76.380000 182.635000 77.180000 183.435000 ;
      RECT 76.380000 184.255000 77.180000 185.055000 ;
      RECT 76.380000 185.875000 77.180000 186.675000 ;
      RECT 76.380000 187.495000 77.180000 188.295000 ;
      RECT 76.380000 189.115000 77.180000 189.915000 ;
      RECT 76.380000 190.735000 77.180000 191.535000 ;
      RECT 76.380000 192.355000 77.180000 193.155000 ;
      RECT 76.380000 193.975000 77.180000 194.775000 ;
      RECT 76.380000 195.595000 77.180000 196.395000 ;
      RECT 76.380000 197.215000 77.180000 198.015000 ;
      RECT 76.380000 198.835000 77.180000 199.635000 ;
      RECT 76.385000  37.145000 77.185000  37.945000 ;
      RECT 76.385000  38.975000 77.185000  39.775000 ;
      RECT 76.385000  58.645000 77.185000  59.445000 ;
      RECT 76.385000  61.475000 77.185000  62.275000 ;
      RECT 77.975000   9.295000 78.775000  10.095000 ;
      RECT 77.975000  12.325000 78.775000  13.125000 ;
      RECT 77.975000  20.195000 78.775000  20.995000 ;
      RECT 77.975000  23.225000 78.775000  24.025000 ;
      RECT 77.975000  41.995000 78.775000  42.795000 ;
      RECT 77.975000  45.025000 78.775000  45.825000 ;
      RECT 77.980000   2.450000 78.780000   3.250000 ;
      RECT 77.980000   4.360000 78.780000   5.160000 ;
      RECT 77.980000   6.270000 78.780000   7.070000 ;
      RECT 77.980000  15.345000 78.780000  16.145000 ;
      RECT 77.980000  17.175000 78.780000  17.975000 ;
      RECT 77.980000  26.245000 78.780000  27.045000 ;
      RECT 77.980000  29.275000 78.780000  30.075000 ;
      RECT 77.980000  32.295000 78.780000  33.095000 ;
      RECT 77.980000  34.125000 78.780000  34.925000 ;
      RECT 77.980000  51.835000 78.780000  52.635000 ;
      RECT 77.980000  64.495000 78.780000  65.295000 ;
      RECT 77.980000  67.325000 78.780000  68.125000 ;
      RECT 77.980000  70.350000 78.780000  71.150000 ;
      RECT 77.980000  72.030000 78.780000  72.830000 ;
      RECT 77.980000  73.710000 78.780000  74.510000 ;
      RECT 77.980000  75.390000 78.780000  76.190000 ;
      RECT 77.980000  77.070000 78.780000  77.870000 ;
      RECT 77.980000  78.750000 78.780000  79.550000 ;
      RECT 77.980000  80.430000 78.780000  81.230000 ;
      RECT 77.980000  82.110000 78.780000  82.910000 ;
      RECT 77.980000  83.790000 78.780000  84.590000 ;
      RECT 77.980000  85.470000 78.780000  86.270000 ;
      RECT 77.980000  87.150000 78.780000  87.950000 ;
      RECT 77.980000  88.830000 78.780000  89.630000 ;
      RECT 77.980000  90.510000 78.780000  91.310000 ;
      RECT 77.980000  92.190000 78.780000  92.990000 ;
      RECT 77.980000  93.870000 78.780000  94.670000 ;
      RECT 77.980000 176.155000 78.780000 176.955000 ;
      RECT 77.980000 177.775000 78.780000 178.575000 ;
      RECT 77.980000 179.395000 78.780000 180.195000 ;
      RECT 77.980000 181.015000 78.780000 181.815000 ;
      RECT 77.980000 182.635000 78.780000 183.435000 ;
      RECT 77.980000 184.255000 78.780000 185.055000 ;
      RECT 77.980000 185.875000 78.780000 186.675000 ;
      RECT 77.980000 187.495000 78.780000 188.295000 ;
      RECT 77.980000 189.115000 78.780000 189.915000 ;
      RECT 77.980000 190.735000 78.780000 191.535000 ;
      RECT 77.980000 192.355000 78.780000 193.155000 ;
      RECT 77.980000 193.975000 78.780000 194.775000 ;
      RECT 77.980000 195.595000 78.780000 196.395000 ;
      RECT 77.980000 197.215000 78.780000 198.015000 ;
      RECT 77.980000 198.835000 78.780000 199.635000 ;
      RECT 77.985000  37.145000 78.785000  37.945000 ;
      RECT 77.985000  38.975000 78.785000  39.775000 ;
      RECT 77.985000  58.645000 78.785000  59.445000 ;
      RECT 77.985000  61.475000 78.785000  62.275000 ;
  END
END sky130_fd_io__overlay_gpiov2
END LIBRARY
