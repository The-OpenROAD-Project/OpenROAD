module dual_spm (clk,
    rstn,
    x,
    y,
    a);
 input clk;
 input rstn;
 input x;
 output y;
 input [31:0] a;

 wire y_iso;

 spm spm_inst_0 (.clk(clk),
    .rst(rstn),
    .x(x),
    .y(y_iso),
    .a({a[31],
    a[30],
    a[29],
    a[28],
    a[27],
    a[26],
    a[25],
    a[24],
    a[23],
    a[22],
    a[21],
    a[20],
    a[19],
    a[18],
    a[17],
    a[16],
    a[15],
    a[14],
    a[13],
    a[12],
    a[11],
    a[10],
    a[9],
    a[8],
    a[7],
    a[6],
    a[5],
    a[4],
    a[3],
    a[2],
    a[1],
    a[0]}));
 spm spm_inst_1 (.clk(clk),
    .rst(rstn),
    .x(y_iso),
    .y(y),
    .a({a[31],
    a[30],
    a[29],
    a[28],
    a[27],
    a[26],
    a[25],
    a[24],
    a[23],
    a[22],
    a[21],
    a[20],
    a[19],
    a[18],
    a[17],
    a[16],
    a[15],
    a[14],
    a[13],
    a[12],
    a[11],
    a[10],
    a[9],
    a[8],
    a[7],
    a[6],
    a[5],
    a[4],
    a[3],
    a[2],
    a[1],
    a[0]}));
endmodule
