VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.1 ;

SITE site1
  CLASS CORE ;
  SIZE 50 BY 20 ;
END site1

MACRO bidir
 SIZE 50 BY 20 ;
 PIN IO DIRECTION INOUT ; END IO
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END bidir

END LIBRARY
