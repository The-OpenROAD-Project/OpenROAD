module test_no_clk ();

 INV_X1 inv1 (.ZN(a));
 INV_X1 inv2 (.A(a));

endmodule
