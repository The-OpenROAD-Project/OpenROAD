# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_io__overlay_vssa_hvc
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 200 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 1.270000 56.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 53.125000 75.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 1.270000 51.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 48.365000 75.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 8.885000 1.270000 13.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 8.885000 75.000000 13.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 8.985000 1.270000 13.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 8.985000 75.000000 13.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2.035000 1.270000 7.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 2.035000 75.000000 7.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 2.135000 1.270000 7.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 2.135000 75.000000 7.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 14.935000 0.965000 18.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035000 14.935000 75.000000 18.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 15.035000 0.965000 18.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 15.035000 75.000000 18.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 19.785000 1.270000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 70.035000 1.270000 95.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 19.785000 75.000000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 70.035000 75.000000 95.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 19.885000 1.270000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 70.035000 1.270000 94.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 19.885000 75.000000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 70.035000 75.000000 94.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 64.085000 1.270000 68.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 64.085000 75.000000 68.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 64.185000 1.270000 68.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 64.185000 75.000000 68.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.495000 51.650000 24.395000 52.820000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 47.740000 24.395000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 56.410000 24.395000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.970000 36.740000 24.395000 40.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390000 36.740000 74.290000 40.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390000 47.740000 74.290000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390000 51.650000 74.290000 52.820000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390000 56.410000 74.290000 56.730000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 36.735000 24.370000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 47.735000 24.370000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 51.645000 24.370000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 56.405000 24.370000 56.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.415000 36.735000 75.000000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.415000 47.735000 75.000000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.415000 51.645000 75.000000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.415000 56.405000 75.000000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 36.840000 1.270000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 47.735000 1.270000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 36.840000 75.000000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 47.735000 75.000000 56.735000 ;
    END
    PORT
      LAYER via3 ;
        RECT  0.585000 51.715000  0.785000 51.915000 ;
        RECT  0.585000 52.135000  0.785000 52.335000 ;
        RECT  0.585000 52.555000  0.785000 52.755000 ;
        RECT  0.620000 47.800000  0.820000 48.000000 ;
        RECT  0.620000 56.470000  0.820000 56.670000 ;
        RECT  0.995000 51.715000  1.195000 51.915000 ;
        RECT  0.995000 52.135000  1.195000 52.335000 ;
        RECT  0.995000 52.555000  1.195000 52.755000 ;
        RECT  1.025000 47.800000  1.225000 48.000000 ;
        RECT  1.025000 56.470000  1.225000 56.670000 ;
        RECT  1.060000 36.820000  1.260000 37.020000 ;
        RECT  1.060000 37.260000  1.260000 37.460000 ;
        RECT  1.060000 37.700000  1.260000 37.900000 ;
        RECT  1.060000 38.140000  1.260000 38.340000 ;
        RECT  1.060000 38.580000  1.260000 38.780000 ;
        RECT  1.060000 39.020000  1.260000 39.220000 ;
        RECT  1.060000 39.460000  1.260000 39.660000 ;
        RECT  1.060000 39.900000  1.260000 40.100000 ;
        RECT  1.405000 51.715000  1.605000 51.915000 ;
        RECT  1.405000 52.135000  1.605000 52.335000 ;
        RECT  1.405000 52.555000  1.605000 52.755000 ;
        RECT  1.430000 47.800000  1.630000 48.000000 ;
        RECT  1.430000 56.470000  1.630000 56.670000 ;
        RECT  1.465000 36.820000  1.665000 37.020000 ;
        RECT  1.465000 37.260000  1.665000 37.460000 ;
        RECT  1.465000 37.700000  1.665000 37.900000 ;
        RECT  1.465000 38.140000  1.665000 38.340000 ;
        RECT  1.465000 38.580000  1.665000 38.780000 ;
        RECT  1.465000 39.020000  1.665000 39.220000 ;
        RECT  1.465000 39.460000  1.665000 39.660000 ;
        RECT  1.465000 39.900000  1.665000 40.100000 ;
        RECT  1.815000 51.715000  2.015000 51.915000 ;
        RECT  1.815000 52.135000  2.015000 52.335000 ;
        RECT  1.815000 52.555000  2.015000 52.755000 ;
        RECT  1.835000 47.800000  2.035000 48.000000 ;
        RECT  1.835000 56.470000  2.035000 56.670000 ;
        RECT  1.870000 36.820000  2.070000 37.020000 ;
        RECT  1.870000 37.260000  2.070000 37.460000 ;
        RECT  1.870000 37.700000  2.070000 37.900000 ;
        RECT  1.870000 38.140000  2.070000 38.340000 ;
        RECT  1.870000 38.580000  2.070000 38.780000 ;
        RECT  1.870000 39.020000  2.070000 39.220000 ;
        RECT  1.870000 39.460000  2.070000 39.660000 ;
        RECT  1.870000 39.900000  2.070000 40.100000 ;
        RECT  2.225000 51.715000  2.425000 51.915000 ;
        RECT  2.225000 52.135000  2.425000 52.335000 ;
        RECT  2.225000 52.555000  2.425000 52.755000 ;
        RECT  2.240000 47.800000  2.440000 48.000000 ;
        RECT  2.240000 56.470000  2.440000 56.670000 ;
        RECT  2.275000 36.820000  2.475000 37.020000 ;
        RECT  2.275000 37.260000  2.475000 37.460000 ;
        RECT  2.275000 37.700000  2.475000 37.900000 ;
        RECT  2.275000 38.140000  2.475000 38.340000 ;
        RECT  2.275000 38.580000  2.475000 38.780000 ;
        RECT  2.275000 39.020000  2.475000 39.220000 ;
        RECT  2.275000 39.460000  2.475000 39.660000 ;
        RECT  2.275000 39.900000  2.475000 40.100000 ;
        RECT  2.635000 51.715000  2.835000 51.915000 ;
        RECT  2.635000 52.135000  2.835000 52.335000 ;
        RECT  2.635000 52.555000  2.835000 52.755000 ;
        RECT  2.645000 47.800000  2.845000 48.000000 ;
        RECT  2.645000 56.470000  2.845000 56.670000 ;
        RECT  2.680000 36.820000  2.880000 37.020000 ;
        RECT  2.680000 37.260000  2.880000 37.460000 ;
        RECT  2.680000 37.700000  2.880000 37.900000 ;
        RECT  2.680000 38.140000  2.880000 38.340000 ;
        RECT  2.680000 38.580000  2.880000 38.780000 ;
        RECT  2.680000 39.020000  2.880000 39.220000 ;
        RECT  2.680000 39.460000  2.880000 39.660000 ;
        RECT  2.680000 39.900000  2.880000 40.100000 ;
        RECT  3.045000 51.715000  3.245000 51.915000 ;
        RECT  3.045000 52.135000  3.245000 52.335000 ;
        RECT  3.045000 52.555000  3.245000 52.755000 ;
        RECT  3.050000 47.800000  3.250000 48.000000 ;
        RECT  3.050000 56.470000  3.250000 56.670000 ;
        RECT  3.085000 36.820000  3.285000 37.020000 ;
        RECT  3.085000 37.260000  3.285000 37.460000 ;
        RECT  3.085000 37.700000  3.285000 37.900000 ;
        RECT  3.085000 38.140000  3.285000 38.340000 ;
        RECT  3.085000 38.580000  3.285000 38.780000 ;
        RECT  3.085000 39.020000  3.285000 39.220000 ;
        RECT  3.085000 39.460000  3.285000 39.660000 ;
        RECT  3.085000 39.900000  3.285000 40.100000 ;
        RECT  3.450000 51.715000  3.650000 51.915000 ;
        RECT  3.450000 52.135000  3.650000 52.335000 ;
        RECT  3.450000 52.555000  3.650000 52.755000 ;
        RECT  3.455000 47.800000  3.655000 48.000000 ;
        RECT  3.455000 56.470000  3.655000 56.670000 ;
        RECT  3.490000 36.820000  3.690000 37.020000 ;
        RECT  3.490000 37.260000  3.690000 37.460000 ;
        RECT  3.490000 37.700000  3.690000 37.900000 ;
        RECT  3.490000 38.140000  3.690000 38.340000 ;
        RECT  3.490000 38.580000  3.690000 38.780000 ;
        RECT  3.490000 39.020000  3.690000 39.220000 ;
        RECT  3.490000 39.460000  3.690000 39.660000 ;
        RECT  3.490000 39.900000  3.690000 40.100000 ;
        RECT  3.855000 51.715000  4.055000 51.915000 ;
        RECT  3.855000 52.135000  4.055000 52.335000 ;
        RECT  3.855000 52.555000  4.055000 52.755000 ;
        RECT  3.860000 47.800000  4.060000 48.000000 ;
        RECT  3.860000 56.470000  4.060000 56.670000 ;
        RECT  3.895000 36.820000  4.095000 37.020000 ;
        RECT  3.895000 37.260000  4.095000 37.460000 ;
        RECT  3.895000 37.700000  4.095000 37.900000 ;
        RECT  3.895000 38.140000  4.095000 38.340000 ;
        RECT  3.895000 38.580000  4.095000 38.780000 ;
        RECT  3.895000 39.020000  4.095000 39.220000 ;
        RECT  3.895000 39.460000  4.095000 39.660000 ;
        RECT  3.895000 39.900000  4.095000 40.100000 ;
        RECT  4.260000 51.715000  4.460000 51.915000 ;
        RECT  4.260000 52.135000  4.460000 52.335000 ;
        RECT  4.260000 52.555000  4.460000 52.755000 ;
        RECT  4.265000 47.800000  4.465000 48.000000 ;
        RECT  4.265000 56.470000  4.465000 56.670000 ;
        RECT  4.300000 36.820000  4.500000 37.020000 ;
        RECT  4.300000 37.260000  4.500000 37.460000 ;
        RECT  4.300000 37.700000  4.500000 37.900000 ;
        RECT  4.300000 38.140000  4.500000 38.340000 ;
        RECT  4.300000 38.580000  4.500000 38.780000 ;
        RECT  4.300000 39.020000  4.500000 39.220000 ;
        RECT  4.300000 39.460000  4.500000 39.660000 ;
        RECT  4.300000 39.900000  4.500000 40.100000 ;
        RECT  4.665000 51.715000  4.865000 51.915000 ;
        RECT  4.665000 52.135000  4.865000 52.335000 ;
        RECT  4.665000 52.555000  4.865000 52.755000 ;
        RECT  4.670000 47.800000  4.870000 48.000000 ;
        RECT  4.670000 56.470000  4.870000 56.670000 ;
        RECT  4.705000 36.820000  4.905000 37.020000 ;
        RECT  4.705000 37.260000  4.905000 37.460000 ;
        RECT  4.705000 37.700000  4.905000 37.900000 ;
        RECT  4.705000 38.140000  4.905000 38.340000 ;
        RECT  4.705000 38.580000  4.905000 38.780000 ;
        RECT  4.705000 39.020000  4.905000 39.220000 ;
        RECT  4.705000 39.460000  4.905000 39.660000 ;
        RECT  4.705000 39.900000  4.905000 40.100000 ;
        RECT  5.070000 51.715000  5.270000 51.915000 ;
        RECT  5.070000 52.135000  5.270000 52.335000 ;
        RECT  5.070000 52.555000  5.270000 52.755000 ;
        RECT  5.075000 47.800000  5.275000 48.000000 ;
        RECT  5.075000 56.470000  5.275000 56.670000 ;
        RECT  5.110000 36.820000  5.310000 37.020000 ;
        RECT  5.110000 37.260000  5.310000 37.460000 ;
        RECT  5.110000 37.700000  5.310000 37.900000 ;
        RECT  5.110000 38.140000  5.310000 38.340000 ;
        RECT  5.110000 38.580000  5.310000 38.780000 ;
        RECT  5.110000 39.020000  5.310000 39.220000 ;
        RECT  5.110000 39.460000  5.310000 39.660000 ;
        RECT  5.110000 39.900000  5.310000 40.100000 ;
        RECT  5.475000 51.715000  5.675000 51.915000 ;
        RECT  5.475000 52.135000  5.675000 52.335000 ;
        RECT  5.475000 52.555000  5.675000 52.755000 ;
        RECT  5.480000 47.800000  5.680000 48.000000 ;
        RECT  5.480000 56.470000  5.680000 56.670000 ;
        RECT  5.515000 36.820000  5.715000 37.020000 ;
        RECT  5.515000 37.260000  5.715000 37.460000 ;
        RECT  5.515000 37.700000  5.715000 37.900000 ;
        RECT  5.515000 38.140000  5.715000 38.340000 ;
        RECT  5.515000 38.580000  5.715000 38.780000 ;
        RECT  5.515000 39.020000  5.715000 39.220000 ;
        RECT  5.515000 39.460000  5.715000 39.660000 ;
        RECT  5.515000 39.900000  5.715000 40.100000 ;
        RECT  5.880000 51.715000  6.080000 51.915000 ;
        RECT  5.880000 52.135000  6.080000 52.335000 ;
        RECT  5.880000 52.555000  6.080000 52.755000 ;
        RECT  5.885000 47.800000  6.085000 48.000000 ;
        RECT  5.885000 56.470000  6.085000 56.670000 ;
        RECT  5.920000 36.820000  6.120000 37.020000 ;
        RECT  5.920000 37.260000  6.120000 37.460000 ;
        RECT  5.920000 37.700000  6.120000 37.900000 ;
        RECT  5.920000 38.140000  6.120000 38.340000 ;
        RECT  5.920000 38.580000  6.120000 38.780000 ;
        RECT  5.920000 39.020000  6.120000 39.220000 ;
        RECT  5.920000 39.460000  6.120000 39.660000 ;
        RECT  5.920000 39.900000  6.120000 40.100000 ;
        RECT  6.285000 51.715000  6.485000 51.915000 ;
        RECT  6.285000 52.135000  6.485000 52.335000 ;
        RECT  6.285000 52.555000  6.485000 52.755000 ;
        RECT  6.290000 47.800000  6.490000 48.000000 ;
        RECT  6.290000 56.470000  6.490000 56.670000 ;
        RECT  6.325000 36.820000  6.525000 37.020000 ;
        RECT  6.325000 37.260000  6.525000 37.460000 ;
        RECT  6.325000 37.700000  6.525000 37.900000 ;
        RECT  6.325000 38.140000  6.525000 38.340000 ;
        RECT  6.325000 38.580000  6.525000 38.780000 ;
        RECT  6.325000 39.020000  6.525000 39.220000 ;
        RECT  6.325000 39.460000  6.525000 39.660000 ;
        RECT  6.325000 39.900000  6.525000 40.100000 ;
        RECT  6.690000 51.715000  6.890000 51.915000 ;
        RECT  6.690000 52.135000  6.890000 52.335000 ;
        RECT  6.690000 52.555000  6.890000 52.755000 ;
        RECT  6.695000 47.800000  6.895000 48.000000 ;
        RECT  6.695000 56.470000  6.895000 56.670000 ;
        RECT  6.730000 36.820000  6.930000 37.020000 ;
        RECT  6.730000 37.260000  6.930000 37.460000 ;
        RECT  6.730000 37.700000  6.930000 37.900000 ;
        RECT  6.730000 38.140000  6.930000 38.340000 ;
        RECT  6.730000 38.580000  6.930000 38.780000 ;
        RECT  6.730000 39.020000  6.930000 39.220000 ;
        RECT  6.730000 39.460000  6.930000 39.660000 ;
        RECT  6.730000 39.900000  6.930000 40.100000 ;
        RECT  7.095000 51.715000  7.295000 51.915000 ;
        RECT  7.095000 52.135000  7.295000 52.335000 ;
        RECT  7.095000 52.555000  7.295000 52.755000 ;
        RECT  7.100000 47.800000  7.300000 48.000000 ;
        RECT  7.100000 56.470000  7.300000 56.670000 ;
        RECT  7.135000 36.820000  7.335000 37.020000 ;
        RECT  7.135000 37.260000  7.335000 37.460000 ;
        RECT  7.135000 37.700000  7.335000 37.900000 ;
        RECT  7.135000 38.140000  7.335000 38.340000 ;
        RECT  7.135000 38.580000  7.335000 38.780000 ;
        RECT  7.135000 39.020000  7.335000 39.220000 ;
        RECT  7.135000 39.460000  7.335000 39.660000 ;
        RECT  7.135000 39.900000  7.335000 40.100000 ;
        RECT  7.500000 51.715000  7.700000 51.915000 ;
        RECT  7.500000 52.135000  7.700000 52.335000 ;
        RECT  7.500000 52.555000  7.700000 52.755000 ;
        RECT  7.505000 47.800000  7.705000 48.000000 ;
        RECT  7.505000 56.470000  7.705000 56.670000 ;
        RECT  7.540000 36.820000  7.740000 37.020000 ;
        RECT  7.540000 37.260000  7.740000 37.460000 ;
        RECT  7.540000 37.700000  7.740000 37.900000 ;
        RECT  7.540000 38.140000  7.740000 38.340000 ;
        RECT  7.540000 38.580000  7.740000 38.780000 ;
        RECT  7.540000 39.020000  7.740000 39.220000 ;
        RECT  7.540000 39.460000  7.740000 39.660000 ;
        RECT  7.540000 39.900000  7.740000 40.100000 ;
        RECT  7.905000 51.715000  8.105000 51.915000 ;
        RECT  7.905000 52.135000  8.105000 52.335000 ;
        RECT  7.905000 52.555000  8.105000 52.755000 ;
        RECT  7.910000 47.800000  8.110000 48.000000 ;
        RECT  7.910000 56.470000  8.110000 56.670000 ;
        RECT  7.945000 36.820000  8.145000 37.020000 ;
        RECT  7.945000 37.260000  8.145000 37.460000 ;
        RECT  7.945000 37.700000  8.145000 37.900000 ;
        RECT  7.945000 38.140000  8.145000 38.340000 ;
        RECT  7.945000 38.580000  8.145000 38.780000 ;
        RECT  7.945000 39.020000  8.145000 39.220000 ;
        RECT  7.945000 39.460000  8.145000 39.660000 ;
        RECT  7.945000 39.900000  8.145000 40.100000 ;
        RECT  8.310000 51.715000  8.510000 51.915000 ;
        RECT  8.310000 52.135000  8.510000 52.335000 ;
        RECT  8.310000 52.555000  8.510000 52.755000 ;
        RECT  8.315000 47.800000  8.515000 48.000000 ;
        RECT  8.315000 56.470000  8.515000 56.670000 ;
        RECT  8.350000 36.820000  8.550000 37.020000 ;
        RECT  8.350000 37.260000  8.550000 37.460000 ;
        RECT  8.350000 37.700000  8.550000 37.900000 ;
        RECT  8.350000 38.140000  8.550000 38.340000 ;
        RECT  8.350000 38.580000  8.550000 38.780000 ;
        RECT  8.350000 39.020000  8.550000 39.220000 ;
        RECT  8.350000 39.460000  8.550000 39.660000 ;
        RECT  8.350000 39.900000  8.550000 40.100000 ;
        RECT  8.715000 51.715000  8.915000 51.915000 ;
        RECT  8.715000 52.135000  8.915000 52.335000 ;
        RECT  8.715000 52.555000  8.915000 52.755000 ;
        RECT  8.720000 47.800000  8.920000 48.000000 ;
        RECT  8.720000 56.470000  8.920000 56.670000 ;
        RECT  8.755000 36.820000  8.955000 37.020000 ;
        RECT  8.755000 37.260000  8.955000 37.460000 ;
        RECT  8.755000 37.700000  8.955000 37.900000 ;
        RECT  8.755000 38.140000  8.955000 38.340000 ;
        RECT  8.755000 38.580000  8.955000 38.780000 ;
        RECT  8.755000 39.020000  8.955000 39.220000 ;
        RECT  8.755000 39.460000  8.955000 39.660000 ;
        RECT  8.755000 39.900000  8.955000 40.100000 ;
        RECT  9.120000 51.715000  9.320000 51.915000 ;
        RECT  9.120000 52.135000  9.320000 52.335000 ;
        RECT  9.120000 52.555000  9.320000 52.755000 ;
        RECT  9.125000 47.800000  9.325000 48.000000 ;
        RECT  9.125000 56.470000  9.325000 56.670000 ;
        RECT  9.160000 36.820000  9.360000 37.020000 ;
        RECT  9.160000 37.260000  9.360000 37.460000 ;
        RECT  9.160000 37.700000  9.360000 37.900000 ;
        RECT  9.160000 38.140000  9.360000 38.340000 ;
        RECT  9.160000 38.580000  9.360000 38.780000 ;
        RECT  9.160000 39.020000  9.360000 39.220000 ;
        RECT  9.160000 39.460000  9.360000 39.660000 ;
        RECT  9.160000 39.900000  9.360000 40.100000 ;
        RECT  9.525000 51.715000  9.725000 51.915000 ;
        RECT  9.525000 52.135000  9.725000 52.335000 ;
        RECT  9.525000 52.555000  9.725000 52.755000 ;
        RECT  9.530000 47.800000  9.730000 48.000000 ;
        RECT  9.530000 56.470000  9.730000 56.670000 ;
        RECT  9.565000 36.820000  9.765000 37.020000 ;
        RECT  9.565000 37.260000  9.765000 37.460000 ;
        RECT  9.565000 37.700000  9.765000 37.900000 ;
        RECT  9.565000 38.140000  9.765000 38.340000 ;
        RECT  9.565000 38.580000  9.765000 38.780000 ;
        RECT  9.565000 39.020000  9.765000 39.220000 ;
        RECT  9.565000 39.460000  9.765000 39.660000 ;
        RECT  9.565000 39.900000  9.765000 40.100000 ;
        RECT  9.930000 51.715000 10.130000 51.915000 ;
        RECT  9.930000 52.135000 10.130000 52.335000 ;
        RECT  9.930000 52.555000 10.130000 52.755000 ;
        RECT  9.935000 47.800000 10.135000 48.000000 ;
        RECT  9.935000 56.470000 10.135000 56.670000 ;
        RECT  9.970000 36.820000 10.170000 37.020000 ;
        RECT  9.970000 37.260000 10.170000 37.460000 ;
        RECT  9.970000 37.700000 10.170000 37.900000 ;
        RECT  9.970000 38.140000 10.170000 38.340000 ;
        RECT  9.970000 38.580000 10.170000 38.780000 ;
        RECT  9.970000 39.020000 10.170000 39.220000 ;
        RECT  9.970000 39.460000 10.170000 39.660000 ;
        RECT  9.970000 39.900000 10.170000 40.100000 ;
        RECT 10.335000 51.715000 10.535000 51.915000 ;
        RECT 10.335000 52.135000 10.535000 52.335000 ;
        RECT 10.335000 52.555000 10.535000 52.755000 ;
        RECT 10.340000 47.800000 10.540000 48.000000 ;
        RECT 10.340000 56.470000 10.540000 56.670000 ;
        RECT 10.375000 36.820000 10.575000 37.020000 ;
        RECT 10.375000 37.260000 10.575000 37.460000 ;
        RECT 10.375000 37.700000 10.575000 37.900000 ;
        RECT 10.375000 38.140000 10.575000 38.340000 ;
        RECT 10.375000 38.580000 10.575000 38.780000 ;
        RECT 10.375000 39.020000 10.575000 39.220000 ;
        RECT 10.375000 39.460000 10.575000 39.660000 ;
        RECT 10.375000 39.900000 10.575000 40.100000 ;
        RECT 10.740000 51.715000 10.940000 51.915000 ;
        RECT 10.740000 52.135000 10.940000 52.335000 ;
        RECT 10.740000 52.555000 10.940000 52.755000 ;
        RECT 10.745000 47.800000 10.945000 48.000000 ;
        RECT 10.745000 56.470000 10.945000 56.670000 ;
        RECT 10.780000 36.820000 10.980000 37.020000 ;
        RECT 10.780000 37.260000 10.980000 37.460000 ;
        RECT 10.780000 37.700000 10.980000 37.900000 ;
        RECT 10.780000 38.140000 10.980000 38.340000 ;
        RECT 10.780000 38.580000 10.980000 38.780000 ;
        RECT 10.780000 39.020000 10.980000 39.220000 ;
        RECT 10.780000 39.460000 10.980000 39.660000 ;
        RECT 10.780000 39.900000 10.980000 40.100000 ;
        RECT 11.145000 51.715000 11.345000 51.915000 ;
        RECT 11.145000 52.135000 11.345000 52.335000 ;
        RECT 11.145000 52.555000 11.345000 52.755000 ;
        RECT 11.150000 47.800000 11.350000 48.000000 ;
        RECT 11.150000 56.470000 11.350000 56.670000 ;
        RECT 11.185000 36.820000 11.385000 37.020000 ;
        RECT 11.185000 37.260000 11.385000 37.460000 ;
        RECT 11.185000 37.700000 11.385000 37.900000 ;
        RECT 11.185000 38.140000 11.385000 38.340000 ;
        RECT 11.185000 38.580000 11.385000 38.780000 ;
        RECT 11.185000 39.020000 11.385000 39.220000 ;
        RECT 11.185000 39.460000 11.385000 39.660000 ;
        RECT 11.185000 39.900000 11.385000 40.100000 ;
        RECT 11.550000 51.715000 11.750000 51.915000 ;
        RECT 11.550000 52.135000 11.750000 52.335000 ;
        RECT 11.550000 52.555000 11.750000 52.755000 ;
        RECT 11.555000 47.800000 11.755000 48.000000 ;
        RECT 11.555000 56.470000 11.755000 56.670000 ;
        RECT 11.590000 36.820000 11.790000 37.020000 ;
        RECT 11.590000 37.260000 11.790000 37.460000 ;
        RECT 11.590000 37.700000 11.790000 37.900000 ;
        RECT 11.590000 38.140000 11.790000 38.340000 ;
        RECT 11.590000 38.580000 11.790000 38.780000 ;
        RECT 11.590000 39.020000 11.790000 39.220000 ;
        RECT 11.590000 39.460000 11.790000 39.660000 ;
        RECT 11.590000 39.900000 11.790000 40.100000 ;
        RECT 11.955000 51.715000 12.155000 51.915000 ;
        RECT 11.955000 52.135000 12.155000 52.335000 ;
        RECT 11.955000 52.555000 12.155000 52.755000 ;
        RECT 11.960000 47.800000 12.160000 48.000000 ;
        RECT 11.960000 56.470000 12.160000 56.670000 ;
        RECT 11.995000 36.820000 12.195000 37.020000 ;
        RECT 11.995000 37.260000 12.195000 37.460000 ;
        RECT 11.995000 37.700000 12.195000 37.900000 ;
        RECT 11.995000 38.140000 12.195000 38.340000 ;
        RECT 11.995000 38.580000 12.195000 38.780000 ;
        RECT 11.995000 39.020000 12.195000 39.220000 ;
        RECT 11.995000 39.460000 12.195000 39.660000 ;
        RECT 11.995000 39.900000 12.195000 40.100000 ;
        RECT 12.360000 51.715000 12.560000 51.915000 ;
        RECT 12.360000 52.135000 12.560000 52.335000 ;
        RECT 12.360000 52.555000 12.560000 52.755000 ;
        RECT 12.365000 47.800000 12.565000 48.000000 ;
        RECT 12.365000 56.470000 12.565000 56.670000 ;
        RECT 12.400000 36.820000 12.600000 37.020000 ;
        RECT 12.400000 37.260000 12.600000 37.460000 ;
        RECT 12.400000 37.700000 12.600000 37.900000 ;
        RECT 12.400000 38.140000 12.600000 38.340000 ;
        RECT 12.400000 38.580000 12.600000 38.780000 ;
        RECT 12.400000 39.020000 12.600000 39.220000 ;
        RECT 12.400000 39.460000 12.600000 39.660000 ;
        RECT 12.400000 39.900000 12.600000 40.100000 ;
        RECT 12.765000 51.715000 12.965000 51.915000 ;
        RECT 12.765000 52.135000 12.965000 52.335000 ;
        RECT 12.765000 52.555000 12.965000 52.755000 ;
        RECT 12.770000 47.800000 12.970000 48.000000 ;
        RECT 12.770000 56.470000 12.970000 56.670000 ;
        RECT 12.805000 36.820000 13.005000 37.020000 ;
        RECT 12.805000 37.260000 13.005000 37.460000 ;
        RECT 12.805000 37.700000 13.005000 37.900000 ;
        RECT 12.805000 38.140000 13.005000 38.340000 ;
        RECT 12.805000 38.580000 13.005000 38.780000 ;
        RECT 12.805000 39.020000 13.005000 39.220000 ;
        RECT 12.805000 39.460000 13.005000 39.660000 ;
        RECT 12.805000 39.900000 13.005000 40.100000 ;
        RECT 13.170000 51.715000 13.370000 51.915000 ;
        RECT 13.170000 52.135000 13.370000 52.335000 ;
        RECT 13.170000 52.555000 13.370000 52.755000 ;
        RECT 13.175000 47.800000 13.375000 48.000000 ;
        RECT 13.175000 56.470000 13.375000 56.670000 ;
        RECT 13.210000 36.820000 13.410000 37.020000 ;
        RECT 13.210000 37.260000 13.410000 37.460000 ;
        RECT 13.210000 37.700000 13.410000 37.900000 ;
        RECT 13.210000 38.140000 13.410000 38.340000 ;
        RECT 13.210000 38.580000 13.410000 38.780000 ;
        RECT 13.210000 39.020000 13.410000 39.220000 ;
        RECT 13.210000 39.460000 13.410000 39.660000 ;
        RECT 13.210000 39.900000 13.410000 40.100000 ;
        RECT 13.575000 51.715000 13.775000 51.915000 ;
        RECT 13.575000 52.135000 13.775000 52.335000 ;
        RECT 13.575000 52.555000 13.775000 52.755000 ;
        RECT 13.580000 47.800000 13.780000 48.000000 ;
        RECT 13.580000 56.470000 13.780000 56.670000 ;
        RECT 13.615000 36.820000 13.815000 37.020000 ;
        RECT 13.615000 37.260000 13.815000 37.460000 ;
        RECT 13.615000 37.700000 13.815000 37.900000 ;
        RECT 13.615000 38.140000 13.815000 38.340000 ;
        RECT 13.615000 38.580000 13.815000 38.780000 ;
        RECT 13.615000 39.020000 13.815000 39.220000 ;
        RECT 13.615000 39.460000 13.815000 39.660000 ;
        RECT 13.615000 39.900000 13.815000 40.100000 ;
        RECT 13.980000 51.715000 14.180000 51.915000 ;
        RECT 13.980000 52.135000 14.180000 52.335000 ;
        RECT 13.980000 52.555000 14.180000 52.755000 ;
        RECT 13.985000 47.800000 14.185000 48.000000 ;
        RECT 13.985000 56.470000 14.185000 56.670000 ;
        RECT 14.020000 36.820000 14.220000 37.020000 ;
        RECT 14.020000 37.260000 14.220000 37.460000 ;
        RECT 14.020000 37.700000 14.220000 37.900000 ;
        RECT 14.020000 38.140000 14.220000 38.340000 ;
        RECT 14.020000 38.580000 14.220000 38.780000 ;
        RECT 14.020000 39.020000 14.220000 39.220000 ;
        RECT 14.020000 39.460000 14.220000 39.660000 ;
        RECT 14.020000 39.900000 14.220000 40.100000 ;
        RECT 14.385000 51.715000 14.585000 51.915000 ;
        RECT 14.385000 52.135000 14.585000 52.335000 ;
        RECT 14.385000 52.555000 14.585000 52.755000 ;
        RECT 14.390000 47.800000 14.590000 48.000000 ;
        RECT 14.390000 56.470000 14.590000 56.670000 ;
        RECT 14.425000 36.820000 14.625000 37.020000 ;
        RECT 14.425000 37.260000 14.625000 37.460000 ;
        RECT 14.425000 37.700000 14.625000 37.900000 ;
        RECT 14.425000 38.140000 14.625000 38.340000 ;
        RECT 14.425000 38.580000 14.625000 38.780000 ;
        RECT 14.425000 39.020000 14.625000 39.220000 ;
        RECT 14.425000 39.460000 14.625000 39.660000 ;
        RECT 14.425000 39.900000 14.625000 40.100000 ;
        RECT 14.790000 51.715000 14.990000 51.915000 ;
        RECT 14.790000 52.135000 14.990000 52.335000 ;
        RECT 14.790000 52.555000 14.990000 52.755000 ;
        RECT 14.795000 47.800000 14.995000 48.000000 ;
        RECT 14.795000 56.470000 14.995000 56.670000 ;
        RECT 14.830000 36.820000 15.030000 37.020000 ;
        RECT 14.830000 37.260000 15.030000 37.460000 ;
        RECT 14.830000 37.700000 15.030000 37.900000 ;
        RECT 14.830000 38.140000 15.030000 38.340000 ;
        RECT 14.830000 38.580000 15.030000 38.780000 ;
        RECT 14.830000 39.020000 15.030000 39.220000 ;
        RECT 14.830000 39.460000 15.030000 39.660000 ;
        RECT 14.830000 39.900000 15.030000 40.100000 ;
        RECT 15.195000 51.715000 15.395000 51.915000 ;
        RECT 15.195000 52.135000 15.395000 52.335000 ;
        RECT 15.195000 52.555000 15.395000 52.755000 ;
        RECT 15.200000 47.800000 15.400000 48.000000 ;
        RECT 15.200000 56.470000 15.400000 56.670000 ;
        RECT 15.235000 36.820000 15.435000 37.020000 ;
        RECT 15.235000 37.260000 15.435000 37.460000 ;
        RECT 15.235000 37.700000 15.435000 37.900000 ;
        RECT 15.235000 38.140000 15.435000 38.340000 ;
        RECT 15.235000 38.580000 15.435000 38.780000 ;
        RECT 15.235000 39.020000 15.435000 39.220000 ;
        RECT 15.235000 39.460000 15.435000 39.660000 ;
        RECT 15.235000 39.900000 15.435000 40.100000 ;
        RECT 15.600000 51.715000 15.800000 51.915000 ;
        RECT 15.600000 52.135000 15.800000 52.335000 ;
        RECT 15.600000 52.555000 15.800000 52.755000 ;
        RECT 15.605000 47.800000 15.805000 48.000000 ;
        RECT 15.605000 56.470000 15.805000 56.670000 ;
        RECT 15.640000 36.820000 15.840000 37.020000 ;
        RECT 15.640000 37.260000 15.840000 37.460000 ;
        RECT 15.640000 37.700000 15.840000 37.900000 ;
        RECT 15.640000 38.140000 15.840000 38.340000 ;
        RECT 15.640000 38.580000 15.840000 38.780000 ;
        RECT 15.640000 39.020000 15.840000 39.220000 ;
        RECT 15.640000 39.460000 15.840000 39.660000 ;
        RECT 15.640000 39.900000 15.840000 40.100000 ;
        RECT 16.005000 51.715000 16.205000 51.915000 ;
        RECT 16.005000 52.135000 16.205000 52.335000 ;
        RECT 16.005000 52.555000 16.205000 52.755000 ;
        RECT 16.010000 47.800000 16.210000 48.000000 ;
        RECT 16.010000 56.470000 16.210000 56.670000 ;
        RECT 16.045000 36.820000 16.245000 37.020000 ;
        RECT 16.045000 37.260000 16.245000 37.460000 ;
        RECT 16.045000 37.700000 16.245000 37.900000 ;
        RECT 16.045000 38.140000 16.245000 38.340000 ;
        RECT 16.045000 38.580000 16.245000 38.780000 ;
        RECT 16.045000 39.020000 16.245000 39.220000 ;
        RECT 16.045000 39.460000 16.245000 39.660000 ;
        RECT 16.045000 39.900000 16.245000 40.100000 ;
        RECT 16.410000 51.715000 16.610000 51.915000 ;
        RECT 16.410000 52.135000 16.610000 52.335000 ;
        RECT 16.410000 52.555000 16.610000 52.755000 ;
        RECT 16.415000 47.800000 16.615000 48.000000 ;
        RECT 16.415000 56.470000 16.615000 56.670000 ;
        RECT 16.450000 36.820000 16.650000 37.020000 ;
        RECT 16.450000 37.260000 16.650000 37.460000 ;
        RECT 16.450000 37.700000 16.650000 37.900000 ;
        RECT 16.450000 38.140000 16.650000 38.340000 ;
        RECT 16.450000 38.580000 16.650000 38.780000 ;
        RECT 16.450000 39.020000 16.650000 39.220000 ;
        RECT 16.450000 39.460000 16.650000 39.660000 ;
        RECT 16.450000 39.900000 16.650000 40.100000 ;
        RECT 16.815000 51.715000 17.015000 51.915000 ;
        RECT 16.815000 52.135000 17.015000 52.335000 ;
        RECT 16.815000 52.555000 17.015000 52.755000 ;
        RECT 16.820000 47.800000 17.020000 48.000000 ;
        RECT 16.820000 56.470000 17.020000 56.670000 ;
        RECT 16.855000 36.820000 17.055000 37.020000 ;
        RECT 16.855000 37.260000 17.055000 37.460000 ;
        RECT 16.855000 37.700000 17.055000 37.900000 ;
        RECT 16.855000 38.140000 17.055000 38.340000 ;
        RECT 16.855000 38.580000 17.055000 38.780000 ;
        RECT 16.855000 39.020000 17.055000 39.220000 ;
        RECT 16.855000 39.460000 17.055000 39.660000 ;
        RECT 16.855000 39.900000 17.055000 40.100000 ;
        RECT 17.220000 51.715000 17.420000 51.915000 ;
        RECT 17.220000 52.135000 17.420000 52.335000 ;
        RECT 17.220000 52.555000 17.420000 52.755000 ;
        RECT 17.225000 47.800000 17.425000 48.000000 ;
        RECT 17.225000 56.470000 17.425000 56.670000 ;
        RECT 17.260000 36.820000 17.460000 37.020000 ;
        RECT 17.260000 37.260000 17.460000 37.460000 ;
        RECT 17.260000 37.700000 17.460000 37.900000 ;
        RECT 17.260000 38.140000 17.460000 38.340000 ;
        RECT 17.260000 38.580000 17.460000 38.780000 ;
        RECT 17.260000 39.020000 17.460000 39.220000 ;
        RECT 17.260000 39.460000 17.460000 39.660000 ;
        RECT 17.260000 39.900000 17.460000 40.100000 ;
        RECT 17.625000 51.715000 17.825000 51.915000 ;
        RECT 17.625000 52.135000 17.825000 52.335000 ;
        RECT 17.625000 52.555000 17.825000 52.755000 ;
        RECT 17.630000 47.800000 17.830000 48.000000 ;
        RECT 17.630000 56.470000 17.830000 56.670000 ;
        RECT 17.665000 36.820000 17.865000 37.020000 ;
        RECT 17.665000 37.260000 17.865000 37.460000 ;
        RECT 17.665000 37.700000 17.865000 37.900000 ;
        RECT 17.665000 38.140000 17.865000 38.340000 ;
        RECT 17.665000 38.580000 17.865000 38.780000 ;
        RECT 17.665000 39.020000 17.865000 39.220000 ;
        RECT 17.665000 39.460000 17.865000 39.660000 ;
        RECT 17.665000 39.900000 17.865000 40.100000 ;
        RECT 18.030000 51.715000 18.230000 51.915000 ;
        RECT 18.030000 52.135000 18.230000 52.335000 ;
        RECT 18.030000 52.555000 18.230000 52.755000 ;
        RECT 18.035000 47.800000 18.235000 48.000000 ;
        RECT 18.035000 56.470000 18.235000 56.670000 ;
        RECT 18.070000 36.820000 18.270000 37.020000 ;
        RECT 18.070000 37.260000 18.270000 37.460000 ;
        RECT 18.070000 37.700000 18.270000 37.900000 ;
        RECT 18.070000 38.140000 18.270000 38.340000 ;
        RECT 18.070000 38.580000 18.270000 38.780000 ;
        RECT 18.070000 39.020000 18.270000 39.220000 ;
        RECT 18.070000 39.460000 18.270000 39.660000 ;
        RECT 18.070000 39.900000 18.270000 40.100000 ;
        RECT 18.435000 51.715000 18.635000 51.915000 ;
        RECT 18.435000 52.135000 18.635000 52.335000 ;
        RECT 18.435000 52.555000 18.635000 52.755000 ;
        RECT 18.440000 47.800000 18.640000 48.000000 ;
        RECT 18.440000 56.470000 18.640000 56.670000 ;
        RECT 18.475000 36.820000 18.675000 37.020000 ;
        RECT 18.475000 37.260000 18.675000 37.460000 ;
        RECT 18.475000 37.700000 18.675000 37.900000 ;
        RECT 18.475000 38.140000 18.675000 38.340000 ;
        RECT 18.475000 38.580000 18.675000 38.780000 ;
        RECT 18.475000 39.020000 18.675000 39.220000 ;
        RECT 18.475000 39.460000 18.675000 39.660000 ;
        RECT 18.475000 39.900000 18.675000 40.100000 ;
        RECT 18.840000 51.715000 19.040000 51.915000 ;
        RECT 18.840000 52.135000 19.040000 52.335000 ;
        RECT 18.840000 52.555000 19.040000 52.755000 ;
        RECT 18.845000 47.800000 19.045000 48.000000 ;
        RECT 18.845000 56.470000 19.045000 56.670000 ;
        RECT 18.880000 36.820000 19.080000 37.020000 ;
        RECT 18.880000 37.260000 19.080000 37.460000 ;
        RECT 18.880000 37.700000 19.080000 37.900000 ;
        RECT 18.880000 38.140000 19.080000 38.340000 ;
        RECT 18.880000 38.580000 19.080000 38.780000 ;
        RECT 18.880000 39.020000 19.080000 39.220000 ;
        RECT 18.880000 39.460000 19.080000 39.660000 ;
        RECT 18.880000 39.900000 19.080000 40.100000 ;
        RECT 19.245000 51.715000 19.445000 51.915000 ;
        RECT 19.245000 52.135000 19.445000 52.335000 ;
        RECT 19.245000 52.555000 19.445000 52.755000 ;
        RECT 19.250000 47.800000 19.450000 48.000000 ;
        RECT 19.250000 56.470000 19.450000 56.670000 ;
        RECT 19.285000 36.820000 19.485000 37.020000 ;
        RECT 19.285000 37.260000 19.485000 37.460000 ;
        RECT 19.285000 37.700000 19.485000 37.900000 ;
        RECT 19.285000 38.140000 19.485000 38.340000 ;
        RECT 19.285000 38.580000 19.485000 38.780000 ;
        RECT 19.285000 39.020000 19.485000 39.220000 ;
        RECT 19.285000 39.460000 19.485000 39.660000 ;
        RECT 19.285000 39.900000 19.485000 40.100000 ;
        RECT 19.650000 51.715000 19.850000 51.915000 ;
        RECT 19.650000 52.135000 19.850000 52.335000 ;
        RECT 19.650000 52.555000 19.850000 52.755000 ;
        RECT 19.655000 47.800000 19.855000 48.000000 ;
        RECT 19.655000 56.470000 19.855000 56.670000 ;
        RECT 19.690000 36.820000 19.890000 37.020000 ;
        RECT 19.690000 37.260000 19.890000 37.460000 ;
        RECT 19.690000 37.700000 19.890000 37.900000 ;
        RECT 19.690000 38.140000 19.890000 38.340000 ;
        RECT 19.690000 38.580000 19.890000 38.780000 ;
        RECT 19.690000 39.020000 19.890000 39.220000 ;
        RECT 19.690000 39.460000 19.890000 39.660000 ;
        RECT 19.690000 39.900000 19.890000 40.100000 ;
        RECT 20.055000 51.715000 20.255000 51.915000 ;
        RECT 20.055000 52.135000 20.255000 52.335000 ;
        RECT 20.055000 52.555000 20.255000 52.755000 ;
        RECT 20.060000 47.800000 20.260000 48.000000 ;
        RECT 20.060000 56.470000 20.260000 56.670000 ;
        RECT 20.095000 36.820000 20.295000 37.020000 ;
        RECT 20.095000 37.260000 20.295000 37.460000 ;
        RECT 20.095000 37.700000 20.295000 37.900000 ;
        RECT 20.095000 38.140000 20.295000 38.340000 ;
        RECT 20.095000 38.580000 20.295000 38.780000 ;
        RECT 20.095000 39.020000 20.295000 39.220000 ;
        RECT 20.095000 39.460000 20.295000 39.660000 ;
        RECT 20.095000 39.900000 20.295000 40.100000 ;
        RECT 20.460000 51.715000 20.660000 51.915000 ;
        RECT 20.460000 52.135000 20.660000 52.335000 ;
        RECT 20.460000 52.555000 20.660000 52.755000 ;
        RECT 20.465000 47.800000 20.665000 48.000000 ;
        RECT 20.465000 56.470000 20.665000 56.670000 ;
        RECT 20.500000 36.820000 20.700000 37.020000 ;
        RECT 20.500000 37.260000 20.700000 37.460000 ;
        RECT 20.500000 37.700000 20.700000 37.900000 ;
        RECT 20.500000 38.140000 20.700000 38.340000 ;
        RECT 20.500000 38.580000 20.700000 38.780000 ;
        RECT 20.500000 39.020000 20.700000 39.220000 ;
        RECT 20.500000 39.460000 20.700000 39.660000 ;
        RECT 20.500000 39.900000 20.700000 40.100000 ;
        RECT 20.865000 51.715000 21.065000 51.915000 ;
        RECT 20.865000 52.135000 21.065000 52.335000 ;
        RECT 20.865000 52.555000 21.065000 52.755000 ;
        RECT 20.870000 47.800000 21.070000 48.000000 ;
        RECT 20.870000 56.470000 21.070000 56.670000 ;
        RECT 20.905000 36.820000 21.105000 37.020000 ;
        RECT 20.905000 37.260000 21.105000 37.460000 ;
        RECT 20.905000 37.700000 21.105000 37.900000 ;
        RECT 20.905000 38.140000 21.105000 38.340000 ;
        RECT 20.905000 38.580000 21.105000 38.780000 ;
        RECT 20.905000 39.020000 21.105000 39.220000 ;
        RECT 20.905000 39.460000 21.105000 39.660000 ;
        RECT 20.905000 39.900000 21.105000 40.100000 ;
        RECT 21.270000 51.715000 21.470000 51.915000 ;
        RECT 21.270000 52.135000 21.470000 52.335000 ;
        RECT 21.270000 52.555000 21.470000 52.755000 ;
        RECT 21.275000 47.800000 21.475000 48.000000 ;
        RECT 21.275000 56.470000 21.475000 56.670000 ;
        RECT 21.305000 36.820000 21.505000 37.020000 ;
        RECT 21.305000 37.260000 21.505000 37.460000 ;
        RECT 21.305000 37.700000 21.505000 37.900000 ;
        RECT 21.305000 38.140000 21.505000 38.340000 ;
        RECT 21.305000 38.580000 21.505000 38.780000 ;
        RECT 21.305000 39.020000 21.505000 39.220000 ;
        RECT 21.305000 39.460000 21.505000 39.660000 ;
        RECT 21.305000 39.900000 21.505000 40.100000 ;
        RECT 21.675000 51.715000 21.875000 51.915000 ;
        RECT 21.675000 52.135000 21.875000 52.335000 ;
        RECT 21.675000 52.555000 21.875000 52.755000 ;
        RECT 21.680000 47.800000 21.880000 48.000000 ;
        RECT 21.680000 56.470000 21.880000 56.670000 ;
        RECT 21.705000 36.820000 21.905000 37.020000 ;
        RECT 21.705000 37.260000 21.905000 37.460000 ;
        RECT 21.705000 37.700000 21.905000 37.900000 ;
        RECT 21.705000 38.140000 21.905000 38.340000 ;
        RECT 21.705000 38.580000 21.905000 38.780000 ;
        RECT 21.705000 39.020000 21.905000 39.220000 ;
        RECT 21.705000 39.460000 21.905000 39.660000 ;
        RECT 21.705000 39.900000 21.905000 40.100000 ;
        RECT 22.080000 51.715000 22.280000 51.915000 ;
        RECT 22.080000 52.135000 22.280000 52.335000 ;
        RECT 22.080000 52.555000 22.280000 52.755000 ;
        RECT 22.085000 47.800000 22.285000 48.000000 ;
        RECT 22.085000 56.470000 22.285000 56.670000 ;
        RECT 22.105000 36.820000 22.305000 37.020000 ;
        RECT 22.105000 37.260000 22.305000 37.460000 ;
        RECT 22.105000 37.700000 22.305000 37.900000 ;
        RECT 22.105000 38.140000 22.305000 38.340000 ;
        RECT 22.105000 38.580000 22.305000 38.780000 ;
        RECT 22.105000 39.020000 22.305000 39.220000 ;
        RECT 22.105000 39.460000 22.305000 39.660000 ;
        RECT 22.105000 39.900000 22.305000 40.100000 ;
        RECT 22.485000 51.715000 22.685000 51.915000 ;
        RECT 22.485000 52.135000 22.685000 52.335000 ;
        RECT 22.485000 52.555000 22.685000 52.755000 ;
        RECT 22.490000 47.800000 22.690000 48.000000 ;
        RECT 22.490000 56.470000 22.690000 56.670000 ;
        RECT 22.505000 36.820000 22.705000 37.020000 ;
        RECT 22.505000 37.260000 22.705000 37.460000 ;
        RECT 22.505000 37.700000 22.705000 37.900000 ;
        RECT 22.505000 38.140000 22.705000 38.340000 ;
        RECT 22.505000 38.580000 22.705000 38.780000 ;
        RECT 22.505000 39.020000 22.705000 39.220000 ;
        RECT 22.505000 39.460000 22.705000 39.660000 ;
        RECT 22.505000 39.900000 22.705000 40.100000 ;
        RECT 22.890000 51.715000 23.090000 51.915000 ;
        RECT 22.890000 52.135000 23.090000 52.335000 ;
        RECT 22.890000 52.555000 23.090000 52.755000 ;
        RECT 22.895000 47.800000 23.095000 48.000000 ;
        RECT 22.895000 56.470000 23.095000 56.670000 ;
        RECT 22.905000 36.820000 23.105000 37.020000 ;
        RECT 22.905000 37.260000 23.105000 37.460000 ;
        RECT 22.905000 37.700000 23.105000 37.900000 ;
        RECT 22.905000 38.140000 23.105000 38.340000 ;
        RECT 22.905000 38.580000 23.105000 38.780000 ;
        RECT 22.905000 39.020000 23.105000 39.220000 ;
        RECT 22.905000 39.460000 23.105000 39.660000 ;
        RECT 22.905000 39.900000 23.105000 40.100000 ;
        RECT 23.295000 51.715000 23.495000 51.915000 ;
        RECT 23.295000 52.135000 23.495000 52.335000 ;
        RECT 23.295000 52.555000 23.495000 52.755000 ;
        RECT 23.300000 47.800000 23.500000 48.000000 ;
        RECT 23.300000 56.470000 23.500000 56.670000 ;
        RECT 23.305000 36.820000 23.505000 37.020000 ;
        RECT 23.305000 37.260000 23.505000 37.460000 ;
        RECT 23.305000 37.700000 23.505000 37.900000 ;
        RECT 23.305000 38.140000 23.505000 38.340000 ;
        RECT 23.305000 38.580000 23.505000 38.780000 ;
        RECT 23.305000 39.020000 23.505000 39.220000 ;
        RECT 23.305000 39.460000 23.505000 39.660000 ;
        RECT 23.305000 39.900000 23.505000 40.100000 ;
        RECT 23.700000 51.715000 23.900000 51.915000 ;
        RECT 23.700000 52.135000 23.900000 52.335000 ;
        RECT 23.700000 52.555000 23.900000 52.755000 ;
        RECT 23.705000 36.820000 23.905000 37.020000 ;
        RECT 23.705000 37.260000 23.905000 37.460000 ;
        RECT 23.705000 37.700000 23.905000 37.900000 ;
        RECT 23.705000 38.140000 23.905000 38.340000 ;
        RECT 23.705000 38.580000 23.905000 38.780000 ;
        RECT 23.705000 39.020000 23.905000 39.220000 ;
        RECT 23.705000 39.460000 23.905000 39.660000 ;
        RECT 23.705000 39.900000 23.905000 40.100000 ;
        RECT 23.705000 47.800000 23.905000 48.000000 ;
        RECT 23.705000 56.470000 23.905000 56.670000 ;
        RECT 24.105000 36.820000 24.305000 37.020000 ;
        RECT 24.105000 37.260000 24.305000 37.460000 ;
        RECT 24.105000 37.700000 24.305000 37.900000 ;
        RECT 24.105000 38.140000 24.305000 38.340000 ;
        RECT 24.105000 38.580000 24.305000 38.780000 ;
        RECT 24.105000 39.020000 24.305000 39.220000 ;
        RECT 24.105000 39.460000 24.305000 39.660000 ;
        RECT 24.105000 39.900000 24.305000 40.100000 ;
        RECT 24.105000 47.800000 24.305000 48.000000 ;
        RECT 24.105000 51.715000 24.305000 51.915000 ;
        RECT 24.105000 52.135000 24.305000 52.335000 ;
        RECT 24.105000 52.555000 24.305000 52.755000 ;
        RECT 24.105000 56.470000 24.305000 56.670000 ;
        RECT 50.480000 36.820000 50.680000 37.020000 ;
        RECT 50.480000 37.260000 50.680000 37.460000 ;
        RECT 50.480000 37.700000 50.680000 37.900000 ;
        RECT 50.480000 38.140000 50.680000 38.340000 ;
        RECT 50.480000 38.580000 50.680000 38.780000 ;
        RECT 50.480000 39.020000 50.680000 39.220000 ;
        RECT 50.480000 39.460000 50.680000 39.660000 ;
        RECT 50.480000 39.900000 50.680000 40.100000 ;
        RECT 50.480000 47.800000 50.680000 48.000000 ;
        RECT 50.480000 51.715000 50.680000 51.915000 ;
        RECT 50.480000 52.135000 50.680000 52.335000 ;
        RECT 50.480000 52.555000 50.680000 52.755000 ;
        RECT 50.480000 56.470000 50.680000 56.670000 ;
        RECT 50.885000 47.800000 51.085000 48.000000 ;
        RECT 50.885000 56.470000 51.085000 56.670000 ;
        RECT 50.890000 36.820000 51.090000 37.020000 ;
        RECT 50.890000 37.260000 51.090000 37.460000 ;
        RECT 50.890000 37.700000 51.090000 37.900000 ;
        RECT 50.890000 38.140000 51.090000 38.340000 ;
        RECT 50.890000 38.580000 51.090000 38.780000 ;
        RECT 50.890000 39.020000 51.090000 39.220000 ;
        RECT 50.890000 39.460000 51.090000 39.660000 ;
        RECT 50.890000 39.900000 51.090000 40.100000 ;
        RECT 50.890000 51.715000 51.090000 51.915000 ;
        RECT 50.890000 52.135000 51.090000 52.335000 ;
        RECT 50.890000 52.555000 51.090000 52.755000 ;
        RECT 51.290000 47.800000 51.490000 48.000000 ;
        RECT 51.290000 56.470000 51.490000 56.670000 ;
        RECT 51.300000 36.820000 51.500000 37.020000 ;
        RECT 51.300000 37.260000 51.500000 37.460000 ;
        RECT 51.300000 37.700000 51.500000 37.900000 ;
        RECT 51.300000 38.140000 51.500000 38.340000 ;
        RECT 51.300000 38.580000 51.500000 38.780000 ;
        RECT 51.300000 39.020000 51.500000 39.220000 ;
        RECT 51.300000 39.460000 51.500000 39.660000 ;
        RECT 51.300000 39.900000 51.500000 40.100000 ;
        RECT 51.300000 51.715000 51.500000 51.915000 ;
        RECT 51.300000 52.135000 51.500000 52.335000 ;
        RECT 51.300000 52.555000 51.500000 52.755000 ;
        RECT 51.695000 47.800000 51.895000 48.000000 ;
        RECT 51.695000 56.470000 51.895000 56.670000 ;
        RECT 51.710000 36.820000 51.910000 37.020000 ;
        RECT 51.710000 37.260000 51.910000 37.460000 ;
        RECT 51.710000 37.700000 51.910000 37.900000 ;
        RECT 51.710000 38.140000 51.910000 38.340000 ;
        RECT 51.710000 38.580000 51.910000 38.780000 ;
        RECT 51.710000 39.020000 51.910000 39.220000 ;
        RECT 51.710000 39.460000 51.910000 39.660000 ;
        RECT 51.710000 39.900000 51.910000 40.100000 ;
        RECT 51.710000 51.715000 51.910000 51.915000 ;
        RECT 51.710000 52.135000 51.910000 52.335000 ;
        RECT 51.710000 52.555000 51.910000 52.755000 ;
        RECT 52.100000 47.800000 52.300000 48.000000 ;
        RECT 52.100000 56.470000 52.300000 56.670000 ;
        RECT 52.120000 36.820000 52.320000 37.020000 ;
        RECT 52.120000 37.260000 52.320000 37.460000 ;
        RECT 52.120000 37.700000 52.320000 37.900000 ;
        RECT 52.120000 38.140000 52.320000 38.340000 ;
        RECT 52.120000 38.580000 52.320000 38.780000 ;
        RECT 52.120000 39.020000 52.320000 39.220000 ;
        RECT 52.120000 39.460000 52.320000 39.660000 ;
        RECT 52.120000 39.900000 52.320000 40.100000 ;
        RECT 52.120000 51.715000 52.320000 51.915000 ;
        RECT 52.120000 52.135000 52.320000 52.335000 ;
        RECT 52.120000 52.555000 52.320000 52.755000 ;
        RECT 52.505000 47.800000 52.705000 48.000000 ;
        RECT 52.505000 56.470000 52.705000 56.670000 ;
        RECT 52.530000 36.820000 52.730000 37.020000 ;
        RECT 52.530000 37.260000 52.730000 37.460000 ;
        RECT 52.530000 37.700000 52.730000 37.900000 ;
        RECT 52.530000 38.140000 52.730000 38.340000 ;
        RECT 52.530000 38.580000 52.730000 38.780000 ;
        RECT 52.530000 39.020000 52.730000 39.220000 ;
        RECT 52.530000 39.460000 52.730000 39.660000 ;
        RECT 52.530000 39.900000 52.730000 40.100000 ;
        RECT 52.530000 51.715000 52.730000 51.915000 ;
        RECT 52.530000 52.135000 52.730000 52.335000 ;
        RECT 52.530000 52.555000 52.730000 52.755000 ;
        RECT 52.910000 47.800000 53.110000 48.000000 ;
        RECT 52.910000 56.470000 53.110000 56.670000 ;
        RECT 52.940000 36.820000 53.140000 37.020000 ;
        RECT 52.940000 37.260000 53.140000 37.460000 ;
        RECT 52.940000 37.700000 53.140000 37.900000 ;
        RECT 52.940000 38.140000 53.140000 38.340000 ;
        RECT 52.940000 38.580000 53.140000 38.780000 ;
        RECT 52.940000 39.020000 53.140000 39.220000 ;
        RECT 52.940000 39.460000 53.140000 39.660000 ;
        RECT 52.940000 39.900000 53.140000 40.100000 ;
        RECT 52.940000 51.715000 53.140000 51.915000 ;
        RECT 52.940000 52.135000 53.140000 52.335000 ;
        RECT 52.940000 52.555000 53.140000 52.755000 ;
        RECT 53.315000 47.800000 53.515000 48.000000 ;
        RECT 53.315000 56.470000 53.515000 56.670000 ;
        RECT 53.345000 36.820000 53.545000 37.020000 ;
        RECT 53.345000 37.260000 53.545000 37.460000 ;
        RECT 53.345000 37.700000 53.545000 37.900000 ;
        RECT 53.345000 38.140000 53.545000 38.340000 ;
        RECT 53.345000 38.580000 53.545000 38.780000 ;
        RECT 53.345000 39.020000 53.545000 39.220000 ;
        RECT 53.345000 39.460000 53.545000 39.660000 ;
        RECT 53.345000 39.900000 53.545000 40.100000 ;
        RECT 53.345000 51.715000 53.545000 51.915000 ;
        RECT 53.345000 52.135000 53.545000 52.335000 ;
        RECT 53.345000 52.555000 53.545000 52.755000 ;
        RECT 53.720000 47.800000 53.920000 48.000000 ;
        RECT 53.720000 56.470000 53.920000 56.670000 ;
        RECT 53.750000 36.820000 53.950000 37.020000 ;
        RECT 53.750000 37.260000 53.950000 37.460000 ;
        RECT 53.750000 37.700000 53.950000 37.900000 ;
        RECT 53.750000 38.140000 53.950000 38.340000 ;
        RECT 53.750000 38.580000 53.950000 38.780000 ;
        RECT 53.750000 39.020000 53.950000 39.220000 ;
        RECT 53.750000 39.460000 53.950000 39.660000 ;
        RECT 53.750000 39.900000 53.950000 40.100000 ;
        RECT 53.750000 51.715000 53.950000 51.915000 ;
        RECT 53.750000 52.135000 53.950000 52.335000 ;
        RECT 53.750000 52.555000 53.950000 52.755000 ;
        RECT 54.125000 47.800000 54.325000 48.000000 ;
        RECT 54.125000 56.470000 54.325000 56.670000 ;
        RECT 54.155000 36.820000 54.355000 37.020000 ;
        RECT 54.155000 37.260000 54.355000 37.460000 ;
        RECT 54.155000 37.700000 54.355000 37.900000 ;
        RECT 54.155000 38.140000 54.355000 38.340000 ;
        RECT 54.155000 38.580000 54.355000 38.780000 ;
        RECT 54.155000 39.020000 54.355000 39.220000 ;
        RECT 54.155000 39.460000 54.355000 39.660000 ;
        RECT 54.155000 39.900000 54.355000 40.100000 ;
        RECT 54.155000 51.715000 54.355000 51.915000 ;
        RECT 54.155000 52.135000 54.355000 52.335000 ;
        RECT 54.155000 52.555000 54.355000 52.755000 ;
        RECT 54.530000 47.800000 54.730000 48.000000 ;
        RECT 54.530000 56.470000 54.730000 56.670000 ;
        RECT 54.560000 36.820000 54.760000 37.020000 ;
        RECT 54.560000 37.260000 54.760000 37.460000 ;
        RECT 54.560000 37.700000 54.760000 37.900000 ;
        RECT 54.560000 38.140000 54.760000 38.340000 ;
        RECT 54.560000 38.580000 54.760000 38.780000 ;
        RECT 54.560000 39.020000 54.760000 39.220000 ;
        RECT 54.560000 39.460000 54.760000 39.660000 ;
        RECT 54.560000 39.900000 54.760000 40.100000 ;
        RECT 54.560000 51.715000 54.760000 51.915000 ;
        RECT 54.560000 52.135000 54.760000 52.335000 ;
        RECT 54.560000 52.555000 54.760000 52.755000 ;
        RECT 54.935000 47.800000 55.135000 48.000000 ;
        RECT 54.935000 56.470000 55.135000 56.670000 ;
        RECT 54.965000 36.820000 55.165000 37.020000 ;
        RECT 54.965000 37.260000 55.165000 37.460000 ;
        RECT 54.965000 37.700000 55.165000 37.900000 ;
        RECT 54.965000 38.140000 55.165000 38.340000 ;
        RECT 54.965000 38.580000 55.165000 38.780000 ;
        RECT 54.965000 39.020000 55.165000 39.220000 ;
        RECT 54.965000 39.460000 55.165000 39.660000 ;
        RECT 54.965000 39.900000 55.165000 40.100000 ;
        RECT 54.965000 51.715000 55.165000 51.915000 ;
        RECT 54.965000 52.135000 55.165000 52.335000 ;
        RECT 54.965000 52.555000 55.165000 52.755000 ;
        RECT 55.340000 47.800000 55.540000 48.000000 ;
        RECT 55.340000 56.470000 55.540000 56.670000 ;
        RECT 55.370000 36.820000 55.570000 37.020000 ;
        RECT 55.370000 37.260000 55.570000 37.460000 ;
        RECT 55.370000 37.700000 55.570000 37.900000 ;
        RECT 55.370000 38.140000 55.570000 38.340000 ;
        RECT 55.370000 38.580000 55.570000 38.780000 ;
        RECT 55.370000 39.020000 55.570000 39.220000 ;
        RECT 55.370000 39.460000 55.570000 39.660000 ;
        RECT 55.370000 39.900000 55.570000 40.100000 ;
        RECT 55.370000 51.715000 55.570000 51.915000 ;
        RECT 55.370000 52.135000 55.570000 52.335000 ;
        RECT 55.370000 52.555000 55.570000 52.755000 ;
        RECT 55.745000 47.800000 55.945000 48.000000 ;
        RECT 55.745000 56.470000 55.945000 56.670000 ;
        RECT 55.775000 36.820000 55.975000 37.020000 ;
        RECT 55.775000 37.260000 55.975000 37.460000 ;
        RECT 55.775000 37.700000 55.975000 37.900000 ;
        RECT 55.775000 38.140000 55.975000 38.340000 ;
        RECT 55.775000 38.580000 55.975000 38.780000 ;
        RECT 55.775000 39.020000 55.975000 39.220000 ;
        RECT 55.775000 39.460000 55.975000 39.660000 ;
        RECT 55.775000 39.900000 55.975000 40.100000 ;
        RECT 55.775000 51.715000 55.975000 51.915000 ;
        RECT 55.775000 52.135000 55.975000 52.335000 ;
        RECT 55.775000 52.555000 55.975000 52.755000 ;
        RECT 56.150000 47.800000 56.350000 48.000000 ;
        RECT 56.150000 56.470000 56.350000 56.670000 ;
        RECT 56.180000 36.820000 56.380000 37.020000 ;
        RECT 56.180000 37.260000 56.380000 37.460000 ;
        RECT 56.180000 37.700000 56.380000 37.900000 ;
        RECT 56.180000 38.140000 56.380000 38.340000 ;
        RECT 56.180000 38.580000 56.380000 38.780000 ;
        RECT 56.180000 39.020000 56.380000 39.220000 ;
        RECT 56.180000 39.460000 56.380000 39.660000 ;
        RECT 56.180000 39.900000 56.380000 40.100000 ;
        RECT 56.180000 51.715000 56.380000 51.915000 ;
        RECT 56.180000 52.135000 56.380000 52.335000 ;
        RECT 56.180000 52.555000 56.380000 52.755000 ;
        RECT 56.555000 47.800000 56.755000 48.000000 ;
        RECT 56.555000 56.470000 56.755000 56.670000 ;
        RECT 56.585000 36.820000 56.785000 37.020000 ;
        RECT 56.585000 37.260000 56.785000 37.460000 ;
        RECT 56.585000 37.700000 56.785000 37.900000 ;
        RECT 56.585000 38.140000 56.785000 38.340000 ;
        RECT 56.585000 38.580000 56.785000 38.780000 ;
        RECT 56.585000 39.020000 56.785000 39.220000 ;
        RECT 56.585000 39.460000 56.785000 39.660000 ;
        RECT 56.585000 39.900000 56.785000 40.100000 ;
        RECT 56.585000 51.715000 56.785000 51.915000 ;
        RECT 56.585000 52.135000 56.785000 52.335000 ;
        RECT 56.585000 52.555000 56.785000 52.755000 ;
        RECT 56.960000 47.800000 57.160000 48.000000 ;
        RECT 56.960000 56.470000 57.160000 56.670000 ;
        RECT 56.990000 36.820000 57.190000 37.020000 ;
        RECT 56.990000 37.260000 57.190000 37.460000 ;
        RECT 56.990000 37.700000 57.190000 37.900000 ;
        RECT 56.990000 38.140000 57.190000 38.340000 ;
        RECT 56.990000 38.580000 57.190000 38.780000 ;
        RECT 56.990000 39.020000 57.190000 39.220000 ;
        RECT 56.990000 39.460000 57.190000 39.660000 ;
        RECT 56.990000 39.900000 57.190000 40.100000 ;
        RECT 56.990000 51.715000 57.190000 51.915000 ;
        RECT 56.990000 52.135000 57.190000 52.335000 ;
        RECT 56.990000 52.555000 57.190000 52.755000 ;
        RECT 57.365000 47.800000 57.565000 48.000000 ;
        RECT 57.365000 56.470000 57.565000 56.670000 ;
        RECT 57.395000 36.820000 57.595000 37.020000 ;
        RECT 57.395000 37.260000 57.595000 37.460000 ;
        RECT 57.395000 37.700000 57.595000 37.900000 ;
        RECT 57.395000 38.140000 57.595000 38.340000 ;
        RECT 57.395000 38.580000 57.595000 38.780000 ;
        RECT 57.395000 39.020000 57.595000 39.220000 ;
        RECT 57.395000 39.460000 57.595000 39.660000 ;
        RECT 57.395000 39.900000 57.595000 40.100000 ;
        RECT 57.395000 51.715000 57.595000 51.915000 ;
        RECT 57.395000 52.135000 57.595000 52.335000 ;
        RECT 57.395000 52.555000 57.595000 52.755000 ;
        RECT 57.770000 47.800000 57.970000 48.000000 ;
        RECT 57.770000 56.470000 57.970000 56.670000 ;
        RECT 57.800000 36.820000 58.000000 37.020000 ;
        RECT 57.800000 37.260000 58.000000 37.460000 ;
        RECT 57.800000 37.700000 58.000000 37.900000 ;
        RECT 57.800000 38.140000 58.000000 38.340000 ;
        RECT 57.800000 38.580000 58.000000 38.780000 ;
        RECT 57.800000 39.020000 58.000000 39.220000 ;
        RECT 57.800000 39.460000 58.000000 39.660000 ;
        RECT 57.800000 39.900000 58.000000 40.100000 ;
        RECT 57.800000 51.715000 58.000000 51.915000 ;
        RECT 57.800000 52.135000 58.000000 52.335000 ;
        RECT 57.800000 52.555000 58.000000 52.755000 ;
        RECT 58.175000 47.800000 58.375000 48.000000 ;
        RECT 58.175000 56.470000 58.375000 56.670000 ;
        RECT 58.205000 36.820000 58.405000 37.020000 ;
        RECT 58.205000 37.260000 58.405000 37.460000 ;
        RECT 58.205000 37.700000 58.405000 37.900000 ;
        RECT 58.205000 38.140000 58.405000 38.340000 ;
        RECT 58.205000 38.580000 58.405000 38.780000 ;
        RECT 58.205000 39.020000 58.405000 39.220000 ;
        RECT 58.205000 39.460000 58.405000 39.660000 ;
        RECT 58.205000 39.900000 58.405000 40.100000 ;
        RECT 58.205000 51.715000 58.405000 51.915000 ;
        RECT 58.205000 52.135000 58.405000 52.335000 ;
        RECT 58.205000 52.555000 58.405000 52.755000 ;
        RECT 58.580000 47.800000 58.780000 48.000000 ;
        RECT 58.580000 56.470000 58.780000 56.670000 ;
        RECT 58.610000 36.820000 58.810000 37.020000 ;
        RECT 58.610000 37.260000 58.810000 37.460000 ;
        RECT 58.610000 37.700000 58.810000 37.900000 ;
        RECT 58.610000 38.140000 58.810000 38.340000 ;
        RECT 58.610000 38.580000 58.810000 38.780000 ;
        RECT 58.610000 39.020000 58.810000 39.220000 ;
        RECT 58.610000 39.460000 58.810000 39.660000 ;
        RECT 58.610000 39.900000 58.810000 40.100000 ;
        RECT 58.610000 51.715000 58.810000 51.915000 ;
        RECT 58.610000 52.135000 58.810000 52.335000 ;
        RECT 58.610000 52.555000 58.810000 52.755000 ;
        RECT 58.985000 47.800000 59.185000 48.000000 ;
        RECT 58.985000 56.470000 59.185000 56.670000 ;
        RECT 59.015000 36.820000 59.215000 37.020000 ;
        RECT 59.015000 37.260000 59.215000 37.460000 ;
        RECT 59.015000 37.700000 59.215000 37.900000 ;
        RECT 59.015000 38.140000 59.215000 38.340000 ;
        RECT 59.015000 38.580000 59.215000 38.780000 ;
        RECT 59.015000 39.020000 59.215000 39.220000 ;
        RECT 59.015000 39.460000 59.215000 39.660000 ;
        RECT 59.015000 39.900000 59.215000 40.100000 ;
        RECT 59.015000 51.715000 59.215000 51.915000 ;
        RECT 59.015000 52.135000 59.215000 52.335000 ;
        RECT 59.015000 52.555000 59.215000 52.755000 ;
        RECT 59.390000 47.800000 59.590000 48.000000 ;
        RECT 59.390000 56.470000 59.590000 56.670000 ;
        RECT 59.420000 36.820000 59.620000 37.020000 ;
        RECT 59.420000 37.260000 59.620000 37.460000 ;
        RECT 59.420000 37.700000 59.620000 37.900000 ;
        RECT 59.420000 38.140000 59.620000 38.340000 ;
        RECT 59.420000 38.580000 59.620000 38.780000 ;
        RECT 59.420000 39.020000 59.620000 39.220000 ;
        RECT 59.420000 39.460000 59.620000 39.660000 ;
        RECT 59.420000 39.900000 59.620000 40.100000 ;
        RECT 59.420000 51.715000 59.620000 51.915000 ;
        RECT 59.420000 52.135000 59.620000 52.335000 ;
        RECT 59.420000 52.555000 59.620000 52.755000 ;
        RECT 59.795000 47.800000 59.995000 48.000000 ;
        RECT 59.795000 56.470000 59.995000 56.670000 ;
        RECT 59.825000 36.820000 60.025000 37.020000 ;
        RECT 59.825000 37.260000 60.025000 37.460000 ;
        RECT 59.825000 37.700000 60.025000 37.900000 ;
        RECT 59.825000 38.140000 60.025000 38.340000 ;
        RECT 59.825000 38.580000 60.025000 38.780000 ;
        RECT 59.825000 39.020000 60.025000 39.220000 ;
        RECT 59.825000 39.460000 60.025000 39.660000 ;
        RECT 59.825000 39.900000 60.025000 40.100000 ;
        RECT 59.825000 51.715000 60.025000 51.915000 ;
        RECT 59.825000 52.135000 60.025000 52.335000 ;
        RECT 59.825000 52.555000 60.025000 52.755000 ;
        RECT 60.200000 47.800000 60.400000 48.000000 ;
        RECT 60.200000 56.470000 60.400000 56.670000 ;
        RECT 60.230000 36.820000 60.430000 37.020000 ;
        RECT 60.230000 37.260000 60.430000 37.460000 ;
        RECT 60.230000 37.700000 60.430000 37.900000 ;
        RECT 60.230000 38.140000 60.430000 38.340000 ;
        RECT 60.230000 38.580000 60.430000 38.780000 ;
        RECT 60.230000 39.020000 60.430000 39.220000 ;
        RECT 60.230000 39.460000 60.430000 39.660000 ;
        RECT 60.230000 39.900000 60.430000 40.100000 ;
        RECT 60.230000 51.715000 60.430000 51.915000 ;
        RECT 60.230000 52.135000 60.430000 52.335000 ;
        RECT 60.230000 52.555000 60.430000 52.755000 ;
        RECT 60.605000 47.800000 60.805000 48.000000 ;
        RECT 60.605000 56.470000 60.805000 56.670000 ;
        RECT 60.635000 36.820000 60.835000 37.020000 ;
        RECT 60.635000 37.260000 60.835000 37.460000 ;
        RECT 60.635000 37.700000 60.835000 37.900000 ;
        RECT 60.635000 38.140000 60.835000 38.340000 ;
        RECT 60.635000 38.580000 60.835000 38.780000 ;
        RECT 60.635000 39.020000 60.835000 39.220000 ;
        RECT 60.635000 39.460000 60.835000 39.660000 ;
        RECT 60.635000 39.900000 60.835000 40.100000 ;
        RECT 60.635000 51.715000 60.835000 51.915000 ;
        RECT 60.635000 52.135000 60.835000 52.335000 ;
        RECT 60.635000 52.555000 60.835000 52.755000 ;
        RECT 61.010000 47.800000 61.210000 48.000000 ;
        RECT 61.010000 56.470000 61.210000 56.670000 ;
        RECT 61.040000 36.820000 61.240000 37.020000 ;
        RECT 61.040000 37.260000 61.240000 37.460000 ;
        RECT 61.040000 37.700000 61.240000 37.900000 ;
        RECT 61.040000 38.140000 61.240000 38.340000 ;
        RECT 61.040000 38.580000 61.240000 38.780000 ;
        RECT 61.040000 39.020000 61.240000 39.220000 ;
        RECT 61.040000 39.460000 61.240000 39.660000 ;
        RECT 61.040000 39.900000 61.240000 40.100000 ;
        RECT 61.040000 51.715000 61.240000 51.915000 ;
        RECT 61.040000 52.135000 61.240000 52.335000 ;
        RECT 61.040000 52.555000 61.240000 52.755000 ;
        RECT 61.415000 47.800000 61.615000 48.000000 ;
        RECT 61.415000 56.470000 61.615000 56.670000 ;
        RECT 61.445000 36.820000 61.645000 37.020000 ;
        RECT 61.445000 37.260000 61.645000 37.460000 ;
        RECT 61.445000 37.700000 61.645000 37.900000 ;
        RECT 61.445000 38.140000 61.645000 38.340000 ;
        RECT 61.445000 38.580000 61.645000 38.780000 ;
        RECT 61.445000 39.020000 61.645000 39.220000 ;
        RECT 61.445000 39.460000 61.645000 39.660000 ;
        RECT 61.445000 39.900000 61.645000 40.100000 ;
        RECT 61.445000 51.715000 61.645000 51.915000 ;
        RECT 61.445000 52.135000 61.645000 52.335000 ;
        RECT 61.445000 52.555000 61.645000 52.755000 ;
        RECT 61.820000 47.800000 62.020000 48.000000 ;
        RECT 61.820000 56.470000 62.020000 56.670000 ;
        RECT 61.850000 36.820000 62.050000 37.020000 ;
        RECT 61.850000 37.260000 62.050000 37.460000 ;
        RECT 61.850000 37.700000 62.050000 37.900000 ;
        RECT 61.850000 38.140000 62.050000 38.340000 ;
        RECT 61.850000 38.580000 62.050000 38.780000 ;
        RECT 61.850000 39.020000 62.050000 39.220000 ;
        RECT 61.850000 39.460000 62.050000 39.660000 ;
        RECT 61.850000 39.900000 62.050000 40.100000 ;
        RECT 61.850000 51.715000 62.050000 51.915000 ;
        RECT 61.850000 52.135000 62.050000 52.335000 ;
        RECT 61.850000 52.555000 62.050000 52.755000 ;
        RECT 62.225000 47.800000 62.425000 48.000000 ;
        RECT 62.225000 56.470000 62.425000 56.670000 ;
        RECT 62.255000 36.820000 62.455000 37.020000 ;
        RECT 62.255000 37.260000 62.455000 37.460000 ;
        RECT 62.255000 37.700000 62.455000 37.900000 ;
        RECT 62.255000 38.140000 62.455000 38.340000 ;
        RECT 62.255000 38.580000 62.455000 38.780000 ;
        RECT 62.255000 39.020000 62.455000 39.220000 ;
        RECT 62.255000 39.460000 62.455000 39.660000 ;
        RECT 62.255000 39.900000 62.455000 40.100000 ;
        RECT 62.255000 51.715000 62.455000 51.915000 ;
        RECT 62.255000 52.135000 62.455000 52.335000 ;
        RECT 62.255000 52.555000 62.455000 52.755000 ;
        RECT 62.630000 47.800000 62.830000 48.000000 ;
        RECT 62.630000 56.470000 62.830000 56.670000 ;
        RECT 62.660000 36.820000 62.860000 37.020000 ;
        RECT 62.660000 37.260000 62.860000 37.460000 ;
        RECT 62.660000 37.700000 62.860000 37.900000 ;
        RECT 62.660000 38.140000 62.860000 38.340000 ;
        RECT 62.660000 38.580000 62.860000 38.780000 ;
        RECT 62.660000 39.020000 62.860000 39.220000 ;
        RECT 62.660000 39.460000 62.860000 39.660000 ;
        RECT 62.660000 39.900000 62.860000 40.100000 ;
        RECT 62.660000 51.715000 62.860000 51.915000 ;
        RECT 62.660000 52.135000 62.860000 52.335000 ;
        RECT 62.660000 52.555000 62.860000 52.755000 ;
        RECT 63.035000 47.800000 63.235000 48.000000 ;
        RECT 63.035000 56.470000 63.235000 56.670000 ;
        RECT 63.065000 36.820000 63.265000 37.020000 ;
        RECT 63.065000 37.260000 63.265000 37.460000 ;
        RECT 63.065000 37.700000 63.265000 37.900000 ;
        RECT 63.065000 38.140000 63.265000 38.340000 ;
        RECT 63.065000 38.580000 63.265000 38.780000 ;
        RECT 63.065000 39.020000 63.265000 39.220000 ;
        RECT 63.065000 39.460000 63.265000 39.660000 ;
        RECT 63.065000 39.900000 63.265000 40.100000 ;
        RECT 63.065000 51.715000 63.265000 51.915000 ;
        RECT 63.065000 52.135000 63.265000 52.335000 ;
        RECT 63.065000 52.555000 63.265000 52.755000 ;
        RECT 63.440000 47.800000 63.640000 48.000000 ;
        RECT 63.440000 56.470000 63.640000 56.670000 ;
        RECT 63.470000 36.820000 63.670000 37.020000 ;
        RECT 63.470000 37.260000 63.670000 37.460000 ;
        RECT 63.470000 37.700000 63.670000 37.900000 ;
        RECT 63.470000 38.140000 63.670000 38.340000 ;
        RECT 63.470000 38.580000 63.670000 38.780000 ;
        RECT 63.470000 39.020000 63.670000 39.220000 ;
        RECT 63.470000 39.460000 63.670000 39.660000 ;
        RECT 63.470000 39.900000 63.670000 40.100000 ;
        RECT 63.470000 51.715000 63.670000 51.915000 ;
        RECT 63.470000 52.135000 63.670000 52.335000 ;
        RECT 63.470000 52.555000 63.670000 52.755000 ;
        RECT 63.845000 47.800000 64.045000 48.000000 ;
        RECT 63.845000 56.470000 64.045000 56.670000 ;
        RECT 63.875000 36.820000 64.075000 37.020000 ;
        RECT 63.875000 37.260000 64.075000 37.460000 ;
        RECT 63.875000 37.700000 64.075000 37.900000 ;
        RECT 63.875000 38.140000 64.075000 38.340000 ;
        RECT 63.875000 38.580000 64.075000 38.780000 ;
        RECT 63.875000 39.020000 64.075000 39.220000 ;
        RECT 63.875000 39.460000 64.075000 39.660000 ;
        RECT 63.875000 39.900000 64.075000 40.100000 ;
        RECT 63.875000 51.715000 64.075000 51.915000 ;
        RECT 63.875000 52.135000 64.075000 52.335000 ;
        RECT 63.875000 52.555000 64.075000 52.755000 ;
        RECT 64.250000 47.800000 64.450000 48.000000 ;
        RECT 64.250000 56.470000 64.450000 56.670000 ;
        RECT 64.280000 36.820000 64.480000 37.020000 ;
        RECT 64.280000 37.260000 64.480000 37.460000 ;
        RECT 64.280000 37.700000 64.480000 37.900000 ;
        RECT 64.280000 38.140000 64.480000 38.340000 ;
        RECT 64.280000 38.580000 64.480000 38.780000 ;
        RECT 64.280000 39.020000 64.480000 39.220000 ;
        RECT 64.280000 39.460000 64.480000 39.660000 ;
        RECT 64.280000 39.900000 64.480000 40.100000 ;
        RECT 64.280000 51.715000 64.480000 51.915000 ;
        RECT 64.280000 52.135000 64.480000 52.335000 ;
        RECT 64.280000 52.555000 64.480000 52.755000 ;
        RECT 64.655000 47.800000 64.855000 48.000000 ;
        RECT 64.655000 56.470000 64.855000 56.670000 ;
        RECT 64.685000 36.820000 64.885000 37.020000 ;
        RECT 64.685000 37.260000 64.885000 37.460000 ;
        RECT 64.685000 37.700000 64.885000 37.900000 ;
        RECT 64.685000 38.140000 64.885000 38.340000 ;
        RECT 64.685000 38.580000 64.885000 38.780000 ;
        RECT 64.685000 39.020000 64.885000 39.220000 ;
        RECT 64.685000 39.460000 64.885000 39.660000 ;
        RECT 64.685000 39.900000 64.885000 40.100000 ;
        RECT 64.685000 51.715000 64.885000 51.915000 ;
        RECT 64.685000 52.135000 64.885000 52.335000 ;
        RECT 64.685000 52.555000 64.885000 52.755000 ;
        RECT 65.060000 47.800000 65.260000 48.000000 ;
        RECT 65.060000 56.470000 65.260000 56.670000 ;
        RECT 65.090000 36.820000 65.290000 37.020000 ;
        RECT 65.090000 37.260000 65.290000 37.460000 ;
        RECT 65.090000 37.700000 65.290000 37.900000 ;
        RECT 65.090000 38.140000 65.290000 38.340000 ;
        RECT 65.090000 38.580000 65.290000 38.780000 ;
        RECT 65.090000 39.020000 65.290000 39.220000 ;
        RECT 65.090000 39.460000 65.290000 39.660000 ;
        RECT 65.090000 39.900000 65.290000 40.100000 ;
        RECT 65.090000 51.715000 65.290000 51.915000 ;
        RECT 65.090000 52.135000 65.290000 52.335000 ;
        RECT 65.090000 52.555000 65.290000 52.755000 ;
        RECT 65.465000 47.800000 65.665000 48.000000 ;
        RECT 65.465000 56.470000 65.665000 56.670000 ;
        RECT 65.495000 36.820000 65.695000 37.020000 ;
        RECT 65.495000 37.260000 65.695000 37.460000 ;
        RECT 65.495000 37.700000 65.695000 37.900000 ;
        RECT 65.495000 38.140000 65.695000 38.340000 ;
        RECT 65.495000 38.580000 65.695000 38.780000 ;
        RECT 65.495000 39.020000 65.695000 39.220000 ;
        RECT 65.495000 39.460000 65.695000 39.660000 ;
        RECT 65.495000 39.900000 65.695000 40.100000 ;
        RECT 65.495000 51.715000 65.695000 51.915000 ;
        RECT 65.495000 52.135000 65.695000 52.335000 ;
        RECT 65.495000 52.555000 65.695000 52.755000 ;
        RECT 65.870000 47.800000 66.070000 48.000000 ;
        RECT 65.870000 56.470000 66.070000 56.670000 ;
        RECT 65.900000 36.820000 66.100000 37.020000 ;
        RECT 65.900000 37.260000 66.100000 37.460000 ;
        RECT 65.900000 37.700000 66.100000 37.900000 ;
        RECT 65.900000 38.140000 66.100000 38.340000 ;
        RECT 65.900000 38.580000 66.100000 38.780000 ;
        RECT 65.900000 39.020000 66.100000 39.220000 ;
        RECT 65.900000 39.460000 66.100000 39.660000 ;
        RECT 65.900000 39.900000 66.100000 40.100000 ;
        RECT 65.900000 51.715000 66.100000 51.915000 ;
        RECT 65.900000 52.135000 66.100000 52.335000 ;
        RECT 65.900000 52.555000 66.100000 52.755000 ;
        RECT 66.275000 47.800000 66.475000 48.000000 ;
        RECT 66.275000 56.470000 66.475000 56.670000 ;
        RECT 66.305000 36.820000 66.505000 37.020000 ;
        RECT 66.305000 37.260000 66.505000 37.460000 ;
        RECT 66.305000 37.700000 66.505000 37.900000 ;
        RECT 66.305000 38.140000 66.505000 38.340000 ;
        RECT 66.305000 38.580000 66.505000 38.780000 ;
        RECT 66.305000 39.020000 66.505000 39.220000 ;
        RECT 66.305000 39.460000 66.505000 39.660000 ;
        RECT 66.305000 39.900000 66.505000 40.100000 ;
        RECT 66.305000 51.715000 66.505000 51.915000 ;
        RECT 66.305000 52.135000 66.505000 52.335000 ;
        RECT 66.305000 52.555000 66.505000 52.755000 ;
        RECT 66.680000 47.800000 66.880000 48.000000 ;
        RECT 66.680000 56.470000 66.880000 56.670000 ;
        RECT 66.710000 36.820000 66.910000 37.020000 ;
        RECT 66.710000 37.260000 66.910000 37.460000 ;
        RECT 66.710000 37.700000 66.910000 37.900000 ;
        RECT 66.710000 38.140000 66.910000 38.340000 ;
        RECT 66.710000 38.580000 66.910000 38.780000 ;
        RECT 66.710000 39.020000 66.910000 39.220000 ;
        RECT 66.710000 39.460000 66.910000 39.660000 ;
        RECT 66.710000 39.900000 66.910000 40.100000 ;
        RECT 66.710000 51.715000 66.910000 51.915000 ;
        RECT 66.710000 52.135000 66.910000 52.335000 ;
        RECT 66.710000 52.555000 66.910000 52.755000 ;
        RECT 67.085000 47.800000 67.285000 48.000000 ;
        RECT 67.085000 56.470000 67.285000 56.670000 ;
        RECT 67.115000 36.820000 67.315000 37.020000 ;
        RECT 67.115000 37.260000 67.315000 37.460000 ;
        RECT 67.115000 37.700000 67.315000 37.900000 ;
        RECT 67.115000 38.140000 67.315000 38.340000 ;
        RECT 67.115000 38.580000 67.315000 38.780000 ;
        RECT 67.115000 39.020000 67.315000 39.220000 ;
        RECT 67.115000 39.460000 67.315000 39.660000 ;
        RECT 67.115000 39.900000 67.315000 40.100000 ;
        RECT 67.115000 51.715000 67.315000 51.915000 ;
        RECT 67.115000 52.135000 67.315000 52.335000 ;
        RECT 67.115000 52.555000 67.315000 52.755000 ;
        RECT 67.490000 47.800000 67.690000 48.000000 ;
        RECT 67.490000 56.470000 67.690000 56.670000 ;
        RECT 67.520000 36.820000 67.720000 37.020000 ;
        RECT 67.520000 37.260000 67.720000 37.460000 ;
        RECT 67.520000 37.700000 67.720000 37.900000 ;
        RECT 67.520000 38.140000 67.720000 38.340000 ;
        RECT 67.520000 38.580000 67.720000 38.780000 ;
        RECT 67.520000 39.020000 67.720000 39.220000 ;
        RECT 67.520000 39.460000 67.720000 39.660000 ;
        RECT 67.520000 39.900000 67.720000 40.100000 ;
        RECT 67.520000 51.715000 67.720000 51.915000 ;
        RECT 67.520000 52.135000 67.720000 52.335000 ;
        RECT 67.520000 52.555000 67.720000 52.755000 ;
        RECT 67.895000 47.800000 68.095000 48.000000 ;
        RECT 67.895000 56.470000 68.095000 56.670000 ;
        RECT 67.925000 36.820000 68.125000 37.020000 ;
        RECT 67.925000 37.260000 68.125000 37.460000 ;
        RECT 67.925000 37.700000 68.125000 37.900000 ;
        RECT 67.925000 38.140000 68.125000 38.340000 ;
        RECT 67.925000 38.580000 68.125000 38.780000 ;
        RECT 67.925000 39.020000 68.125000 39.220000 ;
        RECT 67.925000 39.460000 68.125000 39.660000 ;
        RECT 67.925000 39.900000 68.125000 40.100000 ;
        RECT 67.925000 51.715000 68.125000 51.915000 ;
        RECT 67.925000 52.135000 68.125000 52.335000 ;
        RECT 67.925000 52.555000 68.125000 52.755000 ;
        RECT 68.300000 47.800000 68.500000 48.000000 ;
        RECT 68.300000 56.470000 68.500000 56.670000 ;
        RECT 68.330000 36.820000 68.530000 37.020000 ;
        RECT 68.330000 37.260000 68.530000 37.460000 ;
        RECT 68.330000 37.700000 68.530000 37.900000 ;
        RECT 68.330000 38.140000 68.530000 38.340000 ;
        RECT 68.330000 38.580000 68.530000 38.780000 ;
        RECT 68.330000 39.020000 68.530000 39.220000 ;
        RECT 68.330000 39.460000 68.530000 39.660000 ;
        RECT 68.330000 39.900000 68.530000 40.100000 ;
        RECT 68.330000 51.715000 68.530000 51.915000 ;
        RECT 68.330000 52.135000 68.530000 52.335000 ;
        RECT 68.330000 52.555000 68.530000 52.755000 ;
        RECT 68.705000 47.800000 68.905000 48.000000 ;
        RECT 68.705000 56.470000 68.905000 56.670000 ;
        RECT 68.735000 36.820000 68.935000 37.020000 ;
        RECT 68.735000 37.260000 68.935000 37.460000 ;
        RECT 68.735000 37.700000 68.935000 37.900000 ;
        RECT 68.735000 38.140000 68.935000 38.340000 ;
        RECT 68.735000 38.580000 68.935000 38.780000 ;
        RECT 68.735000 39.020000 68.935000 39.220000 ;
        RECT 68.735000 39.460000 68.935000 39.660000 ;
        RECT 68.735000 39.900000 68.935000 40.100000 ;
        RECT 68.735000 51.715000 68.935000 51.915000 ;
        RECT 68.735000 52.135000 68.935000 52.335000 ;
        RECT 68.735000 52.555000 68.935000 52.755000 ;
        RECT 69.110000 47.800000 69.310000 48.000000 ;
        RECT 69.110000 56.470000 69.310000 56.670000 ;
        RECT 69.140000 36.820000 69.340000 37.020000 ;
        RECT 69.140000 37.260000 69.340000 37.460000 ;
        RECT 69.140000 37.700000 69.340000 37.900000 ;
        RECT 69.140000 38.140000 69.340000 38.340000 ;
        RECT 69.140000 38.580000 69.340000 38.780000 ;
        RECT 69.140000 39.020000 69.340000 39.220000 ;
        RECT 69.140000 39.460000 69.340000 39.660000 ;
        RECT 69.140000 39.900000 69.340000 40.100000 ;
        RECT 69.140000 51.715000 69.340000 51.915000 ;
        RECT 69.140000 52.135000 69.340000 52.335000 ;
        RECT 69.140000 52.555000 69.340000 52.755000 ;
        RECT 69.515000 47.800000 69.715000 48.000000 ;
        RECT 69.515000 56.470000 69.715000 56.670000 ;
        RECT 69.545000 36.820000 69.745000 37.020000 ;
        RECT 69.545000 37.260000 69.745000 37.460000 ;
        RECT 69.545000 37.700000 69.745000 37.900000 ;
        RECT 69.545000 38.140000 69.745000 38.340000 ;
        RECT 69.545000 38.580000 69.745000 38.780000 ;
        RECT 69.545000 39.020000 69.745000 39.220000 ;
        RECT 69.545000 39.460000 69.745000 39.660000 ;
        RECT 69.545000 39.900000 69.745000 40.100000 ;
        RECT 69.545000 51.715000 69.745000 51.915000 ;
        RECT 69.545000 52.135000 69.745000 52.335000 ;
        RECT 69.545000 52.555000 69.745000 52.755000 ;
        RECT 69.920000 47.800000 70.120000 48.000000 ;
        RECT 69.920000 56.470000 70.120000 56.670000 ;
        RECT 69.950000 36.820000 70.150000 37.020000 ;
        RECT 69.950000 37.260000 70.150000 37.460000 ;
        RECT 69.950000 37.700000 70.150000 37.900000 ;
        RECT 69.950000 38.140000 70.150000 38.340000 ;
        RECT 69.950000 38.580000 70.150000 38.780000 ;
        RECT 69.950000 39.020000 70.150000 39.220000 ;
        RECT 69.950000 39.460000 70.150000 39.660000 ;
        RECT 69.950000 39.900000 70.150000 40.100000 ;
        RECT 69.950000 51.715000 70.150000 51.915000 ;
        RECT 69.950000 52.135000 70.150000 52.335000 ;
        RECT 69.950000 52.555000 70.150000 52.755000 ;
        RECT 70.325000 47.800000 70.525000 48.000000 ;
        RECT 70.325000 56.470000 70.525000 56.670000 ;
        RECT 70.355000 36.820000 70.555000 37.020000 ;
        RECT 70.355000 37.260000 70.555000 37.460000 ;
        RECT 70.355000 37.700000 70.555000 37.900000 ;
        RECT 70.355000 38.140000 70.555000 38.340000 ;
        RECT 70.355000 38.580000 70.555000 38.780000 ;
        RECT 70.355000 39.020000 70.555000 39.220000 ;
        RECT 70.355000 39.460000 70.555000 39.660000 ;
        RECT 70.355000 39.900000 70.555000 40.100000 ;
        RECT 70.355000 51.715000 70.555000 51.915000 ;
        RECT 70.355000 52.135000 70.555000 52.335000 ;
        RECT 70.355000 52.555000 70.555000 52.755000 ;
        RECT 70.730000 47.800000 70.930000 48.000000 ;
        RECT 70.730000 56.470000 70.930000 56.670000 ;
        RECT 70.760000 36.820000 70.960000 37.020000 ;
        RECT 70.760000 37.260000 70.960000 37.460000 ;
        RECT 70.760000 37.700000 70.960000 37.900000 ;
        RECT 70.760000 38.140000 70.960000 38.340000 ;
        RECT 70.760000 38.580000 70.960000 38.780000 ;
        RECT 70.760000 39.020000 70.960000 39.220000 ;
        RECT 70.760000 39.460000 70.960000 39.660000 ;
        RECT 70.760000 39.900000 70.960000 40.100000 ;
        RECT 70.760000 51.715000 70.960000 51.915000 ;
        RECT 70.760000 52.135000 70.960000 52.335000 ;
        RECT 70.760000 52.555000 70.960000 52.755000 ;
        RECT 71.135000 47.800000 71.335000 48.000000 ;
        RECT 71.135000 56.470000 71.335000 56.670000 ;
        RECT 71.165000 36.820000 71.365000 37.020000 ;
        RECT 71.165000 37.260000 71.365000 37.460000 ;
        RECT 71.165000 37.700000 71.365000 37.900000 ;
        RECT 71.165000 38.140000 71.365000 38.340000 ;
        RECT 71.165000 38.580000 71.365000 38.780000 ;
        RECT 71.165000 39.020000 71.365000 39.220000 ;
        RECT 71.165000 39.460000 71.365000 39.660000 ;
        RECT 71.165000 39.900000 71.365000 40.100000 ;
        RECT 71.165000 51.715000 71.365000 51.915000 ;
        RECT 71.165000 52.135000 71.365000 52.335000 ;
        RECT 71.165000 52.555000 71.365000 52.755000 ;
        RECT 71.540000 47.800000 71.740000 48.000000 ;
        RECT 71.540000 56.470000 71.740000 56.670000 ;
        RECT 71.570000 36.820000 71.770000 37.020000 ;
        RECT 71.570000 37.260000 71.770000 37.460000 ;
        RECT 71.570000 37.700000 71.770000 37.900000 ;
        RECT 71.570000 38.140000 71.770000 38.340000 ;
        RECT 71.570000 38.580000 71.770000 38.780000 ;
        RECT 71.570000 39.020000 71.770000 39.220000 ;
        RECT 71.570000 39.460000 71.770000 39.660000 ;
        RECT 71.570000 39.900000 71.770000 40.100000 ;
        RECT 71.570000 51.715000 71.770000 51.915000 ;
        RECT 71.570000 52.135000 71.770000 52.335000 ;
        RECT 71.570000 52.555000 71.770000 52.755000 ;
        RECT 71.950000 47.800000 72.150000 48.000000 ;
        RECT 71.950000 56.470000 72.150000 56.670000 ;
        RECT 71.975000 36.820000 72.175000 37.020000 ;
        RECT 71.975000 37.260000 72.175000 37.460000 ;
        RECT 71.975000 37.700000 72.175000 37.900000 ;
        RECT 71.975000 38.140000 72.175000 38.340000 ;
        RECT 71.975000 38.580000 72.175000 38.780000 ;
        RECT 71.975000 39.020000 72.175000 39.220000 ;
        RECT 71.975000 39.460000 72.175000 39.660000 ;
        RECT 71.975000 39.900000 72.175000 40.100000 ;
        RECT 71.975000 51.715000 72.175000 51.915000 ;
        RECT 71.975000 52.135000 72.175000 52.335000 ;
        RECT 71.975000 52.555000 72.175000 52.755000 ;
        RECT 72.360000 47.800000 72.560000 48.000000 ;
        RECT 72.360000 56.470000 72.560000 56.670000 ;
        RECT 72.380000 36.820000 72.580000 37.020000 ;
        RECT 72.380000 37.260000 72.580000 37.460000 ;
        RECT 72.380000 37.700000 72.580000 37.900000 ;
        RECT 72.380000 38.140000 72.580000 38.340000 ;
        RECT 72.380000 38.580000 72.580000 38.780000 ;
        RECT 72.380000 39.020000 72.580000 39.220000 ;
        RECT 72.380000 39.460000 72.580000 39.660000 ;
        RECT 72.380000 39.900000 72.580000 40.100000 ;
        RECT 72.380000 51.715000 72.580000 51.915000 ;
        RECT 72.380000 52.135000 72.580000 52.335000 ;
        RECT 72.380000 52.555000 72.580000 52.755000 ;
        RECT 72.770000 47.800000 72.970000 48.000000 ;
        RECT 72.770000 56.470000 72.970000 56.670000 ;
        RECT 72.785000 36.820000 72.985000 37.020000 ;
        RECT 72.785000 37.260000 72.985000 37.460000 ;
        RECT 72.785000 37.700000 72.985000 37.900000 ;
        RECT 72.785000 38.140000 72.985000 38.340000 ;
        RECT 72.785000 38.580000 72.985000 38.780000 ;
        RECT 72.785000 39.020000 72.985000 39.220000 ;
        RECT 72.785000 39.460000 72.985000 39.660000 ;
        RECT 72.785000 39.900000 72.985000 40.100000 ;
        RECT 72.785000 51.715000 72.985000 51.915000 ;
        RECT 72.785000 52.135000 72.985000 52.335000 ;
        RECT 72.785000 52.555000 72.985000 52.755000 ;
        RECT 73.180000 47.800000 73.380000 48.000000 ;
        RECT 73.180000 56.470000 73.380000 56.670000 ;
        RECT 73.190000 36.820000 73.390000 37.020000 ;
        RECT 73.190000 37.260000 73.390000 37.460000 ;
        RECT 73.190000 37.700000 73.390000 37.900000 ;
        RECT 73.190000 38.140000 73.390000 38.340000 ;
        RECT 73.190000 38.580000 73.390000 38.780000 ;
        RECT 73.190000 39.020000 73.390000 39.220000 ;
        RECT 73.190000 39.460000 73.390000 39.660000 ;
        RECT 73.190000 39.900000 73.390000 40.100000 ;
        RECT 73.190000 51.715000 73.390000 51.915000 ;
        RECT 73.190000 52.135000 73.390000 52.335000 ;
        RECT 73.190000 52.555000 73.390000 52.755000 ;
        RECT 73.590000 47.800000 73.790000 48.000000 ;
        RECT 73.590000 56.470000 73.790000 56.670000 ;
        RECT 73.595000 36.820000 73.795000 37.020000 ;
        RECT 73.595000 37.260000 73.795000 37.460000 ;
        RECT 73.595000 37.700000 73.795000 37.900000 ;
        RECT 73.595000 38.140000 73.795000 38.340000 ;
        RECT 73.595000 38.580000 73.795000 38.780000 ;
        RECT 73.595000 39.020000 73.795000 39.220000 ;
        RECT 73.595000 39.460000 73.795000 39.660000 ;
        RECT 73.595000 39.900000 73.795000 40.100000 ;
        RECT 73.595000 51.715000 73.795000 51.915000 ;
        RECT 73.595000 52.135000 73.795000 52.335000 ;
        RECT 73.595000 52.555000 73.795000 52.755000 ;
        RECT 74.000000 36.820000 74.200000 37.020000 ;
        RECT 74.000000 37.260000 74.200000 37.460000 ;
        RECT 74.000000 37.700000 74.200000 37.900000 ;
        RECT 74.000000 38.140000 74.200000 38.340000 ;
        RECT 74.000000 38.580000 74.200000 38.780000 ;
        RECT 74.000000 39.020000 74.200000 39.220000 ;
        RECT 74.000000 39.460000 74.200000 39.660000 ;
        RECT 74.000000 39.900000 74.200000 40.100000 ;
        RECT 74.000000 47.800000 74.200000 48.000000 ;
        RECT 74.000000 51.715000 74.200000 51.915000 ;
        RECT 74.000000 52.135000 74.200000 52.335000 ;
        RECT 74.000000 52.555000 74.200000 52.755000 ;
        RECT 74.000000 56.470000 74.200000 56.670000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 41.585000 1.270000 46.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 41.585000 75.000000 46.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 41.685000 1.270000 46.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 41.685000 75.000000 46.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 25.835000 1.270000 30.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 25.835000 75.000000 30.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 25.935000 1.270000 30.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 25.935000 75.000000 30.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 58.235000 1.270000 62.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 58.235000 75.000000 62.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 58.335000 1.270000 62.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 58.335000 75.000000 62.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 31.885000 1.270000 35.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 31.885000 75.000000 35.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 31.985000 1.270000 35.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 31.985000 75.000000 35.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met1 ;
      RECT 0.000000 0.000000 75.000000 200.000000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 75.000000 200.000000 ;
    LAYER met3 ;
      RECT  0.000000  0.000000 75.000000  36.340000 ;
      RECT  0.000000 36.340000  0.570000  40.580000 ;
      RECT  0.000000 40.580000 75.000000  47.340000 ;
      RECT  0.000000 48.460000 24.795000  51.250000 ;
      RECT  0.000000 53.220000 24.795000  56.010000 ;
      RECT  0.000000 57.130000 75.000000 200.000000 ;
      RECT 24.795000 36.340000 49.990000  40.580000 ;
      RECT 24.795000 47.340000 49.990000  57.130000 ;
      RECT 49.990000 48.460000 75.000000  51.250000 ;
      RECT 49.990000 53.220000 75.000000  56.010000 ;
      RECT 74.690000 36.340000 75.000000  40.580000 ;
      RECT 74.690000 47.340000 75.000000  48.460000 ;
      RECT 74.690000 51.250000 75.000000  53.220000 ;
      RECT 74.690000 56.010000 75.000000  57.130000 ;
    LAYER met4 ;
      RECT  0.000000   0.000000  1.670000   1.635000 ;
      RECT  0.000000   7.885000  1.670000   8.485000 ;
      RECT  0.000000  13.935000  1.365000  14.535000 ;
      RECT  0.000000  18.785000  1.365000  19.385000 ;
      RECT  0.000000  24.835000  1.670000  25.435000 ;
      RECT  0.000000  30.885000  1.670000  31.485000 ;
      RECT  0.000000  35.735000  1.670000  36.335000 ;
      RECT  0.000000  40.585000  1.670000  41.185000 ;
      RECT  0.000000  46.635000  1.670000  47.335000 ;
      RECT  0.000000  57.135000  1.670000  57.835000 ;
      RECT  0.000000  63.085000  1.670000  63.685000 ;
      RECT  0.000000  68.935000  1.670000  69.635000 ;
      RECT  0.000000  95.400000 75.000000 175.385000 ;
      RECT  1.365000  13.935000 73.635000  19.385000 ;
      RECT  1.670000   0.000000 73.330000  13.935000 ;
      RECT  1.670000  19.385000 73.330000  36.335000 ;
      RECT  1.670000  40.585000 73.330000  47.335000 ;
      RECT  1.670000  48.465000 24.770000  51.245000 ;
      RECT  1.670000  53.225000 24.770000  56.005000 ;
      RECT  1.670000  57.135000 73.330000  95.400000 ;
      RECT  1.670000 175.385000 73.330000 200.000000 ;
      RECT 24.770000  36.335000 50.015000  40.585000 ;
      RECT 24.770000  47.335000 50.015000  57.135000 ;
      RECT 50.015000  48.465000 73.330000  51.245000 ;
      RECT 50.015000  53.225000 73.330000  56.005000 ;
      RECT 73.330000   0.000000 75.000000   1.635000 ;
      RECT 73.330000   7.885000 75.000000   8.485000 ;
      RECT 73.330000  24.835000 75.000000  25.435000 ;
      RECT 73.330000  30.885000 75.000000  31.485000 ;
      RECT 73.330000  35.735000 75.000000  36.335000 ;
      RECT 73.330000  40.585000 75.000000  41.185000 ;
      RECT 73.330000  46.635000 75.000000  47.335000 ;
      RECT 73.330000  57.135000 75.000000  57.835000 ;
      RECT 73.330000  63.085000 75.000000  63.685000 ;
      RECT 73.330000  68.935000 75.000000  69.635000 ;
      RECT 73.635000  13.935000 75.000000  14.535000 ;
      RECT 73.635000  18.785000 75.000000  19.385000 ;
    LAYER met5 ;
      RECT 0.000000   0.000000 75.000000   1.335000 ;
      RECT 0.000000  95.785000 75.000000 174.985000 ;
      RECT 1.765000  14.235000 73.235000  19.085000 ;
      RECT 2.070000   1.335000 72.930000  14.235000 ;
      RECT 2.070000  19.085000 72.930000  95.785000 ;
      RECT 2.070000 174.985000 72.930000 200.000000 ;
  END
END sky130_fd_io__overlay_vssa_hvc
END LIBRARY
