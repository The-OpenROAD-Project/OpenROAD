VERSION 5.8 ;

#USEMINSPACING OBS OFF ;
#BUSBITCHARS "[]" ;

# UNITS
# YBASE MICRON 1000 ;
# END UNITS

SITE IOSITE
  SYMMETRY Y ;
  CLASS PAD ;
  SIZE    1.000 BY 140.000 ;
END IOSITE

MACRO DUMMY_BUMP
  CLASS PAD AREAIO ;
  ORIGIN 0 0 ;
  SIZE 45 BY 45 ;
  SYMMETRY X Y R90 ;
  PIN PAD
    DIRECTION INOUT ;
    PORT
      LAYER metal10 ;
        RECT 0.0 0.0 45.0 45.0 ;
    END
  END PAD
END DUMMY_BUMP

MACRO PADCELL_SIG_V
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN PADCELL_SIG_V 0 0 ;
  SIZE 25.0 BY 140 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE ;
  PIN PAD 
    USE SIGNAL ;
    DIRECTION INOUT ;
    PORT
      CLASS BUMP ;
      LAYER metal10 ;
        RECT 15.0 53.0 20.0 58.0 ;
    END
  END PAD
  PIN A
    USE SIGNAL ;
    DIRECTION INPUT ;
    PORT
      CLASS CORE ;
      LAYER metal4 ;
        RECT 13.170 139.900 13.330 140.000 ;
      LAYER metal5 ; 
        RECT 13.170 139.900 13.330 140.000 ;
      LAYER metal6 ; 
        RECT 13.170 139.900 13.330 140.000 ;
      LAYER metal7 ; 
        RECT 13.170 139.900 13.330 140.000 ;
      LAYER metal8 ;
        RECT 13.170 139.900 13.330 140.000 ;
    END
  END A
  PIN Y
    USE SIGNAL ;
    DIRECTION OUTPUT ;
    PORT
      CLASS CORE ;
      LAYER metal4 ;
        RECT 23.936 139.900 24.096 140.000 ;
      LAYER metal5 ;
        RECT 23.936 139.900 24.096 140.000 ;
      LAYER metal6 ;
        RECT 23.936 139.900 24.096 140.000 ;
      LAYER metal7 ;
        RECT 23.936 139.900 24.096 140.000 ;
      LAYER metal8 ;
        RECT 23.936 139.900 24.096 140.000 ;
    END
  END Y
  PIN PU
    USE SIGNAL ;
    DIRECTION OUTPUT ;
    PORT
      CLASS CORE ;
      LAYER metal4 ;
        RECT 15.170 139.900 15.330 140.000 ;
      LAYER metal5 ;
        RECT 15.170 139.900 15.330 140.000 ;
      LAYER metal6 ;
        RECT 15.170 139.900 15.330 140.000 ;
      LAYER metal7 ;
        RECT 15.170 139.900 15.330 140.000 ;
      LAYER metal8 ;
        RECT 15.170 139.900 15.330 140.000 ;
    END
  END PU
  PIN OE
    USE SIGNAL ;
    DIRECTION OUTPUT ;
    PORT
      CLASS CORE ;
      LAYER metal4 ;
        RECT 15.170 139.900 15.330 140.000 ;
      LAYER metal5 ;
        RECT 15.170 139.900 15.330 140.000 ;
      LAYER metal6 ;
        RECT 15.170 139.900 15.330 140.000 ;
      LAYER metal7 ;
        RECT 15.170 139.900 15.330 140.000 ;
      LAYER metal8 ;
        RECT 15.170 139.900 15.330 140.000 ;
    END
  END OE
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 2.0 25.0 4.0 ;
    END
  END DVSS
  PIN VDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 14.0 25.0 16.0 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 10.0 25.0 12.0 ;
    END
  END VSS
  PIN DVDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 6.0 25.0 8.0 ;
    END
  END DVDD
END PADCELL_SIG_V

MACRO PADCELL_SIG_H
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 25.0 BY 140 ;
  SYMMETRY X Y R90 ;
  PIN PAD 
    DIRECTION INOUT ;
    PORT
      LAYER metal10 ;
        RECT 15.0 53.0 20.0 58.0 ;
    END
  END PAD
  PIN A
    USE SIGNAL ;
    DIRECTION INPUT ;
    PORT
      CLASS CORE ;
      LAYER metal4 ;
        RECT 13.170 139.900 13.330 140.000 ;
      LAYER metal5 ; 
        RECT 13.170 139.900 13.330 140.000 ;
      LAYER metal6 ; 
        RECT 13.170 139.900 13.330 140.000 ;
      LAYER metal7 ; 
        RECT 13.170 139.900 13.330 140.000 ;
      LAYER metal8 ;
        RECT 13.170 139.900 13.330 140.000 ;
    END
  END A
  PIN Y
    USE SIGNAL ;
    DIRECTION OUTPUT ;
    PORT
      CLASS CORE ;
      LAYER metal4 ;
        RECT 23.936 139.900 24.096 140.000 ;
      LAYER metal5 ; 
        RECT 23.936 139.900 24.096 140.000 ;
      LAYER metal6 ; 
        RECT 23.936 139.900 24.096 140.000 ;
      LAYER metal7 ; 
        RECT 23.936 139.900 24.096 140.000 ;
      LAYER metal8 ; 
        RECT 23.936 139.900 24.096 140.000 ;
    END
  END Y
  PIN PU
    USE SIGNAL ;
    DIRECTION OUTPUT ;
    PORT
      CLASS CORE ;
      LAYER metal4 ;
        RECT 15.170 139.900 15.330 140.000 ;
      LAYER metal5 ;
        RECT 15.170 139.900 15.330 140.000 ;
      LAYER metal6 ;
        RECT 15.170 139.900 15.330 140.000 ;
      LAYER metal7 ;
        RECT 15.170 139.900 15.330 140.000 ;
      LAYER metal8 ;
        RECT 15.170 139.900 15.330 140.000 ;
    END
  END PU
  PIN OE
    USE SIGNAL ;
    DIRECTION OUTPUT ;
    PORT
      CLASS CORE ;
      LAYER metal4 ;
        RECT 15.170 139.900 15.330 140.000 ;
      LAYER metal5 ;
        RECT 15.170 139.900 15.330 140.000 ;
      LAYER metal6 ;
        RECT 15.170 139.900 15.330 140.000 ;
      LAYER metal7 ;
        RECT 15.170 139.900 15.330 140.000 ;
      LAYER metal8 ;
        RECT 15.170 139.900 15.330 140.000 ;
    END
  END OE
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 2.0 25.0 4.0 ;
    END
  END DVSS
  PIN VDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 14.0 25.0 16.0 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 10.0 25.0 12.0 ;
    END
  END VSS
  PIN DVDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 6.0 25.0 8.0 ;
    END
  END DVDD
END PADCELL_SIG_H

MACRO PADCELL_VDD_V
  CLASS PAD AREAIO ;
  ORIGIN 0 0 ;
  SIZE 25.0 BY 140 ;
  SYMMETRY X Y R90 ;
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 2.0 25.0 4.0 ;
    END
  END DVSS
  PIN VDD
    USE POWER ;
    PORT
      CLASS BUMP ;
      LAYER metal10 ;
        RECT 15.0 53.0 20.0 58.0 ;
    END
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 14.0 25.0 16.0 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 10.0 25.0 12.0 ;
    END
  END VSS
  PIN DVDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 6.0 25.0 8.0 ;
    END
  END DVDD
END PADCELL_VDD_V

MACRO PADCELL_VDD_H
  CLASS PAD AREAIO ;
  ORIGIN 0 0 ;
  SIZE 25.0 BY 140 ;
  SYMMETRY X Y R90 ;
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 2.0 25.0 4.0 ;
    END
  END DVSS
  PIN VDD
    USE POWER ;
    PORT
      CLASS BUMP ;
      LAYER metal10 ;
        RECT 15.0 53.0 20.0 58.0 ;
    END
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 14.0 25.0 16.0 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 10.0 25.0 12.0 ;
    END
  END VSS
  PIN DVDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 6.0 25.0 8.0 ;
    END
  END DVDD
END PADCELL_VDD_H

MACRO PADCELL_VSS_H
  CLASS PAD AREAIO ;
  ORIGIN 0 0 ;
  SIZE 25.0 BY 140 ;
  SYMMETRY X Y R90 ;
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 2.0 25.0 4.0 ;
    END
  END DVSS
  PIN VDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 14.0 25.0 16.0 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      CLASS BUMP ;
      LAYER metal10 ;
        RECT 15.0 53.0 20.0 58.0 ;
    END
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 10.0 25.0 12.0 ;
    END
  END VSS
  PIN DVDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 6.0 25.0 8.0 ;
    END
  END DVDD
END PADCELL_VSS_H

MACRO PADCELL_VSS_V
  CLASS PAD AREAIO ;
  ORIGIN 0 0 ;
  SIZE 25.0 BY 140 ;
  SYMMETRY X Y R90 ;
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 2.0 25.0 4.0 ;
    END
  END DVSS
  PIN VDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 14.0 25.0 16.0 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      CLASS BUMP ;
      LAYER metal10 ;
        RECT 15.0 53.0 20.0 58.0 ;
    END
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 10.0 25.0 12.0 ;
    END
  END VSS
  PIN DVDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 6.0 25.0 8.0 ;
    END
  END DVDD
END PADCELL_VSS_V

MACRO PADCELL_VDDIO_H
  CLASS PAD AREAIO ;
  ORIGIN 0 0 ;
  SIZE 25.0 BY 140 ;
  SYMMETRY X Y R90 ;
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 2.0 25.0 4.0 ;
    END
  END DVSS
  PIN VDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 14.0 25.0 16.0 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 10.0 25.0 12.0 ;
    END
  END VSS
  PIN DVDD
    USE POWER ;
    PORT
      CLASS BUMP ;
      LAYER metal10 ;
        RECT 15.0 53.0 20.0 58.0 ;
    END
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 6.0 25.0 8.0 ;
    END
  END DVDD
END PADCELL_VDDIO_H

MACRO PADCELL_VDDIO_V
  CLASS PAD AREAIO ;
  ORIGIN 0 0 ;
  SIZE 25.0 BY 140 ;
  SYMMETRY X Y R90 ;
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 2.0 25.0 4.0 ;
    END
  END DVSS
  PIN VDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 14.0 25.0 16.0 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 10.0 25.0 12.0 ;
    END
  END VSS
  PIN DVDD
    USE POWER ;
    PORT
      CLASS BUMP ;
      LAYER metal10 ;
        RECT 15.0 53.0 20.0 58.0 ;
    END
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 6.0 25.0 8.0 ;
    END
  END DVDD
END PADCELL_VDDIO_V

MACRO PADCELL_VSSIO_H
  CLASS PAD AREAIO ;
  ORIGIN 0 0 ;
  SIZE 25.0 BY 140 ;
  SYMMETRY X Y R90 ;
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      CLASS BUMP ;
      LAYER metal10 ;
        RECT 15.0 53.0 20.0 58.0 ;
    END
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 2.0 25.0 4.0 ;
    END
  END DVSS
  PIN VDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 14.0 25.0 16.0 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 10.0 25.0 12.0 ;
    END
  END VSS
  PIN DVDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 6.0 25.0 8.0 ;
    END
  END DVDD
END PADCELL_VSSIO_H

MACRO PADCELL_VSSIO_V
  CLASS PAD AREAIO ;
  ORIGIN 0 0 ;
  SIZE 25.0 BY 140 ;
  SYMMETRY X Y R90 ;
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      CLASS BUMP ;
      LAYER metal10 ;
        RECT 15.0 53.0 20.0 58.0 ;
    END
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 2.0 25.0 4.0 ;
    END
  END DVSS
  PIN VDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 14.0 25.0 16.0 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 10.0 25.0 12.0 ;
    END
  END VSS
  PIN DVDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 6.0 25.0 8.0 ;
    END
  END DVDD
END PADCELL_VSSIO_V

MACRO PAD_CORNER
  CLASS ENDCAP BOTTOMLEFT ;
  ORIGIN 0 0 ;
  SIZE 140 BY 140 ;
  SYMMETRY X Y R90 ;
END PAD_CORNER

MACRO PAD_FILL1_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  SIZE 1 BY 140 ;
  SYMMETRY X Y R90 ;
  PIN DVSS
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 2.0 1.0 4.0 ;
    END
  END DVSS
  PIN VDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 14.0 1.0 16.0 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 10.0 1.0 12.0 ;
    END
  END VSS
  PIN DVDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 6.0 1.0 8.0 ;
    END
  END DVDD
END PAD_FILL1_V

MACRO PAD_FILL5_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  SIZE 5 BY 140 ;
  SYMMETRY X Y R90 ;
  PIN DVSS
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 2.0 5.0 4.0 ;
    END
  END DVSS
  PIN VDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 14.0 5.0 16.0 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 10.0 5.0 12.0 ;
    END
  END VSS
  PIN DVDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 6.0 5.0 8.0 ;
    END
  END DVDD
END PAD_FILL5_V

MACRO PAD_FILL1_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  SIZE 140 BY 1 ;
  SYMMETRY X Y R90 ;
  PIN DVSS
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 2.0 0.0 4.0 1.0 ;
    END
  END DVSS
  PIN VDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 14.0 0.0 16.0 1.0 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 10.0 0.0 12.0 1.0 ;
    END
  END VSS
  PIN DVDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 6.0 0.0 8.0 1.0 ;
    END
  END DVDD
END PAD_FILL1_H

MACRO PAD_FILL5_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  SIZE 140 BY 5 ;
  SYMMETRY X Y R90 ;
  PIN DVSS
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 2.0 0.0 4.0 5.0 ;
    END
  END DVSS
  PIN VDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 14.0 0.0 16.0 5.0 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 10.0 0.0 12.0 5.0 ;
    END
  END VSS
  PIN DVDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 6.0 0.0 8.0 5.0 ;
    END
  END DVDD
END PAD_FILL5_H

MACRO PADCELL_PWRDET_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  SIZE 5 BY 140 ;
  SYMMETRY X Y R90 ;
  PIN DVSS
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 2.0 5.0 4.0 ;
    END
  END DVSS
  PIN VDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 14.0 5.0 16.0 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 10.0 5.0 12.0 ;
    END
  END VSS
  PIN DVDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 6.0 5.0 8.0 ;
    END
  END DVDD
END PADCELL_PWRDET_V

MACRO PADCELL_PWRDET_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  SIZE 5 BY 140 ;
  SYMMETRY X Y R90 ;
  PIN DVSS
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 2.0 5.0 4.0 ;
    END
  END DVSS
  PIN VDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 14.0 5.0 16.0 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 10.0 5.0 12.0 ;
    END
  END VSS
  PIN DVDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 6.0 5.0 8.0 ;
    END
  END DVDD
END PADCELL_PWRDET_H

MACRO PADCELL_CBRK_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  SIZE 5 BY 140 ;
  SYMMETRY X Y R90 ;
  PIN DVSS
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 2.0 5.0 4.0 ;
    END
  END DVSS
  PIN VDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 14.0 5.0 16.0 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 10.0 5.0 12.0 ;
    END
  END VSS
  PIN DVDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 6.0 5.0 8.0 ;
    END
  END DVDD
END PADCELL_CBRK_V

MACRO PADCELL_CBRK_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  SIZE 5 BY 140 ;
  SYMMETRY X Y R90 ;
  PIN DVSS
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 2.0 5.0 4.0 ;
    END
  END DVSS
  PIN VDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 14.0 5.0 16.0 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 10.0 5.0 12.0 ;
    END
  END VSS
  PIN DVDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 6.0 5.0 8.0 ;
    END
  END DVDD
END PADCELL_CBRK_H

MACRO PADCELL_FBRK_V
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  SIZE 5 BY 140 ;
  SYMMETRY X Y R90 ;
  PIN DVSS
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 2.0 5.0 4.0 ;
    END
  END DVSS
  PIN VDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 14.0 5.0 16.0 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 10.0 5.0 12.0 ;
    END
  END VSS
  PIN DVDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 0.0 6.0 5.0 8.0 ;
    END
  END DVDD
END PADCELL_FBRK_V

MACRO PADCELL_FBRK_H
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  SIZE 5 BY 140 ;
  SYMMETRY X Y R90 ;
  PIN DVSS
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 2.0 0.0 4.0 5.0 ;
    END
  END DVSS
  PIN VDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 14.0 0.0 16.0 5.0 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 10.0 0.0 12.0 5.0 ;
    END
  END VSS
  PIN DVDD
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal9 ;
        RECT 6.0 0.0 8.0 5.0 ;
    END
  END DVDD
END PADCELL_FBRK_H

END LIBRARY
