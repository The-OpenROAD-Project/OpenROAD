VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MANUFACTURINGGRID 0.0025 ;

LAYER metal1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.19 ;
  WIDTH 0.065 ;
END metal1

LAYER via1
  TYPE CUT ;
  SPACING 0.075 ;
END via1

LAYER metal2
  TYPE ROUTING ;
  MASK 2 ;
  DIRECTION VERTICAL ;
  PITCH 0.19 ;
  WIDTH 0.07 ;
END metal2

LAYER via2
  TYPE CUT ;
  SPACING 0.085 ;
END via2

LAYER metal3
  TYPE ROUTING ;
  MASK 3 ;
  DIRECTION HORIZONTAL ;
  PITCH 0.19 ;
  WIDTH 0.07 ;
END metal3
