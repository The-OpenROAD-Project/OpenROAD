module Element (clock,
    io_lsbIns_1,
    io_lsbIns_2,
    io_lsbIns_3,
    io_lsbOuts_0,
    io_lsbOuts_1,
    io_lsbOuts_2,
    io_lsbOuts_3,
    io_ins_down,
    io_ins_left,
    io_ins_right,
    io_ins_up,
    io_outs_down,
    io_outs_left,
    io_outs_right,
    io_outs_up);
 input clock;
 input io_lsbIns_1;
 input io_lsbIns_2;
 input io_lsbIns_3;
 output io_lsbOuts_0;
 output io_lsbOuts_1;
 output io_lsbOuts_2;
 output io_lsbOuts_3;
 input [63:0] io_ins_down;
 input [63:0] io_ins_left;
 input [63:0] io_ins_right;
 input [63:0] io_ins_up;
 output [63:0] io_outs_down;
 output [63:0] io_outs_left;
 output [63:0] io_outs_right;
 output [63:0] io_outs_up;

 wire clknet_leaf_32_clock;
 wire clknet_leaf_30_clock;
 wire clknet_leaf_29_clock;
 wire clknet_leaf_28_clock;
 wire clknet_leaf_21_clock;
 wire clknet_leaf_20_clock;
 wire clknet_leaf_14_clock;
 wire clknet_leaf_13_clock;
 wire clknet_leaf_12_clock;
 wire clknet_leaf_11_clock;
 wire clknet_leaf_9_clock;
 wire clknet_leaf_7_clock;
 wire clknet_leaf_5_clock;
 wire clknet_leaf_4_clock;
 wire clknet_leaf_3_clock;
 wire \_io_outs_up_mult_io_o[0] ;
 wire \_io_outs_up_mult_io_o[1] ;
 wire \_io_outs_up_mult_io_o[2] ;
 wire \_io_outs_up_mult_io_o[3] ;
 wire \_io_outs_up_mult_io_o[4] ;
 wire \_io_outs_up_mult_io_o[5] ;
 wire \_io_outs_up_mult_io_o[6] ;
 wire \_io_outs_up_mult_io_o[7] ;
 wire \_io_outs_up_mult_io_o[8] ;
 wire \_io_outs_up_mult_io_o[9] ;
 wire \_io_outs_up_mult_io_o[10] ;
 wire \_io_outs_up_mult_io_o[11] ;
 wire \_io_outs_up_mult_io_o[12] ;
 wire \_io_outs_up_mult_io_o[13] ;
 wire \_io_outs_up_mult_io_o[14] ;
 wire \_io_outs_up_mult_io_o[15] ;
 wire \_io_outs_up_mult_io_o[16] ;
 wire \_io_outs_up_mult_io_o[17] ;
 wire \_io_outs_up_mult_io_o[18] ;
 wire \_io_outs_up_mult_io_o[19] ;
 wire \_io_outs_up_mult_io_o[20] ;
 wire \_io_outs_up_mult_io_o[21] ;
 wire \_io_outs_up_mult_io_o[22] ;
 wire \_io_outs_up_mult_io_o[23] ;
 wire \_io_outs_up_mult_io_o[24] ;
 wire \_io_outs_up_mult_io_o[25] ;
 wire \_io_outs_up_mult_io_o[26] ;
 wire \_io_outs_up_mult_io_o[27] ;
 wire \_io_outs_up_mult_io_o[28] ;
 wire \_io_outs_up_mult_io_o[29] ;
 wire \_io_outs_up_mult_io_o[30] ;
 wire \_io_outs_up_mult_io_o[31] ;
 wire \_io_outs_right_mult_io_o[0] ;
 wire \_io_outs_right_mult_io_o[1] ;
 wire \_io_outs_right_mult_io_o[2] ;
 wire \_io_outs_right_mult_io_o[3] ;
 wire \_io_outs_right_mult_io_o[4] ;
 wire \_io_outs_right_mult_io_o[5] ;
 wire \_io_outs_right_mult_io_o[6] ;
 wire \_io_outs_right_mult_io_o[7] ;
 wire \_io_outs_right_mult_io_o[8] ;
 wire \_io_outs_right_mult_io_o[9] ;
 wire \_io_outs_right_mult_io_o[10] ;
 wire \_io_outs_right_mult_io_o[11] ;
 wire \_io_outs_right_mult_io_o[12] ;
 wire \_io_outs_right_mult_io_o[13] ;
 wire \_io_outs_right_mult_io_o[14] ;
 wire \_io_outs_right_mult_io_o[15] ;
 wire \_io_outs_right_mult_io_o[16] ;
 wire \_io_outs_right_mult_io_o[17] ;
 wire \_io_outs_right_mult_io_o[18] ;
 wire \_io_outs_right_mult_io_o[19] ;
 wire \_io_outs_right_mult_io_o[20] ;
 wire \_io_outs_right_mult_io_o[21] ;
 wire \_io_outs_right_mult_io_o[22] ;
 wire \_io_outs_right_mult_io_o[23] ;
 wire \_io_outs_right_mult_io_o[24] ;
 wire \_io_outs_right_mult_io_o[25] ;
 wire \_io_outs_right_mult_io_o[26] ;
 wire \_io_outs_right_mult_io_o[27] ;
 wire \_io_outs_right_mult_io_o[28] ;
 wire \_io_outs_right_mult_io_o[29] ;
 wire \_io_outs_right_mult_io_o[30] ;
 wire \_io_outs_right_mult_io_o[31] ;
 wire \REG_2[0] ;
 wire \REG_2[1] ;
 wire \REG_2[2] ;
 wire \REG_2[3] ;
 wire \REG_2[4] ;
 wire \REG_2[5] ;
 wire \REG_2[6] ;
 wire \REG_2[7] ;
 wire \REG_2[8] ;
 wire \REG_2[9] ;
 wire \REG_2[10] ;
 wire \REG_2[11] ;
 wire \REG_2[12] ;
 wire \REG_2[13] ;
 wire \REG_2[14] ;
 wire \REG_2[15] ;
 wire \REG_2[16] ;
 wire \REG_2[17] ;
 wire \REG_2[18] ;
 wire \REG_2[19] ;
 wire \REG_2[20] ;
 wire \REG_2[21] ;
 wire \REG_2[22] ;
 wire \REG_2[23] ;
 wire \REG_2[24] ;
 wire \REG_2[25] ;
 wire \REG_2[26] ;
 wire \REG_2[27] ;
 wire \REG_2[28] ;
 wire \REG_2[29] ;
 wire \REG_2[30] ;
 wire \REG_2[31] ;
 wire \_io_outs_left_mult_io_o[0] ;
 wire \_io_outs_left_mult_io_o[1] ;
 wire \_io_outs_left_mult_io_o[2] ;
 wire \_io_outs_left_mult_io_o[3] ;
 wire \_io_outs_left_mult_io_o[4] ;
 wire \_io_outs_left_mult_io_o[5] ;
 wire \_io_outs_left_mult_io_o[6] ;
 wire \_io_outs_left_mult_io_o[7] ;
 wire \_io_outs_left_mult_io_o[8] ;
 wire \_io_outs_left_mult_io_o[9] ;
 wire \_io_outs_left_mult_io_o[10] ;
 wire \_io_outs_left_mult_io_o[11] ;
 wire \_io_outs_left_mult_io_o[12] ;
 wire \_io_outs_left_mult_io_o[13] ;
 wire \_io_outs_left_mult_io_o[14] ;
 wire \_io_outs_left_mult_io_o[15] ;
 wire \_io_outs_left_mult_io_o[16] ;
 wire \_io_outs_left_mult_io_o[17] ;
 wire \_io_outs_left_mult_io_o[18] ;
 wire \_io_outs_left_mult_io_o[19] ;
 wire \_io_outs_left_mult_io_o[20] ;
 wire \_io_outs_left_mult_io_o[21] ;
 wire \_io_outs_left_mult_io_o[22] ;
 wire \_io_outs_left_mult_io_o[23] ;
 wire \_io_outs_left_mult_io_o[24] ;
 wire \_io_outs_left_mult_io_o[25] ;
 wire \_io_outs_left_mult_io_o[26] ;
 wire \_io_outs_left_mult_io_o[27] ;
 wire \_io_outs_left_mult_io_o[28] ;
 wire \_io_outs_left_mult_io_o[29] ;
 wire \_io_outs_left_mult_io_o[30] ;
 wire \_io_outs_left_mult_io_o[31] ;
 wire \REG[0] ;
 wire \REG[1] ;
 wire \REG[2] ;
 wire \REG[3] ;
 wire \REG[4] ;
 wire \REG[5] ;
 wire \REG[6] ;
 wire \REG[7] ;
 wire \REG[8] ;
 wire \REG[9] ;
 wire \REG[10] ;
 wire \REG[11] ;
 wire \REG[12] ;
 wire \REG[13] ;
 wire \REG[14] ;
 wire \REG[15] ;
 wire \REG[16] ;
 wire \REG[17] ;
 wire \REG[18] ;
 wire \REG[19] ;
 wire \REG[20] ;
 wire \REG[21] ;
 wire \REG[22] ;
 wire \REG[23] ;
 wire \REG[24] ;
 wire \REG[25] ;
 wire \REG[26] ;
 wire \REG[27] ;
 wire \REG[28] ;
 wire \REG[29] ;
 wire \REG[30] ;
 wire \REG[31] ;
 wire \_io_outs_down_mult_io_o[0] ;
 wire \_io_outs_down_mult_io_o[1] ;
 wire \_io_outs_down_mult_io_o[2] ;
 wire \_io_outs_down_mult_io_o[3] ;
 wire \_io_outs_down_mult_io_o[4] ;
 wire \_io_outs_down_mult_io_o[5] ;
 wire \_io_outs_down_mult_io_o[6] ;
 wire \_io_outs_down_mult_io_o[7] ;
 wire \_io_outs_down_mult_io_o[8] ;
 wire \_io_outs_down_mult_io_o[9] ;
 wire \_io_outs_down_mult_io_o[10] ;
 wire \_io_outs_down_mult_io_o[11] ;
 wire \_io_outs_down_mult_io_o[12] ;
 wire \_io_outs_down_mult_io_o[13] ;
 wire \_io_outs_down_mult_io_o[14] ;
 wire \_io_outs_down_mult_io_o[15] ;
 wire \_io_outs_down_mult_io_o[16] ;
 wire \_io_outs_down_mult_io_o[17] ;
 wire \_io_outs_down_mult_io_o[18] ;
 wire \_io_outs_down_mult_io_o[19] ;
 wire \_io_outs_down_mult_io_o[20] ;
 wire \_io_outs_down_mult_io_o[21] ;
 wire \_io_outs_down_mult_io_o[22] ;
 wire \_io_outs_down_mult_io_o[23] ;
 wire \_io_outs_down_mult_io_o[24] ;
 wire \_io_outs_down_mult_io_o[25] ;
 wire \_io_outs_down_mult_io_o[26] ;
 wire \_io_outs_down_mult_io_o[27] ;
 wire \_io_outs_down_mult_io_o[28] ;
 wire \_io_outs_down_mult_io_o[29] ;
 wire \_io_outs_down_mult_io_o[30] ;
 wire \_io_outs_down_mult_io_o[31] ;
 wire \REG_4[0] ;
 wire \REG_4[1] ;
 wire \REG_4[2] ;
 wire \REG_4[3] ;
 wire \REG_4[4] ;
 wire \REG_4[5] ;
 wire \REG_4[6] ;
 wire \REG_4[7] ;
 wire \REG_4[8] ;
 wire \REG_4[9] ;
 wire \REG_4[10] ;
 wire \REG_4[11] ;
 wire \REG_4[12] ;
 wire \REG_4[13] ;
 wire \REG_4[14] ;
 wire \REG_4[15] ;
 wire \REG_4[16] ;
 wire \REG_4[17] ;
 wire \REG_4[18] ;
 wire \REG_4[19] ;
 wire \REG_4[20] ;
 wire \REG_4[21] ;
 wire \REG_4[22] ;
 wire \REG_4[23] ;
 wire \REG_4[24] ;
 wire \REG_4[25] ;
 wire \REG_4[26] ;
 wire \REG_4[27] ;
 wire \REG_4[28] ;
 wire \REG_4[29] ;
 wire \REG_4[30] ;
 wire \REG_4[31] ;
 wire \REG_1[0] ;
 wire \REG_1[1] ;
 wire \REG_1[2] ;
 wire \REG_1[3] ;
 wire \REG_1[4] ;
 wire \REG_1[5] ;
 wire \REG_1[6] ;
 wire \REG_1[7] ;
 wire \REG_1[8] ;
 wire \REG_1[9] ;
 wire \REG_1[10] ;
 wire \REG_1[11] ;
 wire \REG_1[12] ;
 wire \REG_1[13] ;
 wire \REG_1[14] ;
 wire \REG_1[15] ;
 wire \REG_1[16] ;
 wire \REG_1[17] ;
 wire \REG_1[18] ;
 wire \REG_1[19] ;
 wire \REG_1[20] ;
 wire \REG_1[21] ;
 wire \REG_1[22] ;
 wire \REG_1[23] ;
 wire \REG_1[24] ;
 wire \REG_1[25] ;
 wire \REG_1[26] ;
 wire \REG_1[27] ;
 wire \REG_1[28] ;
 wire \REG_1[29] ;
 wire \REG_1[30] ;
 wire \REG_1[31] ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire net369;
 wire net368;
 wire net367;
 wire net366;
 wire net365;
 wire net364;
 wire net363;
 wire net362;
 wire net361;
 wire net360;
 wire net359;
 wire net358;
 wire net357;
 wire net356;
 wire net355;
 wire net354;
 wire net353;
 wire net352;
 wire net351;
 wire net350;
 wire net349;
 wire net348;
 wire net375;
 wire net374;
 wire net373;
 wire net372;
 wire net371;
 wire net370;
 wire net341;
 wire net340;
 wire net339;
 wire net338;
 wire net337;
 wire net336;
 wire net335;
 wire net334;
 wire net333;
 wire net332;
 wire net331;
 wire net330;
 wire net329;
 wire net328;
 wire net327;
 wire net326;
 wire net325;
 wire net324;
 wire net323;
 wire net322;
 wire net321;
 wire net320;
 wire net347;
 wire net346;
 wire net345;
 wire net344;
 wire net343;
 wire net342;
 wire net313;
 wire net312;
 wire net311;
 wire net310;
 wire net309;
 wire net308;
 wire net307;
 wire net306;
 wire net305;
 wire net304;
 wire net303;
 wire net302;
 wire net301;
 wire net300;
 wire net299;
 wire net298;
 wire net297;
 wire net296;
 wire net295;
 wire net294;
 wire net293;
 wire net292;
 wire net319;
 wire net318;
 wire net317;
 wire net316;
 wire net315;
 wire net314;
 wire net285;
 wire net284;
 wire net283;
 wire net282;
 wire net281;
 wire net280;
 wire net279;
 wire net278;
 wire net277;
 wire net276;
 wire net275;
 wire net274;
 wire net273;
 wire net272;
 wire net271;
 wire net270;
 wire net269;
 wire net268;
 wire net267;
 wire net266;
 wire net265;
 wire net264;
 wire net291;
 wire net290;
 wire net289;
 wire net288;
 wire net287;
 wire net286;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire clknet_leaf_0_clock;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net392;
 wire net391;
 wire net390;
 wire net389;
 wire net388;
 wire net387;
 wire net386;
 wire net385;
 wire net384;
 wire net383;
 wire net382;
 wire net381;
 wire net380;
 wire net379;
 wire net378;
 wire net377;
 wire net376;
 wire clknet_leaf_1_clock;
 wire clknet_leaf_2_clock;
 wire clknet_leaf_6_clock;
 wire clknet_leaf_8_clock;
 wire clknet_leaf_10_clock;
 wire clknet_leaf_15_clock;
 wire clknet_leaf_16_clock;
 wire clknet_leaf_17_clock;
 wire clknet_leaf_18_clock;
 wire clknet_leaf_19_clock;
 wire clknet_leaf_22_clock;
 wire clknet_leaf_23_clock;
 wire clknet_leaf_24_clock;
 wire clknet_leaf_25_clock;
 wire clknet_leaf_26_clock;
 wire clknet_leaf_27_clock;
 wire clknet_leaf_31_clock;
 wire clknet_leaf_33_clock;
 wire clknet_0_clock;
 wire clknet_2_0__leaf_clock;
 wire clknet_2_1__leaf_clock;
 wire clknet_2_2__leaf_clock;
 wire clknet_2_3__leaf_clock;

 BUFx2_ASAP7_75t_R clkload24 (.A(clknet_leaf_15_clock));
 BUFx2_ASAP7_75t_R clkload23 (.A(clknet_leaf_13_clock));
 BUFx4f_ASAP7_75t_R clkload22 (.A(clknet_leaf_12_clock));
 BUFx2_ASAP7_75t_R clkload21 (.A(clknet_leaf_11_clock));
 BUFx4f_ASAP7_75t_R clkload20 (.A(clknet_leaf_10_clock));
 BUFx2_ASAP7_75t_R clkload19 (.A(clknet_leaf_7_clock));
 BUFx2_ASAP7_75t_R clkload18 (.A(clknet_leaf_6_clock));
 BUFx4f_ASAP7_75t_R clkload17 (.A(clknet_leaf_5_clock));
 BUFx2_ASAP7_75t_R clkload16 (.A(clknet_leaf_4_clock));
 BUFx2_ASAP7_75t_R clkload15 (.A(clknet_leaf_29_clock));
 BUFx2_ASAP7_75t_R clkload14 (.A(clknet_leaf_27_clock));
 BUFx2_ASAP7_75t_R clkload13 (.A(clknet_leaf_25_clock));
 BUFx2_ASAP7_75t_R clkload12 (.A(clknet_leaf_24_clock));
 BUFx2_ASAP7_75t_R clkload11 (.A(clknet_leaf_23_clock));
 BUFx4f_ASAP7_75t_R clkload10 (.A(clknet_leaf_22_clock));
 BUFx4f_ASAP7_75t_R clkload9 (.A(clknet_leaf_21_clock));
 BUFx24_ASAP7_75t_R clkload8 (.A(clknet_leaf_33_clock));
 BUFx2_ASAP7_75t_R clkload7 (.A(clknet_leaf_32_clock));
 BUFx4f_ASAP7_75t_R clkload6 (.A(clknet_leaf_31_clock));
 BUFx2_ASAP7_75t_R clkload5 (.A(clknet_leaf_3_clock));
 BUFx4f_ASAP7_75t_R clkload4 (.A(clknet_leaf_2_clock));
 BUFx2_ASAP7_75t_R clkload3 (.A(clknet_leaf_1_clock));
 BUFx4f_ASAP7_75t_R clkload2 (.A(clknet_leaf_0_clock));
 BUFx8_ASAP7_75t_R clkload1 (.A(clknet_2_3__leaf_clock));
 BUFx8_ASAP7_75t_R clkload0 (.A(clknet_2_0__leaf_clock));
 BUFx4_ASAP7_75t_R clkbuf_2_3__f_clock (.A(clknet_0_clock),
    .Y(clknet_2_3__leaf_clock));
 BUFx4_ASAP7_75t_R clkbuf_2_2__f_clock (.A(clknet_0_clock),
    .Y(clknet_2_2__leaf_clock));
 BUFx4_ASAP7_75t_R clkbuf_2_1__f_clock (.A(clknet_0_clock),
    .Y(clknet_2_1__leaf_clock));
 BUFx4_ASAP7_75t_R clkbuf_2_0__f_clock (.A(clknet_0_clock),
    .Y(clknet_2_0__leaf_clock));
 BUFx4_ASAP7_75t_R clkbuf_0_clock (.A(clock),
    .Y(clknet_0_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_33_clock (.A(clknet_2_0__leaf_clock),
    .Y(clknet_leaf_33_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_32_clock (.A(clknet_2_0__leaf_clock),
    .Y(clknet_leaf_32_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_31_clock (.A(clknet_2_0__leaf_clock),
    .Y(clknet_leaf_31_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_30_clock (.A(clknet_2_0__leaf_clock),
    .Y(clknet_leaf_30_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_29_clock (.A(clknet_2_1__leaf_clock),
    .Y(clknet_leaf_29_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_28_clock (.A(clknet_2_1__leaf_clock),
    .Y(clknet_leaf_28_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_27_clock (.A(clknet_2_1__leaf_clock),
    .Y(clknet_leaf_27_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_26_clock (.A(clknet_2_1__leaf_clock),
    .Y(clknet_leaf_26_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_25_clock (.A(clknet_2_1__leaf_clock),
    .Y(clknet_leaf_25_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_24_clock (.A(clknet_2_1__leaf_clock),
    .Y(clknet_leaf_24_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_23_clock (.A(clknet_2_1__leaf_clock),
    .Y(clknet_leaf_23_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_22_clock (.A(clknet_2_1__leaf_clock),
    .Y(clknet_leaf_22_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_21_clock (.A(clknet_2_1__leaf_clock),
    .Y(clknet_leaf_21_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_20_clock (.A(clknet_2_3__leaf_clock),
    .Y(clknet_leaf_20_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_19_clock (.A(clknet_2_3__leaf_clock),
    .Y(clknet_leaf_19_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_18_clock (.A(clknet_2_3__leaf_clock),
    .Y(clknet_leaf_18_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_17_clock (.A(clknet_2_3__leaf_clock),
    .Y(clknet_leaf_17_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_16_clock (.A(clknet_2_3__leaf_clock),
    .Y(clknet_leaf_16_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_15_clock (.A(clknet_2_3__leaf_clock),
    .Y(clknet_leaf_15_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_14_clock (.A(clknet_2_3__leaf_clock),
    .Y(clknet_leaf_14_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_13_clock (.A(clknet_2_3__leaf_clock),
    .Y(clknet_leaf_13_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_12_clock (.A(clknet_2_2__leaf_clock),
    .Y(clknet_leaf_12_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_11_clock (.A(clknet_2_2__leaf_clock),
    .Y(clknet_leaf_11_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_10_clock (.A(clknet_2_2__leaf_clock),
    .Y(clknet_leaf_10_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_9_clock (.A(clknet_2_2__leaf_clock),
    .Y(clknet_leaf_9_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_8_clock (.A(clknet_2_2__leaf_clock),
    .Y(clknet_leaf_8_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_7_clock (.A(clknet_2_2__leaf_clock),
    .Y(clknet_leaf_7_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_6_clock (.A(clknet_2_2__leaf_clock),
    .Y(clknet_leaf_6_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_5_clock (.A(clknet_2_2__leaf_clock),
    .Y(clknet_leaf_5_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_4_clock (.A(clknet_2_2__leaf_clock),
    .Y(clknet_leaf_4_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_3_clock (.A(clknet_2_0__leaf_clock),
    .Y(clknet_leaf_3_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_2_clock (.A(clknet_2_0__leaf_clock),
    .Y(clknet_leaf_2_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_1_clock (.A(clknet_2_0__leaf_clock),
    .Y(clknet_leaf_1_clock));
 BUFx8_ASAP7_75t_R clkbuf_leaf_0_clock (.A(clknet_2_0__leaf_clock),
    .Y(clknet_leaf_0_clock));
 BUFx2_ASAP7_75t_R output529 (.A(net524),
    .Y(io_outs_up[9]));
 BUFx2_ASAP7_75t_R output528 (.A(net523),
    .Y(io_outs_up[8]));
 BUFx2_ASAP7_75t_R output527 (.A(net522),
    .Y(io_outs_up[7]));
 BUFx2_ASAP7_75t_R output526 (.A(net521),
    .Y(io_outs_up[6]));
 BUFx2_ASAP7_75t_R output525 (.A(net520),
    .Y(io_outs_up[5]));
 BUFx2_ASAP7_75t_R output524 (.A(net519),
    .Y(io_outs_up[4]));
 BUFx2_ASAP7_75t_R output523 (.A(net518),
    .Y(io_outs_up[3]));
 BUFx2_ASAP7_75t_R output522 (.A(net517),
    .Y(io_outs_up[31]));
 BUFx2_ASAP7_75t_R output521 (.A(net516),
    .Y(io_outs_up[30]));
 BUFx2_ASAP7_75t_R output520 (.A(net515),
    .Y(io_outs_up[2]));
 BUFx2_ASAP7_75t_R output519 (.A(net514),
    .Y(io_outs_up[29]));
 BUFx2_ASAP7_75t_R output518 (.A(net513),
    .Y(io_outs_up[28]));
 BUFx2_ASAP7_75t_R output517 (.A(net512),
    .Y(io_outs_up[27]));
 BUFx2_ASAP7_75t_R output516 (.A(net511),
    .Y(io_outs_up[26]));
 BUFx2_ASAP7_75t_R output515 (.A(net510),
    .Y(io_outs_up[25]));
 BUFx2_ASAP7_75t_R output514 (.A(net509),
    .Y(io_outs_up[24]));
 BUFx2_ASAP7_75t_R output513 (.A(net508),
    .Y(io_outs_up[23]));
 BUFx2_ASAP7_75t_R output512 (.A(net507),
    .Y(io_outs_up[22]));
 BUFx2_ASAP7_75t_R output511 (.A(net506),
    .Y(io_outs_up[21]));
 BUFx2_ASAP7_75t_R output510 (.A(net505),
    .Y(io_outs_up[20]));
 BUFx2_ASAP7_75t_R output509 (.A(net504),
    .Y(io_outs_up[1]));
 BUFx2_ASAP7_75t_R output508 (.A(net503),
    .Y(io_outs_up[19]));
 BUFx2_ASAP7_75t_R output507 (.A(net502),
    .Y(io_outs_up[18]));
 BUFx2_ASAP7_75t_R output506 (.A(net501),
    .Y(io_outs_up[17]));
 BUFx2_ASAP7_75t_R output505 (.A(net500),
    .Y(io_outs_up[16]));
 BUFx2_ASAP7_75t_R output504 (.A(net499),
    .Y(io_outs_up[15]));
 BUFx2_ASAP7_75t_R output503 (.A(net498),
    .Y(io_outs_up[14]));
 BUFx2_ASAP7_75t_R output502 (.A(net497),
    .Y(io_outs_up[13]));
 BUFx2_ASAP7_75t_R output501 (.A(net496),
    .Y(io_outs_up[12]));
 BUFx2_ASAP7_75t_R output500 (.A(net495),
    .Y(io_outs_up[11]));
 BUFx2_ASAP7_75t_R output499 (.A(net494),
    .Y(io_outs_up[10]));
 BUFx2_ASAP7_75t_R output498 (.A(net493),
    .Y(io_outs_up[0]));
 BUFx2_ASAP7_75t_R output497 (.A(net492),
    .Y(io_outs_right[9]));
 BUFx2_ASAP7_75t_R output496 (.A(net491),
    .Y(io_outs_right[8]));
 BUFx2_ASAP7_75t_R output495 (.A(net490),
    .Y(io_outs_right[7]));
 BUFx2_ASAP7_75t_R output494 (.A(net489),
    .Y(io_outs_right[6]));
 BUFx2_ASAP7_75t_R output493 (.A(net488),
    .Y(io_outs_right[5]));
 BUFx2_ASAP7_75t_R output492 (.A(net487),
    .Y(io_outs_right[4]));
 BUFx2_ASAP7_75t_R output491 (.A(net486),
    .Y(io_outs_right[3]));
 BUFx2_ASAP7_75t_R output490 (.A(net485),
    .Y(io_outs_right[31]));
 BUFx2_ASAP7_75t_R output489 (.A(net484),
    .Y(io_outs_right[30]));
 BUFx2_ASAP7_75t_R output488 (.A(net483),
    .Y(io_outs_right[2]));
 BUFx2_ASAP7_75t_R output487 (.A(net482),
    .Y(io_outs_right[29]));
 BUFx2_ASAP7_75t_R output486 (.A(net481),
    .Y(io_outs_right[28]));
 BUFx2_ASAP7_75t_R output485 (.A(net480),
    .Y(io_outs_right[27]));
 BUFx2_ASAP7_75t_R output484 (.A(net479),
    .Y(io_outs_right[26]));
 BUFx2_ASAP7_75t_R output483 (.A(net478),
    .Y(io_outs_right[25]));
 BUFx2_ASAP7_75t_R output482 (.A(net477),
    .Y(io_outs_right[24]));
 BUFx2_ASAP7_75t_R output481 (.A(net476),
    .Y(io_outs_right[23]));
 BUFx2_ASAP7_75t_R output480 (.A(net475),
    .Y(io_outs_right[22]));
 BUFx2_ASAP7_75t_R output479 (.A(net474),
    .Y(io_outs_right[21]));
 BUFx2_ASAP7_75t_R output478 (.A(net473),
    .Y(io_outs_right[20]));
 BUFx2_ASAP7_75t_R output477 (.A(net472),
    .Y(io_outs_right[1]));
 BUFx2_ASAP7_75t_R output476 (.A(net471),
    .Y(io_outs_right[19]));
 BUFx2_ASAP7_75t_R output475 (.A(net470),
    .Y(io_outs_right[18]));
 BUFx2_ASAP7_75t_R output474 (.A(net469),
    .Y(io_outs_right[17]));
 BUFx2_ASAP7_75t_R output473 (.A(net468),
    .Y(io_outs_right[16]));
 BUFx2_ASAP7_75t_R output472 (.A(net467),
    .Y(io_outs_right[15]));
 BUFx2_ASAP7_75t_R output471 (.A(net466),
    .Y(io_outs_right[14]));
 BUFx2_ASAP7_75t_R output470 (.A(net465),
    .Y(io_outs_right[13]));
 BUFx2_ASAP7_75t_R output469 (.A(net464),
    .Y(io_outs_right[12]));
 BUFx2_ASAP7_75t_R output468 (.A(net463),
    .Y(io_outs_right[11]));
 BUFx2_ASAP7_75t_R output467 (.A(net462),
    .Y(io_outs_right[10]));
 BUFx2_ASAP7_75t_R output466 (.A(net461),
    .Y(io_outs_right[0]));
 BUFx2_ASAP7_75t_R output465 (.A(net460),
    .Y(io_outs_left[9]));
 BUFx2_ASAP7_75t_R output464 (.A(net459),
    .Y(io_outs_left[8]));
 BUFx2_ASAP7_75t_R output463 (.A(net458),
    .Y(io_outs_left[7]));
 BUFx2_ASAP7_75t_R output462 (.A(net457),
    .Y(io_outs_left[6]));
 BUFx2_ASAP7_75t_R output461 (.A(net456),
    .Y(io_outs_left[5]));
 BUFx2_ASAP7_75t_R output460 (.A(net455),
    .Y(io_outs_left[4]));
 BUFx2_ASAP7_75t_R output459 (.A(net454),
    .Y(io_outs_left[3]));
 BUFx2_ASAP7_75t_R output458 (.A(net453),
    .Y(io_outs_left[31]));
 BUFx2_ASAP7_75t_R output457 (.A(net452),
    .Y(io_outs_left[30]));
 BUFx2_ASAP7_75t_R output456 (.A(net451),
    .Y(io_outs_left[2]));
 BUFx2_ASAP7_75t_R output455 (.A(net450),
    .Y(io_outs_left[29]));
 BUFx2_ASAP7_75t_R output454 (.A(net449),
    .Y(io_outs_left[28]));
 BUFx2_ASAP7_75t_R output453 (.A(net448),
    .Y(io_outs_left[27]));
 BUFx2_ASAP7_75t_R output452 (.A(net447),
    .Y(io_outs_left[26]));
 BUFx2_ASAP7_75t_R output451 (.A(net446),
    .Y(io_outs_left[25]));
 BUFx2_ASAP7_75t_R output450 (.A(net445),
    .Y(io_outs_left[24]));
 BUFx2_ASAP7_75t_R output449 (.A(net444),
    .Y(io_outs_left[23]));
 BUFx2_ASAP7_75t_R output448 (.A(net443),
    .Y(io_outs_left[22]));
 BUFx2_ASAP7_75t_R output447 (.A(net442),
    .Y(io_outs_left[21]));
 BUFx2_ASAP7_75t_R output446 (.A(net441),
    .Y(io_outs_left[20]));
 BUFx2_ASAP7_75t_R output445 (.A(net440),
    .Y(io_outs_left[1]));
 BUFx2_ASAP7_75t_R output444 (.A(net439),
    .Y(io_outs_left[19]));
 BUFx2_ASAP7_75t_R output443 (.A(net438),
    .Y(io_outs_left[18]));
 BUFx2_ASAP7_75t_R output442 (.A(net437),
    .Y(io_outs_left[17]));
 BUFx2_ASAP7_75t_R output441 (.A(net436),
    .Y(io_outs_left[16]));
 BUFx2_ASAP7_75t_R output440 (.A(net435),
    .Y(io_outs_left[15]));
 BUFx2_ASAP7_75t_R output439 (.A(net434),
    .Y(io_outs_left[14]));
 BUFx2_ASAP7_75t_R output438 (.A(net433),
    .Y(io_outs_left[13]));
 BUFx2_ASAP7_75t_R output437 (.A(net432),
    .Y(io_outs_left[12]));
 BUFx2_ASAP7_75t_R output436 (.A(net431),
    .Y(io_outs_left[11]));
 BUFx2_ASAP7_75t_R output435 (.A(net430),
    .Y(io_outs_left[10]));
 BUFx2_ASAP7_75t_R output434 (.A(net396),
    .Y(io_outs_left[0]));
 BUFx2_ASAP7_75t_R output433 (.A(net428),
    .Y(io_outs_down[9]));
 BUFx2_ASAP7_75t_R output432 (.A(net427),
    .Y(io_outs_down[8]));
 BUFx2_ASAP7_75t_R output431 (.A(net426),
    .Y(io_outs_down[7]));
 BUFx2_ASAP7_75t_R output430 (.A(net425),
    .Y(io_outs_down[6]));
 BUFx2_ASAP7_75t_R output429 (.A(net424),
    .Y(io_outs_down[5]));
 BUFx2_ASAP7_75t_R output428 (.A(net423),
    .Y(io_outs_down[4]));
 BUFx2_ASAP7_75t_R output427 (.A(net422),
    .Y(io_outs_down[3]));
 BUFx2_ASAP7_75t_R output426 (.A(net421),
    .Y(io_outs_down[31]));
 BUFx2_ASAP7_75t_R output425 (.A(net420),
    .Y(io_outs_down[30]));
 BUFx2_ASAP7_75t_R output424 (.A(net419),
    .Y(io_outs_down[2]));
 BUFx2_ASAP7_75t_R output423 (.A(net418),
    .Y(io_outs_down[29]));
 BUFx2_ASAP7_75t_R output422 (.A(net417),
    .Y(io_outs_down[28]));
 BUFx2_ASAP7_75t_R output421 (.A(net416),
    .Y(io_outs_down[27]));
 BUFx2_ASAP7_75t_R output420 (.A(net415),
    .Y(io_outs_down[26]));
 BUFx2_ASAP7_75t_R output419 (.A(net414),
    .Y(io_outs_down[25]));
 BUFx2_ASAP7_75t_R output418 (.A(net413),
    .Y(io_outs_down[24]));
 BUFx2_ASAP7_75t_R output417 (.A(net412),
    .Y(io_outs_down[23]));
 BUFx2_ASAP7_75t_R output416 (.A(net411),
    .Y(io_outs_down[22]));
 BUFx2_ASAP7_75t_R output415 (.A(net410),
    .Y(io_outs_down[21]));
 BUFx2_ASAP7_75t_R output414 (.A(net409),
    .Y(io_outs_down[20]));
 BUFx2_ASAP7_75t_R output413 (.A(net408),
    .Y(io_outs_down[1]));
 BUFx2_ASAP7_75t_R output412 (.A(net407),
    .Y(io_outs_down[19]));
 BUFx2_ASAP7_75t_R output411 (.A(net406),
    .Y(io_outs_down[18]));
 BUFx2_ASAP7_75t_R output410 (.A(net405),
    .Y(io_outs_down[17]));
 BUFx2_ASAP7_75t_R output409 (.A(net404),
    .Y(io_outs_down[16]));
 BUFx2_ASAP7_75t_R output408 (.A(net403),
    .Y(io_outs_down[15]));
 BUFx2_ASAP7_75t_R output407 (.A(net402),
    .Y(io_outs_down[14]));
 BUFx2_ASAP7_75t_R output406 (.A(net401),
    .Y(io_outs_down[13]));
 BUFx2_ASAP7_75t_R output405 (.A(net400),
    .Y(io_outs_down[12]));
 BUFx2_ASAP7_75t_R output404 (.A(net399),
    .Y(io_outs_down[11]));
 BUFx2_ASAP7_75t_R output403 (.A(net398),
    .Y(io_outs_down[10]));
 BUFx2_ASAP7_75t_R output402 (.A(net397),
    .Y(io_outs_down[0]));
 BUFx2_ASAP7_75t_R output401 (.A(net396),
    .Y(io_lsbOuts_3));
 BUFx2_ASAP7_75t_R output400 (.A(net395),
    .Y(io_lsbOuts_2));
 BUFx2_ASAP7_75t_R output399 (.A(net394),
    .Y(io_lsbOuts_1));
 BUFx2_ASAP7_75t_R output398 (.A(net393),
    .Y(io_lsbOuts_0));
 BUFx2_ASAP7_75t_R input397 (.A(io_lsbIns_2),
    .Y(net392));
 BUFx2_ASAP7_75t_R input396 (.A(io_ins_up[9]),
    .Y(net391));
 BUFx2_ASAP7_75t_R input395 (.A(io_ins_up[8]),
    .Y(net390));
 BUFx2_ASAP7_75t_R input394 (.A(io_ins_up[7]),
    .Y(net389));
 BUFx2_ASAP7_75t_R input393 (.A(io_ins_up[6]),
    .Y(net388));
 BUFx2_ASAP7_75t_R input392 (.A(io_ins_up[5]),
    .Y(net387));
 BUFx2_ASAP7_75t_R input391 (.A(io_ins_up[4]),
    .Y(net386));
 BUFx2_ASAP7_75t_R input390 (.A(io_ins_up[3]),
    .Y(net385));
 BUFx2_ASAP7_75t_R input389 (.A(io_ins_up[31]),
    .Y(net384));
 BUFx2_ASAP7_75t_R input388 (.A(io_ins_up[30]),
    .Y(net383));
 BUFx2_ASAP7_75t_R input387 (.A(io_ins_up[2]),
    .Y(net382));
 BUFx2_ASAP7_75t_R input386 (.A(io_ins_up[29]),
    .Y(net381));
 BUFx2_ASAP7_75t_R input385 (.A(io_ins_up[28]),
    .Y(net380));
 BUFx2_ASAP7_75t_R input384 (.A(io_ins_up[27]),
    .Y(net379));
 BUFx2_ASAP7_75t_R input383 (.A(io_ins_up[26]),
    .Y(net378));
 BUFx2_ASAP7_75t_R input382 (.A(io_ins_up[25]),
    .Y(net377));
 BUFx2_ASAP7_75t_R input381 (.A(io_ins_up[24]),
    .Y(net376));
 BUFx2_ASAP7_75t_R input380 (.A(io_ins_up[23]),
    .Y(net375));
 BUFx2_ASAP7_75t_R input379 (.A(io_ins_up[22]),
    .Y(net374));
 BUFx2_ASAP7_75t_R input378 (.A(io_ins_up[21]),
    .Y(net373));
 BUFx2_ASAP7_75t_R input377 (.A(io_ins_up[20]),
    .Y(net372));
 BUFx2_ASAP7_75t_R input376 (.A(io_ins_up[1]),
    .Y(net371));
 BUFx2_ASAP7_75t_R input375 (.A(io_ins_up[19]),
    .Y(net370));
 BUFx2_ASAP7_75t_R input374 (.A(io_ins_up[18]),
    .Y(net369));
 BUFx2_ASAP7_75t_R input373 (.A(io_ins_up[17]),
    .Y(net368));
 BUFx2_ASAP7_75t_R input372 (.A(io_ins_up[16]),
    .Y(net367));
 BUFx2_ASAP7_75t_R input371 (.A(io_ins_up[15]),
    .Y(net366));
 BUFx2_ASAP7_75t_R input370 (.A(io_ins_up[14]),
    .Y(net365));
 BUFx2_ASAP7_75t_R input369 (.A(io_ins_up[13]),
    .Y(net364));
 BUFx2_ASAP7_75t_R input368 (.A(io_ins_up[12]),
    .Y(net363));
 BUFx2_ASAP7_75t_R input367 (.A(io_ins_up[11]),
    .Y(net362));
 BUFx2_ASAP7_75t_R input366 (.A(io_ins_up[10]),
    .Y(net361));
 BUFx2_ASAP7_75t_R input365 (.A(io_ins_up[0]),
    .Y(net360));
 BUFx2_ASAP7_75t_R input364 (.A(io_ins_right[9]),
    .Y(net359));
 BUFx2_ASAP7_75t_R input363 (.A(io_ins_right[8]),
    .Y(net358));
 BUFx2_ASAP7_75t_R input362 (.A(io_ins_right[7]),
    .Y(net357));
 BUFx2_ASAP7_75t_R input361 (.A(io_ins_right[6]),
    .Y(net356));
 BUFx2_ASAP7_75t_R input360 (.A(io_ins_right[5]),
    .Y(net355));
 BUFx2_ASAP7_75t_R input359 (.A(io_ins_right[4]),
    .Y(net354));
 BUFx2_ASAP7_75t_R input358 (.A(io_ins_right[3]),
    .Y(net353));
 BUFx2_ASAP7_75t_R input357 (.A(io_ins_right[31]),
    .Y(net352));
 BUFx2_ASAP7_75t_R input356 (.A(io_ins_right[30]),
    .Y(net351));
 BUFx2_ASAP7_75t_R input355 (.A(io_ins_right[2]),
    .Y(net350));
 BUFx2_ASAP7_75t_R input354 (.A(io_ins_right[29]),
    .Y(net349));
 BUFx2_ASAP7_75t_R input353 (.A(io_ins_right[28]),
    .Y(net348));
 BUFx2_ASAP7_75t_R input352 (.A(io_ins_right[27]),
    .Y(net347));
 BUFx2_ASAP7_75t_R input351 (.A(io_ins_right[26]),
    .Y(net346));
 BUFx2_ASAP7_75t_R input350 (.A(io_ins_right[25]),
    .Y(net345));
 BUFx2_ASAP7_75t_R input349 (.A(io_ins_right[24]),
    .Y(net344));
 BUFx2_ASAP7_75t_R input348 (.A(io_ins_right[23]),
    .Y(net343));
 BUFx2_ASAP7_75t_R input347 (.A(io_ins_right[22]),
    .Y(net342));
 BUFx2_ASAP7_75t_R input346 (.A(io_ins_right[21]),
    .Y(net341));
 BUFx2_ASAP7_75t_R input345 (.A(io_ins_right[20]),
    .Y(net340));
 BUFx2_ASAP7_75t_R input344 (.A(io_ins_right[1]),
    .Y(net339));
 BUFx2_ASAP7_75t_R input343 (.A(io_ins_right[19]),
    .Y(net338));
 BUFx2_ASAP7_75t_R input342 (.A(io_ins_right[18]),
    .Y(net337));
 BUFx2_ASAP7_75t_R input341 (.A(io_ins_right[17]),
    .Y(net336));
 BUFx2_ASAP7_75t_R input340 (.A(io_ins_right[16]),
    .Y(net335));
 BUFx2_ASAP7_75t_R input339 (.A(io_ins_right[15]),
    .Y(net334));
 BUFx2_ASAP7_75t_R input338 (.A(io_ins_right[14]),
    .Y(net333));
 BUFx2_ASAP7_75t_R input337 (.A(io_ins_right[13]),
    .Y(net332));
 BUFx2_ASAP7_75t_R input336 (.A(io_ins_right[12]),
    .Y(net331));
 BUFx2_ASAP7_75t_R input335 (.A(io_ins_right[11]),
    .Y(net330));
 BUFx2_ASAP7_75t_R input334 (.A(io_ins_right[10]),
    .Y(net329));
 BUFx2_ASAP7_75t_R input333 (.A(io_ins_right[0]),
    .Y(net328));
 BUFx2_ASAP7_75t_R input332 (.A(io_ins_left[9]),
    .Y(net327));
 BUFx2_ASAP7_75t_R input331 (.A(io_ins_left[8]),
    .Y(net326));
 BUFx2_ASAP7_75t_R input330 (.A(io_ins_left[7]),
    .Y(net325));
 BUFx2_ASAP7_75t_R input329 (.A(io_ins_left[6]),
    .Y(net324));
 BUFx2_ASAP7_75t_R input328 (.A(io_ins_left[5]),
    .Y(net323));
 BUFx2_ASAP7_75t_R input327 (.A(io_ins_left[4]),
    .Y(net322));
 BUFx2_ASAP7_75t_R input326 (.A(io_ins_left[3]),
    .Y(net321));
 BUFx2_ASAP7_75t_R input325 (.A(io_ins_left[31]),
    .Y(net320));
 BUFx2_ASAP7_75t_R input324 (.A(io_ins_left[30]),
    .Y(net319));
 BUFx2_ASAP7_75t_R input323 (.A(io_ins_left[2]),
    .Y(net318));
 BUFx2_ASAP7_75t_R input322 (.A(io_ins_left[29]),
    .Y(net317));
 BUFx2_ASAP7_75t_R input321 (.A(io_ins_left[28]),
    .Y(net316));
 BUFx2_ASAP7_75t_R input320 (.A(io_ins_left[27]),
    .Y(net315));
 BUFx2_ASAP7_75t_R input319 (.A(io_ins_left[26]),
    .Y(net314));
 BUFx2_ASAP7_75t_R input318 (.A(io_ins_left[25]),
    .Y(net313));
 BUFx2_ASAP7_75t_R input317 (.A(io_ins_left[24]),
    .Y(net312));
 BUFx2_ASAP7_75t_R input316 (.A(io_ins_left[23]),
    .Y(net311));
 BUFx2_ASAP7_75t_R input315 (.A(io_ins_left[22]),
    .Y(net310));
 BUFx2_ASAP7_75t_R input314 (.A(io_ins_left[21]),
    .Y(net309));
 BUFx2_ASAP7_75t_R input313 (.A(io_ins_left[20]),
    .Y(net308));
 BUFx2_ASAP7_75t_R input312 (.A(io_ins_left[1]),
    .Y(net307));
 BUFx2_ASAP7_75t_R input311 (.A(io_ins_left[19]),
    .Y(net306));
 BUFx2_ASAP7_75t_R input310 (.A(io_ins_left[18]),
    .Y(net305));
 BUFx2_ASAP7_75t_R input309 (.A(io_ins_left[17]),
    .Y(net304));
 BUFx2_ASAP7_75t_R input308 (.A(io_ins_left[16]),
    .Y(net303));
 BUFx2_ASAP7_75t_R input307 (.A(io_ins_left[15]),
    .Y(net302));
 BUFx2_ASAP7_75t_R input306 (.A(io_ins_left[14]),
    .Y(net301));
 BUFx2_ASAP7_75t_R input305 (.A(io_ins_left[13]),
    .Y(net300));
 BUFx2_ASAP7_75t_R input304 (.A(io_ins_left[12]),
    .Y(net299));
 BUFx2_ASAP7_75t_R input303 (.A(io_ins_left[11]),
    .Y(net298));
 BUFx2_ASAP7_75t_R input302 (.A(io_ins_left[10]),
    .Y(net297));
 BUFx2_ASAP7_75t_R input301 (.A(io_ins_left[0]),
    .Y(net296));
 BUFx2_ASAP7_75t_R input300 (.A(io_ins_down[9]),
    .Y(net295));
 BUFx2_ASAP7_75t_R input299 (.A(io_ins_down[8]),
    .Y(net294));
 BUFx2_ASAP7_75t_R input298 (.A(io_ins_down[7]),
    .Y(net293));
 BUFx2_ASAP7_75t_R input297 (.A(io_ins_down[6]),
    .Y(net292));
 BUFx2_ASAP7_75t_R input296 (.A(io_ins_down[5]),
    .Y(net291));
 BUFx2_ASAP7_75t_R input295 (.A(io_ins_down[4]),
    .Y(net290));
 BUFx2_ASAP7_75t_R input294 (.A(io_ins_down[3]),
    .Y(net289));
 BUFx2_ASAP7_75t_R input293 (.A(io_ins_down[31]),
    .Y(net288));
 BUFx2_ASAP7_75t_R input292 (.A(io_ins_down[30]),
    .Y(net287));
 BUFx2_ASAP7_75t_R input291 (.A(io_ins_down[2]),
    .Y(net286));
 BUFx2_ASAP7_75t_R input290 (.A(io_ins_down[29]),
    .Y(net285));
 BUFx2_ASAP7_75t_R input289 (.A(io_ins_down[28]),
    .Y(net284));
 BUFx2_ASAP7_75t_R input288 (.A(io_ins_down[27]),
    .Y(net283));
 BUFx2_ASAP7_75t_R input287 (.A(io_ins_down[26]),
    .Y(net282));
 BUFx2_ASAP7_75t_R input286 (.A(io_ins_down[25]),
    .Y(net281));
 BUFx2_ASAP7_75t_R input285 (.A(io_ins_down[24]),
    .Y(net280));
 BUFx2_ASAP7_75t_R input284 (.A(io_ins_down[23]),
    .Y(net279));
 BUFx2_ASAP7_75t_R input283 (.A(io_ins_down[22]),
    .Y(net278));
 BUFx2_ASAP7_75t_R input282 (.A(io_ins_down[21]),
    .Y(net277));
 BUFx2_ASAP7_75t_R input281 (.A(io_ins_down[20]),
    .Y(net276));
 BUFx2_ASAP7_75t_R input280 (.A(io_ins_down[1]),
    .Y(net275));
 BUFx2_ASAP7_75t_R input279 (.A(io_ins_down[19]),
    .Y(net274));
 BUFx2_ASAP7_75t_R input278 (.A(io_ins_down[18]),
    .Y(net273));
 BUFx2_ASAP7_75t_R input277 (.A(io_ins_down[17]),
    .Y(net272));
 BUFx2_ASAP7_75t_R input276 (.A(io_ins_down[16]),
    .Y(net271));
 BUFx2_ASAP7_75t_R input275 (.A(io_ins_down[15]),
    .Y(net270));
 BUFx2_ASAP7_75t_R input274 (.A(io_ins_down[14]),
    .Y(net269));
 BUFx2_ASAP7_75t_R input273 (.A(io_ins_down[13]),
    .Y(net268));
 BUFx2_ASAP7_75t_R input272 (.A(io_ins_down[12]),
    .Y(net267));
 BUFx2_ASAP7_75t_R input271 (.A(io_ins_down[11]),
    .Y(net266));
 BUFx2_ASAP7_75t_R input270 (.A(io_ins_down[10]),
    .Y(net265));
 BUFx2_ASAP7_75t_R input269 (.A(io_ins_down[0]),
    .Y(net264));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_55_Left_111 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_Left_110 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_Left_109 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_Left_108 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_Left_107 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_Left_106 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_Left_105 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_Left_104 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Left_103 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Left_102 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Left_101 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Left_100 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Left_99 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Left_98 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Left_97 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Left_96 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Left_95 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Left_94 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Left_93 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Left_92 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Left_91 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Left_90 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Left_89 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Left_88 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Left_87 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Left_86 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Left_85 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Left_84 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Left_83 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Left_82 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Left_81 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Left_80 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Left_79 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Left_78 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Left_77 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Left_76 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Left_75 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Left_74 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Left_73 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Left_72 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Left_71 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Left_70 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Left_69 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Left_68 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Left_67 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Left_66 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Left_65 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Left_64 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Left_63 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Left_62 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Left_61 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Left_60 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Left_59 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Left_58 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Left_57 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Left_56 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Right_0 ();
 TIELOx1_ASAP7_75t_R _646__128 (.L(io_outs_up[63]));
 TIELOx1_ASAP7_75t_R _645__127 (.L(io_outs_up[62]));
 TIELOx1_ASAP7_75t_R _644__126 (.L(io_outs_up[61]));
 TIELOx1_ASAP7_75t_R _643__125 (.L(io_outs_up[60]));
 TIELOx1_ASAP7_75t_R _642__124 (.L(io_outs_up[59]));
 TIELOx1_ASAP7_75t_R _641__123 (.L(io_outs_up[58]));
 TIELOx1_ASAP7_75t_R _640__122 (.L(io_outs_up[57]));
 TIELOx1_ASAP7_75t_R _639__121 (.L(io_outs_up[56]));
 TIELOx1_ASAP7_75t_R _638__120 (.L(io_outs_up[55]));
 TIELOx1_ASAP7_75t_R _637__119 (.L(io_outs_up[54]));
 TIELOx1_ASAP7_75t_R _636__118 (.L(io_outs_up[53]));
 TIELOx1_ASAP7_75t_R _635__117 (.L(io_outs_up[52]));
 TIELOx1_ASAP7_75t_R _634__116 (.L(io_outs_up[51]));
 TIELOx1_ASAP7_75t_R _633__115 (.L(io_outs_up[50]));
 TIELOx1_ASAP7_75t_R _632__114 (.L(io_outs_up[49]));
 TIELOx1_ASAP7_75t_R _631__113 (.L(io_outs_up[48]));
 TIELOx1_ASAP7_75t_R _630__112 (.L(io_outs_up[47]));
 TIELOx1_ASAP7_75t_R _629__111 (.L(io_outs_up[46]));
 TIELOx1_ASAP7_75t_R _628__110 (.L(io_outs_up[45]));
 TIELOx1_ASAP7_75t_R _627__109 (.L(io_outs_up[44]));
 TIELOx1_ASAP7_75t_R _626__108 (.L(io_outs_up[43]));
 TIELOx1_ASAP7_75t_R _625__107 (.L(io_outs_up[42]));
 TIELOx1_ASAP7_75t_R _624__106 (.L(io_outs_up[41]));
 TIELOx1_ASAP7_75t_R _623__105 (.L(io_outs_up[40]));
 TIELOx1_ASAP7_75t_R _622__104 (.L(io_outs_up[39]));
 TIELOx1_ASAP7_75t_R _621__103 (.L(io_outs_up[38]));
 TIELOx1_ASAP7_75t_R _620__102 (.L(io_outs_up[37]));
 TIELOx1_ASAP7_75t_R _619__101 (.L(io_outs_up[36]));
 TIELOx1_ASAP7_75t_R _618__100 (.L(io_outs_up[35]));
 TIELOx1_ASAP7_75t_R _617__99 (.L(io_outs_up[34]));
 TIELOx1_ASAP7_75t_R _616__98 (.L(io_outs_up[33]));
 TIELOx1_ASAP7_75t_R _615__97 (.L(io_outs_up[32]));
 TIELOx1_ASAP7_75t_R _614__96 (.L(io_outs_right[63]));
 TIELOx1_ASAP7_75t_R _613__95 (.L(io_outs_right[62]));
 TIELOx1_ASAP7_75t_R _612__94 (.L(io_outs_right[61]));
 TIELOx1_ASAP7_75t_R _611__93 (.L(io_outs_right[60]));
 TIELOx1_ASAP7_75t_R _610__92 (.L(io_outs_right[59]));
 TIELOx1_ASAP7_75t_R _609__91 (.L(io_outs_right[58]));
 TIELOx1_ASAP7_75t_R _608__90 (.L(io_outs_right[57]));
 TIELOx1_ASAP7_75t_R _607__89 (.L(io_outs_right[56]));
 TIELOx1_ASAP7_75t_R _606__88 (.L(io_outs_right[55]));
 TIELOx1_ASAP7_75t_R _605__87 (.L(io_outs_right[54]));
 TIELOx1_ASAP7_75t_R _604__86 (.L(io_outs_right[53]));
 TIELOx1_ASAP7_75t_R _603__85 (.L(io_outs_right[52]));
 TIELOx1_ASAP7_75t_R _602__84 (.L(io_outs_right[51]));
 TIELOx1_ASAP7_75t_R _601__83 (.L(io_outs_right[50]));
 TIELOx1_ASAP7_75t_R _600__82 (.L(io_outs_right[49]));
 TIELOx1_ASAP7_75t_R _599__81 (.L(io_outs_right[48]));
 TIELOx1_ASAP7_75t_R _598__80 (.L(io_outs_right[47]));
 TIELOx1_ASAP7_75t_R _597__79 (.L(io_outs_right[46]));
 TIELOx1_ASAP7_75t_R _596__78 (.L(io_outs_right[45]));
 TIELOx1_ASAP7_75t_R _595__77 (.L(io_outs_right[44]));
 TIELOx1_ASAP7_75t_R _594__76 (.L(io_outs_right[43]));
 TIELOx1_ASAP7_75t_R _593__75 (.L(io_outs_right[42]));
 TIELOx1_ASAP7_75t_R _592__74 (.L(io_outs_right[41]));
 TIELOx1_ASAP7_75t_R _591__73 (.L(io_outs_right[40]));
 TIELOx1_ASAP7_75t_R _590__72 (.L(io_outs_right[39]));
 TIELOx1_ASAP7_75t_R _589__71 (.L(io_outs_right[38]));
 TIELOx1_ASAP7_75t_R _588__70 (.L(io_outs_right[37]));
 TIELOx1_ASAP7_75t_R _587__69 (.L(io_outs_right[36]));
 TIELOx1_ASAP7_75t_R _586__68 (.L(io_outs_right[35]));
 TIELOx1_ASAP7_75t_R _585__67 (.L(io_outs_right[34]));
 TIELOx1_ASAP7_75t_R _584__66 (.L(io_outs_right[33]));
 TIELOx1_ASAP7_75t_R _583__65 (.L(io_outs_right[32]));
 TIELOx1_ASAP7_75t_R _582__64 (.L(io_outs_left[63]));
 TIELOx1_ASAP7_75t_R _581__63 (.L(io_outs_left[62]));
 TIELOx1_ASAP7_75t_R _580__62 (.L(io_outs_left[61]));
 TIELOx1_ASAP7_75t_R _579__61 (.L(io_outs_left[60]));
 TIELOx1_ASAP7_75t_R _578__60 (.L(io_outs_left[59]));
 TIELOx1_ASAP7_75t_R _577__59 (.L(io_outs_left[58]));
 TIELOx1_ASAP7_75t_R _576__58 (.L(io_outs_left[57]));
 TIELOx1_ASAP7_75t_R _575__57 (.L(io_outs_left[56]));
 TIELOx1_ASAP7_75t_R _574__56 (.L(io_outs_left[55]));
 TIELOx1_ASAP7_75t_R _573__55 (.L(io_outs_left[54]));
 TIELOx1_ASAP7_75t_R _572__54 (.L(io_outs_left[53]));
 TIELOx1_ASAP7_75t_R _571__53 (.L(io_outs_left[52]));
 TIELOx1_ASAP7_75t_R _570__52 (.L(io_outs_left[51]));
 TIELOx1_ASAP7_75t_R _569__51 (.L(io_outs_left[50]));
 TIELOx1_ASAP7_75t_R _568__50 (.L(io_outs_left[49]));
 TIELOx1_ASAP7_75t_R _567__49 (.L(io_outs_left[48]));
 TIELOx1_ASAP7_75t_R _566__48 (.L(io_outs_left[47]));
 TIELOx1_ASAP7_75t_R _565__47 (.L(io_outs_left[46]));
 TIELOx1_ASAP7_75t_R _564__46 (.L(io_outs_left[45]));
 TIELOx1_ASAP7_75t_R _563__45 (.L(io_outs_left[44]));
 TIELOx1_ASAP7_75t_R _562__44 (.L(io_outs_left[43]));
 TIELOx1_ASAP7_75t_R _561__43 (.L(io_outs_left[42]));
 TIELOx1_ASAP7_75t_R _560__42 (.L(io_outs_left[41]));
 TIELOx1_ASAP7_75t_R _559__41 (.L(io_outs_left[40]));
 TIELOx1_ASAP7_75t_R _558__40 (.L(io_outs_left[39]));
 TIELOx1_ASAP7_75t_R _557__39 (.L(io_outs_left[38]));
 TIELOx1_ASAP7_75t_R _556__38 (.L(io_outs_left[37]));
 TIELOx1_ASAP7_75t_R _555__37 (.L(io_outs_left[36]));
 TIELOx1_ASAP7_75t_R _554__36 (.L(io_outs_left[35]));
 TIELOx1_ASAP7_75t_R _553__35 (.L(io_outs_left[34]));
 TIELOx1_ASAP7_75t_R _552__34 (.L(io_outs_left[33]));
 TIELOx1_ASAP7_75t_R _551__33 (.L(io_outs_left[32]));
 TIELOx1_ASAP7_75t_R _549__32 (.L(io_outs_down[63]));
 TIELOx1_ASAP7_75t_R _548__31 (.L(io_outs_down[62]));
 TIELOx1_ASAP7_75t_R _547__30 (.L(io_outs_down[61]));
 TIELOx1_ASAP7_75t_R _546__29 (.L(io_outs_down[60]));
 TIELOx1_ASAP7_75t_R _545__28 (.L(io_outs_down[59]));
 TIELOx1_ASAP7_75t_R _544__27 (.L(io_outs_down[58]));
 TIELOx1_ASAP7_75t_R _543__26 (.L(io_outs_down[57]));
 TIELOx1_ASAP7_75t_R _542__25 (.L(io_outs_down[56]));
 TIELOx1_ASAP7_75t_R _541__24 (.L(io_outs_down[55]));
 TIELOx1_ASAP7_75t_R _540__23 (.L(io_outs_down[54]));
 TIELOx1_ASAP7_75t_R _539__22 (.L(io_outs_down[53]));
 TIELOx1_ASAP7_75t_R _538__21 (.L(io_outs_down[52]));
 TIELOx1_ASAP7_75t_R _537__20 (.L(io_outs_down[51]));
 TIELOx1_ASAP7_75t_R _536__19 (.L(io_outs_down[50]));
 TIELOx1_ASAP7_75t_R _535__18 (.L(io_outs_down[49]));
 TIELOx1_ASAP7_75t_R _534__17 (.L(io_outs_down[48]));
 TIELOx1_ASAP7_75t_R _533__16 (.L(io_outs_down[47]));
 TIELOx1_ASAP7_75t_R _532__15 (.L(io_outs_down[46]));
 TIELOx1_ASAP7_75t_R _531__14 (.L(io_outs_down[45]));
 TIELOx1_ASAP7_75t_R _530__13 (.L(io_outs_down[44]));
 TIELOx1_ASAP7_75t_R _529__12 (.L(io_outs_down[43]));
 TIELOx1_ASAP7_75t_R _528__11 (.L(io_outs_down[42]));
 TIELOx1_ASAP7_75t_R _527__10 (.L(io_outs_down[41]));
 TIELOx1_ASAP7_75t_R _526__9 (.L(io_outs_down[40]));
 TIELOx1_ASAP7_75t_R _525__8 (.L(io_outs_down[39]));
 TIELOx1_ASAP7_75t_R _524__7 (.L(io_outs_down[38]));
 TIELOx1_ASAP7_75t_R _523__6 (.L(io_outs_down[37]));
 TIELOx1_ASAP7_75t_R _522__5 (.L(io_outs_down[36]));
 TIELOx1_ASAP7_75t_R _521__4 (.L(io_outs_down[35]));
 TIELOx1_ASAP7_75t_R _520__3 (.L(io_outs_down[34]));
 TIELOx1_ASAP7_75t_R _519__2 (.L(io_outs_down[33]));
 TIELOx1_ASAP7_75t_R _518__1 (.L(io_outs_down[32]));
 DFFHQNx1_ASAP7_75t_R \REG[0]$_DFF_P_  (.CLK(clknet_leaf_13_clock),
    .D(net264),
    .QN(_001_));
 DFFHQNx1_ASAP7_75t_R \REG[10]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(net265),
    .QN(_002_));
 DFFHQNx1_ASAP7_75t_R \REG[11]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(net266),
    .QN(_003_));
 DFFHQNx1_ASAP7_75t_R \REG[12]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net267),
    .QN(_004_));
 DFFHQNx1_ASAP7_75t_R \REG[13]$_DFF_P_  (.CLK(clknet_leaf_9_clock),
    .D(net268),
    .QN(_005_));
 DFFHQNx1_ASAP7_75t_R \REG[14]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(net269),
    .QN(_006_));
 DFFHQNx1_ASAP7_75t_R \REG[15]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(net270),
    .QN(_007_));
 DFFHQNx1_ASAP7_75t_R \REG[16]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(net271),
    .QN(_008_));
 DFFHQNx1_ASAP7_75t_R \REG[17]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(net272),
    .QN(_009_));
 DFFHQNx1_ASAP7_75t_R \REG[18]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net273),
    .QN(_010_));
 DFFHQNx1_ASAP7_75t_R \REG[19]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(net274),
    .QN(_011_));
 DFFHQNx1_ASAP7_75t_R \REG[1]$_DFF_P_  (.CLK(clknet_leaf_11_clock),
    .D(net275),
    .QN(_012_));
 DFFHQNx1_ASAP7_75t_R \REG[20]$_DFF_P_  (.CLK(clknet_leaf_14_clock),
    .D(net276),
    .QN(_013_));
 DFFHQNx1_ASAP7_75t_R \REG[21]$_DFF_P_  (.CLK(clknet_leaf_9_clock),
    .D(net277),
    .QN(_014_));
 DFFHQNx1_ASAP7_75t_R \REG[22]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net278),
    .QN(_015_));
 DFFHQNx1_ASAP7_75t_R \REG[23]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(net279),
    .QN(_016_));
 DFFHQNx1_ASAP7_75t_R \REG[24]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(net280),
    .QN(_017_));
 DFFHQNx1_ASAP7_75t_R \REG[25]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(net281),
    .QN(_018_));
 DFFHQNx1_ASAP7_75t_R \REG[26]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(net282),
    .QN(_019_));
 DFFHQNx1_ASAP7_75t_R \REG[27]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net283),
    .QN(_020_));
 DFFHQNx1_ASAP7_75t_R \REG[28]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(net284),
    .QN(_021_));
 DFFHQNx1_ASAP7_75t_R \REG[29]$_DFF_P_  (.CLK(clknet_leaf_14_clock),
    .D(net285),
    .QN(_022_));
 DFFHQNx1_ASAP7_75t_R \REG[2]$_DFF_P_  (.CLK(clknet_leaf_11_clock),
    .D(net286),
    .QN(_023_));
 DFFHQNx1_ASAP7_75t_R \REG[30]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(net287),
    .QN(_024_));
 DFFHQNx1_ASAP7_75t_R \REG[31]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(net288),
    .QN(_025_));
 DFFHQNx1_ASAP7_75t_R \REG[3]$_DFF_P_  (.CLK(clknet_leaf_11_clock),
    .D(net289),
    .QN(_026_));
 DFFHQNx1_ASAP7_75t_R \REG[4]$_DFF_P_  (.CLK(clknet_leaf_14_clock),
    .D(net290),
    .QN(_027_));
 DFFHQNx1_ASAP7_75t_R \REG[5]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net291),
    .QN(_028_));
 DFFHQNx1_ASAP7_75t_R \REG[6]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(net292),
    .QN(_029_));
 DFFHQNx1_ASAP7_75t_R \REG[7]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(net293),
    .QN(_030_));
 DFFHQNx1_ASAP7_75t_R \REG[8]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(net294),
    .QN(_031_));
 DFFHQNx1_ASAP7_75t_R \REG[9]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(net295),
    .QN(_032_));
 DFFHQNx1_ASAP7_75t_R \REG_1[0]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(net296),
    .QN(_033_));
 DFFHQNx1_ASAP7_75t_R \REG_1[10]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(net297),
    .QN(_034_));
 DFFHQNx1_ASAP7_75t_R \REG_1[11]$_DFF_P_  (.CLK(clknet_leaf_23_clock),
    .D(net298),
    .QN(_035_));
 DFFHQNx1_ASAP7_75t_R \REG_1[12]$_DFF_P_  (.CLK(clknet_leaf_23_clock),
    .D(net299),
    .QN(_036_));
 DFFHQNx1_ASAP7_75t_R \REG_1[13]$_DFF_P_  (.CLK(clknet_leaf_25_clock),
    .D(net300),
    .QN(_037_));
 DFFHQNx1_ASAP7_75t_R \REG_1[14]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(net301),
    .QN(_038_));
 DFFHQNx1_ASAP7_75t_R \REG_1[15]$_DFF_P_  (.CLK(clknet_leaf_24_clock),
    .D(net302),
    .QN(_039_));
 DFFHQNx1_ASAP7_75t_R \REG_1[16]$_DFF_P_  (.CLK(clknet_leaf_24_clock),
    .D(net303),
    .QN(_040_));
 DFFHQNx1_ASAP7_75t_R \REG_1[17]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(net304),
    .QN(_041_));
 DFFHQNx1_ASAP7_75t_R \REG_1[18]$_DFF_P_  (.CLK(clknet_leaf_23_clock),
    .D(net305),
    .QN(_042_));
 DFFHQNx1_ASAP7_75t_R \REG_1[19]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(net306),
    .QN(_043_));
 DFFHQNx1_ASAP7_75t_R \REG_1[1]$_DFF_P_  (.CLK(clknet_leaf_20_clock),
    .D(net307),
    .QN(_044_));
 DFFHQNx1_ASAP7_75t_R \REG_1[20]$_DFF_P_  (.CLK(clknet_leaf_23_clock),
    .D(net308),
    .QN(_045_));
 DFFHQNx1_ASAP7_75t_R \REG_1[21]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(net309),
    .QN(_046_));
 DFFHQNx1_ASAP7_75t_R \REG_1[22]$_DFF_P_  (.CLK(clknet_leaf_25_clock),
    .D(net310),
    .QN(_047_));
 DFFHQNx1_ASAP7_75t_R \REG_1[23]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(net311),
    .QN(_048_));
 DFFHQNx1_ASAP7_75t_R \REG_1[24]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(net312),
    .QN(_049_));
 DFFHQNx1_ASAP7_75t_R \REG_1[25]$_DFF_P_  (.CLK(clknet_leaf_23_clock),
    .D(net313),
    .QN(_050_));
 DFFHQNx1_ASAP7_75t_R \REG_1[26]$_DFF_P_  (.CLK(clknet_leaf_24_clock),
    .D(net314),
    .QN(_051_));
 DFFHQNx1_ASAP7_75t_R \REG_1[27]$_DFF_P_  (.CLK(clknet_leaf_23_clock),
    .D(net315),
    .QN(_052_));
 DFFHQNx1_ASAP7_75t_R \REG_1[28]$_DFF_P_  (.CLK(clknet_leaf_24_clock),
    .D(net316),
    .QN(_053_));
 DFFHQNx1_ASAP7_75t_R \REG_1[29]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(net317),
    .QN(_054_));
 DFFHQNx1_ASAP7_75t_R \REG_1[2]$_DFF_P_  (.CLK(clknet_leaf_20_clock),
    .D(net318),
    .QN(_055_));
 DFFHQNx1_ASAP7_75t_R \REG_1[30]$_DFF_P_  (.CLK(clknet_leaf_24_clock),
    .D(net319),
    .QN(_056_));
 DFFHQNx1_ASAP7_75t_R \REG_1[31]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(net320),
    .QN(_057_));
 DFFHQNx1_ASAP7_75t_R \REG_1[3]$_DFF_P_  (.CLK(clknet_leaf_20_clock),
    .D(net321),
    .QN(_058_));
 DFFHQNx1_ASAP7_75t_R \REG_1[4]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(net322),
    .QN(_059_));
 DFFHQNx1_ASAP7_75t_R \REG_1[5]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(net323),
    .QN(_060_));
 DFFHQNx1_ASAP7_75t_R \REG_1[6]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(net324),
    .QN(_061_));
 DFFHQNx1_ASAP7_75t_R \REG_1[7]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(net325),
    .QN(_062_));
 DFFHQNx1_ASAP7_75t_R \REG_1[8]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(net326),
    .QN(_063_));
 DFFHQNx1_ASAP7_75t_R \REG_1[9]$_DFF_P_  (.CLK(clknet_leaf_24_clock),
    .D(net327),
    .QN(_064_));
 DFFHQNx1_ASAP7_75t_R \REG_2[0]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(net328),
    .QN(_065_));
 DFFHQNx1_ASAP7_75t_R \REG_2[10]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(net329),
    .QN(_066_));
 DFFHQNx1_ASAP7_75t_R \REG_2[11]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(net330),
    .QN(_067_));
 DFFHQNx1_ASAP7_75t_R \REG_2[12]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(net331),
    .QN(_068_));
 DFFHQNx1_ASAP7_75t_R \REG_2[13]$_DFF_P_  (.CLK(clknet_leaf_3_clock),
    .D(net332),
    .QN(_069_));
 DFFHQNx1_ASAP7_75t_R \REG_2[14]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(net333),
    .QN(_070_));
 DFFHQNx1_ASAP7_75t_R \REG_2[15]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(net334),
    .QN(_071_));
 DFFHQNx1_ASAP7_75t_R \REG_2[16]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(net335),
    .QN(_072_));
 DFFHQNx1_ASAP7_75t_R \REG_2[17]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(net336),
    .QN(_073_));
 DFFHQNx1_ASAP7_75t_R \REG_2[18]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(net337),
    .QN(_074_));
 DFFHQNx1_ASAP7_75t_R \REG_2[19]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(net338),
    .QN(_075_));
 DFFHQNx1_ASAP7_75t_R \REG_2[1]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(net339),
    .QN(_076_));
 DFFHQNx1_ASAP7_75t_R \REG_2[20]$_DFF_P_  (.CLK(clknet_leaf_3_clock),
    .D(net340),
    .QN(_077_));
 DFFHQNx1_ASAP7_75t_R \REG_2[21]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(net341),
    .QN(_078_));
 DFFHQNx1_ASAP7_75t_R \REG_2[22]$_DFF_P_  (.CLK(clknet_leaf_33_clock),
    .D(net342),
    .QN(_079_));
 DFFHQNx1_ASAP7_75t_R \REG_2[23]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(net343),
    .QN(_080_));
 DFFHQNx1_ASAP7_75t_R \REG_2[24]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(net344),
    .QN(_081_));
 DFFHQNx1_ASAP7_75t_R \REG_2[25]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(net345),
    .QN(_082_));
 DFFHQNx1_ASAP7_75t_R \REG_2[26]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(net346),
    .QN(_083_));
 DFFHQNx1_ASAP7_75t_R \REG_2[27]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(net347),
    .QN(_084_));
 DFFHQNx1_ASAP7_75t_R \REG_2[28]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(net348),
    .QN(_085_));
 DFFHQNx1_ASAP7_75t_R \REG_2[29]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(net349),
    .QN(_086_));
 DFFHQNx1_ASAP7_75t_R \REG_2[2]$_DFF_P_  (.CLK(clknet_leaf_5_clock),
    .D(net350),
    .QN(_087_));
 DFFHQNx1_ASAP7_75t_R \REG_2[30]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(net351),
    .QN(_088_));
 DFFHQNx1_ASAP7_75t_R \REG_2[31]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(net352),
    .QN(_089_));
 DFFHQNx1_ASAP7_75t_R \REG_2[3]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(net353),
    .QN(_090_));
 DFFHQNx1_ASAP7_75t_R \REG_2[4]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(net354),
    .QN(_091_));
 DFFHQNx1_ASAP7_75t_R \REG_2[5]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(net355),
    .QN(_092_));
 DFFHQNx1_ASAP7_75t_R \REG_2[6]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(net356),
    .QN(_093_));
 DFFHQNx1_ASAP7_75t_R \REG_2[7]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(net357),
    .QN(_094_));
 DFFHQNx1_ASAP7_75t_R \REG_2[8]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(net358),
    .QN(_095_));
 DFFHQNx1_ASAP7_75t_R \REG_2[9]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(net359),
    .QN(_096_));
 DFFHQNx1_ASAP7_75t_R \REG_4[0]$_DFF_P_  (.CLK(clknet_leaf_28_clock),
    .D(net360),
    .QN(_097_));
 DFFHQNx1_ASAP7_75t_R \REG_4[10]$_DFF_P_  (.CLK(clknet_leaf_25_clock),
    .D(net361),
    .QN(_098_));
 DFFHQNx1_ASAP7_75t_R \REG_4[11]$_DFF_P_  (.CLK(clknet_leaf_25_clock),
    .D(net362),
    .QN(_099_));
 DFFHQNx1_ASAP7_75t_R \REG_4[12]$_DFF_P_  (.CLK(clknet_leaf_25_clock),
    .D(net363),
    .QN(_100_));
 DFFHQNx1_ASAP7_75t_R \REG_4[13]$_DFF_P_  (.CLK(clknet_leaf_31_clock),
    .D(net364),
    .QN(_101_));
 DFFHQNx1_ASAP7_75t_R \REG_4[14]$_DFF_P_  (.CLK(clknet_leaf_26_clock),
    .D(net365),
    .QN(_102_));
 DFFHQNx1_ASAP7_75t_R \REG_4[15]$_DFF_P_  (.CLK(clknet_leaf_25_clock),
    .D(net366),
    .QN(_103_));
 DFFHQNx1_ASAP7_75t_R \REG_4[16]$_DFF_P_  (.CLK(clknet_leaf_26_clock),
    .D(net367),
    .QN(_104_));
 DFFHQNx1_ASAP7_75t_R \REG_4[17]$_DFF_P_  (.CLK(clknet_leaf_31_clock),
    .D(net368),
    .QN(_105_));
 DFFHQNx1_ASAP7_75t_R \REG_4[18]$_DFF_P_  (.CLK(clknet_leaf_25_clock),
    .D(net369),
    .QN(_106_));
 DFFHQNx1_ASAP7_75t_R \REG_4[19]$_DFF_P_  (.CLK(clknet_leaf_31_clock),
    .D(net370),
    .QN(_107_));
 DFFHQNx1_ASAP7_75t_R \REG_4[1]$_DFF_P_  (.CLK(clknet_leaf_32_clock),
    .D(net371),
    .QN(_108_));
 DFFHQNx1_ASAP7_75t_R \REG_4[20]$_DFF_P_  (.CLK(clknet_leaf_27_clock),
    .D(net372),
    .QN(_109_));
 DFFHQNx1_ASAP7_75t_R \REG_4[21]$_DFF_P_  (.CLK(clknet_leaf_33_clock),
    .D(net373),
    .QN(_110_));
 DFFHQNx1_ASAP7_75t_R \REG_4[22]$_DFF_P_  (.CLK(clknet_leaf_27_clock),
    .D(net374),
    .QN(_111_));
 DFFHQNx1_ASAP7_75t_R \REG_4[23]$_DFF_P_  (.CLK(clknet_leaf_31_clock),
    .D(net375),
    .QN(_112_));
 DFFHQNx1_ASAP7_75t_R \REG_4[24]$_DFF_P_  (.CLK(clknet_leaf_26_clock),
    .D(net376),
    .QN(_113_));
 DFFHQNx1_ASAP7_75t_R \REG_4[25]$_DFF_P_  (.CLK(clknet_leaf_31_clock),
    .D(net377),
    .QN(_114_));
 DFFHQNx1_ASAP7_75t_R \REG_4[26]$_DFF_P_  (.CLK(clknet_leaf_26_clock),
    .D(net378),
    .QN(_115_));
 DFFHQNx1_ASAP7_75t_R \REG_4[27]$_DFF_P_  (.CLK(clknet_leaf_33_clock),
    .D(net379),
    .QN(_116_));
 DFFHQNx1_ASAP7_75t_R \REG_4[28]$_DFF_P_  (.CLK(clknet_leaf_26_clock),
    .D(net380),
    .QN(_117_));
 DFFHQNx1_ASAP7_75t_R \REG_4[29]$_DFF_P_  (.CLK(clknet_leaf_27_clock),
    .D(net381),
    .QN(_118_));
 DFFHQNx1_ASAP7_75t_R \REG_4[2]$_DFF_P_  (.CLK(clknet_leaf_32_clock),
    .D(net382),
    .QN(_119_));
 DFFHQNx1_ASAP7_75t_R \REG_4[30]$_DFF_P_  (.CLK(clknet_leaf_32_clock),
    .D(net383),
    .QN(_120_));
 DFFHQNx1_ASAP7_75t_R \REG_4[31]$_DFF_P_  (.CLK(clknet_leaf_32_clock),
    .D(net384),
    .QN(_121_));
 DFFHQNx1_ASAP7_75t_R \REG_4[3]$_DFF_P_  (.CLK(clknet_leaf_22_clock),
    .D(net385),
    .QN(_122_));
 DFFHQNx1_ASAP7_75t_R \REG_4[4]$_DFF_P_  (.CLK(clknet_leaf_27_clock),
    .D(net386),
    .QN(_123_));
 DFFHQNx1_ASAP7_75t_R \REG_4[5]$_DFF_P_  (.CLK(clknet_leaf_33_clock),
    .D(net387),
    .QN(_124_));
 DFFHQNx1_ASAP7_75t_R \REG_4[6]$_DFF_P_  (.CLK(clknet_leaf_25_clock),
    .D(net388),
    .QN(_125_));
 DFFHQNx1_ASAP7_75t_R \REG_4[7]$_DFF_P_  (.CLK(clknet_leaf_26_clock),
    .D(net389),
    .QN(_126_));
 DFFHQNx1_ASAP7_75t_R \REG_4[8]$_DFF_P_  (.CLK(clknet_leaf_31_clock),
    .D(net390),
    .QN(_127_));
 DFFHQNx1_ASAP7_75t_R \REG_4[9]$_DFF_P_  (.CLK(clknet_leaf_27_clock),
    .D(net391),
    .QN(_128_));
 DFFHQNx1_ASAP7_75t_R \REG_8$_DFF_P_  (.CLK(clknet_leaf_9_clock),
    .D(net392),
    .QN(_129_));
 INVx3_ASAP7_75t_R _258_ (.A(_000_),
    .Y(net524));
 INVx3_ASAP7_75t_R _259_ (.A(_001_),
    .Y(\REG[0] ));
 INVx3_ASAP7_75t_R _260_ (.A(_002_),
    .Y(\REG[10] ));
 INVx3_ASAP7_75t_R _261_ (.A(_003_),
    .Y(\REG[11] ));
 INVx3_ASAP7_75t_R _262_ (.A(_004_),
    .Y(\REG[12] ));
 INVx3_ASAP7_75t_R _263_ (.A(_005_),
    .Y(\REG[13] ));
 INVx3_ASAP7_75t_R _264_ (.A(_006_),
    .Y(\REG[14] ));
 INVx3_ASAP7_75t_R _265_ (.A(_007_),
    .Y(\REG[15] ));
 INVx3_ASAP7_75t_R _266_ (.A(_008_),
    .Y(\REG[16] ));
 INVx3_ASAP7_75t_R _267_ (.A(_009_),
    .Y(\REG[17] ));
 INVx3_ASAP7_75t_R _268_ (.A(_010_),
    .Y(\REG[18] ));
 INVx3_ASAP7_75t_R _269_ (.A(_011_),
    .Y(\REG[19] ));
 INVx3_ASAP7_75t_R _270_ (.A(_012_),
    .Y(\REG[1] ));
 INVx3_ASAP7_75t_R _271_ (.A(_013_),
    .Y(\REG[20] ));
 INVx3_ASAP7_75t_R _272_ (.A(_014_),
    .Y(\REG[21] ));
 INVx3_ASAP7_75t_R _273_ (.A(_015_),
    .Y(\REG[22] ));
 INVx3_ASAP7_75t_R _274_ (.A(_016_),
    .Y(\REG[23] ));
 INVx3_ASAP7_75t_R _275_ (.A(_017_),
    .Y(\REG[24] ));
 INVx3_ASAP7_75t_R _276_ (.A(_018_),
    .Y(\REG[25] ));
 INVx3_ASAP7_75t_R _277_ (.A(_019_),
    .Y(\REG[26] ));
 INVx3_ASAP7_75t_R _278_ (.A(_020_),
    .Y(\REG[27] ));
 INVx3_ASAP7_75t_R _279_ (.A(_021_),
    .Y(\REG[28] ));
 INVx3_ASAP7_75t_R _280_ (.A(_022_),
    .Y(\REG[29] ));
 INVx3_ASAP7_75t_R _281_ (.A(_023_),
    .Y(\REG[2] ));
 INVx3_ASAP7_75t_R _282_ (.A(_024_),
    .Y(\REG[30] ));
 INVx3_ASAP7_75t_R _283_ (.A(_025_),
    .Y(\REG[31] ));
 INVx3_ASAP7_75t_R _284_ (.A(_026_),
    .Y(\REG[3] ));
 INVx3_ASAP7_75t_R _285_ (.A(_027_),
    .Y(\REG[4] ));
 INVx3_ASAP7_75t_R _286_ (.A(_028_),
    .Y(\REG[5] ));
 INVx3_ASAP7_75t_R _287_ (.A(_029_),
    .Y(\REG[6] ));
 INVx3_ASAP7_75t_R _288_ (.A(_030_),
    .Y(\REG[7] ));
 INVx3_ASAP7_75t_R _289_ (.A(_031_),
    .Y(\REG[8] ));
 INVx3_ASAP7_75t_R _290_ (.A(_032_),
    .Y(\REG[9] ));
 INVx3_ASAP7_75t_R _291_ (.A(_033_),
    .Y(\REG_1[0] ));
 INVx3_ASAP7_75t_R _292_ (.A(_034_),
    .Y(\REG_1[10] ));
 INVx3_ASAP7_75t_R _293_ (.A(_035_),
    .Y(\REG_1[11] ));
 INVx3_ASAP7_75t_R _294_ (.A(_036_),
    .Y(\REG_1[12] ));
 INVx3_ASAP7_75t_R _295_ (.A(_037_),
    .Y(\REG_1[13] ));
 INVx3_ASAP7_75t_R _296_ (.A(_038_),
    .Y(\REG_1[14] ));
 INVx3_ASAP7_75t_R _297_ (.A(_039_),
    .Y(\REG_1[15] ));
 INVx3_ASAP7_75t_R _298_ (.A(_040_),
    .Y(\REG_1[16] ));
 INVx3_ASAP7_75t_R _299_ (.A(_041_),
    .Y(\REG_1[17] ));
 INVx3_ASAP7_75t_R _300_ (.A(_042_),
    .Y(\REG_1[18] ));
 INVx3_ASAP7_75t_R _301_ (.A(_043_),
    .Y(\REG_1[19] ));
 INVx3_ASAP7_75t_R _302_ (.A(_044_),
    .Y(\REG_1[1] ));
 INVx3_ASAP7_75t_R _303_ (.A(_045_),
    .Y(\REG_1[20] ));
 INVx3_ASAP7_75t_R _304_ (.A(_046_),
    .Y(\REG_1[21] ));
 INVx3_ASAP7_75t_R _305_ (.A(_047_),
    .Y(\REG_1[22] ));
 INVx3_ASAP7_75t_R _306_ (.A(_048_),
    .Y(\REG_1[23] ));
 INVx3_ASAP7_75t_R _307_ (.A(_049_),
    .Y(\REG_1[24] ));
 INVx3_ASAP7_75t_R _308_ (.A(_050_),
    .Y(\REG_1[25] ));
 INVx3_ASAP7_75t_R _309_ (.A(_051_),
    .Y(\REG_1[26] ));
 INVx3_ASAP7_75t_R _310_ (.A(_052_),
    .Y(\REG_1[27] ));
 INVx3_ASAP7_75t_R _311_ (.A(_053_),
    .Y(\REG_1[28] ));
 INVx3_ASAP7_75t_R _312_ (.A(_054_),
    .Y(\REG_1[29] ));
 INVx3_ASAP7_75t_R _313_ (.A(_055_),
    .Y(\REG_1[2] ));
 INVx3_ASAP7_75t_R _314_ (.A(_056_),
    .Y(\REG_1[30] ));
 INVx3_ASAP7_75t_R _315_ (.A(_057_),
    .Y(\REG_1[31] ));
 INVx3_ASAP7_75t_R _316_ (.A(_058_),
    .Y(\REG_1[3] ));
 INVx3_ASAP7_75t_R _317_ (.A(_059_),
    .Y(\REG_1[4] ));
 INVx3_ASAP7_75t_R _318_ (.A(_060_),
    .Y(\REG_1[5] ));
 INVx3_ASAP7_75t_R _319_ (.A(_061_),
    .Y(\REG_1[6] ));
 INVx3_ASAP7_75t_R _320_ (.A(_062_),
    .Y(\REG_1[7] ));
 INVx3_ASAP7_75t_R _321_ (.A(_063_),
    .Y(\REG_1[8] ));
 INVx3_ASAP7_75t_R _322_ (.A(_064_),
    .Y(\REG_1[9] ));
 INVx3_ASAP7_75t_R _323_ (.A(_065_),
    .Y(\REG_2[0] ));
 INVx3_ASAP7_75t_R _324_ (.A(_066_),
    .Y(\REG_2[10] ));
 INVx3_ASAP7_75t_R _325_ (.A(_067_),
    .Y(\REG_2[11] ));
 INVx3_ASAP7_75t_R _326_ (.A(_068_),
    .Y(\REG_2[12] ));
 INVx3_ASAP7_75t_R _327_ (.A(_069_),
    .Y(\REG_2[13] ));
 INVx3_ASAP7_75t_R _328_ (.A(_070_),
    .Y(\REG_2[14] ));
 INVx3_ASAP7_75t_R _329_ (.A(_071_),
    .Y(\REG_2[15] ));
 INVx3_ASAP7_75t_R _330_ (.A(_072_),
    .Y(\REG_2[16] ));
 INVx3_ASAP7_75t_R _331_ (.A(_073_),
    .Y(\REG_2[17] ));
 INVx3_ASAP7_75t_R _332_ (.A(_074_),
    .Y(\REG_2[18] ));
 INVx3_ASAP7_75t_R _333_ (.A(_075_),
    .Y(\REG_2[19] ));
 INVx3_ASAP7_75t_R _334_ (.A(_076_),
    .Y(\REG_2[1] ));
 INVx3_ASAP7_75t_R _335_ (.A(_077_),
    .Y(\REG_2[20] ));
 INVx3_ASAP7_75t_R _336_ (.A(_078_),
    .Y(\REG_2[21] ));
 INVx3_ASAP7_75t_R _337_ (.A(_079_),
    .Y(\REG_2[22] ));
 INVx3_ASAP7_75t_R _338_ (.A(_080_),
    .Y(\REG_2[23] ));
 INVx3_ASAP7_75t_R _339_ (.A(_081_),
    .Y(\REG_2[24] ));
 INVx3_ASAP7_75t_R _340_ (.A(_082_),
    .Y(\REG_2[25] ));
 INVx3_ASAP7_75t_R _341_ (.A(_083_),
    .Y(\REG_2[26] ));
 INVx3_ASAP7_75t_R _342_ (.A(_084_),
    .Y(\REG_2[27] ));
 INVx3_ASAP7_75t_R _343_ (.A(_085_),
    .Y(\REG_2[28] ));
 INVx3_ASAP7_75t_R _344_ (.A(_086_),
    .Y(\REG_2[29] ));
 INVx3_ASAP7_75t_R _345_ (.A(_087_),
    .Y(\REG_2[2] ));
 INVx3_ASAP7_75t_R _346_ (.A(_088_),
    .Y(\REG_2[30] ));
 INVx3_ASAP7_75t_R _347_ (.A(_089_),
    .Y(\REG_2[31] ));
 INVx3_ASAP7_75t_R _348_ (.A(_090_),
    .Y(\REG_2[3] ));
 INVx3_ASAP7_75t_R _349_ (.A(_091_),
    .Y(\REG_2[4] ));
 INVx3_ASAP7_75t_R _350_ (.A(_092_),
    .Y(\REG_2[5] ));
 INVx3_ASAP7_75t_R _351_ (.A(_093_),
    .Y(\REG_2[6] ));
 INVx3_ASAP7_75t_R _352_ (.A(_094_),
    .Y(\REG_2[7] ));
 INVx3_ASAP7_75t_R _353_ (.A(_095_),
    .Y(\REG_2[8] ));
 INVx3_ASAP7_75t_R _354_ (.A(_096_),
    .Y(\REG_2[9] ));
 INVx3_ASAP7_75t_R _355_ (.A(_097_),
    .Y(\REG_4[0] ));
 INVx3_ASAP7_75t_R _356_ (.A(_098_),
    .Y(\REG_4[10] ));
 INVx3_ASAP7_75t_R _357_ (.A(_099_),
    .Y(\REG_4[11] ));
 INVx3_ASAP7_75t_R _358_ (.A(_100_),
    .Y(\REG_4[12] ));
 INVx3_ASAP7_75t_R _359_ (.A(_101_),
    .Y(\REG_4[13] ));
 INVx3_ASAP7_75t_R _360_ (.A(_102_),
    .Y(\REG_4[14] ));
 INVx3_ASAP7_75t_R _361_ (.A(_103_),
    .Y(\REG_4[15] ));
 INVx3_ASAP7_75t_R _362_ (.A(_104_),
    .Y(\REG_4[16] ));
 INVx3_ASAP7_75t_R _363_ (.A(_105_),
    .Y(\REG_4[17] ));
 INVx3_ASAP7_75t_R _364_ (.A(_106_),
    .Y(\REG_4[18] ));
 INVx3_ASAP7_75t_R _365_ (.A(_107_),
    .Y(\REG_4[19] ));
 INVx3_ASAP7_75t_R _366_ (.A(_108_),
    .Y(\REG_4[1] ));
 INVx3_ASAP7_75t_R _367_ (.A(_109_),
    .Y(\REG_4[20] ));
 INVx3_ASAP7_75t_R _368_ (.A(_110_),
    .Y(\REG_4[21] ));
 INVx3_ASAP7_75t_R _369_ (.A(_111_),
    .Y(\REG_4[22] ));
 INVx3_ASAP7_75t_R _370_ (.A(_112_),
    .Y(\REG_4[23] ));
 INVx3_ASAP7_75t_R _371_ (.A(_113_),
    .Y(\REG_4[24] ));
 INVx3_ASAP7_75t_R _372_ (.A(_114_),
    .Y(\REG_4[25] ));
 INVx3_ASAP7_75t_R _373_ (.A(_115_),
    .Y(\REG_4[26] ));
 INVx3_ASAP7_75t_R _374_ (.A(_116_),
    .Y(\REG_4[27] ));
 INVx3_ASAP7_75t_R _375_ (.A(_117_),
    .Y(\REG_4[28] ));
 INVx3_ASAP7_75t_R _376_ (.A(_118_),
    .Y(\REG_4[29] ));
 INVx3_ASAP7_75t_R _377_ (.A(_119_),
    .Y(\REG_4[2] ));
 INVx3_ASAP7_75t_R _378_ (.A(_120_),
    .Y(\REG_4[30] ));
 INVx3_ASAP7_75t_R _379_ (.A(_121_),
    .Y(\REG_4[31] ));
 INVx3_ASAP7_75t_R _380_ (.A(_122_),
    .Y(\REG_4[3] ));
 INVx3_ASAP7_75t_R _381_ (.A(_123_),
    .Y(\REG_4[4] ));
 INVx3_ASAP7_75t_R _382_ (.A(_124_),
    .Y(\REG_4[5] ));
 INVx3_ASAP7_75t_R _383_ (.A(_125_),
    .Y(\REG_4[6] ));
 INVx3_ASAP7_75t_R _384_ (.A(_126_),
    .Y(\REG_4[7] ));
 INVx3_ASAP7_75t_R _385_ (.A(_127_),
    .Y(\REG_4[8] ));
 INVx3_ASAP7_75t_R _386_ (.A(_128_),
    .Y(\REG_4[9] ));
 INVx3_ASAP7_75t_R _387_ (.A(_129_),
    .Y(net394));
 INVx3_ASAP7_75t_R _388_ (.A(_130_),
    .Y(net397));
 INVx3_ASAP7_75t_R _389_ (.A(_131_),
    .Y(net398));
 INVx3_ASAP7_75t_R _390_ (.A(_132_),
    .Y(net399));
 INVx3_ASAP7_75t_R _391_ (.A(_133_),
    .Y(net400));
 INVx3_ASAP7_75t_R _392_ (.A(_134_),
    .Y(net401));
 INVx3_ASAP7_75t_R _393_ (.A(_135_),
    .Y(net402));
 INVx3_ASAP7_75t_R _394_ (.A(_136_),
    .Y(net403));
 INVx3_ASAP7_75t_R _395_ (.A(_137_),
    .Y(net404));
 INVx3_ASAP7_75t_R _396_ (.A(_138_),
    .Y(net405));
 INVx3_ASAP7_75t_R _397_ (.A(_139_),
    .Y(net406));
 INVx3_ASAP7_75t_R _398_ (.A(_140_),
    .Y(net407));
 INVx3_ASAP7_75t_R _399_ (.A(_141_),
    .Y(net408));
 INVx3_ASAP7_75t_R _400_ (.A(_142_),
    .Y(net409));
 INVx3_ASAP7_75t_R _401_ (.A(_143_),
    .Y(net410));
 INVx3_ASAP7_75t_R _402_ (.A(_144_),
    .Y(net411));
 INVx3_ASAP7_75t_R _403_ (.A(_145_),
    .Y(net412));
 INVx3_ASAP7_75t_R _404_ (.A(_146_),
    .Y(net413));
 INVx3_ASAP7_75t_R _405_ (.A(_147_),
    .Y(net414));
 INVx3_ASAP7_75t_R _406_ (.A(_148_),
    .Y(net415));
 INVx3_ASAP7_75t_R _407_ (.A(_149_),
    .Y(net416));
 INVx3_ASAP7_75t_R _408_ (.A(_150_),
    .Y(net417));
 INVx3_ASAP7_75t_R _409_ (.A(_151_),
    .Y(net418));
 INVx3_ASAP7_75t_R _410_ (.A(_152_),
    .Y(net419));
 INVx3_ASAP7_75t_R _411_ (.A(_153_),
    .Y(net420));
 INVx3_ASAP7_75t_R _412_ (.A(_154_),
    .Y(net421));
 INVx3_ASAP7_75t_R _413_ (.A(_155_),
    .Y(net422));
 INVx3_ASAP7_75t_R _414_ (.A(_156_),
    .Y(net423));
 INVx3_ASAP7_75t_R _415_ (.A(_157_),
    .Y(net424));
 INVx3_ASAP7_75t_R _416_ (.A(_158_),
    .Y(net425));
 INVx3_ASAP7_75t_R _417_ (.A(_159_),
    .Y(net426));
 INVx3_ASAP7_75t_R _418_ (.A(_160_),
    .Y(net427));
 INVx3_ASAP7_75t_R _419_ (.A(_161_),
    .Y(net428));
 INVx3_ASAP7_75t_R _420_ (.A(_162_),
    .Y(net396));
 INVx3_ASAP7_75t_R _421_ (.A(_163_),
    .Y(net430));
 INVx3_ASAP7_75t_R _422_ (.A(_164_),
    .Y(net431));
 INVx3_ASAP7_75t_R _423_ (.A(_165_),
    .Y(net432));
 INVx3_ASAP7_75t_R _424_ (.A(_166_),
    .Y(net433));
 INVx3_ASAP7_75t_R _425_ (.A(_167_),
    .Y(net434));
 INVx3_ASAP7_75t_R _426_ (.A(_168_),
    .Y(net435));
 INVx3_ASAP7_75t_R _427_ (.A(_169_),
    .Y(net436));
 INVx3_ASAP7_75t_R _428_ (.A(_170_),
    .Y(net437));
 INVx3_ASAP7_75t_R _429_ (.A(_171_),
    .Y(net438));
 INVx3_ASAP7_75t_R _430_ (.A(_172_),
    .Y(net439));
 INVx3_ASAP7_75t_R _431_ (.A(_173_),
    .Y(net440));
 INVx3_ASAP7_75t_R _432_ (.A(_174_),
    .Y(net441));
 INVx3_ASAP7_75t_R _433_ (.A(_175_),
    .Y(net442));
 INVx3_ASAP7_75t_R _434_ (.A(_176_),
    .Y(net443));
 INVx3_ASAP7_75t_R _435_ (.A(_177_),
    .Y(net444));
 INVx3_ASAP7_75t_R _436_ (.A(_178_),
    .Y(net445));
 INVx3_ASAP7_75t_R _437_ (.A(_179_),
    .Y(net446));
 INVx3_ASAP7_75t_R _438_ (.A(_180_),
    .Y(net447));
 INVx3_ASAP7_75t_R _439_ (.A(_181_),
    .Y(net448));
 INVx3_ASAP7_75t_R _440_ (.A(_182_),
    .Y(net449));
 INVx3_ASAP7_75t_R _441_ (.A(_183_),
    .Y(net450));
 INVx3_ASAP7_75t_R _442_ (.A(_184_),
    .Y(net451));
 INVx3_ASAP7_75t_R _443_ (.A(_185_),
    .Y(net452));
 INVx3_ASAP7_75t_R _444_ (.A(_186_),
    .Y(net453));
 INVx3_ASAP7_75t_R _445_ (.A(_187_),
    .Y(net454));
 INVx3_ASAP7_75t_R _446_ (.A(_188_),
    .Y(net455));
 INVx3_ASAP7_75t_R _447_ (.A(_189_),
    .Y(net456));
 INVx3_ASAP7_75t_R _448_ (.A(_190_),
    .Y(net457));
 INVx3_ASAP7_75t_R _449_ (.A(_191_),
    .Y(net458));
 INVx3_ASAP7_75t_R _450_ (.A(_192_),
    .Y(net459));
 INVx3_ASAP7_75t_R _451_ (.A(_193_),
    .Y(net460));
 INVx3_ASAP7_75t_R _452_ (.A(_194_),
    .Y(net461));
 INVx3_ASAP7_75t_R _453_ (.A(_195_),
    .Y(net462));
 INVx3_ASAP7_75t_R _454_ (.A(_196_),
    .Y(net463));
 INVx3_ASAP7_75t_R _455_ (.A(_197_),
    .Y(net464));
 INVx3_ASAP7_75t_R _456_ (.A(_198_),
    .Y(net465));
 INVx3_ASAP7_75t_R _457_ (.A(_199_),
    .Y(net466));
 INVx3_ASAP7_75t_R _458_ (.A(_200_),
    .Y(net467));
 INVx3_ASAP7_75t_R _459_ (.A(_201_),
    .Y(net468));
 INVx3_ASAP7_75t_R _460_ (.A(_202_),
    .Y(net469));
 INVx3_ASAP7_75t_R _461_ (.A(_203_),
    .Y(net470));
 INVx3_ASAP7_75t_R _462_ (.A(_204_),
    .Y(net471));
 INVx3_ASAP7_75t_R _463_ (.A(_205_),
    .Y(net472));
 INVx3_ASAP7_75t_R _464_ (.A(_206_),
    .Y(net473));
 INVx3_ASAP7_75t_R _465_ (.A(_207_),
    .Y(net474));
 INVx3_ASAP7_75t_R _466_ (.A(_208_),
    .Y(net475));
 INVx3_ASAP7_75t_R _467_ (.A(_209_),
    .Y(net476));
 INVx3_ASAP7_75t_R _468_ (.A(_210_),
    .Y(net477));
 INVx3_ASAP7_75t_R _469_ (.A(_211_),
    .Y(net478));
 INVx3_ASAP7_75t_R _470_ (.A(_212_),
    .Y(net479));
 INVx3_ASAP7_75t_R _471_ (.A(_213_),
    .Y(net480));
 INVx3_ASAP7_75t_R _472_ (.A(_214_),
    .Y(net481));
 INVx3_ASAP7_75t_R _473_ (.A(_215_),
    .Y(net482));
 INVx3_ASAP7_75t_R _474_ (.A(_216_),
    .Y(net483));
 INVx3_ASAP7_75t_R _475_ (.A(_217_),
    .Y(net484));
 INVx3_ASAP7_75t_R _476_ (.A(_218_),
    .Y(net485));
 INVx3_ASAP7_75t_R _477_ (.A(_219_),
    .Y(net486));
 INVx3_ASAP7_75t_R _478_ (.A(_220_),
    .Y(net487));
 INVx3_ASAP7_75t_R _479_ (.A(_221_),
    .Y(net488));
 INVx3_ASAP7_75t_R _480_ (.A(_222_),
    .Y(net489));
 INVx3_ASAP7_75t_R _481_ (.A(_223_),
    .Y(net490));
 INVx3_ASAP7_75t_R _482_ (.A(_224_),
    .Y(net491));
 INVx3_ASAP7_75t_R _483_ (.A(_225_),
    .Y(net492));
 INVx3_ASAP7_75t_R _484_ (.A(_226_),
    .Y(net493));
 INVx3_ASAP7_75t_R _485_ (.A(_227_),
    .Y(net494));
 INVx3_ASAP7_75t_R _486_ (.A(_228_),
    .Y(net495));
 INVx3_ASAP7_75t_R _487_ (.A(_229_),
    .Y(net496));
 INVx3_ASAP7_75t_R _488_ (.A(_230_),
    .Y(net497));
 INVx3_ASAP7_75t_R _489_ (.A(_231_),
    .Y(net498));
 INVx3_ASAP7_75t_R _490_ (.A(_232_),
    .Y(net499));
 INVx3_ASAP7_75t_R _491_ (.A(_233_),
    .Y(net500));
 INVx3_ASAP7_75t_R _492_ (.A(_234_),
    .Y(net501));
 INVx3_ASAP7_75t_R _493_ (.A(_235_),
    .Y(net502));
 INVx3_ASAP7_75t_R _494_ (.A(_236_),
    .Y(net503));
 INVx3_ASAP7_75t_R _495_ (.A(_237_),
    .Y(net504));
 INVx3_ASAP7_75t_R _496_ (.A(_238_),
    .Y(net505));
 INVx3_ASAP7_75t_R _497_ (.A(_239_),
    .Y(net506));
 INVx3_ASAP7_75t_R _498_ (.A(_240_),
    .Y(net507));
 INVx3_ASAP7_75t_R _499_ (.A(_241_),
    .Y(net508));
 INVx3_ASAP7_75t_R _500_ (.A(_242_),
    .Y(net509));
 INVx3_ASAP7_75t_R _501_ (.A(_243_),
    .Y(net510));
 INVx3_ASAP7_75t_R _502_ (.A(_244_),
    .Y(net511));
 INVx3_ASAP7_75t_R _503_ (.A(_245_),
    .Y(net512));
 INVx3_ASAP7_75t_R _504_ (.A(_246_),
    .Y(net513));
 INVx3_ASAP7_75t_R _505_ (.A(_247_),
    .Y(net514));
 INVx3_ASAP7_75t_R _506_ (.A(_248_),
    .Y(net515));
 INVx3_ASAP7_75t_R _507_ (.A(_249_),
    .Y(net516));
 INVx3_ASAP7_75t_R _508_ (.A(_250_),
    .Y(net517));
 INVx3_ASAP7_75t_R _509_ (.A(_251_),
    .Y(net518));
 INVx3_ASAP7_75t_R _510_ (.A(_252_),
    .Y(net519));
 INVx3_ASAP7_75t_R _511_ (.A(_253_),
    .Y(net520));
 INVx3_ASAP7_75t_R _512_ (.A(_254_),
    .Y(net521));
 INVx3_ASAP7_75t_R _513_ (.A(_255_),
    .Y(net522));
 INVx3_ASAP7_75t_R _514_ (.A(_256_),
    .Y(net523));
 BUFx2_ASAP7_75t_R _516_ (.A(io_lsbIns_1),
    .Y(net393));
 BUFx2_ASAP7_75t_R _517_ (.A(io_lsbIns_3),
    .Y(net395));
 DFFHQNx1_ASAP7_75t_R \io_outs_down_REG[0]$_DFF_P_  (.CLK(clknet_leaf_28_clock),
    .D(\_io_outs_down_mult_io_o[0] ),
    .QN(_130_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down_REG[10]$_DFF_P_  (.CLK(clknet_leaf_27_clock),
    .D(\_io_outs_down_mult_io_o[10] ),
    .QN(_131_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down_REG[11]$_DFF_P_  (.CLK(clknet_leaf_26_clock),
    .D(\_io_outs_down_mult_io_o[11] ),
    .QN(_132_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down_REG[12]$_DFF_P_  (.CLK(clknet_leaf_32_clock),
    .D(\_io_outs_down_mult_io_o[12] ),
    .QN(_133_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down_REG[13]$_DFF_P_  (.CLK(clknet_leaf_33_clock),
    .D(\_io_outs_down_mult_io_o[13] ),
    .QN(_134_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down_REG[14]$_DFF_P_  (.CLK(clknet_leaf_27_clock),
    .D(\_io_outs_down_mult_io_o[14] ),
    .QN(_135_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down_REG[15]$_DFF_P_  (.CLK(clknet_leaf_27_clock),
    .D(\_io_outs_down_mult_io_o[15] ),
    .QN(_136_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down_REG[16]$_DFF_P_  (.CLK(clknet_leaf_26_clock),
    .D(\_io_outs_down_mult_io_o[16] ),
    .QN(_137_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down_REG[17]$_DFF_P_  (.CLK(clknet_leaf_27_clock),
    .D(\_io_outs_down_mult_io_o[17] ),
    .QN(_138_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down_REG[18]$_DFF_P_  (.CLK(clknet_leaf_32_clock),
    .D(\_io_outs_down_mult_io_o[18] ),
    .QN(_139_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down_REG[19]$_DFF_P_  (.CLK(clknet_leaf_26_clock),
    .D(\_io_outs_down_mult_io_o[19] ),
    .QN(_140_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down_REG[1]$_DFF_P_  (.CLK(clknet_leaf_32_clock),
    .D(\_io_outs_down_mult_io_o[1] ),
    .QN(_141_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down_REG[20]$_DFF_P_  (.CLK(clknet_leaf_31_clock),
    .D(\_io_outs_down_mult_io_o[20] ),
    .QN(_142_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down_REG[21]$_DFF_P_  (.CLK(clknet_leaf_32_clock),
    .D(\_io_outs_down_mult_io_o[21] ),
    .QN(_143_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down_REG[22]$_DFF_P_  (.CLK(clknet_leaf_32_clock),
    .D(\_io_outs_down_mult_io_o[22] ),
    .QN(_144_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down_REG[23]$_DFF_P_  (.CLK(clknet_leaf_26_clock),
    .D(\_io_outs_down_mult_io_o[23] ),
    .QN(_145_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down_REG[24]$_DFF_P_  (.CLK(clknet_leaf_28_clock),
    .D(\_io_outs_down_mult_io_o[24] ),
    .QN(_146_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down_REG[25]$_DFF_P_  (.CLK(clknet_leaf_25_clock),
    .D(\_io_outs_down_mult_io_o[25] ),
    .QN(_147_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down_REG[26]$_DFF_P_  (.CLK(clknet_leaf_27_clock),
    .D(\_io_outs_down_mult_io_o[26] ),
    .QN(_148_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down_REG[27]$_DFF_P_  (.CLK(clknet_leaf_32_clock),
    .D(\_io_outs_down_mult_io_o[27] ),
    .QN(_149_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down_REG[28]$_DFF_P_  (.CLK(clknet_leaf_26_clock),
    .D(\_io_outs_down_mult_io_o[28] ),
    .QN(_150_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down_REG[29]$_DFF_P_  (.CLK(clknet_leaf_31_clock),
    .D(\_io_outs_down_mult_io_o[29] ),
    .QN(_151_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down_REG[2]$_DFF_P_  (.CLK(clknet_leaf_30_clock),
    .D(\_io_outs_down_mult_io_o[2] ),
    .QN(_152_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down_REG[30]$_DFF_P_  (.CLK(clknet_leaf_33_clock),
    .D(\_io_outs_down_mult_io_o[30] ),
    .QN(_153_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down_REG[31]$_DFF_P_  (.CLK(clknet_leaf_28_clock),
    .D(\_io_outs_down_mult_io_o[31] ),
    .QN(_154_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down_REG[3]$_DFF_P_  (.CLK(clknet_leaf_31_clock),
    .D(\_io_outs_down_mult_io_o[3] ),
    .QN(_155_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down_REG[4]$_DFF_P_  (.CLK(clknet_leaf_27_clock),
    .D(\_io_outs_down_mult_io_o[4] ),
    .QN(_156_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down_REG[5]$_DFF_P_  (.CLK(clknet_leaf_31_clock),
    .D(\_io_outs_down_mult_io_o[5] ),
    .QN(_157_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down_REG[6]$_DFF_P_  (.CLK(clknet_leaf_26_clock),
    .D(\_io_outs_down_mult_io_o[6] ),
    .QN(_158_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down_REG[7]$_DFF_P_  (.CLK(clknet_leaf_33_clock),
    .D(\_io_outs_down_mult_io_o[7] ),
    .QN(_159_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down_REG[8]$_DFF_P_  (.CLK(clknet_leaf_28_clock),
    .D(\_io_outs_down_mult_io_o[8] ),
    .QN(_160_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down_REG[9]$_DFF_P_  (.CLK(clknet_leaf_25_clock),
    .D(\_io_outs_down_mult_io_o[9] ),
    .QN(_161_));
 DFFHQNx1_ASAP7_75t_R \io_outs_left_REG[0]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(\_io_outs_left_mult_io_o[0] ),
    .QN(_162_));
 DFFHQNx1_ASAP7_75t_R \io_outs_left_REG[10]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(\_io_outs_left_mult_io_o[10] ),
    .QN(_163_));
 DFFHQNx1_ASAP7_75t_R \io_outs_left_REG[11]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(\_io_outs_left_mult_io_o[11] ),
    .QN(_164_));
 DFFHQNx1_ASAP7_75t_R \io_outs_left_REG[12]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(\_io_outs_left_mult_io_o[12] ),
    .QN(_165_));
 DFFHQNx1_ASAP7_75t_R \io_outs_left_REG[13]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(\_io_outs_left_mult_io_o[13] ),
    .QN(_166_));
 DFFHQNx1_ASAP7_75t_R \io_outs_left_REG[14]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(\_io_outs_left_mult_io_o[14] ),
    .QN(_167_));
 DFFHQNx1_ASAP7_75t_R \io_outs_left_REG[15]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(\_io_outs_left_mult_io_o[15] ),
    .QN(_168_));
 DFFHQNx1_ASAP7_75t_R \io_outs_left_REG[16]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(\_io_outs_left_mult_io_o[16] ),
    .QN(_169_));
 DFFHQNx1_ASAP7_75t_R \io_outs_left_REG[17]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(\_io_outs_left_mult_io_o[17] ),
    .QN(_170_));
 DFFHQNx1_ASAP7_75t_R \io_outs_left_REG[18]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(\_io_outs_left_mult_io_o[18] ),
    .QN(_171_));
 DFFHQNx1_ASAP7_75t_R \io_outs_left_REG[19]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(\_io_outs_left_mult_io_o[19] ),
    .QN(_172_));
 DFFHQNx1_ASAP7_75t_R \io_outs_left_REG[1]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(\_io_outs_left_mult_io_o[1] ),
    .QN(_173_));
 DFFHQNx1_ASAP7_75t_R \io_outs_left_REG[20]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(\_io_outs_left_mult_io_o[20] ),
    .QN(_174_));
 DFFHQNx1_ASAP7_75t_R \io_outs_left_REG[21]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(\_io_outs_left_mult_io_o[21] ),
    .QN(_175_));
 DFFHQNx1_ASAP7_75t_R \io_outs_left_REG[22]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(\_io_outs_left_mult_io_o[22] ),
    .QN(_176_));
 DFFHQNx1_ASAP7_75t_R \io_outs_left_REG[23]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(\_io_outs_left_mult_io_o[23] ),
    .QN(_177_));
 DFFHQNx1_ASAP7_75t_R \io_outs_left_REG[24]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(\_io_outs_left_mult_io_o[24] ),
    .QN(_178_));
 DFFHQNx1_ASAP7_75t_R \io_outs_left_REG[25]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(\_io_outs_left_mult_io_o[25] ),
    .QN(_179_));
 DFFHQNx1_ASAP7_75t_R \io_outs_left_REG[26]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(\_io_outs_left_mult_io_o[26] ),
    .QN(_180_));
 DFFHQNx1_ASAP7_75t_R \io_outs_left_REG[27]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(\_io_outs_left_mult_io_o[27] ),
    .QN(_181_));
 DFFHQNx1_ASAP7_75t_R \io_outs_left_REG[28]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(\_io_outs_left_mult_io_o[28] ),
    .QN(_182_));
 DFFHQNx1_ASAP7_75t_R \io_outs_left_REG[29]$_DFF_P_  (.CLK(clknet_leaf_5_clock),
    .D(\_io_outs_left_mult_io_o[29] ),
    .QN(_183_));
 DFFHQNx1_ASAP7_75t_R \io_outs_left_REG[2]$_DFF_P_  (.CLK(clknet_leaf_5_clock),
    .D(\_io_outs_left_mult_io_o[2] ),
    .QN(_184_));
 DFFHQNx1_ASAP7_75t_R \io_outs_left_REG[30]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(\_io_outs_left_mult_io_o[30] ),
    .QN(_185_));
 DFFHQNx1_ASAP7_75t_R \io_outs_left_REG[31]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(\_io_outs_left_mult_io_o[31] ),
    .QN(_186_));
 DFFHQNx1_ASAP7_75t_R \io_outs_left_REG[3]$_DFF_P_  (.CLK(clknet_leaf_9_clock),
    .D(\_io_outs_left_mult_io_o[3] ),
    .QN(_187_));
 DFFHQNx1_ASAP7_75t_R \io_outs_left_REG[4]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(\_io_outs_left_mult_io_o[4] ),
    .QN(_188_));
 DFFHQNx1_ASAP7_75t_R \io_outs_left_REG[5]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(\_io_outs_left_mult_io_o[5] ),
    .QN(_189_));
 DFFHQNx1_ASAP7_75t_R \io_outs_left_REG[6]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(\_io_outs_left_mult_io_o[6] ),
    .QN(_190_));
 DFFHQNx1_ASAP7_75t_R \io_outs_left_REG[7]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(\_io_outs_left_mult_io_o[7] ),
    .QN(_191_));
 DFFHQNx1_ASAP7_75t_R \io_outs_left_REG[8]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(\_io_outs_left_mult_io_o[8] ),
    .QN(_192_));
 DFFHQNx1_ASAP7_75t_R \io_outs_left_REG[9]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(\_io_outs_left_mult_io_o[9] ),
    .QN(_193_));
 DFFHQNx1_ASAP7_75t_R \io_outs_right_REG[0]$_DFF_P_  (.CLK(clknet_leaf_20_clock),
    .D(\_io_outs_right_mult_io_o[0] ),
    .QN(_194_));
 DFFHQNx1_ASAP7_75t_R \io_outs_right_REG[10]$_DFF_P_  (.CLK(clknet_leaf_22_clock),
    .D(\_io_outs_right_mult_io_o[10] ),
    .QN(_195_));
 DFFHQNx1_ASAP7_75t_R \io_outs_right_REG[11]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(\_io_outs_right_mult_io_o[11] ),
    .QN(_196_));
 DFFHQNx1_ASAP7_75t_R \io_outs_right_REG[12]$_DFF_P_  (.CLK(clknet_leaf_22_clock),
    .D(\_io_outs_right_mult_io_o[12] ),
    .QN(_197_));
 DFFHQNx1_ASAP7_75t_R \io_outs_right_REG[13]$_DFF_P_  (.CLK(clknet_leaf_22_clock),
    .D(\_io_outs_right_mult_io_o[13] ),
    .QN(_198_));
 DFFHQNx1_ASAP7_75t_R \io_outs_right_REG[14]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(\_io_outs_right_mult_io_o[14] ),
    .QN(_199_));
 DFFHQNx1_ASAP7_75t_R \io_outs_right_REG[15]$_DFF_P_  (.CLK(clknet_leaf_23_clock),
    .D(\_io_outs_right_mult_io_o[15] ),
    .QN(_200_));
 DFFHQNx1_ASAP7_75t_R \io_outs_right_REG[16]$_DFF_P_  (.CLK(clknet_leaf_23_clock),
    .D(\_io_outs_right_mult_io_o[16] ),
    .QN(_201_));
 DFFHQNx1_ASAP7_75t_R \io_outs_right_REG[17]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(\_io_outs_right_mult_io_o[17] ),
    .QN(_202_));
 DFFHQNx1_ASAP7_75t_R \io_outs_right_REG[18]$_DFF_P_  (.CLK(clknet_leaf_23_clock),
    .D(\_io_outs_right_mult_io_o[18] ),
    .QN(_203_));
 DFFHQNx1_ASAP7_75t_R \io_outs_right_REG[19]$_DFF_P_  (.CLK(clknet_leaf_24_clock),
    .D(\_io_outs_right_mult_io_o[19] ),
    .QN(_204_));
 DFFHQNx1_ASAP7_75t_R \io_outs_right_REG[1]$_DFF_P_  (.CLK(clknet_leaf_22_clock),
    .D(\_io_outs_right_mult_io_o[1] ),
    .QN(_205_));
 DFFHQNx1_ASAP7_75t_R \io_outs_right_REG[20]$_DFF_P_  (.CLK(clknet_leaf_22_clock),
    .D(\_io_outs_right_mult_io_o[20] ),
    .QN(_206_));
 DFFHQNx1_ASAP7_75t_R \io_outs_right_REG[21]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(\_io_outs_right_mult_io_o[21] ),
    .QN(_207_));
 DFFHQNx1_ASAP7_75t_R \io_outs_right_REG[22]$_DFF_P_  (.CLK(clknet_leaf_25_clock),
    .D(\_io_outs_right_mult_io_o[22] ),
    .QN(_208_));
 DFFHQNx1_ASAP7_75t_R \io_outs_right_REG[23]$_DFF_P_  (.CLK(clknet_leaf_22_clock),
    .D(\_io_outs_right_mult_io_o[23] ),
    .QN(_209_));
 DFFHQNx1_ASAP7_75t_R \io_outs_right_REG[24]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(\_io_outs_right_mult_io_o[24] ),
    .QN(_210_));
 DFFHQNx1_ASAP7_75t_R \io_outs_right_REG[25]$_DFF_P_  (.CLK(clknet_leaf_24_clock),
    .D(\_io_outs_right_mult_io_o[25] ),
    .QN(_211_));
 DFFHQNx1_ASAP7_75t_R \io_outs_right_REG[26]$_DFF_P_  (.CLK(clknet_leaf_23_clock),
    .D(\_io_outs_right_mult_io_o[26] ),
    .QN(_212_));
 DFFHQNx1_ASAP7_75t_R \io_outs_right_REG[27]$_DFF_P_  (.CLK(clknet_leaf_24_clock),
    .D(\_io_outs_right_mult_io_o[27] ),
    .QN(_213_));
 DFFHQNx1_ASAP7_75t_R \io_outs_right_REG[28]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(\_io_outs_right_mult_io_o[28] ),
    .QN(_214_));
 DFFHQNx1_ASAP7_75t_R \io_outs_right_REG[29]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(\_io_outs_right_mult_io_o[29] ),
    .QN(_215_));
 DFFHQNx1_ASAP7_75t_R \io_outs_right_REG[2]$_DFF_P_  (.CLK(clknet_leaf_22_clock),
    .D(\_io_outs_right_mult_io_o[2] ),
    .QN(_216_));
 DFFHQNx1_ASAP7_75t_R \io_outs_right_REG[30]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(\_io_outs_right_mult_io_o[30] ),
    .QN(_217_));
 DFFHQNx1_ASAP7_75t_R \io_outs_right_REG[31]$_DFF_P_  (.CLK(clknet_leaf_22_clock),
    .D(\_io_outs_right_mult_io_o[31] ),
    .QN(_218_));
 DFFHQNx1_ASAP7_75t_R \io_outs_right_REG[3]$_DFF_P_  (.CLK(clknet_leaf_22_clock),
    .D(\_io_outs_right_mult_io_o[3] ),
    .QN(_219_));
 DFFHQNx1_ASAP7_75t_R \io_outs_right_REG[4]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(\_io_outs_right_mult_io_o[4] ),
    .QN(_220_));
 DFFHQNx1_ASAP7_75t_R \io_outs_right_REG[5]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(\_io_outs_right_mult_io_o[5] ),
    .QN(_221_));
 DFFHQNx1_ASAP7_75t_R \io_outs_right_REG[6]$_DFF_P_  (.CLK(clknet_leaf_24_clock),
    .D(\_io_outs_right_mult_io_o[6] ),
    .QN(_222_));
 DFFHQNx1_ASAP7_75t_R \io_outs_right_REG[7]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(\_io_outs_right_mult_io_o[7] ),
    .QN(_223_));
 DFFHQNx1_ASAP7_75t_R \io_outs_right_REG[8]$_DFF_P_  (.CLK(clknet_leaf_23_clock),
    .D(\_io_outs_right_mult_io_o[8] ),
    .QN(_224_));
 DFFHQNx1_ASAP7_75t_R \io_outs_right_REG[9]$_DFF_P_  (.CLK(clknet_leaf_24_clock),
    .D(\_io_outs_right_mult_io_o[9] ),
    .QN(_225_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up_REG[0]$_DFF_P_  (.CLK(clknet_leaf_14_clock),
    .D(\_io_outs_up_mult_io_o[0] ),
    .QN(_226_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up_REG[10]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(\_io_outs_up_mult_io_o[10] ),
    .QN(_227_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up_REG[11]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(\_io_outs_up_mult_io_o[11] ),
    .QN(_228_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up_REG[12]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(\_io_outs_up_mult_io_o[12] ),
    .QN(_229_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up_REG[13]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(\_io_outs_up_mult_io_o[13] ),
    .QN(_230_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up_REG[14]$_DFF_P_  (.CLK(clknet_leaf_13_clock),
    .D(\_io_outs_up_mult_io_o[14] ),
    .QN(_231_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up_REG[15]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(\_io_outs_up_mult_io_o[15] ),
    .QN(_232_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up_REG[16]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(\_io_outs_up_mult_io_o[16] ),
    .QN(_233_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up_REG[17]$_DFF_P_  (.CLK(clknet_leaf_9_clock),
    .D(\_io_outs_up_mult_io_o[17] ),
    .QN(_234_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up_REG[18]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(\_io_outs_up_mult_io_o[18] ),
    .QN(_235_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up_REG[19]$_DFF_P_  (.CLK(clknet_leaf_9_clock),
    .D(\_io_outs_up_mult_io_o[19] ),
    .QN(_236_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up_REG[1]$_DFF_P_  (.CLK(clknet_leaf_9_clock),
    .D(\_io_outs_up_mult_io_o[1] ),
    .QN(_237_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up_REG[20]$_DFF_P_  (.CLK(clknet_leaf_14_clock),
    .D(\_io_outs_up_mult_io_o[20] ),
    .QN(_238_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up_REG[21]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(\_io_outs_up_mult_io_o[21] ),
    .QN(_239_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up_REG[22]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(\_io_outs_up_mult_io_o[22] ),
    .QN(_240_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up_REG[23]$_DFF_P_  (.CLK(clknet_leaf_9_clock),
    .D(\_io_outs_up_mult_io_o[23] ),
    .QN(_241_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up_REG[24]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(\_io_outs_up_mult_io_o[24] ),
    .QN(_242_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up_REG[25]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(\_io_outs_up_mult_io_o[25] ),
    .QN(_243_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up_REG[26]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(\_io_outs_up_mult_io_o[26] ),
    .QN(_244_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up_REG[27]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(\_io_outs_up_mult_io_o[27] ),
    .QN(_245_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up_REG[28]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(\_io_outs_up_mult_io_o[28] ),
    .QN(_246_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up_REG[29]$_DFF_P_  (.CLK(clknet_leaf_14_clock),
    .D(\_io_outs_up_mult_io_o[29] ),
    .QN(_247_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up_REG[2]$_DFF_P_  (.CLK(clknet_leaf_14_clock),
    .D(\_io_outs_up_mult_io_o[2] ),
    .QN(_248_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up_REG[30]$_DFF_P_  (.CLK(clknet_leaf_9_clock),
    .D(\_io_outs_up_mult_io_o[30] ),
    .QN(_249_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up_REG[31]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(\_io_outs_up_mult_io_o[31] ),
    .QN(_250_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up_REG[3]$_DFF_P_  (.CLK(clknet_leaf_13_clock),
    .D(\_io_outs_up_mult_io_o[3] ),
    .QN(_251_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up_REG[4]$_DFF_P_  (.CLK(clknet_leaf_14_clock),
    .D(\_io_outs_up_mult_io_o[4] ),
    .QN(_252_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up_REG[5]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(\_io_outs_up_mult_io_o[5] ),
    .QN(_253_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up_REG[6]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(\_io_outs_up_mult_io_o[6] ),
    .QN(_254_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up_REG[7]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(\_io_outs_up_mult_io_o[7] ),
    .QN(_255_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up_REG[8]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(\_io_outs_up_mult_io_o[8] ),
    .QN(_256_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up_REG[9]$_DFF_P_  (.CLK(clknet_leaf_14_clock),
    .D(\_io_outs_up_mult_io_o[9] ),
    .QN(_000_));
 Multiplier io_outs_down_mult (.clknet_leaf_32_clock_i(clknet_leaf_32_clock),
    .clknet_leaf_30_clock_i(clknet_leaf_30_clock),
    .clknet_leaf_29_clock_i(clknet_leaf_29_clock),
    .clknet_leaf_28_clock_i(clknet_leaf_28_clock),
    .clknet_leaf_12_clock_i(clknet_leaf_12_clock),
    .clknet_leaf_4_clock_i(clknet_leaf_4_clock),
    .clknet_leaf_3_clock_i(clknet_leaf_3_clock),
    .io_a({\REG_1[31] ,
    \REG_1[30] ,
    \REG_1[29] ,
    \REG_1[28] ,
    \REG_1[27] ,
    \REG_1[26] ,
    \REG_1[25] ,
    \REG_1[24] ,
    \REG_1[23] ,
    \REG_1[22] ,
    \REG_1[21] ,
    \REG_1[20] ,
    \REG_1[19] ,
    \REG_1[18] ,
    \REG_1[17] ,
    \REG_1[16] ,
    \REG_1[15] ,
    \REG_1[14] ,
    \REG_1[13] ,
    \REG_1[12] ,
    \REG_1[11] ,
    \REG_1[10] ,
    \REG_1[9] ,
    \REG_1[8] ,
    \REG_1[7] ,
    \REG_1[6] ,
    \REG_1[5] ,
    \REG_1[4] ,
    \REG_1[3] ,
    \REG_1[2] ,
    \REG_1[1] ,
    \REG_1[0] }),
    .io_b({\REG_4[31] ,
    \REG_4[30] ,
    \REG_4[29] ,
    \REG_4[28] ,
    \REG_4[27] ,
    \REG_4[26] ,
    \REG_4[25] ,
    \REG_4[24] ,
    \REG_4[23] ,
    \REG_4[22] ,
    \REG_4[21] ,
    \REG_4[20] ,
    \REG_4[19] ,
    \REG_4[18] ,
    \REG_4[17] ,
    \REG_4[16] ,
    \REG_4[15] ,
    \REG_4[14] ,
    \REG_4[13] ,
    \REG_4[12] ,
    \REG_4[11] ,
    \REG_4[10] ,
    \REG_4[9] ,
    \REG_4[8] ,
    \REG_4[7] ,
    \REG_4[6] ,
    \REG_4[5] ,
    \REG_4[4] ,
    \REG_4[3] ,
    \REG_4[2] ,
    \REG_4[1] ,
    \REG_4[0] }),
    .io_o({\_io_outs_down_mult_io_o[31] ,
    \_io_outs_down_mult_io_o[30] ,
    \_io_outs_down_mult_io_o[29] ,
    \_io_outs_down_mult_io_o[28] ,
    \_io_outs_down_mult_io_o[27] ,
    \_io_outs_down_mult_io_o[26] ,
    \_io_outs_down_mult_io_o[25] ,
    \_io_outs_down_mult_io_o[24] ,
    \_io_outs_down_mult_io_o[23] ,
    \_io_outs_down_mult_io_o[22] ,
    \_io_outs_down_mult_io_o[21] ,
    \_io_outs_down_mult_io_o[20] ,
    \_io_outs_down_mult_io_o[19] ,
    \_io_outs_down_mult_io_o[18] ,
    \_io_outs_down_mult_io_o[17] ,
    \_io_outs_down_mult_io_o[16] ,
    \_io_outs_down_mult_io_o[15] ,
    \_io_outs_down_mult_io_o[14] ,
    \_io_outs_down_mult_io_o[13] ,
    \_io_outs_down_mult_io_o[12] ,
    \_io_outs_down_mult_io_o[11] ,
    \_io_outs_down_mult_io_o[10] ,
    \_io_outs_down_mult_io_o[9] ,
    \_io_outs_down_mult_io_o[8] ,
    \_io_outs_down_mult_io_o[7] ,
    \_io_outs_down_mult_io_o[6] ,
    \_io_outs_down_mult_io_o[5] ,
    \_io_outs_down_mult_io_o[4] ,
    \_io_outs_down_mult_io_o[3] ,
    \_io_outs_down_mult_io_o[2] ,
    \_io_outs_down_mult_io_o[1] ,
    \_io_outs_down_mult_io_o[0] }));
 Multiplier_io_outs_left_mult io_outs_left_mult (.clknet_leaf_21_clock_i(clknet_leaf_21_clock),
    .clknet_leaf_20_clock_i(clknet_leaf_20_clock),
    .clknet_leaf_13_clock_i(clknet_leaf_13_clock),
    .clknet_leaf_12_clock_i(clknet_leaf_12_clock),
    .clknet_leaf_7_clock_i(clknet_leaf_7_clock),
    .clknet_leaf_5_clock_i(clknet_leaf_5_clock),
    .io_a({\REG[31] ,
    \REG[30] ,
    \REG[29] ,
    \REG[28] ,
    \REG[27] ,
    \REG[26] ,
    \REG[25] ,
    \REG[24] ,
    \REG[23] ,
    \REG[22] ,
    \REG[21] ,
    \REG[20] ,
    \REG[19] ,
    \REG[18] ,
    \REG[17] ,
    \REG[16] ,
    \REG[15] ,
    \REG[14] ,
    \REG[13] ,
    \REG[12] ,
    \REG[11] ,
    \REG[10] ,
    \REG[9] ,
    \REG[8] ,
    \REG[7] ,
    \REG[6] ,
    \REG[5] ,
    \REG[4] ,
    \REG[3] ,
    \REG[2] ,
    \REG[1] ,
    \REG[0] }),
    .io_b({\REG_1[31] ,
    \REG_1[30] ,
    \REG_1[29] ,
    \REG_1[28] ,
    \REG_1[27] ,
    \REG_1[26] ,
    \REG_1[25] ,
    \REG_1[24] ,
    \REG_1[23] ,
    \REG_1[22] ,
    \REG_1[21] ,
    \REG_1[20] ,
    \REG_1[19] ,
    \REG_1[18] ,
    \REG_1[17] ,
    \REG_1[16] ,
    \REG_1[15] ,
    \REG_1[14] ,
    \REG_1[13] ,
    \REG_1[12] ,
    \REG_1[11] ,
    \REG_1[10] ,
    \REG_1[9] ,
    \REG_1[8] ,
    \REG_1[7] ,
    \REG_1[6] ,
    \REG_1[5] ,
    \REG_1[4] ,
    \REG_1[3] ,
    \REG_1[2] ,
    \REG_1[1] ,
    \REG_1[0] }),
    .io_o({\_io_outs_left_mult_io_o[31] ,
    \_io_outs_left_mult_io_o[30] ,
    \_io_outs_left_mult_io_o[29] ,
    \_io_outs_left_mult_io_o[28] ,
    \_io_outs_left_mult_io_o[27] ,
    \_io_outs_left_mult_io_o[26] ,
    \_io_outs_left_mult_io_o[25] ,
    \_io_outs_left_mult_io_o[24] ,
    \_io_outs_left_mult_io_o[23] ,
    \_io_outs_left_mult_io_o[22] ,
    \_io_outs_left_mult_io_o[21] ,
    \_io_outs_left_mult_io_o[20] ,
    \_io_outs_left_mult_io_o[19] ,
    \_io_outs_left_mult_io_o[18] ,
    \_io_outs_left_mult_io_o[17] ,
    \_io_outs_left_mult_io_o[16] ,
    \_io_outs_left_mult_io_o[15] ,
    \_io_outs_left_mult_io_o[14] ,
    \_io_outs_left_mult_io_o[13] ,
    \_io_outs_left_mult_io_o[12] ,
    \_io_outs_left_mult_io_o[11] ,
    \_io_outs_left_mult_io_o[10] ,
    \_io_outs_left_mult_io_o[9] ,
    \_io_outs_left_mult_io_o[8] ,
    \_io_outs_left_mult_io_o[7] ,
    \_io_outs_left_mult_io_o[6] ,
    \_io_outs_left_mult_io_o[5] ,
    \_io_outs_left_mult_io_o[4] ,
    \_io_outs_left_mult_io_o[3] ,
    \_io_outs_left_mult_io_o[2] ,
    \_io_outs_left_mult_io_o[1] ,
    \_io_outs_left_mult_io_o[0] }));
 Multiplier_io_outs_right_mult io_outs_right_mult (.clknet_leaf_30_clock_i(clknet_leaf_30_clock),
    .clknet_leaf_29_clock_i(clknet_leaf_29_clock),
    .clknet_leaf_21_clock_i(clknet_leaf_21_clock),
    .clknet_leaf_5_clock_i(clknet_leaf_5_clock),
    .clknet_leaf_4_clock_i(clknet_leaf_4_clock),
    .clknet_leaf_3_clock_i(clknet_leaf_3_clock),
    .io_a({\REG_4[31] ,
    \REG_4[30] ,
    \REG_4[29] ,
    \REG_4[28] ,
    \REG_4[27] ,
    \REG_4[26] ,
    \REG_4[25] ,
    \REG_4[24] ,
    \REG_4[23] ,
    \REG_4[22] ,
    \REG_4[21] ,
    \REG_4[20] ,
    \REG_4[19] ,
    \REG_4[18] ,
    \REG_4[17] ,
    \REG_4[16] ,
    \REG_4[15] ,
    \REG_4[14] ,
    \REG_4[13] ,
    \REG_4[12] ,
    \REG_4[11] ,
    \REG_4[10] ,
    \REG_4[9] ,
    \REG_4[8] ,
    \REG_4[7] ,
    \REG_4[6] ,
    \REG_4[5] ,
    \REG_4[4] ,
    \REG_4[3] ,
    \REG_4[2] ,
    \REG_4[1] ,
    \REG_4[0] }),
    .io_b({\REG_2[31] ,
    \REG_2[30] ,
    \REG_2[29] ,
    \REG_2[28] ,
    \REG_2[27] ,
    \REG_2[26] ,
    \REG_2[25] ,
    \REG_2[24] ,
    \REG_2[23] ,
    \REG_2[22] ,
    \REG_2[21] ,
    \REG_2[20] ,
    \REG_2[19] ,
    \REG_2[18] ,
    \REG_2[17] ,
    \REG_2[16] ,
    \REG_2[15] ,
    \REG_2[14] ,
    \REG_2[13] ,
    \REG_2[12] ,
    \REG_2[11] ,
    \REG_2[10] ,
    \REG_2[9] ,
    \REG_2[8] ,
    \REG_2[7] ,
    \REG_2[6] ,
    \REG_2[5] ,
    \REG_2[4] ,
    \REG_2[3] ,
    \REG_2[2] ,
    \REG_2[1] ,
    \REG_2[0] }),
    .io_o({\_io_outs_right_mult_io_o[31] ,
    \_io_outs_right_mult_io_o[30] ,
    \_io_outs_right_mult_io_o[29] ,
    \_io_outs_right_mult_io_o[28] ,
    \_io_outs_right_mult_io_o[27] ,
    \_io_outs_right_mult_io_o[26] ,
    \_io_outs_right_mult_io_o[25] ,
    \_io_outs_right_mult_io_o[24] ,
    \_io_outs_right_mult_io_o[23] ,
    \_io_outs_right_mult_io_o[22] ,
    \_io_outs_right_mult_io_o[21] ,
    \_io_outs_right_mult_io_o[20] ,
    \_io_outs_right_mult_io_o[19] ,
    \_io_outs_right_mult_io_o[18] ,
    \_io_outs_right_mult_io_o[17] ,
    \_io_outs_right_mult_io_o[16] ,
    \_io_outs_right_mult_io_o[15] ,
    \_io_outs_right_mult_io_o[14] ,
    \_io_outs_right_mult_io_o[13] ,
    \_io_outs_right_mult_io_o[12] ,
    \_io_outs_right_mult_io_o[11] ,
    \_io_outs_right_mult_io_o[10] ,
    \_io_outs_right_mult_io_o[9] ,
    \_io_outs_right_mult_io_o[8] ,
    \_io_outs_right_mult_io_o[7] ,
    \_io_outs_right_mult_io_o[6] ,
    \_io_outs_right_mult_io_o[5] ,
    \_io_outs_right_mult_io_o[4] ,
    \_io_outs_right_mult_io_o[3] ,
    \_io_outs_right_mult_io_o[2] ,
    \_io_outs_right_mult_io_o[1] ,
    \_io_outs_right_mult_io_o[0] }));
 Multiplier_io_outs_up_mult io_outs_up_mult (.clknet_leaf_14_clock_i(clknet_leaf_14_clock),
    .clknet_leaf_13_clock_i(clknet_leaf_13_clock),
    .clknet_leaf_11_clock_i(clknet_leaf_11_clock),
    .clknet_leaf_9_clock_i(clknet_leaf_9_clock),
    .clknet_leaf_7_clock_i(clknet_leaf_7_clock),
    .clknet_leaf_5_clock_i(clknet_leaf_5_clock),
    .clknet_leaf_4_clock_i(clknet_leaf_4_clock),
    .clknet_leaf_3_clock_i(clknet_leaf_3_clock),
    .io_a({\REG_2[31] ,
    \REG_2[30] ,
    \REG_2[29] ,
    \REG_2[28] ,
    \REG_2[27] ,
    \REG_2[26] ,
    \REG_2[25] ,
    \REG_2[24] ,
    \REG_2[23] ,
    \REG_2[22] ,
    \REG_2[21] ,
    \REG_2[20] ,
    \REG_2[19] ,
    \REG_2[18] ,
    \REG_2[17] ,
    \REG_2[16] ,
    \REG_2[15] ,
    \REG_2[14] ,
    \REG_2[13] ,
    \REG_2[12] ,
    \REG_2[11] ,
    \REG_2[10] ,
    \REG_2[9] ,
    \REG_2[8] ,
    \REG_2[7] ,
    \REG_2[6] ,
    \REG_2[5] ,
    \REG_2[4] ,
    \REG_2[3] ,
    \REG_2[2] ,
    \REG_2[1] ,
    \REG_2[0] }),
    .io_b({\REG[31] ,
    \REG[30] ,
    \REG[29] ,
    \REG[28] ,
    \REG[27] ,
    \REG[26] ,
    \REG[25] ,
    \REG[24] ,
    \REG[23] ,
    \REG[22] ,
    \REG[21] ,
    \REG[20] ,
    \REG[19] ,
    \REG[18] ,
    \REG[17] ,
    \REG[16] ,
    \REG[15] ,
    \REG[14] ,
    \REG[13] ,
    \REG[12] ,
    \REG[11] ,
    \REG[10] ,
    \REG[9] ,
    \REG[8] ,
    \REG[7] ,
    \REG[6] ,
    \REG[5] ,
    \REG[4] ,
    \REG[3] ,
    \REG[2] ,
    \REG[1] ,
    \REG[0] }),
    .io_o({\_io_outs_up_mult_io_o[31] ,
    \_io_outs_up_mult_io_o[30] ,
    \_io_outs_up_mult_io_o[29] ,
    \_io_outs_up_mult_io_o[28] ,
    \_io_outs_up_mult_io_o[27] ,
    \_io_outs_up_mult_io_o[26] ,
    \_io_outs_up_mult_io_o[25] ,
    \_io_outs_up_mult_io_o[24] ,
    \_io_outs_up_mult_io_o[23] ,
    \_io_outs_up_mult_io_o[22] ,
    \_io_outs_up_mult_io_o[21] ,
    \_io_outs_up_mult_io_o[20] ,
    \_io_outs_up_mult_io_o[19] ,
    \_io_outs_up_mult_io_o[18] ,
    \_io_outs_up_mult_io_o[17] ,
    \_io_outs_up_mult_io_o[16] ,
    \_io_outs_up_mult_io_o[15] ,
    \_io_outs_up_mult_io_o[14] ,
    \_io_outs_up_mult_io_o[13] ,
    \_io_outs_up_mult_io_o[12] ,
    \_io_outs_up_mult_io_o[11] ,
    \_io_outs_up_mult_io_o[10] ,
    \_io_outs_up_mult_io_o[9] ,
    \_io_outs_up_mult_io_o[8] ,
    \_io_outs_up_mult_io_o[7] ,
    \_io_outs_up_mult_io_o[6] ,
    \_io_outs_up_mult_io_o[5] ,
    \_io_outs_up_mult_io_o[4] ,
    \_io_outs_up_mult_io_o[3] ,
    \_io_outs_up_mult_io_o[2] ,
    \_io_outs_up_mult_io_o[1] ,
    \_io_outs_up_mult_io_o[0] }));
endmodule
module Multiplier (clknet_leaf_32_clock_i,
    clknet_leaf_30_clock_i,
    clknet_leaf_29_clock_i,
    clknet_leaf_28_clock_i,
    clknet_leaf_12_clock_i,
    clknet_leaf_4_clock_i,
    clknet_leaf_3_clock_i,
    io_a,
    io_b,
    io_o);
 input clknet_leaf_32_clock_i;
 input clknet_leaf_30_clock_i;
 input clknet_leaf_29_clock_i;
 input clknet_leaf_28_clock_i;
 input clknet_leaf_12_clock_i;
 input clknet_leaf_4_clock_i;
 input clknet_leaf_3_clock_i;
 input [31:0] io_a;
 input [31:0] io_b;
 output [31:0] io_o;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire \mod.$1 ;
 wire \mod.$2 ;
 wire \mod.$3 ;
 wire \mod.$4 ;
 wire \mod.$5 ;
 wire \mod.$54 ;
 wire \mod.$55 ;
 wire \mod.$56 ;
 wire \mod.$57 ;
 wire \mod.$6 ;
 wire \mod.a_registered[0] ;
 wire \mod.a_registered[1] ;
 wire \mod.a_registered[2] ;
 wire \mod.a_registered[3] ;
 wire \mod.b_registered[0] ;
 wire \mod.b_registered[1] ;
 wire \mod.b_registered[2] ;
 wire \mod.b_registered[3] ;
 wire \mod.booth_b0_m0 ;
 wire \mod.booth_b0_m1 ;
 wire \mod.booth_b0_m2 ;
 wire \mod.booth_b0_m3 ;
 wire \mod.booth_b2_m0 ;
 wire \mod.booth_b2_m1 ;
 wire \mod.c ;
 wire \mod.con$4400 ;
 wire \mod.con$4402 ;
 wire \mod.final_a_registered[0] ;
 wire \mod.final_a_registered[1] ;
 wire \mod.final_a_registered[2] ;
 wire \mod.final_a_registered[3] ;
 wire \mod.final_adder.$signal ;
 wire \mod.final_adder.$signal$10 ;
 wire \mod.final_adder.$signal$263 ;
 wire \mod.final_adder.$signal$264 ;
 wire \mod.final_adder.$signal$265 ;
 wire \mod.final_adder.$signal$6 ;
 wire \mod.final_adder.$signal$8 ;
 wire \mod.final_adder.con ;
 wire \mod.final_adder.con$137 ;
 wire \mod.final_adder.con$139 ;
 wire \mod.final_adder.con$141 ;
 wire \mod.final_adder.g_new ;
 wire \mod.final_adder.g_new$477 ;
 wire \mod.final_adder.sn ;
 wire \mod.final_adder.sn$138 ;
 wire \mod.final_adder.sn$140 ;
 wire \mod.final_adder.sn$142 ;
 wire \mod.final_b_registered[0] ;
 wire \mod.final_b_registered[2] ;
 wire \mod.final_b_registered[3] ;
 wire \mod.pp_row0_0 ;
 wire \mod.pp_row0_1 ;
 wire \mod.pp_row1_0 ;
 wire \mod.pp_row2_0 ;
 wire \mod.pp_row2_1 ;
 wire \mod.pp_row2_2 ;
 wire \mod.pp_row3_0 ;
 wire \mod.pp_row3_1 ;
 wire \mod.s ;
 wire \mod.s$1260 ;
 wire \mod.sel_0 ;
 wire \mod.sel_0$1365 ;
 wire \mod.sel_1 ;
 wire \mod.sel_1$1366 ;
 wire \mod.sn$4401 ;
 wire \mod.sn$4403 ;
 wire \mod.t ;
 wire \mod.t$1976 ;
 wire \mod.t$1977 ;
 wire \mod.t$1978 ;
 wire \mod.t$2009 ;
 wire \mod.t$2010 ;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;

 TIELOx1_ASAP7_75t_R \mod.final_adder.U$375_163  (.L(net161));
 TIELOx1_ASAP7_75t_R \mod.final_adder.U$3_162  (.L(net160));
 TIELOx1_ASAP7_75t_R \mod.U$603_161  (.L(net159));
 TIELOx1_ASAP7_75t_R \mod.U$531_160  (.L(net158));
 TIELOx1_ASAP7_75t_R \mod.U$530_159  (.L(net157));
 TIELOx1_ASAP7_75t_R \mod.U$529_158  (.L(net156));
 TIELOx1_ASAP7_75t_R \mod.U$526_157  (.L(net155));
 TIELOx1_ASAP7_75t_R _83__156 (.L(io_o[31]));
 TIELOx1_ASAP7_75t_R _82__155 (.L(io_o[30]));
 TIELOx1_ASAP7_75t_R _81__154 (.L(io_o[29]));
 TIELOx1_ASAP7_75t_R _80__153 (.L(io_o[28]));
 TIELOx1_ASAP7_75t_R _79__152 (.L(io_o[27]));
 TIELOx1_ASAP7_75t_R _78__151 (.L(io_o[26]));
 TIELOx1_ASAP7_75t_R _77__150 (.L(io_o[25]));
 TIELOx1_ASAP7_75t_R _76__149 (.L(io_o[24]));
 TIELOx1_ASAP7_75t_R _75__148 (.L(io_o[23]));
 TIELOx1_ASAP7_75t_R _74__147 (.L(io_o[22]));
 TIELOx1_ASAP7_75t_R _73__146 (.L(io_o[21]));
 TIELOx1_ASAP7_75t_R _72__145 (.L(io_o[20]));
 TIELOx1_ASAP7_75t_R _71__144 (.L(io_o[19]));
 TIELOx1_ASAP7_75t_R _70__143 (.L(io_o[18]));
 TIELOx1_ASAP7_75t_R _69__142 (.L(io_o[17]));
 TIELOx1_ASAP7_75t_R _68__141 (.L(io_o[16]));
 TIELOx1_ASAP7_75t_R _67__140 (.L(io_o[15]));
 TIELOx1_ASAP7_75t_R _66__139 (.L(io_o[14]));
 TIELOx1_ASAP7_75t_R _65__138 (.L(io_o[13]));
 TIELOx1_ASAP7_75t_R _64__137 (.L(io_o[12]));
 TIELOx1_ASAP7_75t_R _63__136 (.L(io_o[11]));
 TIELOx1_ASAP7_75t_R _62__135 (.L(io_o[10]));
 TIELOx1_ASAP7_75t_R _61__134 (.L(io_o[9]));
 TIELOx1_ASAP7_75t_R _60__133 (.L(io_o[8]));
 TIELOx1_ASAP7_75t_R _59__132 (.L(io_o[7]));
 TIELOx1_ASAP7_75t_R _58__131 (.L(io_o[6]));
 TIELOx1_ASAP7_75t_R _57__130 (.L(io_o[5]));
 TIELOx1_ASAP7_75t_R _56__129 (.L(io_o[4]));
 INVx3_ASAP7_75t_R _28_ (.A(_00_),
    .Y(\mod.pp_row3_1 ));
 INVx3_ASAP7_75t_R _29_ (.A(_01_),
    .Y(\mod.a_registered[0] ));
 INVx3_ASAP7_75t_R _30_ (.A(_02_),
    .Y(\mod.a_registered[1] ));
 INVx3_ASAP7_75t_R _31_ (.A(_03_),
    .Y(\mod.a_registered[2] ));
 INVx3_ASAP7_75t_R _32_ (.A(_04_),
    .Y(\mod.a_registered[3] ));
 INVx3_ASAP7_75t_R _33_ (.A(_05_),
    .Y(\mod.b_registered[0] ));
 INVx3_ASAP7_75t_R _34_ (.A(_06_),
    .Y(\mod.b_registered[1] ));
 INVx3_ASAP7_75t_R _35_ (.A(_07_),
    .Y(\mod.b_registered[2] ));
 INVx3_ASAP7_75t_R _36_ (.A(_08_),
    .Y(\mod.b_registered[3] ));
 INVx3_ASAP7_75t_R _37_ (.A(_09_),
    .Y(\mod.final_a_registered[0] ));
 INVx3_ASAP7_75t_R _38_ (.A(_10_),
    .Y(\mod.final_a_registered[1] ));
 INVx3_ASAP7_75t_R _39_ (.A(_11_),
    .Y(\mod.final_a_registered[2] ));
 INVx3_ASAP7_75t_R _40_ (.A(_12_),
    .Y(\mod.final_a_registered[3] ));
 INVx3_ASAP7_75t_R _41_ (.A(_13_),
    .Y(\mod.final_b_registered[0] ));
 INVx3_ASAP7_75t_R _42_ (.A(_14_),
    .Y(\mod.final_b_registered[2] ));
 INVx3_ASAP7_75t_R _43_ (.A(_15_),
    .Y(\mod.final_b_registered[3] ));
 INVx3_ASAP7_75t_R _44_ (.A(_16_),
    .Y(io_o[0]));
 INVx3_ASAP7_75t_R _45_ (.A(_17_),
    .Y(io_o[1]));
 INVx3_ASAP7_75t_R _46_ (.A(_18_),
    .Y(io_o[2]));
 INVx3_ASAP7_75t_R _47_ (.A(_19_),
    .Y(io_o[3]));
 INVx3_ASAP7_75t_R _48_ (.A(_20_),
    .Y(\mod.pp_row0_0 ));
 INVx3_ASAP7_75t_R _49_ (.A(_21_),
    .Y(\mod.pp_row0_1 ));
 INVx3_ASAP7_75t_R _50_ (.A(_22_),
    .Y(\mod.pp_row1_0 ));
 INVx3_ASAP7_75t_R _51_ (.A(_23_),
    .Y(\mod.pp_row2_0 ));
 INVx3_ASAP7_75t_R _52_ (.A(_24_),
    .Y(\mod.pp_row2_1 ));
 INVx3_ASAP7_75t_R _53_ (.A(_25_),
    .Y(\mod.pp_row2_2 ));
 INVx3_ASAP7_75t_R _54_ (.A(_26_),
    .Y(\mod.pp_row3_0 ));
 INVx1_ASAP7_75t_R \mod.U$2674  (.A(\mod.con$4400 ),
    .Y(\mod.c ));
 INVx1_ASAP7_75t_R \mod.U$2675  (.A(\mod.sn$4401 ),
    .Y(\mod.s ));
 INVx1_ASAP7_75t_R \mod.U$2677  (.A(\mod.sn$4403 ),
    .Y(\mod.s$1260 ));
 INVx1_ASAP7_75t_R \mod.U$526  (.A(net155),
    .Y(\mod.$1 ));
 INVx1_ASAP7_75t_R \mod.U$527  (.A(\mod.a_registered[0] ),
    .Y(\mod.$2 ));
 INVx1_ASAP7_75t_R \mod.U$528  (.A(\mod.a_registered[1] ),
    .Y(\mod.$3 ));
 AO33x2_ASAP7_75t_R \mod.U$529  (.A1(\mod.$3 ),
    .A2(\mod.a_registered[0] ),
    .A3(net156),
    .B1(\mod.a_registered[1] ),
    .B2(\mod.$2 ),
    .B3(\mod.$1 ),
    .Y(\mod.sel_0 ));
 XOR2x1_ASAP7_75t_R \mod.U$530  (.A(\mod.a_registered[0] ),
    .Y(\mod.sel_1 ),
    .B(net157));
 AO22x1_ASAP7_75t_R \mod.U$531  (.A1(net158),
    .A2(\mod.sel_0 ),
    .B1(\mod.b_registered[0] ),
    .B2(\mod.sel_1 ),
    .Y(\mod.t ));
 XOR2x1_ASAP7_75t_R \mod.U$532  (.A(\mod.t ),
    .Y(\mod.booth_b0_m0 ),
    .B(\mod.a_registered[1] ));
 AO22x1_ASAP7_75t_R \mod.U$533  (.A1(\mod.b_registered[0] ),
    .A2(\mod.sel_0 ),
    .B1(\mod.b_registered[1] ),
    .B2(\mod.sel_1 ),
    .Y(\mod.t$1976 ));
 XOR2x1_ASAP7_75t_R \mod.U$534  (.A(\mod.t$1976 ),
    .Y(\mod.booth_b0_m1 ),
    .B(\mod.a_registered[1] ));
 AO22x1_ASAP7_75t_R \mod.U$535  (.A1(\mod.b_registered[1] ),
    .A2(\mod.sel_0 ),
    .B1(\mod.b_registered[2] ),
    .B2(\mod.sel_1 ),
    .Y(\mod.t$1977 ));
 XOR2x1_ASAP7_75t_R \mod.U$536  (.A(\mod.t$1977 ),
    .Y(\mod.booth_b0_m2 ),
    .B(\mod.a_registered[1] ));
 AO22x1_ASAP7_75t_R \mod.U$537  (.A1(\mod.b_registered[2] ),
    .A2(\mod.sel_0 ),
    .B1(\mod.b_registered[3] ),
    .B2(\mod.sel_1 ),
    .Y(\mod.t$1978 ));
 XOR2x1_ASAP7_75t_R \mod.U$538  (.A(\mod.t$1978 ),
    .Y(\mod.booth_b0_m3 ),
    .B(\mod.a_registered[1] ));
 INVx1_ASAP7_75t_R \mod.U$598  (.A(\mod.a_registered[1] ),
    .Y(\mod.$4 ));
 INVx1_ASAP7_75t_R \mod.U$599  (.A(\mod.a_registered[2] ),
    .Y(\mod.$5 ));
 INVx1_ASAP7_75t_R \mod.U$600  (.A(\mod.a_registered[3] ),
    .Y(\mod.$6 ));
 AO33x2_ASAP7_75t_R \mod.U$601  (.A1(\mod.$6 ),
    .A2(\mod.a_registered[2] ),
    .A3(\mod.a_registered[1] ),
    .B1(\mod.a_registered[3] ),
    .B2(\mod.$5 ),
    .B3(\mod.$4 ),
    .Y(\mod.sel_0$1365 ));
 XOR2x1_ASAP7_75t_R \mod.U$602  (.A(\mod.a_registered[2] ),
    .Y(\mod.sel_1$1366 ),
    .B(\mod.a_registered[1] ));
 AO22x1_ASAP7_75t_R \mod.U$603  (.A1(net159),
    .A2(\mod.sel_0$1365 ),
    .B1(\mod.b_registered[0] ),
    .B2(\mod.sel_1$1366 ),
    .Y(\mod.t$2009 ));
 XOR2x1_ASAP7_75t_R \mod.U$604  (.A(\mod.t$2009 ),
    .Y(\mod.booth_b2_m0 ),
    .B(\mod.a_registered[3] ));
 AO22x1_ASAP7_75t_R \mod.U$605  (.A1(\mod.b_registered[0] ),
    .A2(\mod.sel_0$1365 ),
    .B1(\mod.b_registered[1] ),
    .B2(\mod.sel_1$1366 ),
    .Y(\mod.t$2010 ));
 XOR2x1_ASAP7_75t_R \mod.U$606  (.A(\mod.t$2010 ),
    .Y(\mod.booth_b2_m1 ),
    .B(\mod.a_registered[3] ));
 DFFHQNx1_ASAP7_75t_R \mod.a_registered[0]$_DFF_P_  (.CLK(clknet_leaf_4_clock_i),
    .D(io_a[0]),
    .QN(_01_));
 DFFHQNx1_ASAP7_75t_R \mod.a_registered[1]$_DFF_P_  (.CLK(clknet_leaf_12_clock_i),
    .D(io_a[1]),
    .QN(_02_));
 DFFHQNx1_ASAP7_75t_R \mod.a_registered[2]$_DFF_P_  (.CLK(clknet_leaf_4_clock_i),
    .D(io_a[2]),
    .QN(_03_));
 DFFHQNx1_ASAP7_75t_R \mod.a_registered[3]$_DFF_P_  (.CLK(clknet_leaf_29_clock_i),
    .D(io_a[3]),
    .QN(_04_));
 DFFHQNx1_ASAP7_75t_R \mod.b_registered[0]$_DFF_P_  (.CLK(clknet_leaf_3_clock_i),
    .D(io_b[0]),
    .QN(_05_));
 DFFHQNx1_ASAP7_75t_R \mod.b_registered[1]$_DFF_P_  (.CLK(clknet_leaf_3_clock_i),
    .D(io_b[1]),
    .QN(_06_));
 DFFHQNx1_ASAP7_75t_R \mod.b_registered[2]$_DFF_P_  (.CLK(clknet_leaf_3_clock_i),
    .D(io_b[2]),
    .QN(_07_));
 DFFHQNx1_ASAP7_75t_R \mod.b_registered[3]$_DFF_P_  (.CLK(clknet_leaf_3_clock_i),
    .D(io_b[3]),
    .QN(_08_));
 HAxp5_ASAP7_75t_R \mod.dadda_ha_5_2_0  (.A(\mod.pp_row2_0 ),
    .B(\mod.pp_row2_1 ),
    .CON(\mod.con$4400 ),
    .SN(\mod.sn$4401 ));
 HAxp5_ASAP7_75t_R \mod.dadda_ha_5_3_0  (.A(\mod.pp_row3_0 ),
    .B(\mod.pp_row3_1 ),
    .CON(\mod.con$4402 ),
    .SN(\mod.sn$4403 ));
 DFFHQNx1_ASAP7_75t_R \mod.final_a_registered[0]$_DFF_P_  (.CLK(clknet_leaf_30_clock_i),
    .D(\mod.pp_row0_0 ),
    .QN(_09_));
 DFFHQNx1_ASAP7_75t_R \mod.final_a_registered[1]$_DFF_P_  (.CLK(clknet_leaf_30_clock_i),
    .D(\mod.pp_row1_0 ),
    .QN(_10_));
 DFFHQNx1_ASAP7_75t_R \mod.final_a_registered[2]$_DFF_P_  (.CLK(clknet_leaf_28_clock_i),
    .D(\mod.pp_row2_2 ),
    .QN(_11_));
 DFFHQNx1_ASAP7_75t_R \mod.final_a_registered[3]$_DFF_P_  (.CLK(clknet_leaf_28_clock_i),
    .D(\mod.c ),
    .QN(_12_));
 HAxp5_ASAP7_75t_R \mod.final_adder.U$0  (.A(\mod.final_a_registered[0] ),
    .B(\mod.final_b_registered[0] ),
    .CON(\mod.final_adder.con ),
    .SN(\mod.final_adder.sn ));
 INVx1_ASAP7_75t_R \mod.final_adder.U$1  (.A(\mod.final_adder.con ),
    .Y(\mod.final_adder.$signal$263 ));
 INVx1_ASAP7_75t_R \mod.final_adder.U$11  (.A(\mod.final_adder.sn$142 ),
    .Y(\mod.final_adder.$signal$10 ));
 AO21x1_ASAP7_75t_R \mod.final_adder.U$193  (.A1(\mod.final_adder.$signal$6 ),
    .A2(\mod.final_adder.$signal$263 ),
    .B(\mod.final_adder.$signal$264 ),
    .Y(\mod.final_adder.g_new ));
 INVx1_ASAP7_75t_R \mod.final_adder.U$2  (.A(\mod.final_adder.sn ),
    .Y(\mod.final_adder.$signal ));
 HAxp5_ASAP7_75t_R \mod.final_adder.U$3  (.A(\mod.final_a_registered[1] ),
    .B(net160),
    .CON(\mod.final_adder.con$137 ),
    .SN(\mod.final_adder.sn$138 ));
 AO21x1_ASAP7_75t_R \mod.final_adder.U$344  (.A1(\mod.final_adder.$signal$8 ),
    .A2(\mod.final_adder.g_new ),
    .B(\mod.final_adder.$signal$265 ),
    .Y(\mod.final_adder.g_new$477 ));
 XOR2x1_ASAP7_75t_R \mod.final_adder.U$375  (.A(\mod.final_adder.$signal ),
    .Y(\mod.$54 ),
    .B(net161));
 XOR2x1_ASAP7_75t_R \mod.final_adder.U$376  (.A(\mod.final_adder.$signal$6 ),
    .Y(\mod.$55 ),
    .B(\mod.final_adder.$signal$263 ));
 XOR2x1_ASAP7_75t_R \mod.final_adder.U$377  (.A(\mod.final_adder.$signal$8 ),
    .Y(\mod.$56 ),
    .B(\mod.final_adder.g_new ));
 XOR2x1_ASAP7_75t_R \mod.final_adder.U$378  (.A(\mod.final_adder.$signal$10 ),
    .Y(\mod.$57 ),
    .B(\mod.final_adder.g_new$477 ));
 INVx1_ASAP7_75t_R \mod.final_adder.U$4  (.A(\mod.final_adder.con$137 ),
    .Y(\mod.final_adder.$signal$264 ));
 INVx1_ASAP7_75t_R \mod.final_adder.U$5  (.A(\mod.final_adder.sn$138 ),
    .Y(\mod.final_adder.$signal$6 ));
 HAxp5_ASAP7_75t_R \mod.final_adder.U$6  (.A(\mod.final_a_registered[2] ),
    .B(\mod.final_b_registered[2] ),
    .CON(\mod.final_adder.con$139 ),
    .SN(\mod.final_adder.sn$140 ));
 INVx1_ASAP7_75t_R \mod.final_adder.U$7  (.A(\mod.final_adder.con$139 ),
    .Y(\mod.final_adder.$signal$265 ));
 INVx1_ASAP7_75t_R \mod.final_adder.U$8  (.A(\mod.final_adder.sn$140 ),
    .Y(\mod.final_adder.$signal$8 ));
 HAxp5_ASAP7_75t_R \mod.final_adder.U$9  (.A(\mod.final_a_registered[3] ),
    .B(\mod.final_b_registered[3] ),
    .CON(\mod.final_adder.con$141 ),
    .SN(\mod.final_adder.sn$142 ));
 DFFHQNx1_ASAP7_75t_R \mod.final_b_registered[0]$_DFF_P_  (.CLK(clknet_leaf_30_clock_i),
    .D(\mod.pp_row0_1 ),
    .QN(_13_));
 DFFHQNx1_ASAP7_75t_R \mod.final_b_registered[2]$_DFF_P_  (.CLK(clknet_leaf_28_clock_i),
    .D(\mod.s ),
    .QN(_14_));
 DFFHQNx1_ASAP7_75t_R \mod.final_b_registered[3]$_DFF_P_  (.CLK(clknet_leaf_28_clock_i),
    .D(\mod.s$1260 ),
    .QN(_15_));
 DFFHQNx1_ASAP7_75t_R \mod.o[0]$_DFF_P_  (.CLK(clknet_leaf_28_clock_i),
    .D(\mod.$54 ),
    .QN(_16_));
 DFFHQNx1_ASAP7_75t_R \mod.o[1]$_DFF_P_  (.CLK(clknet_leaf_32_clock_i),
    .D(\mod.$55 ),
    .QN(_17_));
 DFFHQNx1_ASAP7_75t_R \mod.o[2]$_DFF_P_  (.CLK(clknet_leaf_30_clock_i),
    .D(\mod.$56 ),
    .QN(_18_));
 DFFHQNx1_ASAP7_75t_R \mod.o[3]$_DFF_P_  (.CLK(clknet_leaf_28_clock_i),
    .D(\mod.$57 ),
    .QN(_19_));
 DFFHQNx1_ASAP7_75t_R \mod.pp_row0_0$_DFF_P_  (.CLK(clknet_leaf_30_clock_i),
    .D(\mod.booth_b0_m0 ),
    .QN(_20_));
 DFFHQNx1_ASAP7_75t_R \mod.pp_row0_1$_DFF_P_  (.CLK(clknet_leaf_30_clock_i),
    .D(\mod.a_registered[1] ),
    .QN(_21_));
 DFFHQNx1_ASAP7_75t_R \mod.pp_row1_0$_DFF_P_  (.CLK(clknet_leaf_30_clock_i),
    .D(\mod.booth_b0_m1 ),
    .QN(_22_));
 DFFHQNx1_ASAP7_75t_R \mod.pp_row2_0$_DFF_P_  (.CLK(clknet_leaf_30_clock_i),
    .D(\mod.booth_b0_m2 ),
    .QN(_23_));
 DFFHQNx1_ASAP7_75t_R \mod.pp_row2_1$_DFF_P_  (.CLK(clknet_leaf_30_clock_i),
    .D(\mod.booth_b2_m0 ),
    .QN(_24_));
 DFFHQNx1_ASAP7_75t_R \mod.pp_row2_2$_DFF_P_  (.CLK(clknet_leaf_28_clock_i),
    .D(\mod.a_registered[3] ),
    .QN(_25_));
 DFFHQNx1_ASAP7_75t_R \mod.pp_row3_0$_DFF_P_  (.CLK(clknet_leaf_30_clock_i),
    .D(\mod.booth_b0_m3 ),
    .QN(_26_));
 DFFHQNx1_ASAP7_75t_R \mod.pp_row3_1$_DFF_P_  (.CLK(clknet_leaf_29_clock_i),
    .D(\mod.booth_b2_m1 ),
    .QN(_00_));
endmodule
module Multiplier_io_outs_left_mult (clknet_leaf_21_clock_i,
    clknet_leaf_20_clock_i,
    clknet_leaf_13_clock_i,
    clknet_leaf_12_clock_i,
    clknet_leaf_7_clock_i,
    clknet_leaf_5_clock_i,
    io_a,
    io_b,
    io_o);
 input clknet_leaf_21_clock_i;
 input clknet_leaf_20_clock_i;
 input clknet_leaf_13_clock_i;
 input clknet_leaf_12_clock_i;
 input clknet_leaf_7_clock_i;
 input clknet_leaf_5_clock_i;
 input [31:0] io_a;
 input [31:0] io_b;
 output [31:0] io_o;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire \mod.$1 ;
 wire \mod.$2 ;
 wire \mod.$3 ;
 wire \mod.$4 ;
 wire \mod.$5 ;
 wire \mod.$54 ;
 wire \mod.$55 ;
 wire \mod.$56 ;
 wire \mod.$57 ;
 wire \mod.$6 ;
 wire \mod.a_registered[0] ;
 wire \mod.a_registered[1] ;
 wire \mod.a_registered[2] ;
 wire \mod.a_registered[3] ;
 wire \mod.b_registered[0] ;
 wire \mod.b_registered[1] ;
 wire \mod.b_registered[2] ;
 wire \mod.b_registered[3] ;
 wire \mod.booth_b0_m0 ;
 wire \mod.booth_b0_m1 ;
 wire \mod.booth_b0_m2 ;
 wire \mod.booth_b0_m3 ;
 wire \mod.booth_b2_m0 ;
 wire \mod.booth_b2_m1 ;
 wire \mod.c ;
 wire \mod.con$4400 ;
 wire \mod.con$4402 ;
 wire \mod.final_a_registered[0] ;
 wire \mod.final_a_registered[1] ;
 wire \mod.final_a_registered[2] ;
 wire \mod.final_a_registered[3] ;
 wire \mod.final_adder.$signal ;
 wire \mod.final_adder.$signal$10 ;
 wire \mod.final_adder.$signal$263 ;
 wire \mod.final_adder.$signal$264 ;
 wire \mod.final_adder.$signal$265 ;
 wire \mod.final_adder.$signal$6 ;
 wire \mod.final_adder.$signal$8 ;
 wire \mod.final_adder.con ;
 wire \mod.final_adder.con$137 ;
 wire \mod.final_adder.con$139 ;
 wire \mod.final_adder.con$141 ;
 wire \mod.final_adder.g_new ;
 wire \mod.final_adder.g_new$477 ;
 wire \mod.final_adder.sn ;
 wire \mod.final_adder.sn$138 ;
 wire \mod.final_adder.sn$140 ;
 wire \mod.final_adder.sn$142 ;
 wire \mod.final_b_registered[0] ;
 wire \mod.final_b_registered[2] ;
 wire \mod.final_b_registered[3] ;
 wire \mod.pp_row0_0 ;
 wire \mod.pp_row0_1 ;
 wire \mod.pp_row1_0 ;
 wire \mod.pp_row2_0 ;
 wire \mod.pp_row2_1 ;
 wire \mod.pp_row2_2 ;
 wire \mod.pp_row3_0 ;
 wire \mod.pp_row3_1 ;
 wire \mod.s ;
 wire \mod.s$1260 ;
 wire \mod.sel_0 ;
 wire \mod.sel_0$1365 ;
 wire \mod.sel_1 ;
 wire \mod.sel_1$1366 ;
 wire \mod.sn$4401 ;
 wire \mod.sn$4403 ;
 wire \mod.t ;
 wire \mod.t$1976 ;
 wire \mod.t$1977 ;
 wire \mod.t$1978 ;
 wire \mod.t$2009 ;
 wire \mod.t$2010 ;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;

 TIELOx1_ASAP7_75t_R \mod.final_adder.U$375_198  (.L(net195));
 TIELOx1_ASAP7_75t_R \mod.final_adder.U$3_197  (.L(net194));
 TIELOx1_ASAP7_75t_R \mod.U$603_196  (.L(net193));
 TIELOx1_ASAP7_75t_R \mod.U$531_195  (.L(net192));
 TIELOx1_ASAP7_75t_R \mod.U$530_194  (.L(net191));
 TIELOx1_ASAP7_75t_R \mod.U$529_193  (.L(net190));
 TIELOx1_ASAP7_75t_R \mod.U$526_192  (.L(net189));
 TIELOx1_ASAP7_75t_R _83__191 (.L(io_o[31]));
 TIELOx1_ASAP7_75t_R _82__190 (.L(io_o[30]));
 TIELOx1_ASAP7_75t_R _81__189 (.L(io_o[29]));
 TIELOx1_ASAP7_75t_R _80__188 (.L(io_o[28]));
 TIELOx1_ASAP7_75t_R _79__187 (.L(io_o[27]));
 TIELOx1_ASAP7_75t_R _78__186 (.L(io_o[26]));
 TIELOx1_ASAP7_75t_R _77__185 (.L(io_o[25]));
 TIELOx1_ASAP7_75t_R _76__184 (.L(io_o[24]));
 TIELOx1_ASAP7_75t_R _75__183 (.L(io_o[23]));
 TIELOx1_ASAP7_75t_R _74__182 (.L(io_o[22]));
 TIELOx1_ASAP7_75t_R _73__181 (.L(io_o[21]));
 TIELOx1_ASAP7_75t_R _72__180 (.L(io_o[20]));
 TIELOx1_ASAP7_75t_R _71__179 (.L(io_o[19]));
 TIELOx1_ASAP7_75t_R _70__178 (.L(io_o[18]));
 TIELOx1_ASAP7_75t_R _69__177 (.L(io_o[17]));
 TIELOx1_ASAP7_75t_R _68__176 (.L(io_o[16]));
 TIELOx1_ASAP7_75t_R _67__175 (.L(io_o[15]));
 TIELOx1_ASAP7_75t_R _66__174 (.L(io_o[14]));
 TIELOx1_ASAP7_75t_R _65__173 (.L(io_o[13]));
 TIELOx1_ASAP7_75t_R _64__172 (.L(io_o[12]));
 TIELOx1_ASAP7_75t_R _63__171 (.L(io_o[11]));
 TIELOx1_ASAP7_75t_R _62__170 (.L(io_o[10]));
 TIELOx1_ASAP7_75t_R _61__169 (.L(io_o[9]));
 TIELOx1_ASAP7_75t_R _60__168 (.L(io_o[8]));
 TIELOx1_ASAP7_75t_R _59__167 (.L(io_o[7]));
 TIELOx1_ASAP7_75t_R _58__166 (.L(io_o[6]));
 TIELOx1_ASAP7_75t_R _57__165 (.L(io_o[5]));
 TIELOx1_ASAP7_75t_R _56__164 (.L(io_o[4]));
 INVx3_ASAP7_75t_R _28_ (.A(_00_),
    .Y(\mod.pp_row3_1 ));
 INVx3_ASAP7_75t_R _29_ (.A(_01_),
    .Y(\mod.a_registered[0] ));
 INVx3_ASAP7_75t_R _30_ (.A(_02_),
    .Y(\mod.a_registered[1] ));
 INVx3_ASAP7_75t_R _31_ (.A(_03_),
    .Y(\mod.a_registered[2] ));
 INVx3_ASAP7_75t_R _32_ (.A(_04_),
    .Y(\mod.a_registered[3] ));
 INVx3_ASAP7_75t_R _33_ (.A(_05_),
    .Y(\mod.b_registered[0] ));
 INVx3_ASAP7_75t_R _34_ (.A(_06_),
    .Y(\mod.b_registered[1] ));
 INVx3_ASAP7_75t_R _35_ (.A(_07_),
    .Y(\mod.b_registered[2] ));
 INVx3_ASAP7_75t_R _36_ (.A(_08_),
    .Y(\mod.b_registered[3] ));
 INVx3_ASAP7_75t_R _37_ (.A(_09_),
    .Y(\mod.final_a_registered[0] ));
 INVx3_ASAP7_75t_R _38_ (.A(_10_),
    .Y(\mod.final_a_registered[1] ));
 INVx3_ASAP7_75t_R _39_ (.A(_11_),
    .Y(\mod.final_a_registered[2] ));
 INVx3_ASAP7_75t_R _40_ (.A(_12_),
    .Y(\mod.final_a_registered[3] ));
 INVx3_ASAP7_75t_R _41_ (.A(_13_),
    .Y(\mod.final_b_registered[0] ));
 INVx3_ASAP7_75t_R _42_ (.A(_14_),
    .Y(\mod.final_b_registered[2] ));
 INVx3_ASAP7_75t_R _43_ (.A(_15_),
    .Y(\mod.final_b_registered[3] ));
 INVx3_ASAP7_75t_R _44_ (.A(_16_),
    .Y(io_o[0]));
 INVx3_ASAP7_75t_R _45_ (.A(_17_),
    .Y(io_o[1]));
 INVx3_ASAP7_75t_R _46_ (.A(_18_),
    .Y(io_o[2]));
 INVx3_ASAP7_75t_R _47_ (.A(_19_),
    .Y(io_o[3]));
 INVx3_ASAP7_75t_R _48_ (.A(_20_),
    .Y(\mod.pp_row0_0 ));
 INVx3_ASAP7_75t_R _49_ (.A(_21_),
    .Y(\mod.pp_row0_1 ));
 INVx3_ASAP7_75t_R _50_ (.A(_22_),
    .Y(\mod.pp_row1_0 ));
 INVx3_ASAP7_75t_R _51_ (.A(_23_),
    .Y(\mod.pp_row2_0 ));
 INVx3_ASAP7_75t_R _52_ (.A(_24_),
    .Y(\mod.pp_row2_1 ));
 INVx3_ASAP7_75t_R _53_ (.A(_25_),
    .Y(\mod.pp_row2_2 ));
 INVx3_ASAP7_75t_R _54_ (.A(_26_),
    .Y(\mod.pp_row3_0 ));
 INVx1_ASAP7_75t_R \mod.U$2674  (.A(\mod.con$4400 ),
    .Y(\mod.c ));
 INVx1_ASAP7_75t_R \mod.U$2675  (.A(\mod.sn$4401 ),
    .Y(\mod.s ));
 INVx1_ASAP7_75t_R \mod.U$2677  (.A(\mod.sn$4403 ),
    .Y(\mod.s$1260 ));
 INVx1_ASAP7_75t_R \mod.U$526  (.A(net189),
    .Y(\mod.$1 ));
 INVx1_ASAP7_75t_R \mod.U$527  (.A(\mod.a_registered[0] ),
    .Y(\mod.$2 ));
 INVx1_ASAP7_75t_R \mod.U$528  (.A(\mod.a_registered[1] ),
    .Y(\mod.$3 ));
 AO33x2_ASAP7_75t_R \mod.U$529  (.A1(\mod.$3 ),
    .A2(\mod.a_registered[0] ),
    .A3(net190),
    .B1(\mod.a_registered[1] ),
    .B2(\mod.$2 ),
    .B3(\mod.$1 ),
    .Y(\mod.sel_0 ));
 XOR2x1_ASAP7_75t_R \mod.U$530  (.A(\mod.a_registered[0] ),
    .Y(\mod.sel_1 ),
    .B(net191));
 AO22x1_ASAP7_75t_R \mod.U$531  (.A1(net192),
    .A2(\mod.sel_0 ),
    .B1(\mod.b_registered[0] ),
    .B2(\mod.sel_1 ),
    .Y(\mod.t ));
 XOR2x1_ASAP7_75t_R \mod.U$532  (.A(\mod.t ),
    .Y(\mod.booth_b0_m0 ),
    .B(\mod.a_registered[1] ));
 AO22x1_ASAP7_75t_R \mod.U$533  (.A1(\mod.b_registered[0] ),
    .A2(\mod.sel_0 ),
    .B1(\mod.b_registered[1] ),
    .B2(\mod.sel_1 ),
    .Y(\mod.t$1976 ));
 XOR2x1_ASAP7_75t_R \mod.U$534  (.A(\mod.t$1976 ),
    .Y(\mod.booth_b0_m1 ),
    .B(\mod.a_registered[1] ));
 AO22x1_ASAP7_75t_R \mod.U$535  (.A1(\mod.b_registered[1] ),
    .A2(\mod.sel_0 ),
    .B1(\mod.b_registered[2] ),
    .B2(\mod.sel_1 ),
    .Y(\mod.t$1977 ));
 XOR2x1_ASAP7_75t_R \mod.U$536  (.A(\mod.t$1977 ),
    .Y(\mod.booth_b0_m2 ),
    .B(\mod.a_registered[1] ));
 AO22x1_ASAP7_75t_R \mod.U$537  (.A1(\mod.b_registered[2] ),
    .A2(\mod.sel_0 ),
    .B1(\mod.b_registered[3] ),
    .B2(\mod.sel_1 ),
    .Y(\mod.t$1978 ));
 XOR2x1_ASAP7_75t_R \mod.U$538  (.A(\mod.t$1978 ),
    .Y(\mod.booth_b0_m3 ),
    .B(\mod.a_registered[1] ));
 INVx1_ASAP7_75t_R \mod.U$598  (.A(\mod.a_registered[1] ),
    .Y(\mod.$4 ));
 INVx1_ASAP7_75t_R \mod.U$599  (.A(\mod.a_registered[2] ),
    .Y(\mod.$5 ));
 INVx1_ASAP7_75t_R \mod.U$600  (.A(\mod.a_registered[3] ),
    .Y(\mod.$6 ));
 AO33x2_ASAP7_75t_R \mod.U$601  (.A1(\mod.$6 ),
    .A2(\mod.a_registered[2] ),
    .A3(\mod.a_registered[1] ),
    .B1(\mod.a_registered[3] ),
    .B2(\mod.$5 ),
    .B3(\mod.$4 ),
    .Y(\mod.sel_0$1365 ));
 XOR2x1_ASAP7_75t_R \mod.U$602  (.A(\mod.a_registered[2] ),
    .Y(\mod.sel_1$1366 ),
    .B(\mod.a_registered[1] ));
 AO22x1_ASAP7_75t_R \mod.U$603  (.A1(net193),
    .A2(\mod.sel_0$1365 ),
    .B1(\mod.b_registered[0] ),
    .B2(\mod.sel_1$1366 ),
    .Y(\mod.t$2009 ));
 XOR2x1_ASAP7_75t_R \mod.U$604  (.A(\mod.t$2009 ),
    .Y(\mod.booth_b2_m0 ),
    .B(\mod.a_registered[3] ));
 AO22x1_ASAP7_75t_R \mod.U$605  (.A1(\mod.b_registered[0] ),
    .A2(\mod.sel_0$1365 ),
    .B1(\mod.b_registered[1] ),
    .B2(\mod.sel_1$1366 ),
    .Y(\mod.t$2010 ));
 XOR2x1_ASAP7_75t_R \mod.U$606  (.A(\mod.t$2010 ),
    .Y(\mod.booth_b2_m1 ),
    .B(\mod.a_registered[3] ));
 DFFHQNx1_ASAP7_75t_R \mod.a_registered[0]$_DFF_P_  (.CLK(clknet_leaf_13_clock_i),
    .D(io_a[0]),
    .QN(_01_));
 DFFHQNx1_ASAP7_75t_R \mod.a_registered[1]$_DFF_P_  (.CLK(clknet_leaf_13_clock_i),
    .D(io_a[1]),
    .QN(_02_));
 DFFHQNx1_ASAP7_75t_R \mod.a_registered[2]$_DFF_P_  (.CLK(clknet_leaf_12_clock_i),
    .D(io_a[2]),
    .QN(_03_));
 DFFHQNx1_ASAP7_75t_R \mod.a_registered[3]$_DFF_P_  (.CLK(clknet_leaf_12_clock_i),
    .D(io_a[3]),
    .QN(_04_));
 DFFHQNx1_ASAP7_75t_R \mod.b_registered[0]$_DFF_P_  (.CLK(clknet_leaf_12_clock_i),
    .D(io_b[0]),
    .QN(_05_));
 DFFHQNx1_ASAP7_75t_R \mod.b_registered[1]$_DFF_P_  (.CLK(clknet_leaf_12_clock_i),
    .D(io_b[1]),
    .QN(_06_));
 DFFHQNx1_ASAP7_75t_R \mod.b_registered[2]$_DFF_P_  (.CLK(clknet_leaf_12_clock_i),
    .D(io_b[2]),
    .QN(_07_));
 DFFHQNx1_ASAP7_75t_R \mod.b_registered[3]$_DFF_P_  (.CLK(clknet_leaf_12_clock_i),
    .D(io_b[3]),
    .QN(_08_));
 HAxp5_ASAP7_75t_R \mod.dadda_ha_5_2_0  (.A(\mod.pp_row2_0 ),
    .B(\mod.pp_row2_1 ),
    .CON(\mod.con$4400 ),
    .SN(\mod.sn$4401 ));
 HAxp5_ASAP7_75t_R \mod.dadda_ha_5_3_0  (.A(\mod.pp_row3_0 ),
    .B(\mod.pp_row3_1 ),
    .CON(\mod.con$4402 ),
    .SN(\mod.sn$4403 ));
 DFFHQNx1_ASAP7_75t_R \mod.final_a_registered[0]$_DFF_P_  (.CLK(clknet_leaf_20_clock_i),
    .D(\mod.pp_row0_0 ),
    .QN(_09_));
 DFFHQNx1_ASAP7_75t_R \mod.final_a_registered[1]$_DFF_P_  (.CLK(clknet_leaf_20_clock_i),
    .D(\mod.pp_row1_0 ),
    .QN(_10_));
 DFFHQNx1_ASAP7_75t_R \mod.final_a_registered[2]$_DFF_P_  (.CLK(clknet_leaf_12_clock_i),
    .D(\mod.pp_row2_2 ),
    .QN(_11_));
 DFFHQNx1_ASAP7_75t_R \mod.final_a_registered[3]$_DFF_P_  (.CLK(clknet_leaf_20_clock_i),
    .D(\mod.c ),
    .QN(_12_));
 HAxp5_ASAP7_75t_R \mod.final_adder.U$0  (.A(\mod.final_a_registered[0] ),
    .B(\mod.final_b_registered[0] ),
    .CON(\mod.final_adder.con ),
    .SN(\mod.final_adder.sn ));
 INVx1_ASAP7_75t_R \mod.final_adder.U$1  (.A(\mod.final_adder.con ),
    .Y(\mod.final_adder.$signal$263 ));
 INVx1_ASAP7_75t_R \mod.final_adder.U$11  (.A(\mod.final_adder.sn$142 ),
    .Y(\mod.final_adder.$signal$10 ));
 AO21x1_ASAP7_75t_R \mod.final_adder.U$193  (.A1(\mod.final_adder.$signal$6 ),
    .A2(\mod.final_adder.$signal$263 ),
    .B(\mod.final_adder.$signal$264 ),
    .Y(\mod.final_adder.g_new ));
 INVx1_ASAP7_75t_R \mod.final_adder.U$2  (.A(\mod.final_adder.sn ),
    .Y(\mod.final_adder.$signal ));
 HAxp5_ASAP7_75t_R \mod.final_adder.U$3  (.A(\mod.final_a_registered[1] ),
    .B(net194),
    .CON(\mod.final_adder.con$137 ),
    .SN(\mod.final_adder.sn$138 ));
 AO21x1_ASAP7_75t_R \mod.final_adder.U$344  (.A1(\mod.final_adder.$signal$8 ),
    .A2(\mod.final_adder.g_new ),
    .B(\mod.final_adder.$signal$265 ),
    .Y(\mod.final_adder.g_new$477 ));
 XOR2x1_ASAP7_75t_R \mod.final_adder.U$375  (.A(\mod.final_adder.$signal ),
    .Y(\mod.$54 ),
    .B(net195));
 XOR2x1_ASAP7_75t_R \mod.final_adder.U$376  (.A(\mod.final_adder.$signal$6 ),
    .Y(\mod.$55 ),
    .B(\mod.final_adder.$signal$263 ));
 XOR2x1_ASAP7_75t_R \mod.final_adder.U$377  (.A(\mod.final_adder.$signal$8 ),
    .Y(\mod.$56 ),
    .B(\mod.final_adder.g_new ));
 XOR2x1_ASAP7_75t_R \mod.final_adder.U$378  (.A(\mod.final_adder.$signal$10 ),
    .Y(\mod.$57 ),
    .B(\mod.final_adder.g_new$477 ));
 INVx1_ASAP7_75t_R \mod.final_adder.U$4  (.A(\mod.final_adder.con$137 ),
    .Y(\mod.final_adder.$signal$264 ));
 INVx1_ASAP7_75t_R \mod.final_adder.U$5  (.A(\mod.final_adder.sn$138 ),
    .Y(\mod.final_adder.$signal$6 ));
 HAxp5_ASAP7_75t_R \mod.final_adder.U$6  (.A(\mod.final_a_registered[2] ),
    .B(\mod.final_b_registered[2] ),
    .CON(\mod.final_adder.con$139 ),
    .SN(\mod.final_adder.sn$140 ));
 INVx1_ASAP7_75t_R \mod.final_adder.U$7  (.A(\mod.final_adder.con$139 ),
    .Y(\mod.final_adder.$signal$265 ));
 INVx1_ASAP7_75t_R \mod.final_adder.U$8  (.A(\mod.final_adder.sn$140 ),
    .Y(\mod.final_adder.$signal$8 ));
 HAxp5_ASAP7_75t_R \mod.final_adder.U$9  (.A(\mod.final_a_registered[3] ),
    .B(\mod.final_b_registered[3] ),
    .CON(\mod.final_adder.con$141 ),
    .SN(\mod.final_adder.sn$142 ));
 DFFHQNx1_ASAP7_75t_R \mod.final_b_registered[0]$_DFF_P_  (.CLK(clknet_leaf_13_clock_i),
    .D(\mod.pp_row0_1 ),
    .QN(_13_));
 DFFHQNx1_ASAP7_75t_R \mod.final_b_registered[2]$_DFF_P_  (.CLK(clknet_leaf_12_clock_i),
    .D(\mod.s ),
    .QN(_14_));
 DFFHQNx1_ASAP7_75t_R \mod.final_b_registered[3]$_DFF_P_  (.CLK(clknet_leaf_20_clock_i),
    .D(\mod.s$1260 ),
    .QN(_15_));
 DFFHQNx1_ASAP7_75t_R \mod.o[0]$_DFF_P_  (.CLK(clknet_leaf_20_clock_i),
    .D(\mod.$54 ),
    .QN(_16_));
 DFFHQNx1_ASAP7_75t_R \mod.o[1]$_DFF_P_  (.CLK(clknet_leaf_7_clock_i),
    .D(\mod.$55 ),
    .QN(_17_));
 DFFHQNx1_ASAP7_75t_R \mod.o[2]$_DFF_P_  (.CLK(clknet_leaf_5_clock_i),
    .D(\mod.$56 ),
    .QN(_18_));
 DFFHQNx1_ASAP7_75t_R \mod.o[3]$_DFF_P_  (.CLK(clknet_leaf_7_clock_i),
    .D(\mod.$57 ),
    .QN(_19_));
 DFFHQNx1_ASAP7_75t_R \mod.pp_row0_0$_DFF_P_  (.CLK(clknet_leaf_20_clock_i),
    .D(\mod.booth_b0_m0 ),
    .QN(_20_));
 DFFHQNx1_ASAP7_75t_R \mod.pp_row0_1$_DFF_P_  (.CLK(clknet_leaf_13_clock_i),
    .D(\mod.a_registered[1] ),
    .QN(_21_));
 DFFHQNx1_ASAP7_75t_R \mod.pp_row1_0$_DFF_P_  (.CLK(clknet_leaf_13_clock_i),
    .D(\mod.booth_b0_m1 ),
    .QN(_22_));
 DFFHQNx1_ASAP7_75t_R \mod.pp_row2_0$_DFF_P_  (.CLK(clknet_leaf_21_clock_i),
    .D(\mod.booth_b0_m2 ),
    .QN(_23_));
 DFFHQNx1_ASAP7_75t_R \mod.pp_row2_1$_DFF_P_  (.CLK(clknet_leaf_21_clock_i),
    .D(\mod.booth_b2_m0 ),
    .QN(_24_));
 DFFHQNx1_ASAP7_75t_R \mod.pp_row2_2$_DFF_P_  (.CLK(clknet_leaf_12_clock_i),
    .D(\mod.a_registered[3] ),
    .QN(_25_));
 DFFHQNx1_ASAP7_75t_R \mod.pp_row3_0$_DFF_P_  (.CLK(clknet_leaf_20_clock_i),
    .D(\mod.booth_b0_m3 ),
    .QN(_26_));
 DFFHQNx1_ASAP7_75t_R \mod.pp_row3_1$_DFF_P_  (.CLK(clknet_leaf_21_clock_i),
    .D(\mod.booth_b2_m1 ),
    .QN(_00_));
endmodule
module Multiplier_io_outs_right_mult (clknet_leaf_30_clock_i,
    clknet_leaf_29_clock_i,
    clknet_leaf_21_clock_i,
    clknet_leaf_5_clock_i,
    clknet_leaf_4_clock_i,
    clknet_leaf_3_clock_i,
    io_a,
    io_b,
    io_o);
 input clknet_leaf_30_clock_i;
 input clknet_leaf_29_clock_i;
 input clknet_leaf_21_clock_i;
 input clknet_leaf_5_clock_i;
 input clknet_leaf_4_clock_i;
 input clknet_leaf_3_clock_i;
 input [31:0] io_a;
 input [31:0] io_b;
 output [31:0] io_o;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire \mod.$1 ;
 wire \mod.$2 ;
 wire \mod.$3 ;
 wire \mod.$4 ;
 wire \mod.$5 ;
 wire \mod.$54 ;
 wire \mod.$55 ;
 wire \mod.$56 ;
 wire \mod.$57 ;
 wire \mod.$6 ;
 wire \mod.a_registered[0] ;
 wire \mod.a_registered[1] ;
 wire \mod.a_registered[2] ;
 wire \mod.a_registered[3] ;
 wire \mod.b_registered[0] ;
 wire \mod.b_registered[1] ;
 wire \mod.b_registered[2] ;
 wire \mod.b_registered[3] ;
 wire \mod.booth_b0_m0 ;
 wire \mod.booth_b0_m1 ;
 wire \mod.booth_b0_m2 ;
 wire \mod.booth_b0_m3 ;
 wire \mod.booth_b2_m0 ;
 wire \mod.booth_b2_m1 ;
 wire \mod.c ;
 wire \mod.con$4400 ;
 wire \mod.con$4402 ;
 wire \mod.final_a_registered[0] ;
 wire \mod.final_a_registered[1] ;
 wire \mod.final_a_registered[2] ;
 wire \mod.final_a_registered[3] ;
 wire \mod.final_adder.$signal ;
 wire \mod.final_adder.$signal$10 ;
 wire \mod.final_adder.$signal$263 ;
 wire \mod.final_adder.$signal$264 ;
 wire \mod.final_adder.$signal$265 ;
 wire \mod.final_adder.$signal$6 ;
 wire \mod.final_adder.$signal$8 ;
 wire \mod.final_adder.con ;
 wire \mod.final_adder.con$137 ;
 wire \mod.final_adder.con$139 ;
 wire \mod.final_adder.con$141 ;
 wire \mod.final_adder.g_new ;
 wire \mod.final_adder.g_new$477 ;
 wire \mod.final_adder.sn ;
 wire \mod.final_adder.sn$138 ;
 wire \mod.final_adder.sn$140 ;
 wire \mod.final_adder.sn$142 ;
 wire \mod.final_b_registered[0] ;
 wire \mod.final_b_registered[2] ;
 wire \mod.final_b_registered[3] ;
 wire \mod.pp_row0_0 ;
 wire \mod.pp_row0_1 ;
 wire \mod.pp_row1_0 ;
 wire \mod.pp_row2_0 ;
 wire \mod.pp_row2_1 ;
 wire \mod.pp_row2_2 ;
 wire \mod.pp_row3_0 ;
 wire \mod.pp_row3_1 ;
 wire \mod.s ;
 wire \mod.s$1260 ;
 wire \mod.sel_0 ;
 wire \mod.sel_0$1365 ;
 wire \mod.sel_1 ;
 wire \mod.sel_1$1366 ;
 wire \mod.sn$4401 ;
 wire \mod.sn$4403 ;
 wire \mod.t ;
 wire \mod.t$1976 ;
 wire \mod.t$1977 ;
 wire \mod.t$1978 ;
 wire \mod.t$2009 ;
 wire \mod.t$2010 ;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;

 TIELOx1_ASAP7_75t_R \mod.final_adder.U$375_233  (.L(net229));
 TIELOx1_ASAP7_75t_R \mod.final_adder.U$3_232  (.L(net228));
 TIELOx1_ASAP7_75t_R \mod.U$603_231  (.L(net227));
 TIELOx1_ASAP7_75t_R \mod.U$531_230  (.L(net226));
 TIELOx1_ASAP7_75t_R \mod.U$530_229  (.L(net225));
 TIELOx1_ASAP7_75t_R \mod.U$529_228  (.L(net224));
 TIELOx1_ASAP7_75t_R \mod.U$526_227  (.L(net223));
 TIELOx1_ASAP7_75t_R _83__226 (.L(io_o[31]));
 TIELOx1_ASAP7_75t_R _82__225 (.L(io_o[30]));
 TIELOx1_ASAP7_75t_R _81__224 (.L(io_o[29]));
 TIELOx1_ASAP7_75t_R _80__223 (.L(io_o[28]));
 TIELOx1_ASAP7_75t_R _79__222 (.L(io_o[27]));
 TIELOx1_ASAP7_75t_R _78__221 (.L(io_o[26]));
 TIELOx1_ASAP7_75t_R _77__220 (.L(io_o[25]));
 TIELOx1_ASAP7_75t_R _76__219 (.L(io_o[24]));
 TIELOx1_ASAP7_75t_R _75__218 (.L(io_o[23]));
 TIELOx1_ASAP7_75t_R _74__217 (.L(io_o[22]));
 TIELOx1_ASAP7_75t_R _73__216 (.L(io_o[21]));
 TIELOx1_ASAP7_75t_R _72__215 (.L(io_o[20]));
 TIELOx1_ASAP7_75t_R _71__214 (.L(io_o[19]));
 TIELOx1_ASAP7_75t_R _70__213 (.L(io_o[18]));
 TIELOx1_ASAP7_75t_R _69__212 (.L(io_o[17]));
 TIELOx1_ASAP7_75t_R _68__211 (.L(io_o[16]));
 TIELOx1_ASAP7_75t_R _67__210 (.L(io_o[15]));
 TIELOx1_ASAP7_75t_R _66__209 (.L(io_o[14]));
 TIELOx1_ASAP7_75t_R _65__208 (.L(io_o[13]));
 TIELOx1_ASAP7_75t_R _64__207 (.L(io_o[12]));
 TIELOx1_ASAP7_75t_R _63__206 (.L(io_o[11]));
 TIELOx1_ASAP7_75t_R _62__205 (.L(io_o[10]));
 TIELOx1_ASAP7_75t_R _61__204 (.L(io_o[9]));
 TIELOx1_ASAP7_75t_R _60__203 (.L(io_o[8]));
 TIELOx1_ASAP7_75t_R _59__202 (.L(io_o[7]));
 TIELOx1_ASAP7_75t_R _58__201 (.L(io_o[6]));
 TIELOx1_ASAP7_75t_R _57__200 (.L(io_o[5]));
 TIELOx1_ASAP7_75t_R _56__199 (.L(io_o[4]));
 INVx3_ASAP7_75t_R _28_ (.A(_00_),
    .Y(\mod.pp_row3_1 ));
 INVx3_ASAP7_75t_R _29_ (.A(_01_),
    .Y(\mod.a_registered[0] ));
 INVx3_ASAP7_75t_R _30_ (.A(_02_),
    .Y(\mod.a_registered[1] ));
 INVx3_ASAP7_75t_R _31_ (.A(_03_),
    .Y(\mod.a_registered[2] ));
 INVx3_ASAP7_75t_R _32_ (.A(_04_),
    .Y(\mod.a_registered[3] ));
 INVx3_ASAP7_75t_R _33_ (.A(_05_),
    .Y(\mod.b_registered[0] ));
 INVx3_ASAP7_75t_R _34_ (.A(_06_),
    .Y(\mod.b_registered[1] ));
 INVx3_ASAP7_75t_R _35_ (.A(_07_),
    .Y(\mod.b_registered[2] ));
 INVx3_ASAP7_75t_R _36_ (.A(_08_),
    .Y(\mod.b_registered[3] ));
 INVx3_ASAP7_75t_R _37_ (.A(_09_),
    .Y(\mod.final_a_registered[0] ));
 INVx3_ASAP7_75t_R _38_ (.A(_10_),
    .Y(\mod.final_a_registered[1] ));
 INVx3_ASAP7_75t_R _39_ (.A(_11_),
    .Y(\mod.final_a_registered[2] ));
 INVx3_ASAP7_75t_R _40_ (.A(_12_),
    .Y(\mod.final_a_registered[3] ));
 INVx3_ASAP7_75t_R _41_ (.A(_13_),
    .Y(\mod.final_b_registered[0] ));
 INVx3_ASAP7_75t_R _42_ (.A(_14_),
    .Y(\mod.final_b_registered[2] ));
 INVx3_ASAP7_75t_R _43_ (.A(_15_),
    .Y(\mod.final_b_registered[3] ));
 INVx3_ASAP7_75t_R _44_ (.A(_16_),
    .Y(io_o[0]));
 INVx3_ASAP7_75t_R _45_ (.A(_17_),
    .Y(io_o[1]));
 INVx3_ASAP7_75t_R _46_ (.A(_18_),
    .Y(io_o[2]));
 INVx3_ASAP7_75t_R _47_ (.A(_19_),
    .Y(io_o[3]));
 INVx3_ASAP7_75t_R _48_ (.A(_20_),
    .Y(\mod.pp_row0_0 ));
 INVx3_ASAP7_75t_R _49_ (.A(_21_),
    .Y(\mod.pp_row0_1 ));
 INVx3_ASAP7_75t_R _50_ (.A(_22_),
    .Y(\mod.pp_row1_0 ));
 INVx3_ASAP7_75t_R _51_ (.A(_23_),
    .Y(\mod.pp_row2_0 ));
 INVx3_ASAP7_75t_R _52_ (.A(_24_),
    .Y(\mod.pp_row2_1 ));
 INVx3_ASAP7_75t_R _53_ (.A(_25_),
    .Y(\mod.pp_row2_2 ));
 INVx3_ASAP7_75t_R _54_ (.A(_26_),
    .Y(\mod.pp_row3_0 ));
 INVx1_ASAP7_75t_R \mod.U$2674  (.A(\mod.con$4400 ),
    .Y(\mod.c ));
 INVx1_ASAP7_75t_R \mod.U$2675  (.A(\mod.sn$4401 ),
    .Y(\mod.s ));
 INVx1_ASAP7_75t_R \mod.U$2677  (.A(\mod.sn$4403 ),
    .Y(\mod.s$1260 ));
 INVx1_ASAP7_75t_R \mod.U$526  (.A(net223),
    .Y(\mod.$1 ));
 INVx1_ASAP7_75t_R \mod.U$527  (.A(\mod.a_registered[0] ),
    .Y(\mod.$2 ));
 INVx1_ASAP7_75t_R \mod.U$528  (.A(\mod.a_registered[1] ),
    .Y(\mod.$3 ));
 AO33x2_ASAP7_75t_R \mod.U$529  (.A1(\mod.$3 ),
    .A2(\mod.a_registered[0] ),
    .A3(net224),
    .B1(\mod.a_registered[1] ),
    .B2(\mod.$2 ),
    .B3(\mod.$1 ),
    .Y(\mod.sel_0 ));
 XOR2x1_ASAP7_75t_R \mod.U$530  (.A(\mod.a_registered[0] ),
    .Y(\mod.sel_1 ),
    .B(net225));
 AO22x1_ASAP7_75t_R \mod.U$531  (.A1(net226),
    .A2(\mod.sel_0 ),
    .B1(\mod.b_registered[0] ),
    .B2(\mod.sel_1 ),
    .Y(\mod.t ));
 XOR2x1_ASAP7_75t_R \mod.U$532  (.A(\mod.t ),
    .Y(\mod.booth_b0_m0 ),
    .B(\mod.a_registered[1] ));
 AO22x1_ASAP7_75t_R \mod.U$533  (.A1(\mod.b_registered[0] ),
    .A2(\mod.sel_0 ),
    .B1(\mod.b_registered[1] ),
    .B2(\mod.sel_1 ),
    .Y(\mod.t$1976 ));
 XOR2x1_ASAP7_75t_R \mod.U$534  (.A(\mod.t$1976 ),
    .Y(\mod.booth_b0_m1 ),
    .B(\mod.a_registered[1] ));
 AO22x1_ASAP7_75t_R \mod.U$535  (.A1(\mod.b_registered[1] ),
    .A2(\mod.sel_0 ),
    .B1(\mod.b_registered[2] ),
    .B2(\mod.sel_1 ),
    .Y(\mod.t$1977 ));
 XOR2x1_ASAP7_75t_R \mod.U$536  (.A(\mod.t$1977 ),
    .Y(\mod.booth_b0_m2 ),
    .B(\mod.a_registered[1] ));
 AO22x1_ASAP7_75t_R \mod.U$537  (.A1(\mod.b_registered[2] ),
    .A2(\mod.sel_0 ),
    .B1(\mod.b_registered[3] ),
    .B2(\mod.sel_1 ),
    .Y(\mod.t$1978 ));
 XOR2x1_ASAP7_75t_R \mod.U$538  (.A(\mod.t$1978 ),
    .Y(\mod.booth_b0_m3 ),
    .B(\mod.a_registered[1] ));
 INVx1_ASAP7_75t_R \mod.U$598  (.A(\mod.a_registered[1] ),
    .Y(\mod.$4 ));
 INVx1_ASAP7_75t_R \mod.U$599  (.A(\mod.a_registered[2] ),
    .Y(\mod.$5 ));
 INVx1_ASAP7_75t_R \mod.U$600  (.A(\mod.a_registered[3] ),
    .Y(\mod.$6 ));
 AO33x2_ASAP7_75t_R \mod.U$601  (.A1(\mod.$6 ),
    .A2(\mod.a_registered[2] ),
    .A3(\mod.a_registered[1] ),
    .B1(\mod.a_registered[3] ),
    .B2(\mod.$5 ),
    .B3(\mod.$4 ),
    .Y(\mod.sel_0$1365 ));
 XOR2x1_ASAP7_75t_R \mod.U$602  (.A(\mod.a_registered[2] ),
    .Y(\mod.sel_1$1366 ),
    .B(\mod.a_registered[1] ));
 AO22x1_ASAP7_75t_R \mod.U$603  (.A1(net227),
    .A2(\mod.sel_0$1365 ),
    .B1(\mod.b_registered[0] ),
    .B2(\mod.sel_1$1366 ),
    .Y(\mod.t$2009 ));
 XOR2x1_ASAP7_75t_R \mod.U$604  (.A(\mod.t$2009 ),
    .Y(\mod.booth_b2_m0 ),
    .B(\mod.a_registered[3] ));
 AO22x1_ASAP7_75t_R \mod.U$605  (.A1(\mod.b_registered[0] ),
    .A2(\mod.sel_0$1365 ),
    .B1(\mod.b_registered[1] ),
    .B2(\mod.sel_1$1366 ),
    .Y(\mod.t$2010 ));
 XOR2x1_ASAP7_75t_R \mod.U$606  (.A(\mod.t$2010 ),
    .Y(\mod.booth_b2_m1 ),
    .B(\mod.a_registered[3] ));
 DFFHQNx1_ASAP7_75t_R \mod.a_registered[0]$_DFF_P_  (.CLK(clknet_leaf_3_clock_i),
    .D(io_a[0]),
    .QN(_01_));
 DFFHQNx1_ASAP7_75t_R \mod.a_registered[1]$_DFF_P_  (.CLK(clknet_leaf_3_clock_i),
    .D(io_a[1]),
    .QN(_02_));
 DFFHQNx1_ASAP7_75t_R \mod.a_registered[2]$_DFF_P_  (.CLK(clknet_leaf_30_clock_i),
    .D(io_a[2]),
    .QN(_03_));
 DFFHQNx1_ASAP7_75t_R \mod.a_registered[3]$_DFF_P_  (.CLK(clknet_leaf_29_clock_i),
    .D(io_a[3]),
    .QN(_04_));
 DFFHQNx1_ASAP7_75t_R \mod.b_registered[0]$_DFF_P_  (.CLK(clknet_leaf_5_clock_i),
    .D(io_b[0]),
    .QN(_05_));
 DFFHQNx1_ASAP7_75t_R \mod.b_registered[1]$_DFF_P_  (.CLK(clknet_leaf_3_clock_i),
    .D(io_b[1]),
    .QN(_06_));
 DFFHQNx1_ASAP7_75t_R \mod.b_registered[2]$_DFF_P_  (.CLK(clknet_leaf_5_clock_i),
    .D(io_b[2]),
    .QN(_07_));
 DFFHQNx1_ASAP7_75t_R \mod.b_registered[3]$_DFF_P_  (.CLK(clknet_leaf_3_clock_i),
    .D(io_b[3]),
    .QN(_08_));
 HAxp5_ASAP7_75t_R \mod.dadda_ha_5_2_0  (.A(\mod.pp_row2_0 ),
    .B(\mod.pp_row2_1 ),
    .CON(\mod.con$4400 ),
    .SN(\mod.sn$4401 ));
 HAxp5_ASAP7_75t_R \mod.dadda_ha_5_3_0  (.A(\mod.pp_row3_0 ),
    .B(\mod.pp_row3_1 ),
    .CON(\mod.con$4402 ),
    .SN(\mod.sn$4403 ));
 DFFHQNx1_ASAP7_75t_R \mod.final_a_registered[0]$_DFF_P_  (.CLK(clknet_leaf_21_clock_i),
    .D(\mod.pp_row0_0 ),
    .QN(_09_));
 DFFHQNx1_ASAP7_75t_R \mod.final_a_registered[1]$_DFF_P_  (.CLK(clknet_leaf_21_clock_i),
    .D(\mod.pp_row1_0 ),
    .QN(_10_));
 DFFHQNx1_ASAP7_75t_R \mod.final_a_registered[2]$_DFF_P_  (.CLK(clknet_leaf_29_clock_i),
    .D(\mod.pp_row2_2 ),
    .QN(_11_));
 DFFHQNx1_ASAP7_75t_R \mod.final_a_registered[3]$_DFF_P_  (.CLK(clknet_leaf_29_clock_i),
    .D(\mod.c ),
    .QN(_12_));
 HAxp5_ASAP7_75t_R \mod.final_adder.U$0  (.A(\mod.final_a_registered[0] ),
    .B(\mod.final_b_registered[0] ),
    .CON(\mod.final_adder.con ),
    .SN(\mod.final_adder.sn ));
 INVx1_ASAP7_75t_R \mod.final_adder.U$1  (.A(\mod.final_adder.con ),
    .Y(\mod.final_adder.$signal$263 ));
 INVx1_ASAP7_75t_R \mod.final_adder.U$11  (.A(\mod.final_adder.sn$142 ),
    .Y(\mod.final_adder.$signal$10 ));
 AO21x1_ASAP7_75t_R \mod.final_adder.U$193  (.A1(\mod.final_adder.$signal$6 ),
    .A2(\mod.final_adder.$signal$263 ),
    .B(\mod.final_adder.$signal$264 ),
    .Y(\mod.final_adder.g_new ));
 INVx1_ASAP7_75t_R \mod.final_adder.U$2  (.A(\mod.final_adder.sn ),
    .Y(\mod.final_adder.$signal ));
 HAxp5_ASAP7_75t_R \mod.final_adder.U$3  (.A(\mod.final_a_registered[1] ),
    .B(net228),
    .CON(\mod.final_adder.con$137 ),
    .SN(\mod.final_adder.sn$138 ));
 AO21x1_ASAP7_75t_R \mod.final_adder.U$344  (.A1(\mod.final_adder.$signal$8 ),
    .A2(\mod.final_adder.g_new ),
    .B(\mod.final_adder.$signal$265 ),
    .Y(\mod.final_adder.g_new$477 ));
 XOR2x1_ASAP7_75t_R \mod.final_adder.U$375  (.A(\mod.final_adder.$signal ),
    .Y(\mod.$54 ),
    .B(net229));
 XOR2x1_ASAP7_75t_R \mod.final_adder.U$376  (.A(\mod.final_adder.$signal$6 ),
    .Y(\mod.$55 ),
    .B(\mod.final_adder.$signal$263 ));
 XOR2x1_ASAP7_75t_R \mod.final_adder.U$377  (.A(\mod.final_adder.$signal$8 ),
    .Y(\mod.$56 ),
    .B(\mod.final_adder.g_new ));
 XOR2x1_ASAP7_75t_R \mod.final_adder.U$378  (.A(\mod.final_adder.$signal$10 ),
    .Y(\mod.$57 ),
    .B(\mod.final_adder.g_new$477 ));
 INVx1_ASAP7_75t_R \mod.final_adder.U$4  (.A(\mod.final_adder.con$137 ),
    .Y(\mod.final_adder.$signal$264 ));
 INVx1_ASAP7_75t_R \mod.final_adder.U$5  (.A(\mod.final_adder.sn$138 ),
    .Y(\mod.final_adder.$signal$6 ));
 HAxp5_ASAP7_75t_R \mod.final_adder.U$6  (.A(\mod.final_a_registered[2] ),
    .B(\mod.final_b_registered[2] ),
    .CON(\mod.final_adder.con$139 ),
    .SN(\mod.final_adder.sn$140 ));
 INVx1_ASAP7_75t_R \mod.final_adder.U$7  (.A(\mod.final_adder.con$139 ),
    .Y(\mod.final_adder.$signal$265 ));
 INVx1_ASAP7_75t_R \mod.final_adder.U$8  (.A(\mod.final_adder.sn$140 ),
    .Y(\mod.final_adder.$signal$8 ));
 HAxp5_ASAP7_75t_R \mod.final_adder.U$9  (.A(\mod.final_a_registered[3] ),
    .B(\mod.final_b_registered[3] ),
    .CON(\mod.final_adder.con$141 ),
    .SN(\mod.final_adder.sn$142 ));
 DFFHQNx1_ASAP7_75t_R \mod.final_b_registered[0]$_DFF_P_  (.CLK(clknet_leaf_21_clock_i),
    .D(\mod.pp_row0_1 ),
    .QN(_13_));
 DFFHQNx1_ASAP7_75t_R \mod.final_b_registered[2]$_DFF_P_  (.CLK(clknet_leaf_29_clock_i),
    .D(\mod.s ),
    .QN(_14_));
 DFFHQNx1_ASAP7_75t_R \mod.final_b_registered[3]$_DFF_P_  (.CLK(clknet_leaf_29_clock_i),
    .D(\mod.s$1260 ),
    .QN(_15_));
 DFFHQNx1_ASAP7_75t_R \mod.o[0]$_DFF_P_  (.CLK(clknet_leaf_21_clock_i),
    .D(\mod.$54 ),
    .QN(_16_));
 DFFHQNx1_ASAP7_75t_R \mod.o[1]$_DFF_P_  (.CLK(clknet_leaf_21_clock_i),
    .D(\mod.$55 ),
    .QN(_17_));
 DFFHQNx1_ASAP7_75t_R \mod.o[2]$_DFF_P_  (.CLK(clknet_leaf_21_clock_i),
    .D(\mod.$56 ),
    .QN(_18_));
 DFFHQNx1_ASAP7_75t_R \mod.o[3]$_DFF_P_  (.CLK(clknet_leaf_21_clock_i),
    .D(\mod.$57 ),
    .QN(_19_));
 DFFHQNx1_ASAP7_75t_R \mod.pp_row0_0$_DFF_P_  (.CLK(clknet_leaf_4_clock_i),
    .D(\mod.booth_b0_m0 ),
    .QN(_20_));
 DFFHQNx1_ASAP7_75t_R \mod.pp_row0_1$_DFF_P_  (.CLK(clknet_leaf_4_clock_i),
    .D(\mod.a_registered[1] ),
    .QN(_21_));
 DFFHQNx1_ASAP7_75t_R \mod.pp_row1_0$_DFF_P_  (.CLK(clknet_leaf_29_clock_i),
    .D(\mod.booth_b0_m1 ),
    .QN(_22_));
 DFFHQNx1_ASAP7_75t_R \mod.pp_row2_0$_DFF_P_  (.CLK(clknet_leaf_29_clock_i),
    .D(\mod.booth_b0_m2 ),
    .QN(_23_));
 DFFHQNx1_ASAP7_75t_R \mod.pp_row2_1$_DFF_P_  (.CLK(clknet_leaf_29_clock_i),
    .D(\mod.booth_b2_m0 ),
    .QN(_24_));
 DFFHQNx1_ASAP7_75t_R \mod.pp_row2_2$_DFF_P_  (.CLK(clknet_leaf_29_clock_i),
    .D(\mod.a_registered[3] ),
    .QN(_25_));
 DFFHQNx1_ASAP7_75t_R \mod.pp_row3_0$_DFF_P_  (.CLK(clknet_leaf_4_clock_i),
    .D(\mod.booth_b0_m3 ),
    .QN(_26_));
 DFFHQNx1_ASAP7_75t_R \mod.pp_row3_1$_DFF_P_  (.CLK(clknet_leaf_4_clock_i),
    .D(\mod.booth_b2_m1 ),
    .QN(_00_));
endmodule
module Multiplier_io_outs_up_mult (clknet_leaf_14_clock_i,
    clknet_leaf_13_clock_i,
    clknet_leaf_11_clock_i,
    clknet_leaf_9_clock_i,
    clknet_leaf_7_clock_i,
    clknet_leaf_5_clock_i,
    clknet_leaf_4_clock_i,
    clknet_leaf_3_clock_i,
    io_a,
    io_b,
    io_o);
 input clknet_leaf_14_clock_i;
 input clknet_leaf_13_clock_i;
 input clknet_leaf_11_clock_i;
 input clknet_leaf_9_clock_i;
 input clknet_leaf_7_clock_i;
 input clknet_leaf_5_clock_i;
 input clknet_leaf_4_clock_i;
 input clknet_leaf_3_clock_i;
 input [31:0] io_a;
 input [31:0] io_b;
 output [31:0] io_o;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire \mod.$1 ;
 wire \mod.$2 ;
 wire \mod.$3 ;
 wire \mod.$4 ;
 wire \mod.$5 ;
 wire \mod.$54 ;
 wire \mod.$55 ;
 wire \mod.$56 ;
 wire \mod.$57 ;
 wire \mod.$6 ;
 wire \mod.a_registered[0] ;
 wire \mod.a_registered[1] ;
 wire \mod.a_registered[2] ;
 wire \mod.a_registered[3] ;
 wire \mod.b_registered[0] ;
 wire \mod.b_registered[1] ;
 wire \mod.b_registered[2] ;
 wire \mod.b_registered[3] ;
 wire \mod.booth_b0_m0 ;
 wire \mod.booth_b0_m1 ;
 wire \mod.booth_b0_m2 ;
 wire \mod.booth_b0_m3 ;
 wire \mod.booth_b2_m0 ;
 wire \mod.booth_b2_m1 ;
 wire \mod.c ;
 wire \mod.con$4400 ;
 wire \mod.con$4402 ;
 wire \mod.final_a_registered[0] ;
 wire \mod.final_a_registered[1] ;
 wire \mod.final_a_registered[2] ;
 wire \mod.final_a_registered[3] ;
 wire \mod.final_adder.$signal ;
 wire \mod.final_adder.$signal$10 ;
 wire \mod.final_adder.$signal$263 ;
 wire \mod.final_adder.$signal$264 ;
 wire \mod.final_adder.$signal$265 ;
 wire \mod.final_adder.$signal$6 ;
 wire \mod.final_adder.$signal$8 ;
 wire \mod.final_adder.con ;
 wire \mod.final_adder.con$137 ;
 wire \mod.final_adder.con$139 ;
 wire \mod.final_adder.con$141 ;
 wire \mod.final_adder.g_new ;
 wire \mod.final_adder.g_new$477 ;
 wire \mod.final_adder.sn ;
 wire \mod.final_adder.sn$138 ;
 wire \mod.final_adder.sn$140 ;
 wire \mod.final_adder.sn$142 ;
 wire \mod.final_b_registered[0] ;
 wire \mod.final_b_registered[2] ;
 wire \mod.final_b_registered[3] ;
 wire \mod.pp_row0_0 ;
 wire \mod.pp_row0_1 ;
 wire \mod.pp_row1_0 ;
 wire \mod.pp_row2_0 ;
 wire \mod.pp_row2_1 ;
 wire \mod.pp_row2_2 ;
 wire \mod.pp_row3_0 ;
 wire \mod.pp_row3_1 ;
 wire \mod.s ;
 wire \mod.s$1260 ;
 wire \mod.sel_0 ;
 wire \mod.sel_0$1365 ;
 wire \mod.sel_1 ;
 wire \mod.sel_1$1366 ;
 wire \mod.sn$4401 ;
 wire \mod.sn$4403 ;
 wire \mod.t ;
 wire \mod.t$1976 ;
 wire \mod.t$1977 ;
 wire \mod.t$1978 ;
 wire \mod.t$2009 ;
 wire \mod.t$2010 ;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;

 TIELOx1_ASAP7_75t_R \mod.final_adder.U$375_268  (.L(net263));
 TIELOx1_ASAP7_75t_R \mod.final_adder.U$3_267  (.L(net262));
 TIELOx1_ASAP7_75t_R \mod.U$603_266  (.L(net261));
 TIELOx1_ASAP7_75t_R \mod.U$531_265  (.L(net260));
 TIELOx1_ASAP7_75t_R \mod.U$530_264  (.L(net259));
 TIELOx1_ASAP7_75t_R \mod.U$529_263  (.L(net258));
 TIELOx1_ASAP7_75t_R \mod.U$526_262  (.L(net257));
 TIELOx1_ASAP7_75t_R _83__261 (.L(io_o[31]));
 TIELOx1_ASAP7_75t_R _82__260 (.L(io_o[30]));
 TIELOx1_ASAP7_75t_R _81__259 (.L(io_o[29]));
 TIELOx1_ASAP7_75t_R _80__258 (.L(io_o[28]));
 TIELOx1_ASAP7_75t_R _79__257 (.L(io_o[27]));
 TIELOx1_ASAP7_75t_R _78__256 (.L(io_o[26]));
 TIELOx1_ASAP7_75t_R _77__255 (.L(io_o[25]));
 TIELOx1_ASAP7_75t_R _76__254 (.L(io_o[24]));
 TIELOx1_ASAP7_75t_R _75__253 (.L(io_o[23]));
 TIELOx1_ASAP7_75t_R _74__252 (.L(io_o[22]));
 TIELOx1_ASAP7_75t_R _73__251 (.L(io_o[21]));
 TIELOx1_ASAP7_75t_R _72__250 (.L(io_o[20]));
 TIELOx1_ASAP7_75t_R _71__249 (.L(io_o[19]));
 TIELOx1_ASAP7_75t_R _70__248 (.L(io_o[18]));
 TIELOx1_ASAP7_75t_R _69__247 (.L(io_o[17]));
 TIELOx1_ASAP7_75t_R _68__246 (.L(io_o[16]));
 TIELOx1_ASAP7_75t_R _67__245 (.L(io_o[15]));
 TIELOx1_ASAP7_75t_R _66__244 (.L(io_o[14]));
 TIELOx1_ASAP7_75t_R _65__243 (.L(io_o[13]));
 TIELOx1_ASAP7_75t_R _64__242 (.L(io_o[12]));
 TIELOx1_ASAP7_75t_R _63__241 (.L(io_o[11]));
 TIELOx1_ASAP7_75t_R _62__240 (.L(io_o[10]));
 TIELOx1_ASAP7_75t_R _61__239 (.L(io_o[9]));
 TIELOx1_ASAP7_75t_R _60__238 (.L(io_o[8]));
 TIELOx1_ASAP7_75t_R _59__237 (.L(io_o[7]));
 TIELOx1_ASAP7_75t_R _58__236 (.L(io_o[6]));
 TIELOx1_ASAP7_75t_R _57__235 (.L(io_o[5]));
 TIELOx1_ASAP7_75t_R _56__234 (.L(io_o[4]));
 INVx3_ASAP7_75t_R _28_ (.A(_00_),
    .Y(\mod.pp_row3_1 ));
 INVx3_ASAP7_75t_R _29_ (.A(_01_),
    .Y(\mod.a_registered[0] ));
 INVx3_ASAP7_75t_R _30_ (.A(_02_),
    .Y(\mod.a_registered[1] ));
 INVx3_ASAP7_75t_R _31_ (.A(_03_),
    .Y(\mod.a_registered[2] ));
 INVx3_ASAP7_75t_R _32_ (.A(_04_),
    .Y(\mod.a_registered[3] ));
 INVx3_ASAP7_75t_R _33_ (.A(_05_),
    .Y(\mod.b_registered[0] ));
 INVx3_ASAP7_75t_R _34_ (.A(_06_),
    .Y(\mod.b_registered[1] ));
 INVx3_ASAP7_75t_R _35_ (.A(_07_),
    .Y(\mod.b_registered[2] ));
 INVx3_ASAP7_75t_R _36_ (.A(_08_),
    .Y(\mod.b_registered[3] ));
 INVx3_ASAP7_75t_R _37_ (.A(_09_),
    .Y(\mod.final_a_registered[0] ));
 INVx3_ASAP7_75t_R _38_ (.A(_10_),
    .Y(\mod.final_a_registered[1] ));
 INVx3_ASAP7_75t_R _39_ (.A(_11_),
    .Y(\mod.final_a_registered[2] ));
 INVx3_ASAP7_75t_R _40_ (.A(_12_),
    .Y(\mod.final_a_registered[3] ));
 INVx3_ASAP7_75t_R _41_ (.A(_13_),
    .Y(\mod.final_b_registered[0] ));
 INVx3_ASAP7_75t_R _42_ (.A(_14_),
    .Y(\mod.final_b_registered[2] ));
 INVx3_ASAP7_75t_R _43_ (.A(_15_),
    .Y(\mod.final_b_registered[3] ));
 INVx3_ASAP7_75t_R _44_ (.A(_16_),
    .Y(io_o[0]));
 INVx3_ASAP7_75t_R _45_ (.A(_17_),
    .Y(io_o[1]));
 INVx3_ASAP7_75t_R _46_ (.A(_18_),
    .Y(io_o[2]));
 INVx3_ASAP7_75t_R _47_ (.A(_19_),
    .Y(io_o[3]));
 INVx3_ASAP7_75t_R _48_ (.A(_20_),
    .Y(\mod.pp_row0_0 ));
 INVx3_ASAP7_75t_R _49_ (.A(_21_),
    .Y(\mod.pp_row0_1 ));
 INVx3_ASAP7_75t_R _50_ (.A(_22_),
    .Y(\mod.pp_row1_0 ));
 INVx3_ASAP7_75t_R _51_ (.A(_23_),
    .Y(\mod.pp_row2_0 ));
 INVx3_ASAP7_75t_R _52_ (.A(_24_),
    .Y(\mod.pp_row2_1 ));
 INVx3_ASAP7_75t_R _53_ (.A(_25_),
    .Y(\mod.pp_row2_2 ));
 INVx3_ASAP7_75t_R _54_ (.A(_26_),
    .Y(\mod.pp_row3_0 ));
 INVx1_ASAP7_75t_R \mod.U$2674  (.A(\mod.con$4400 ),
    .Y(\mod.c ));
 INVx1_ASAP7_75t_R \mod.U$2675  (.A(\mod.sn$4401 ),
    .Y(\mod.s ));
 INVx1_ASAP7_75t_R \mod.U$2677  (.A(\mod.sn$4403 ),
    .Y(\mod.s$1260 ));
 INVx1_ASAP7_75t_R \mod.U$526  (.A(net257),
    .Y(\mod.$1 ));
 INVx1_ASAP7_75t_R \mod.U$527  (.A(\mod.a_registered[0] ),
    .Y(\mod.$2 ));
 INVx1_ASAP7_75t_R \mod.U$528  (.A(\mod.a_registered[1] ),
    .Y(\mod.$3 ));
 AO33x2_ASAP7_75t_R \mod.U$529  (.A1(\mod.$3 ),
    .A2(\mod.a_registered[0] ),
    .A3(net258),
    .B1(\mod.a_registered[1] ),
    .B2(\mod.$2 ),
    .B3(\mod.$1 ),
    .Y(\mod.sel_0 ));
 XOR2x1_ASAP7_75t_R \mod.U$530  (.A(\mod.a_registered[0] ),
    .Y(\mod.sel_1 ),
    .B(net259));
 AO22x1_ASAP7_75t_R \mod.U$531  (.A1(net260),
    .A2(\mod.sel_0 ),
    .B1(\mod.b_registered[0] ),
    .B2(\mod.sel_1 ),
    .Y(\mod.t ));
 XOR2x1_ASAP7_75t_R \mod.U$532  (.A(\mod.t ),
    .Y(\mod.booth_b0_m0 ),
    .B(\mod.a_registered[1] ));
 AO22x1_ASAP7_75t_R \mod.U$533  (.A1(\mod.b_registered[0] ),
    .A2(\mod.sel_0 ),
    .B1(\mod.b_registered[1] ),
    .B2(\mod.sel_1 ),
    .Y(\mod.t$1976 ));
 XOR2x1_ASAP7_75t_R \mod.U$534  (.A(\mod.t$1976 ),
    .Y(\mod.booth_b0_m1 ),
    .B(\mod.a_registered[1] ));
 AO22x1_ASAP7_75t_R \mod.U$535  (.A1(\mod.b_registered[1] ),
    .A2(\mod.sel_0 ),
    .B1(\mod.b_registered[2] ),
    .B2(\mod.sel_1 ),
    .Y(\mod.t$1977 ));
 XOR2x1_ASAP7_75t_R \mod.U$536  (.A(\mod.t$1977 ),
    .Y(\mod.booth_b0_m2 ),
    .B(\mod.a_registered[1] ));
 AO22x1_ASAP7_75t_R \mod.U$537  (.A1(\mod.b_registered[2] ),
    .A2(\mod.sel_0 ),
    .B1(\mod.b_registered[3] ),
    .B2(\mod.sel_1 ),
    .Y(\mod.t$1978 ));
 XOR2x1_ASAP7_75t_R \mod.U$538  (.A(\mod.t$1978 ),
    .Y(\mod.booth_b0_m3 ),
    .B(\mod.a_registered[1] ));
 INVx1_ASAP7_75t_R \mod.U$598  (.A(\mod.a_registered[1] ),
    .Y(\mod.$4 ));
 INVx1_ASAP7_75t_R \mod.U$599  (.A(\mod.a_registered[2] ),
    .Y(\mod.$5 ));
 INVx1_ASAP7_75t_R \mod.U$600  (.A(\mod.a_registered[3] ),
    .Y(\mod.$6 ));
 AO33x2_ASAP7_75t_R \mod.U$601  (.A1(\mod.$6 ),
    .A2(\mod.a_registered[2] ),
    .A3(\mod.a_registered[1] ),
    .B1(\mod.a_registered[3] ),
    .B2(\mod.$5 ),
    .B3(\mod.$4 ),
    .Y(\mod.sel_0$1365 ));
 XOR2x1_ASAP7_75t_R \mod.U$602  (.A(\mod.a_registered[2] ),
    .Y(\mod.sel_1$1366 ),
    .B(\mod.a_registered[1] ));
 AO22x1_ASAP7_75t_R \mod.U$603  (.A1(net261),
    .A2(\mod.sel_0$1365 ),
    .B1(\mod.b_registered[0] ),
    .B2(\mod.sel_1$1366 ),
    .Y(\mod.t$2009 ));
 XOR2x1_ASAP7_75t_R \mod.U$604  (.A(\mod.t$2009 ),
    .Y(\mod.booth_b2_m0 ),
    .B(\mod.a_registered[3] ));
 AO22x1_ASAP7_75t_R \mod.U$605  (.A1(\mod.b_registered[0] ),
    .A2(\mod.sel_0$1365 ),
    .B1(\mod.b_registered[1] ),
    .B2(\mod.sel_1$1366 ),
    .Y(\mod.t$2010 ));
 XOR2x1_ASAP7_75t_R \mod.U$606  (.A(\mod.t$2010 ),
    .Y(\mod.booth_b2_m1 ),
    .B(\mod.a_registered[3] ));
 DFFHQNx1_ASAP7_75t_R \mod.a_registered[0]$_DFF_P_  (.CLK(clknet_leaf_5_clock_i),
    .D(io_a[0]),
    .QN(_01_));
 DFFHQNx1_ASAP7_75t_R \mod.a_registered[1]$_DFF_P_  (.CLK(clknet_leaf_3_clock_i),
    .D(io_a[1]),
    .QN(_02_));
 DFFHQNx1_ASAP7_75t_R \mod.a_registered[2]$_DFF_P_  (.CLK(clknet_leaf_5_clock_i),
    .D(io_a[2]),
    .QN(_03_));
 DFFHQNx1_ASAP7_75t_R \mod.a_registered[3]$_DFF_P_  (.CLK(clknet_leaf_5_clock_i),
    .D(io_a[3]),
    .QN(_04_));
 DFFHQNx1_ASAP7_75t_R \mod.b_registered[0]$_DFF_P_  (.CLK(clknet_leaf_13_clock_i),
    .D(io_b[0]),
    .QN(_05_));
 DFFHQNx1_ASAP7_75t_R \mod.b_registered[1]$_DFF_P_  (.CLK(clknet_leaf_7_clock_i),
    .D(io_b[1]),
    .QN(_06_));
 DFFHQNx1_ASAP7_75t_R \mod.b_registered[2]$_DFF_P_  (.CLK(clknet_leaf_5_clock_i),
    .D(io_b[2]),
    .QN(_07_));
 DFFHQNx1_ASAP7_75t_R \mod.b_registered[3]$_DFF_P_  (.CLK(clknet_leaf_11_clock_i),
    .D(io_b[3]),
    .QN(_08_));
 HAxp5_ASAP7_75t_R \mod.dadda_ha_5_2_0  (.A(\mod.pp_row2_0 ),
    .B(\mod.pp_row2_1 ),
    .CON(\mod.con$4400 ),
    .SN(\mod.sn$4401 ));
 HAxp5_ASAP7_75t_R \mod.dadda_ha_5_3_0  (.A(\mod.pp_row3_0 ),
    .B(\mod.pp_row3_1 ),
    .CON(\mod.con$4402 ),
    .SN(\mod.sn$4403 ));
 DFFHQNx1_ASAP7_75t_R \mod.final_a_registered[0]$_DFF_P_  (.CLK(clknet_leaf_11_clock_i),
    .D(\mod.pp_row0_0 ),
    .QN(_09_));
 DFFHQNx1_ASAP7_75t_R \mod.final_a_registered[1]$_DFF_P_  (.CLK(clknet_leaf_11_clock_i),
    .D(\mod.pp_row1_0 ),
    .QN(_10_));
 DFFHQNx1_ASAP7_75t_R \mod.final_a_registered[2]$_DFF_P_  (.CLK(clknet_leaf_4_clock_i),
    .D(\mod.pp_row2_2 ),
    .QN(_11_));
 DFFHQNx1_ASAP7_75t_R \mod.final_a_registered[3]$_DFF_P_  (.CLK(clknet_leaf_11_clock_i),
    .D(\mod.c ),
    .QN(_12_));
 HAxp5_ASAP7_75t_R \mod.final_adder.U$0  (.A(\mod.final_a_registered[0] ),
    .B(\mod.final_b_registered[0] ),
    .CON(\mod.final_adder.con ),
    .SN(\mod.final_adder.sn ));
 INVx1_ASAP7_75t_R \mod.final_adder.U$1  (.A(\mod.final_adder.con ),
    .Y(\mod.final_adder.$signal$263 ));
 INVx1_ASAP7_75t_R \mod.final_adder.U$11  (.A(\mod.final_adder.sn$142 ),
    .Y(\mod.final_adder.$signal$10 ));
 AO21x1_ASAP7_75t_R \mod.final_adder.U$193  (.A1(\mod.final_adder.$signal$6 ),
    .A2(\mod.final_adder.$signal$263 ),
    .B(\mod.final_adder.$signal$264 ),
    .Y(\mod.final_adder.g_new ));
 INVx1_ASAP7_75t_R \mod.final_adder.U$2  (.A(\mod.final_adder.sn ),
    .Y(\mod.final_adder.$signal ));
 HAxp5_ASAP7_75t_R \mod.final_adder.U$3  (.A(\mod.final_a_registered[1] ),
    .B(net262),
    .CON(\mod.final_adder.con$137 ),
    .SN(\mod.final_adder.sn$138 ));
 AO21x1_ASAP7_75t_R \mod.final_adder.U$344  (.A1(\mod.final_adder.$signal$8 ),
    .A2(\mod.final_adder.g_new ),
    .B(\mod.final_adder.$signal$265 ),
    .Y(\mod.final_adder.g_new$477 ));
 XOR2x1_ASAP7_75t_R \mod.final_adder.U$375  (.A(\mod.final_adder.$signal ),
    .Y(\mod.$54 ),
    .B(net263));
 XOR2x1_ASAP7_75t_R \mod.final_adder.U$376  (.A(\mod.final_adder.$signal$6 ),
    .Y(\mod.$55 ),
    .B(\mod.final_adder.$signal$263 ));
 XOR2x1_ASAP7_75t_R \mod.final_adder.U$377  (.A(\mod.final_adder.$signal$8 ),
    .Y(\mod.$56 ),
    .B(\mod.final_adder.g_new ));
 XOR2x1_ASAP7_75t_R \mod.final_adder.U$378  (.A(\mod.final_adder.$signal$10 ),
    .Y(\mod.$57 ),
    .B(\mod.final_adder.g_new$477 ));
 INVx1_ASAP7_75t_R \mod.final_adder.U$4  (.A(\mod.final_adder.con$137 ),
    .Y(\mod.final_adder.$signal$264 ));
 INVx1_ASAP7_75t_R \mod.final_adder.U$5  (.A(\mod.final_adder.sn$138 ),
    .Y(\mod.final_adder.$signal$6 ));
 HAxp5_ASAP7_75t_R \mod.final_adder.U$6  (.A(\mod.final_a_registered[2] ),
    .B(\mod.final_b_registered[2] ),
    .CON(\mod.final_adder.con$139 ),
    .SN(\mod.final_adder.sn$140 ));
 INVx1_ASAP7_75t_R \mod.final_adder.U$7  (.A(\mod.final_adder.con$139 ),
    .Y(\mod.final_adder.$signal$265 ));
 INVx1_ASAP7_75t_R \mod.final_adder.U$8  (.A(\mod.final_adder.sn$140 ),
    .Y(\mod.final_adder.$signal$8 ));
 HAxp5_ASAP7_75t_R \mod.final_adder.U$9  (.A(\mod.final_a_registered[3] ),
    .B(\mod.final_b_registered[3] ),
    .CON(\mod.final_adder.con$141 ),
    .SN(\mod.final_adder.sn$142 ));
 DFFHQNx1_ASAP7_75t_R \mod.final_b_registered[0]$_DFF_P_  (.CLK(clknet_leaf_9_clock_i),
    .D(\mod.pp_row0_1 ),
    .QN(_13_));
 DFFHQNx1_ASAP7_75t_R \mod.final_b_registered[2]$_DFF_P_  (.CLK(clknet_leaf_11_clock_i),
    .D(\mod.s ),
    .QN(_14_));
 DFFHQNx1_ASAP7_75t_R \mod.final_b_registered[3]$_DFF_P_  (.CLK(clknet_leaf_11_clock_i),
    .D(\mod.s$1260 ),
    .QN(_15_));
 DFFHQNx1_ASAP7_75t_R \mod.o[0]$_DFF_P_  (.CLK(clknet_leaf_14_clock_i),
    .D(\mod.$54 ),
    .QN(_16_));
 DFFHQNx1_ASAP7_75t_R \mod.o[1]$_DFF_P_  (.CLK(clknet_leaf_7_clock_i),
    .D(\mod.$55 ),
    .QN(_17_));
 DFFHQNx1_ASAP7_75t_R \mod.o[2]$_DFF_P_  (.CLK(clknet_leaf_14_clock_i),
    .D(\mod.$56 ),
    .QN(_18_));
 DFFHQNx1_ASAP7_75t_R \mod.o[3]$_DFF_P_  (.CLK(clknet_leaf_13_clock_i),
    .D(\mod.$57 ),
    .QN(_19_));
 DFFHQNx1_ASAP7_75t_R \mod.pp_row0_0$_DFF_P_  (.CLK(clknet_leaf_9_clock_i),
    .D(\mod.booth_b0_m0 ),
    .QN(_20_));
 DFFHQNx1_ASAP7_75t_R \mod.pp_row0_1$_DFF_P_  (.CLK(clknet_leaf_9_clock_i),
    .D(\mod.a_registered[1] ),
    .QN(_21_));
 DFFHQNx1_ASAP7_75t_R \mod.pp_row1_0$_DFF_P_  (.CLK(clknet_leaf_11_clock_i),
    .D(\mod.booth_b0_m1 ),
    .QN(_22_));
 DFFHQNx1_ASAP7_75t_R \mod.pp_row2_0$_DFF_P_  (.CLK(clknet_leaf_11_clock_i),
    .D(\mod.booth_b0_m2 ),
    .QN(_23_));
 DFFHQNx1_ASAP7_75t_R \mod.pp_row2_1$_DFF_P_  (.CLK(clknet_leaf_4_clock_i),
    .D(\mod.booth_b2_m0 ),
    .QN(_24_));
 DFFHQNx1_ASAP7_75t_R \mod.pp_row2_2$_DFF_P_  (.CLK(clknet_leaf_4_clock_i),
    .D(\mod.a_registered[3] ),
    .QN(_25_));
 DFFHQNx1_ASAP7_75t_R \mod.pp_row3_0$_DFF_P_  (.CLK(clknet_leaf_4_clock_i),
    .D(\mod.booth_b0_m3 ),
    .QN(_26_));
 DFFHQNx1_ASAP7_75t_R \mod.pp_row3_1$_DFF_P_  (.CLK(clknet_leaf_4_clock_i),
    .D(\mod.booth_b2_m1 ),
    .QN(_00_));
endmodule
