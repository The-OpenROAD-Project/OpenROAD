# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS

MACRO sky130_fd_sc_hs__a2111o_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.440000 0.840000 0.670000 ;
        RECT 0.510000 0.255000 0.840000 0.440000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.050000 1.500000 2.275000 1.800000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435000 0.255000 1.795000 0.490000 ;
        RECT 1.595000 0.490000 1.795000 0.670000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.005000 0.255000 2.335000 0.490000 ;
        RECT 2.005000 0.490000 2.245000 0.670000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 1.500000 2.775000 1.800000 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.504100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.860000 0.370000 4.195000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.360000  1.940000 0.690000 1.970000 ;
      RECT 0.360000  1.970000 1.630000 2.140000 ;
      RECT 0.360000  2.140000 0.690000 2.980000 ;
      RECT 0.385000  0.840000 0.715000 1.160000 ;
      RECT 0.385000  1.160000 3.115000 1.320000 ;
      RECT 0.385000  1.320000 3.690000 1.330000 ;
      RECT 0.385000  1.330000 0.715000 1.340000 ;
      RECT 0.890000  2.310000 1.100000 3.245000 ;
      RECT 1.095000  0.085000 1.265000 0.660000 ;
      RECT 1.095000  0.660000 1.425000 0.990000 ;
      RECT 1.300000  2.140000 1.630000 2.980000 ;
      RECT 1.715000  0.840000 2.045000 1.160000 ;
      RECT 2.415000  0.660000 2.675000 0.990000 ;
      RECT 2.505000  0.085000 2.675000 0.660000 ;
      RECT 2.530000  1.970000 3.115000 2.140000 ;
      RECT 2.530000  2.140000 2.860000 2.980000 ;
      RECT 2.845000  0.660000 3.115000 1.160000 ;
      RECT 2.945000  1.330000 3.690000 1.650000 ;
      RECT 2.945000  1.650000 3.115000 1.970000 ;
      RECT 3.410000  1.820000 3.660000 3.245000 ;
      RECT 3.435000  0.085000 3.685000 1.150000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__a2111o_1


MACRO sky130_fd_sc_hs__a2111o_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.365000 1.350000 4.695000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.350000 4.195000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.985000 1.350000 3.315000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 1.350000 2.775000 2.890000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.350000 2.275000 1.780000 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.550000 0.860000 2.980000 ;
        RECT 0.690000 0.350000 0.860000 1.550000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.155000  1.820000 0.405000 3.245000 ;
      RECT 0.180000  0.085000 0.510000 1.130000 ;
      RECT 1.030000  1.220000 1.360000 1.550000 ;
      RECT 1.040000  0.085000 1.370000 0.840000 ;
      RECT 1.055000  2.290000 1.385000 3.245000 ;
      RECT 1.190000  1.010000 4.520000 1.180000 ;
      RECT 1.190000  1.180000 1.360000 1.220000 ;
      RECT 1.190000  1.550000 1.360000 1.950000 ;
      RECT 1.190000  1.950000 2.085000 2.120000 ;
      RECT 1.755000  2.120000 2.085000 2.980000 ;
      RECT 1.780000  0.350000 2.030000 1.010000 ;
      RECT 2.210000  0.085000 2.580000 0.840000 ;
      RECT 2.760000  0.350000 3.010000 1.010000 ;
      RECT 3.135000  1.950000 4.545000 2.120000 ;
      RECT 3.135000  2.120000 3.505000 2.980000 ;
      RECT 3.180000  0.085000 3.730000 0.840000 ;
      RECT 3.675000  2.290000 4.045000 3.245000 ;
      RECT 4.190000  0.350000 4.520000 1.010000 ;
      RECT 4.215000  2.120000 4.545000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_hs__a2111o_2
MACRO sky130_fd_sc_hs__a2111o_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.285000 1.450000 7.075000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.245000 1.260000 8.035000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.405000 1.450000 6.115000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.450000 5.155000 1.780000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.385000 1.260000 3.715000 1.780000 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.960000 2.445000 1.130000 ;
        RECT 0.125000 1.130000 0.650000 1.800000 ;
        RECT 0.125000 1.800000 2.065000 1.970000 ;
        RECT 0.835000 1.970000 1.165000 2.980000 ;
        RECT 1.415000 0.350000 1.665000 0.960000 ;
        RECT 1.735000 1.970000 2.065000 2.980000 ;
        RECT 2.195000 0.350000 2.445000 0.960000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.385000  2.140000 0.635000 3.245000 ;
      RECT 0.870000  1.300000 3.215000 1.630000 ;
      RECT 0.905000  0.085000 1.235000 0.790000 ;
      RECT 1.365000  2.140000 1.535000 3.245000 ;
      RECT 1.845000  0.085000 2.015000 0.790000 ;
      RECT 2.265000  1.820000 2.515000 3.245000 ;
      RECT 2.625000  0.085000 2.875000 1.030000 ;
      RECT 2.705000  2.290000 3.035000 2.905000 ;
      RECT 2.705000  2.905000 4.835000 3.075000 ;
      RECT 3.045000  0.350000 3.350000 0.920000 ;
      RECT 3.045000  0.920000 4.220000 1.090000 ;
      RECT 3.045000  1.090000 3.215000 1.300000 ;
      RECT 3.045000  1.630000 3.215000 1.950000 ;
      RECT 3.045000  1.950000 3.405000 2.120000 ;
      RECT 3.235000  2.120000 3.405000 2.735000 ;
      RECT 3.530000  0.085000 3.870000 0.750000 ;
      RECT 3.605000  1.950000 3.935000 2.905000 ;
      RECT 4.050000  0.350000 4.220000 0.920000 ;
      RECT 4.050000  1.090000 4.220000 1.110000 ;
      RECT 4.050000  1.110000 6.770000 1.280000 ;
      RECT 4.135000  1.950000 5.805000 2.120000 ;
      RECT 4.135000  2.120000 4.305000 2.735000 ;
      RECT 4.400000  0.085000 4.740000 0.940000 ;
      RECT 4.505000  2.290000 4.835000 2.905000 ;
      RECT 4.920000  0.350000 5.090000 1.110000 ;
      RECT 5.025000  2.290000 5.305000 2.905000 ;
      RECT 5.025000  2.905000 6.175000 3.075000 ;
      RECT 5.270000  0.085000 5.600000 0.940000 ;
      RECT 5.475000  2.120000 5.805000 2.735000 ;
      RECT 6.005000  1.950000 8.055000 2.120000 ;
      RECT 6.005000  2.120000 6.175000 2.905000 ;
      RECT 6.010000  0.285000 7.120000 0.455000 ;
      RECT 6.010000  0.455000 6.340000 0.940000 ;
      RECT 6.375000  2.290000 6.705000 3.245000 ;
      RECT 6.510000  0.625000 6.770000 1.110000 ;
      RECT 6.905000  2.120000 7.075000 2.980000 ;
      RECT 6.950000  0.455000 7.120000 0.920000 ;
      RECT 6.950000  0.920000 8.060000 1.090000 ;
      RECT 7.275000  2.290000 7.525000 3.245000 ;
      RECT 7.300000  0.085000 7.630000 0.750000 ;
      RECT 7.725000  2.120000 8.055000 2.980000 ;
      RECT 7.810000  0.350000 8.060000 0.920000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_hs__a2111o_4
MACRO sky130_fd_sc_hs__a2111oi_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.350000 2.415000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.625000 1.180000 3.235000 1.550000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.545000 1.350000 1.875000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.350000 1.335000 1.780000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.465000 1.350000 0.835000 1.780000 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  0.722400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.010000 2.180000 1.180000 ;
        RECT 0.125000 1.180000 0.295000 1.950000 ;
        RECT 0.125000 1.950000 1.315000 2.980000 ;
        RECT 0.850000 0.350000 1.100000 1.010000 ;
        RECT 1.850000 0.350000 2.180000 1.010000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.340000  0.085000 0.670000 0.840000 ;
      RECT 1.270000  0.085000 1.680000 0.840000 ;
      RECT 1.695000  1.950000 3.105000 2.120000 ;
      RECT 1.695000  2.120000 2.065000 2.980000 ;
      RECT 2.235000  2.290000 2.605000 3.245000 ;
      RECT 2.750000  0.085000 3.080000 1.010000 ;
      RECT 2.775000  1.820000 3.105000 1.950000 ;
      RECT 2.775000  2.120000 3.105000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__a2111oi_1
MACRO sky130_fd_sc_hs__a2111oi_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.350000 4.675000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.850000 1.350000 5.180000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.180000 3.715000 1.550000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505000 1.350000 2.755000 1.780000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.350000 1.315000 1.780000 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  1.027900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.010000 2.500000 1.180000 ;
        RECT 0.125000 1.180000 0.355000 1.950000 ;
        RECT 0.125000 1.950000 1.085000 2.120000 ;
        RECT 0.755000 2.120000 1.085000 2.735000 ;
        RECT 1.160000 0.350000 1.490000 1.010000 ;
        RECT 2.170000 0.350000 2.500000 0.770000 ;
        RECT 2.170000 0.770000 4.330000 0.975000 ;
        RECT 2.170000 0.975000 2.500000 1.010000 ;
        RECT 4.000000 0.975000 4.330000 1.130000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.305000  2.290000 0.555000 2.905000 ;
      RECT 0.305000  2.905000 2.435000 3.075000 ;
      RECT 0.660000  0.085000 0.990000 0.840000 ;
      RECT 1.285000  1.950000 1.455000 2.905000 ;
      RECT 1.655000  1.950000 3.325000 2.120000 ;
      RECT 1.655000  2.120000 1.985000 2.735000 ;
      RECT 1.660000  0.085000 2.000000 0.840000 ;
      RECT 2.185000  2.290000 2.435000 2.905000 ;
      RECT 2.625000  2.290000 2.905000 2.905000 ;
      RECT 2.625000  2.905000 3.855000 3.075000 ;
      RECT 3.075000  1.820000 3.325000 1.950000 ;
      RECT 3.075000  2.120000 3.325000 2.735000 ;
      RECT 3.525000  1.950000 5.655000 2.120000 ;
      RECT 3.525000  2.120000 3.855000 2.905000 ;
      RECT 3.570000  0.350000 4.680000 0.600000 ;
      RECT 4.055000  2.290000 4.225000 3.245000 ;
      RECT 4.425000  2.120000 4.675000 2.980000 ;
      RECT 4.510000  0.600000 4.680000 1.010000 ;
      RECT 4.510000  1.010000 5.630000 1.180000 ;
      RECT 4.860000  0.085000 5.200000 0.840000 ;
      RECT 4.875000  2.290000 5.205000 3.245000 ;
      RECT 5.380000  0.350000 5.630000 1.010000 ;
      RECT 5.405000  1.820000 5.655000 1.950000 ;
      RECT 5.405000  2.120000 5.655000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_hs__a2111oi_2
MACRO sky130_fd_sc_hs__a2111oi_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.450000 1.350000 8.035000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.205000 1.350000 9.555000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.275000 1.350000 6.075000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.235000 1.350000 3.510000 1.780000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.555000 1.180000 1.905000 1.550000 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  1.708000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.840000 2.640000 1.010000 ;
        RECT 0.125000 1.010000 0.355000 1.720000 ;
        RECT 0.125000 1.720000 1.705000 1.890000 ;
        RECT 0.555000 1.890000 0.885000 2.735000 ;
        RECT 1.455000 1.890000 1.705000 2.735000 ;
        RECT 1.530000 0.330000 1.700000 0.840000 ;
        RECT 2.390000 0.350000 2.640000 0.840000 ;
        RECT 2.390000 1.010000 7.740000 1.130000 ;
        RECT 2.390000 1.130000 6.880000 1.180000 ;
        RECT 4.070000 0.350000 4.320000 0.975000 ;
        RECT 4.070000 0.975000 7.740000 1.010000 ;
        RECT 6.550000 0.770000 6.880000 0.915000 ;
        RECT 6.550000 0.915000 7.740000 0.975000 ;
        RECT 7.410000 0.770000 7.740000 0.915000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.105000  2.060000  0.355000 2.905000 ;
      RECT 0.105000  2.905000  2.235000 3.075000 ;
      RECT 1.020000  0.085000  1.350000 0.670000 ;
      RECT 1.085000  2.060000  1.255000 2.905000 ;
      RECT 1.880000  0.085000  2.210000 0.670000 ;
      RECT 1.905000  1.950000  4.035000 2.120000 ;
      RECT 1.905000  2.120000  2.235000 2.905000 ;
      RECT 2.435000  2.290000  2.685000 2.905000 ;
      RECT 2.435000  2.905000  5.925000 3.075000 ;
      RECT 2.810000  0.085000  3.900000 0.840000 ;
      RECT 2.855000  2.120000  3.085000 2.735000 ;
      RECT 3.255000  2.290000  3.585000 2.905000 ;
      RECT 3.705000  1.820000  4.035000 1.950000 ;
      RECT 3.755000  2.120000  4.035000 2.735000 ;
      RECT 4.245000  1.950000  9.975000 2.120000 ;
      RECT 4.245000  2.120000  4.525000 2.735000 ;
      RECT 4.500000  0.085000  4.830000 0.805000 ;
      RECT 4.695000  2.290000  5.025000 2.905000 ;
      RECT 5.195000  2.120000  5.425000 2.735000 ;
      RECT 5.595000  2.290000  5.925000 2.905000 ;
      RECT 6.120000  0.350000  8.090000 0.600000 ;
      RECT 6.120000  0.600000  6.380000 0.680000 ;
      RECT 6.125000  2.120000  6.295000 2.980000 ;
      RECT 6.495000  2.290000  6.825000 3.245000 ;
      RECT 7.025000  2.120000  7.195000 2.980000 ;
      RECT 7.040000  0.600000  7.250000 0.680000 ;
      RECT 7.395000  2.290000  7.725000 3.245000 ;
      RECT 7.920000  0.600000  8.090000 1.010000 ;
      RECT 7.920000  1.010000  9.890000 1.180000 ;
      RECT 7.925000  2.120000  8.095000 2.980000 ;
      RECT 8.270000  0.085000  8.600000 0.840000 ;
      RECT 8.295000  2.290000  8.545000 3.245000 ;
      RECT 8.745000  2.120000  9.075000 2.980000 ;
      RECT 8.780000  0.350000  8.950000 1.010000 ;
      RECT 9.130000  0.085000  9.460000 0.840000 ;
      RECT 9.275000  2.290000  9.525000 3.245000 ;
      RECT 9.640000  0.350000  9.890000 1.010000 ;
      RECT 9.725000  1.820000  9.975000 1.950000 ;
      RECT 9.725000  2.120000  9.975000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
  END
END sky130_fd_sc_hs__a2111oi_4
MACRO sky130_fd_sc_hs__a211o_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.450000 2.755000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.585000 1.450000 1.835000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 0.255000 2.875000 0.570000 ;
        RECT 2.045000 0.570000 2.275000 0.670000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.385000 0.255000 3.715000 0.670000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.504100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.435000 1.075000 1.130000 ;
        RECT 0.085000 1.130000 0.255000 1.820000 ;
        RECT 0.085000 1.820000 0.435000 2.980000 ;
        RECT 0.825000 0.345000 1.075000 0.435000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.425000  1.400000 1.415000 1.650000 ;
      RECT 0.635000  1.820000 0.885000 3.245000 ;
      RECT 1.245000  1.110000 3.540000 1.280000 ;
      RECT 1.245000  1.280000 1.415000 1.400000 ;
      RECT 1.255000  0.085000 1.705000 0.940000 ;
      RECT 1.355000  1.950000 2.615000 2.120000 ;
      RECT 1.355000  2.120000 1.685000 2.980000 ;
      RECT 1.885000  2.290000 2.085000 3.245000 ;
      RECT 2.280000  0.840000 2.610000 1.080000 ;
      RECT 2.280000  1.080000 3.540000 1.110000 ;
      RECT 2.285000  2.120000 2.615000 2.980000 ;
      RECT 2.780000  0.740000 3.215000 0.910000 ;
      RECT 3.045000  0.085000 3.215000 0.740000 ;
      RECT 3.125000  1.280000 3.540000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__a211o_1
MACRO sky130_fd_sc_hs__a211o_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.260000 2.535000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.545000 1.260000 1.875000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.745000 1.260000 3.235000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405000 1.450000 3.735000 1.780000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.575000 1.010000 0.980000 1.180000 ;
        RECT 0.575000 1.180000 0.835000 2.980000 ;
        RECT 0.810000 0.350000 0.980000 1.010000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.125000  1.820000 0.375000 3.245000 ;
      RECT 0.300000  0.085000 0.630000 0.840000 ;
      RECT 1.005000  1.350000 1.335000 1.680000 ;
      RECT 1.025000  2.290000 1.355000 3.245000 ;
      RECT 1.160000  0.085000 1.330000 0.350000 ;
      RECT 1.160000  0.350000 1.870000 0.750000 ;
      RECT 1.165000  0.920000 3.740000 1.090000 ;
      RECT 1.165000  1.090000 1.335000 1.350000 ;
      RECT 1.165000  1.680000 1.335000 1.950000 ;
      RECT 1.165000  1.950000 3.735000 2.120000 ;
      RECT 1.545000  2.290000 2.865000 2.460000 ;
      RECT 1.545000  2.460000 1.875000 2.980000 ;
      RECT 2.075000  2.630000 2.365000 3.245000 ;
      RECT 2.330000  0.350000 2.700000 0.920000 ;
      RECT 2.535000  2.460000 2.865000 2.980000 ;
      RECT 2.870000  0.085000 3.040000 0.350000 ;
      RECT 2.870000  0.350000 3.310000 0.750000 ;
      RECT 3.405000  2.120000 3.735000 2.980000 ;
      RECT 3.490000  0.350000 3.740000 0.920000 ;
      RECT 3.490000  1.090000 3.740000 1.130000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__a211o_2
MACRO sky130_fd_sc_hs__a211o_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925000 1.450000 6.115000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925000 0.255000 5.320000 0.505000 ;
        RECT 4.925000 0.505000 5.125000 0.670000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.785000 1.470000 3.105000 1.720000 ;
        RECT 2.785000 1.720000 4.515000 1.890000 ;
        RECT 3.965000 1.470000 4.515000 1.720000 ;
        RECT 3.995000 1.890000 4.195000 2.150000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.450000 1.210000 3.780000 1.550000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.675000 1.240000 1.795000 1.410000 ;
        RECT 0.675000 1.410000 0.925000 1.720000 ;
        RECT 0.675000 1.720000 1.905000 1.890000 ;
        RECT 0.675000 1.890000 0.925000 2.980000 ;
        RECT 1.330000 0.350000 1.500000 0.790000 ;
        RECT 1.330000 0.790000 2.370000 0.960000 ;
        RECT 1.330000 0.960000 1.795000 1.240000 ;
        RECT 1.575000 1.890000 1.905000 2.980000 ;
        RECT 2.180000 0.545000 2.370000 0.790000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.200000 0.085000 ;
      RECT 0.000000  3.245000 7.200000 3.415000 ;
      RECT 0.225000  1.820000 0.475000 3.245000 ;
      RECT 0.820000  0.085000 1.150000 1.050000 ;
      RECT 1.125000  2.060000 1.375000 3.245000 ;
      RECT 1.680000  0.085000 2.010000 0.620000 ;
      RECT 1.965000  1.130000 3.280000 1.300000 ;
      RECT 1.965000  1.300000 2.615000 1.550000 ;
      RECT 2.105000  1.820000 2.275000 3.245000 ;
      RECT 2.445000  1.550000 2.615000 2.060000 ;
      RECT 2.445000  2.060000 3.825000 2.230000 ;
      RECT 2.540000  0.085000 2.870000 0.960000 ;
      RECT 2.545000  2.400000 4.710000 2.570000 ;
      RECT 2.545000  2.570000 2.875000 2.780000 ;
      RECT 3.040000  0.450000 3.280000 0.870000 ;
      RECT 3.040000  0.870000 4.245000 1.040000 ;
      RECT 3.040000  1.040000 3.280000 1.130000 ;
      RECT 3.045000  2.740000 4.300000 2.990000 ;
      RECT 3.460000  0.085000 3.790000 0.700000 ;
      RECT 3.960000  0.595000 4.245000 0.870000 ;
      RECT 3.960000  1.040000 4.245000 1.110000 ;
      RECT 3.960000  1.110000 6.055000 1.280000 ;
      RECT 4.420000  2.060000 6.910000 2.120000 ;
      RECT 4.420000  2.120000 5.960000 2.230000 ;
      RECT 4.420000  2.230000 4.710000 2.400000 ;
      RECT 4.425000  0.085000 4.755000 0.940000 ;
      RECT 4.500000  2.570000 4.710000 2.990000 ;
      RECT 4.880000  2.400000 5.555000 3.245000 ;
      RECT 5.295000  0.675000 6.405000 0.845000 ;
      RECT 5.680000  1.950000 6.910000 2.060000 ;
      RECT 5.725000  1.015000 6.055000 1.110000 ;
      RECT 5.725000  2.230000 5.960000 2.980000 ;
      RECT 6.130000  2.290000 6.460000 3.245000 ;
      RECT 6.235000  0.595000 6.405000 0.675000 ;
      RECT 6.235000  0.845000 6.405000 1.275000 ;
      RECT 6.580000  1.940000 6.910000 1.950000 ;
      RECT 6.585000  0.085000 6.915000 1.275000 ;
      RECT 6.630000  2.120000 6.910000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
  END
END sky130_fd_sc_hs__a211o_4
MACRO sky130_fd_sc_hs__a211oi_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.880000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.350000 1.335000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.465000 1.350000 0.835000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.545000 1.350000 1.875000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 1.180000 2.775000 1.550000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.792700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 0.350000 1.500000 0.810000 ;
        RECT 1.085000 0.810000 2.540000 1.010000 ;
        RECT 1.085000 1.010000 2.275000 1.025000 ;
        RECT 1.085000 1.025000 2.215000 1.180000 ;
        RECT 2.045000 1.180000 2.215000 1.820000 ;
        RECT 2.045000 1.820000 2.565000 2.980000 ;
        RECT 2.210000 0.350000 2.540000 0.810000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.880000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.880000 0.085000 ;
      RECT 0.000000  3.245000 2.880000 3.415000 ;
      RECT 0.315000  1.950000 1.635000 2.120000 ;
      RECT 0.315000  2.120000 0.645000 2.980000 ;
      RECT 0.340000  0.085000 0.670000 1.130000 ;
      RECT 0.815000  2.290000 1.135000 3.245000 ;
      RECT 1.305000  2.120000 1.635000 2.980000 ;
      RECT 1.670000  0.085000 2.040000 0.640000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
  END
END sky130_fd_sc_hs__a211oi_1
MACRO sky130_fd_sc_hs__a211oi_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 0.480000 1.550000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.430000 2.275000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.180000 3.715000 1.550000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.180000 4.675000 1.550000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.076000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.650000 0.635000 0.830000 1.090000 ;
        RECT 0.650000 1.090000 2.755000 1.260000 ;
        RECT 2.525000 1.260000 2.755000 1.720000 ;
        RECT 2.525000 1.720000 4.145000 1.890000 ;
        RECT 2.585000 0.840000 3.590000 1.010000 ;
        RECT 2.585000 1.010000 2.755000 1.090000 ;
        RECT 2.960000 0.330000 3.590000 0.840000 ;
        RECT 3.815000 1.890000 4.145000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.105000  1.820000 0.355000 3.245000 ;
      RECT 0.150000  0.255000 1.260000 0.425000 ;
      RECT 0.150000  0.425000 0.480000 1.010000 ;
      RECT 0.555000  1.820000 0.805000 1.950000 ;
      RECT 0.555000  1.950000 2.355000 2.060000 ;
      RECT 0.555000  2.060000 3.245000 2.120000 ;
      RECT 0.555000  2.120000 0.805000 2.980000 ;
      RECT 1.005000  2.290000 1.335000 3.245000 ;
      RECT 1.010000  0.425000 1.260000 0.750000 ;
      RECT 1.010000  0.750000 2.240000 0.920000 ;
      RECT 1.440000  0.085000 1.610000 0.330000 ;
      RECT 1.440000  0.330000 1.810000 0.580000 ;
      RECT 1.535000  2.120000 3.245000 2.230000 ;
      RECT 1.535000  2.230000 1.705000 2.980000 ;
      RECT 1.905000  2.400000 2.235000 3.245000 ;
      RECT 1.990000  0.330000 2.240000 0.750000 ;
      RECT 2.460000  0.085000 2.790000 0.670000 ;
      RECT 2.465000  2.400000 2.795000 2.905000 ;
      RECT 2.465000  2.905000 4.595000 3.075000 ;
      RECT 2.965000  2.230000 3.245000 2.735000 ;
      RECT 3.445000  2.060000 3.615000 2.905000 ;
      RECT 3.760000  0.085000 4.090000 1.010000 ;
      RECT 4.345000  1.820000 4.595000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_hs__a211oi_2
MACRO sky130_fd_sc_hs__a211oi_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505000 1.350000 3.855000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 2.275000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.300000 6.115000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365000 1.350000 7.555000 1.780000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.685800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.570000 0.785000 3.760000 0.960000 ;
        RECT 2.570000 0.960000 6.490000 1.010000 ;
        RECT 2.570000 1.010000 8.515000 1.130000 ;
        RECT 5.380000 0.350000 5.630000 0.960000 ;
        RECT 6.320000 0.350000 6.490000 0.960000 ;
        RECT 6.320000 1.130000 8.515000 1.180000 ;
        RECT 6.795000 1.950000 7.895000 2.120000 ;
        RECT 6.795000 2.120000 6.965000 2.735000 ;
        RECT 7.180000 0.350000 8.515000 1.010000 ;
        RECT 7.695000 2.120000 7.895000 2.735000 ;
        RECT 7.725000 1.180000 8.515000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
      RECT 0.000000  3.245000 8.640000 3.415000 ;
      RECT 0.345000  1.950000 6.145000 2.120000 ;
      RECT 0.345000  2.120000 0.675000 2.980000 ;
      RECT 0.420000  0.350000 0.670000 1.010000 ;
      RECT 0.420000  1.010000 2.390000 1.180000 ;
      RECT 0.850000  0.085000 1.180000 0.840000 ;
      RECT 0.875000  2.290000 1.045000 3.245000 ;
      RECT 1.245000  2.120000 1.495000 2.980000 ;
      RECT 1.360000  0.350000 1.530000 1.010000 ;
      RECT 1.695000  2.290000 2.025000 3.245000 ;
      RECT 1.710000  0.085000 2.040000 0.840000 ;
      RECT 2.220000  0.350000 4.190000 0.615000 ;
      RECT 2.220000  0.615000 2.390000 1.010000 ;
      RECT 2.225000  2.120000 2.395000 2.980000 ;
      RECT 2.595000  2.290000 2.925000 3.245000 ;
      RECT 3.125000  2.120000 3.295000 2.980000 ;
      RECT 3.495000  2.290000 3.825000 3.245000 ;
      RECT 4.025000  1.820000 4.275000 1.950000 ;
      RECT 4.025000  2.120000 4.275000 2.980000 ;
      RECT 4.465000  2.290000 4.795000 2.905000 ;
      RECT 4.465000  2.905000 8.395000 3.075000 ;
      RECT 4.995000  2.120000 5.165000 2.735000 ;
      RECT 5.365000  2.290000 5.695000 2.905000 ;
      RECT 5.810000  0.085000 6.140000 0.790000 ;
      RECT 5.895000  2.120000 6.145000 2.735000 ;
      RECT 6.315000  1.950000 6.595000 2.905000 ;
      RECT 6.670000  0.085000 7.000000 0.840000 ;
      RECT 7.165000  2.290000 7.495000 2.905000 ;
      RECT 8.065000  2.120000 8.395000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
  END
END sky130_fd_sc_hs__a211oi_4
MACRO sky130_fd_sc_hs__a21bo_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.655000 1.450000 1.315000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.255000 0.435000 0.670000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.515000 1.180000 2.845000 1.550000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.504100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.295000 0.350000 3.755000 1.130000 ;
        RECT 3.430000 1.820000 3.755000 2.980000 ;
        RECT 3.585000 1.130000 3.755000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.130000  1.940000 0.460000 1.950000 ;
      RECT 0.130000  1.950000 1.390000 2.120000 ;
      RECT 0.130000  2.120000 0.460000 2.980000 ;
      RECT 0.155000  0.840000 0.775000 1.095000 ;
      RECT 0.155000  1.095000 0.485000 1.340000 ;
      RECT 0.605000  0.085000 0.775000 0.840000 ;
      RECT 0.660000  2.290000 0.860000 3.245000 ;
      RECT 0.945000  0.660000 1.315000 1.110000 ;
      RECT 0.945000  1.110000 1.745000 1.280000 ;
      RECT 1.060000  2.120000 1.390000 2.980000 ;
      RECT 1.485000  0.085000 1.815000 0.930000 ;
      RECT 1.575000  1.280000 1.745000 1.940000 ;
      RECT 1.575000  1.940000 1.760000 2.240000 ;
      RECT 1.575000  2.240000 3.255000 2.410000 ;
      RECT 1.575000  2.410000 1.760000 2.980000 ;
      RECT 1.915000  1.100000 2.245000 1.770000 ;
      RECT 2.075000  0.350000 2.720000 0.940000 ;
      RECT 2.075000  0.940000 2.245000 1.100000 ;
      RECT 2.075000  1.770000 2.245000 1.820000 ;
      RECT 2.075000  1.820000 2.695000 2.070000 ;
      RECT 2.900000  0.085000 3.115000 0.895000 ;
      RECT 2.900000  2.580000 3.230000 3.245000 ;
      RECT 3.085000  1.320000 3.415000 1.650000 ;
      RECT 3.085000  1.650000 3.255000 2.240000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__a21bo_1
MACRO sky130_fd_sc_hs__a21bo_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.725000 1.260000 3.235000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405000 1.450000 3.735000 1.780000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 0.510000 1.550000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.020000 0.840000 1.395000 1.040000 ;
        RECT 1.020000 1.040000 1.190000 1.820000 ;
        RECT 1.020000 1.820000 1.415000 2.070000 ;
        RECT 1.225000 0.350000 1.565000 0.750000 ;
        RECT 1.225000 0.750000 1.395000 0.840000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.120000  1.820000 0.450000 2.240000 ;
      RECT 0.120000  2.240000 1.810000 2.410000 ;
      RECT 0.120000  2.410000 0.450000 2.700000 ;
      RECT 0.270000  0.540000 0.600000 0.840000 ;
      RECT 0.270000  0.840000 0.850000 1.010000 ;
      RECT 0.635000  2.580000 0.965000 3.245000 ;
      RECT 0.680000  1.010000 0.850000 2.240000 ;
      RECT 0.805000  0.085000 1.055000 0.670000 ;
      RECT 1.360000  1.220000 1.735000 1.550000 ;
      RECT 1.535000  2.580000 1.865000 3.245000 ;
      RECT 1.565000  0.920000 2.810000 1.090000 ;
      RECT 1.565000  1.090000 1.735000 1.220000 ;
      RECT 1.605000  1.720000 2.075000 1.890000 ;
      RECT 1.605000  1.890000 1.810000 2.240000 ;
      RECT 1.735000  0.085000 2.310000 0.750000 ;
      RECT 1.905000  1.260000 2.215000 1.590000 ;
      RECT 1.905000  1.590000 2.075000 1.720000 ;
      RECT 2.055000  2.060000 2.415000 2.980000 ;
      RECT 2.245000  1.760000 2.555000 1.930000 ;
      RECT 2.245000  1.930000 2.415000 2.060000 ;
      RECT 2.385000  1.090000 2.555000 1.760000 ;
      RECT 2.480000  0.350000 2.810000 0.920000 ;
      RECT 2.585000  2.100000 3.735000 2.270000 ;
      RECT 2.585000  2.270000 2.755000 2.980000 ;
      RECT 2.955000  2.440000 3.205000 3.245000 ;
      RECT 3.380000  0.085000 3.710000 1.090000 ;
      RECT 3.405000  1.950000 3.735000 2.100000 ;
      RECT 3.405000  2.270000 3.735000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__a21bo_2
MACRO sky130_fd_sc_hs__a21bo_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.450000 5.200000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.935000 0.255000 4.265000 0.670000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.255000 0.625000 0.505000 ;
        RECT 0.125000 0.505000 0.355000 0.670000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.510000 1.420000 1.850000 ;
        RECT 0.605000 1.850000 2.300000 2.100000 ;
        RECT 1.250000 0.480000 1.555000 1.010000 ;
        RECT 1.250000 1.010000 2.415000 1.180000 ;
        RECT 1.250000 1.180000 1.420000 1.510000 ;
        RECT 2.165000 0.480000 2.415000 1.010000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.240000 0.085000 ;
      RECT 0.000000  3.245000 6.240000 3.415000 ;
      RECT 0.105000  0.840000 0.615000 1.275000 ;
      RECT 0.105000  1.275000 0.435000 2.270000 ;
      RECT 0.105000  2.270000 2.640000 2.440000 ;
      RECT 0.105000  2.440000 0.435000 2.980000 ;
      RECT 0.620000  2.610000 0.950000 3.245000 ;
      RECT 0.795000  0.085000 1.045000 1.275000 ;
      RECT 1.520000  2.610000 1.850000 3.245000 ;
      RECT 1.590000  1.350000 2.755000 1.680000 ;
      RECT 1.735000  0.085000 1.985000 0.840000 ;
      RECT 2.420000  2.610000 2.750000 3.245000 ;
      RECT 2.470000  1.850000 3.290000 2.020000 ;
      RECT 2.470000  2.020000 2.640000 2.270000 ;
      RECT 2.585000  1.110000 5.035000 1.280000 ;
      RECT 2.585000  1.280000 2.755000 1.350000 ;
      RECT 2.595000  0.085000 2.845000 0.940000 ;
      RECT 2.940000  2.190000 3.270000 2.905000 ;
      RECT 2.940000  2.905000 4.090000 3.075000 ;
      RECT 2.960000  1.450000 3.290000 1.850000 ;
      RECT 3.085000  0.595000 3.415000 1.110000 ;
      RECT 3.470000  1.280000 3.720000 2.735000 ;
      RECT 3.595000  0.085000 3.765000 0.940000 ;
      RECT 3.920000  1.940000 4.090000 1.950000 ;
      RECT 3.920000  1.950000 5.970000 2.120000 ;
      RECT 3.920000  2.120000 4.090000 2.905000 ;
      RECT 4.290000  2.290000 4.540000 3.245000 ;
      RECT 4.435000  0.255000 5.545000 0.425000 ;
      RECT 4.435000  0.425000 4.605000 0.940000 ;
      RECT 4.740000  2.120000 5.070000 2.980000 ;
      RECT 4.785000  0.595000 5.035000 1.110000 ;
      RECT 5.215000  0.425000 5.545000 1.275000 ;
      RECT 5.270000  2.290000 5.520000 3.245000 ;
      RECT 5.720000  1.940000 5.970000 1.950000 ;
      RECT 5.720000  2.120000 5.970000 2.980000 ;
      RECT 5.725000  0.085000 5.975000 1.275000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
  END
END sky130_fd_sc_hs__a21bo_4
MACRO sky130_fd_sc_hs__a21boi_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.350000 2.295000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505000 1.180000 3.235000 1.550000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.120000 0.255000 0.450000 1.605000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.515200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.920000 1.525000 2.980000 ;
        RECT 1.275000 1.720000 1.875000 1.890000 ;
        RECT 1.275000 1.890000 1.525000 1.920000 ;
        RECT 1.705000 1.010000 2.060000 1.180000 ;
        RECT 1.705000 1.180000 1.875000 1.720000 ;
        RECT 1.810000 0.350000 2.060000 1.010000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.105000  1.775000 0.915000 1.945000 ;
      RECT 0.105000  1.945000 0.435000 2.980000 ;
      RECT 0.620000  0.540000 0.950000 1.050000 ;
      RECT 0.635000  2.115000 0.885000 3.245000 ;
      RECT 0.745000  1.050000 0.950000 1.220000 ;
      RECT 0.745000  1.220000 1.535000 1.550000 ;
      RECT 0.745000  1.550000 0.915000 1.775000 ;
      RECT 1.120000  0.085000 1.630000 0.760000 ;
      RECT 1.120000  0.760000 1.450000 1.050000 ;
      RECT 1.725000  2.060000 2.985000 2.230000 ;
      RECT 1.725000  2.230000 2.020000 2.980000 ;
      RECT 2.190000  2.400000 2.520000 3.245000 ;
      RECT 2.630000  0.085000 2.960000 1.010000 ;
      RECT 2.655000  1.820000 2.985000 2.060000 ;
      RECT 2.690000  2.230000 2.985000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__a21boi_1
MACRO sky130_fd_sc_hs__a21boi_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.485000 1.320000 2.815000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.265000 1.220000 3.715000 1.550000 ;
        RECT 3.485000 1.180000 3.715000 1.220000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.450000 0.475000 1.780000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.750400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.270000 0.350000 1.440000 0.980000 ;
        RECT 1.270000 0.980000 2.900000 1.150000 ;
        RECT 1.615000 1.150000 2.275000 1.410000 ;
        RECT 1.615000 1.410000 1.945000 2.735000 ;
        RECT 2.570000 0.770000 2.900000 0.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.195000  1.950000 0.445000 3.245000 ;
      RECT 0.270000  0.450000 0.520000 1.110000 ;
      RECT 0.270000  1.110000 0.975000 1.280000 ;
      RECT 0.645000  1.940000 0.975000 2.980000 ;
      RECT 0.760000  0.085000 1.090000 0.940000 ;
      RECT 0.805000  1.280000 0.975000 1.320000 ;
      RECT 0.805000  1.320000 1.395000 1.650000 ;
      RECT 0.805000  1.650000 0.975000 1.940000 ;
      RECT 1.165000  1.820000 1.415000 2.905000 ;
      RECT 1.165000  2.905000 2.315000 3.075000 ;
      RECT 1.620000  0.085000 1.950000 0.810000 ;
      RECT 2.115000  1.820000 2.315000 1.950000 ;
      RECT 2.115000  1.950000 3.215000 2.120000 ;
      RECT 2.115000  2.120000 2.315000 2.905000 ;
      RECT 2.140000  0.350000 3.250000 0.600000 ;
      RECT 2.515000  2.290000 2.845000 3.245000 ;
      RECT 3.045000  1.720000 4.215000 1.890000 ;
      RECT 3.045000  1.890000 3.215000 1.950000 ;
      RECT 3.045000  2.120000 3.215000 2.980000 ;
      RECT 3.080000  0.600000 3.250000 0.840000 ;
      RECT 3.080000  0.840000 4.190000 1.010000 ;
      RECT 3.080000  1.010000 3.250000 1.050000 ;
      RECT 3.415000  2.060000 3.765000 3.245000 ;
      RECT 3.430000  0.085000 3.760000 0.670000 ;
      RECT 3.940000  0.350000 4.190000 0.840000 ;
      RECT 3.940000  1.010000 4.190000 1.130000 ;
      RECT 3.965000  1.890000 4.215000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__a21boi_2
MACRO sky130_fd_sc_hs__a21boi_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.430000 1.795000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.365000 1.430000 3.715000 1.780000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.363000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365000 1.490000 7.555000 1.820000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  1.500800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.700000 0.770000 1.810000 0.940000 ;
        RECT 0.700000 0.940000 0.950000 1.130000 ;
        RECT 1.480000 0.940000 1.810000 1.090000 ;
        RECT 1.480000 1.090000 5.720000 1.150000 ;
        RECT 1.480000 1.150000 4.745000 1.260000 ;
        RECT 3.965000 1.260000 4.745000 1.780000 ;
        RECT 4.165000 1.780000 4.745000 1.820000 ;
        RECT 4.165000 1.820000 5.395000 1.990000 ;
        RECT 4.165000 1.990000 4.495000 2.735000 ;
        RECT 4.575000 0.980000 5.720000 1.090000 ;
        RECT 4.610000 0.350000 4.860000 0.980000 ;
        RECT 5.065000 1.990000 5.395000 2.735000 ;
        RECT 5.470000 0.350000 5.720000 0.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.680000 0.085000 ;
      RECT 0.000000  3.245000 7.680000 3.415000 ;
      RECT 0.115000  1.950000 3.995000 2.120000 ;
      RECT 0.115000  2.120000 0.365000 2.980000 ;
      RECT 0.190000  0.350000 2.160000 0.600000 ;
      RECT 0.190000  0.600000 0.520000 1.130000 ;
      RECT 0.565000  2.290000 0.895000 3.245000 ;
      RECT 1.095000  2.120000 1.265000 2.980000 ;
      RECT 1.465000  2.290000 1.795000 3.245000 ;
      RECT 1.990000  0.600000 2.160000 0.750000 ;
      RECT 1.990000  0.750000 3.960000 0.920000 ;
      RECT 1.995000  1.820000 2.165000 1.950000 ;
      RECT 1.995000  2.120000 2.165000 2.980000 ;
      RECT 2.340000  0.085000 2.670000 0.580000 ;
      RECT 2.365000  2.290000 2.615000 3.245000 ;
      RECT 2.815000  2.120000 3.145000 2.980000 ;
      RECT 2.850000  0.510000 3.020000 0.750000 ;
      RECT 3.200000  0.085000 3.530000 0.580000 ;
      RECT 3.345000  2.290000 3.515000 3.245000 ;
      RECT 3.710000  0.510000 3.960000 0.750000 ;
      RECT 3.715000  2.120000 3.995000 2.905000 ;
      RECT 3.715000  2.905000 5.845000 3.075000 ;
      RECT 4.180000  0.085000 4.430000 0.880000 ;
      RECT 4.665000  2.160000 4.895000 2.905000 ;
      RECT 4.915000  1.320000 6.195000 1.650000 ;
      RECT 5.040000  0.085000 5.290000 0.810000 ;
      RECT 5.565000  1.820000 5.845000 2.905000 ;
      RECT 5.900000  0.085000 6.230000 0.980000 ;
      RECT 6.025000  1.150000 6.660000 1.320000 ;
      RECT 6.025000  1.650000 6.195000 1.990000 ;
      RECT 6.025000  1.990000 6.815000 2.160000 ;
      RECT 6.035000  2.330000 6.365000 3.245000 ;
      RECT 6.400000  0.350000 6.660000 1.150000 ;
      RECT 6.535000  2.160000 6.815000 2.980000 ;
      RECT 7.015000  2.100000 7.265000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
  END
END sky130_fd_sc_hs__a21boi_4
MACRO sky130_fd_sc_hs__a21o_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.450000 2.375000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.645000 0.255000 3.235000 0.570000 ;
        RECT 3.005000 0.570000 3.235000 0.670000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.585000 1.450000 1.835000 1.780000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.504100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.980000 1.075000 1.150000 ;
        RECT 0.085000 1.150000 0.255000 1.820000 ;
        RECT 0.085000 1.820000 0.435000 2.980000 ;
        RECT 0.825000 0.670000 1.075000 0.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.425000  1.320000 1.415000 1.650000 ;
      RECT 0.635000  1.820000 0.885000 3.245000 ;
      RECT 1.245000  1.110000 2.135000 1.280000 ;
      RECT 1.245000  1.280000 1.415000 1.320000 ;
      RECT 1.245000  1.650000 1.415000 1.950000 ;
      RECT 1.245000  1.950000 1.605000 2.980000 ;
      RECT 1.255000  0.085000 1.585000 0.940000 ;
      RECT 1.805000  0.660000 2.135000 1.110000 ;
      RECT 1.805000  1.950000 3.065000 2.120000 ;
      RECT 1.805000  2.120000 2.135000 2.980000 ;
      RECT 2.305000  0.085000 2.475000 0.840000 ;
      RECT 2.305000  0.840000 3.040000 1.010000 ;
      RECT 2.335000  2.290000 2.535000 3.245000 ;
      RECT 2.710000  1.010000 3.040000 1.340000 ;
      RECT 2.735000  1.940000 3.065000 1.950000 ;
      RECT 2.735000  2.120000 3.065000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__a21o_1
MACRO sky130_fd_sc_hs__a21o_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.200000 1.180000 2.755000 1.550000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925000 1.180000 3.255000 1.550000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.180000 1.990000 1.535000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.570000 1.550000 0.900000 1.890000 ;
        RECT 0.570000 1.890000 0.850000 2.980000 ;
        RECT 0.725000 0.350000 1.055000 1.050000 ;
        RECT 0.725000 1.050000 0.900000 1.550000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.120000  1.820000 0.370000 3.245000 ;
      RECT 0.295000  0.085000 0.545000 1.130000 ;
      RECT 1.020000  2.045000 1.350000 3.245000 ;
      RECT 1.070000  1.220000 1.395000 1.705000 ;
      RECT 1.070000  1.705000 1.790000 1.875000 ;
      RECT 1.225000  0.085000 1.795000 0.670000 ;
      RECT 1.225000  0.840000 2.295000 1.010000 ;
      RECT 1.225000  1.010000 1.395000 1.220000 ;
      RECT 1.540000  1.875000 1.790000 2.980000 ;
      RECT 1.965000  0.350000 2.295000 0.840000 ;
      RECT 1.990000  1.720000 3.220000 1.890000 ;
      RECT 1.990000  1.890000 2.240000 2.980000 ;
      RECT 2.440000  2.060000 2.770000 3.245000 ;
      RECT 2.865000  0.085000 3.195000 1.010000 ;
      RECT 2.970000  1.890000 3.220000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__a21o_2
MACRO sky130_fd_sc_hs__a21o_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.450000 4.195000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.260000 4.905000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.425000 1.435000 2.755000 1.780000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.960000 1.690000 1.130000 ;
        RECT 0.125000 1.130000 0.355000 1.800000 ;
        RECT 0.125000 1.800000 1.835000 1.970000 ;
        RECT 0.660000 0.350000 0.830000 0.960000 ;
        RECT 0.685000 1.970000 0.855000 2.980000 ;
        RECT 1.440000 0.350000 1.690000 0.960000 ;
        RECT 1.505000 1.970000 1.835000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.150000  0.085000 0.480000 0.790000 ;
      RECT 0.155000  2.140000 0.485000 3.245000 ;
      RECT 0.635000  1.300000 2.205000 1.630000 ;
      RECT 1.010000  0.085000 1.260000 0.790000 ;
      RECT 1.055000  2.140000 1.305000 3.245000 ;
      RECT 1.870000  0.085000 2.120000 0.925000 ;
      RECT 1.870000  1.095000 3.255000 1.110000 ;
      RECT 1.870000  1.110000 4.220000 1.265000 ;
      RECT 1.870000  1.265000 2.205000 1.300000 ;
      RECT 2.035000  1.950000 2.285000 3.245000 ;
      RECT 2.360000  0.450000 2.610000 1.095000 ;
      RECT 2.475000  1.950000 2.725000 2.905000 ;
      RECT 2.475000  2.905000 3.625000 3.075000 ;
      RECT 2.790000  0.085000 3.120000 0.925000 ;
      RECT 2.925000  1.265000 4.220000 1.280000 ;
      RECT 2.925000  1.280000 3.255000 2.735000 ;
      RECT 3.455000  1.950000 5.505000 2.120000 ;
      RECT 3.455000  2.120000 3.625000 2.905000 ;
      RECT 3.460000  0.255000 4.570000 0.425000 ;
      RECT 3.460000  0.425000 3.790000 0.940000 ;
      RECT 3.825000  2.290000 4.075000 3.245000 ;
      RECT 3.960000  0.595000 4.220000 1.110000 ;
      RECT 4.275000  2.120000 4.525000 2.980000 ;
      RECT 4.400000  0.425000 4.570000 0.920000 ;
      RECT 4.400000  0.920000 5.510000 1.090000 ;
      RECT 4.725000  2.290000 5.055000 3.245000 ;
      RECT 4.750000  0.085000 5.080000 0.750000 ;
      RECT 5.255000  1.940000 5.505000 1.950000 ;
      RECT 5.255000  2.120000 5.505000 2.980000 ;
      RECT 5.260000  0.350000 5.510000 0.920000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_hs__a21o_4
MACRO sky130_fd_sc_hs__a21oi_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.920000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.350000 1.050000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.435000 1.550000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.560000 1.190000 1.815000 1.550000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.596600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.920000 0.350000 1.290000 1.010000 ;
        RECT 0.920000 1.010000 1.390000 1.180000 ;
        RECT 1.220000 1.180000 1.390000 1.720000 ;
        RECT 1.220000 1.720000 1.815000 1.890000 ;
        RECT 1.565000 1.890000 1.815000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 1.920000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 1.920000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.920000 0.085000 ;
      RECT 0.000000  3.245000 1.920000 3.415000 ;
      RECT 0.105000  1.820000 0.435000 1.985000 ;
      RECT 0.105000  1.985000 0.955000 2.060000 ;
      RECT 0.105000  2.060000 1.365000 2.230000 ;
      RECT 0.105000  2.230000 0.400000 2.980000 ;
      RECT 0.130000  0.085000 0.460000 1.010000 ;
      RECT 0.570000  2.400000 0.900000 3.245000 ;
      RECT 1.070000  2.230000 1.365000 2.980000 ;
      RECT 1.560000  0.085000 1.790000 1.020000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
  END
END sky130_fd_sc_hs__a21oi_1
MACRO sky130_fd_sc_hs__a21oi_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.350000 3.350000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.180000 2.755000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.435000 0.435000 1.780000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.739300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.350000 0.860000 0.750000 ;
        RECT 0.605000 0.750000 3.180000 0.920000 ;
        RECT 0.605000 0.920000 0.860000 1.550000 ;
        RECT 0.605000 1.550000 1.395000 1.780000 ;
        RECT 1.065000 1.780000 1.395000 2.735000 ;
        RECT 2.930000 0.920000 3.180000 1.130000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.100000  0.085000 0.430000 1.130000 ;
      RECT 0.615000  1.950000 0.895000 2.905000 ;
      RECT 0.615000  2.905000 1.845000 3.075000 ;
      RECT 1.360000  1.090000 1.775000 1.260000 ;
      RECT 1.565000  1.260000 1.775000 1.950000 ;
      RECT 1.565000  1.950000 3.690000 2.120000 ;
      RECT 1.565000  2.290000 3.705000 2.460000 ;
      RECT 1.565000  2.460000 1.845000 2.905000 ;
      RECT 2.000000  0.085000 2.330000 0.580000 ;
      RECT 2.045000  2.630000 2.305000 3.245000 ;
      RECT 2.475000  2.460000 2.805000 2.980000 ;
      RECT 2.500000  0.330000 3.690000 0.580000 ;
      RECT 3.005000  2.630000 3.175000 3.245000 ;
      RECT 3.360000  0.580000 3.690000 1.130000 ;
      RECT 3.375000  2.460000 3.705000 2.980000 ;
      RECT 3.520000  1.130000 3.690000 1.950000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__a21oi_2
MACRO sky130_fd_sc_hs__a21oi_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925000 1.350000 3.935000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.785000 1.350000 2.275000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.235000 1.350000 5.245000 1.780000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.478600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 0.595000 2.780000 0.880000 ;
        RECT 2.525000 0.880000 4.650000 1.010000 ;
        RECT 2.525000 1.010000 5.590000 1.180000 ;
        RECT 2.525000 1.180000 2.755000 1.950000 ;
        RECT 2.525000 1.950000 5.585000 2.120000 ;
        RECT 4.355000 2.120000 4.685000 2.735000 ;
        RECT 4.400000 0.350000 4.650000 0.880000 ;
        RECT 5.255000 2.120000 5.585000 2.735000 ;
        RECT 5.340000 0.350000 5.590000 1.010000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.240000 0.085000 ;
      RECT 0.000000  3.245000 6.240000 3.415000 ;
      RECT 0.305000  1.820000 0.555000 1.950000 ;
      RECT 0.305000  1.950000 2.355000 2.120000 ;
      RECT 0.305000  2.120000 0.555000 2.980000 ;
      RECT 0.380000  0.350000 0.630000 1.010000 ;
      RECT 0.380000  1.010000 2.350000 1.180000 ;
      RECT 0.755000  2.290000 1.005000 3.245000 ;
      RECT 0.810000  0.085000 1.140000 0.840000 ;
      RECT 1.205000  2.120000 1.535000 2.980000 ;
      RECT 1.320000  0.350000 1.490000 1.010000 ;
      RECT 1.670000  0.085000 2.000000 0.840000 ;
      RECT 1.735000  2.290000 1.905000 3.245000 ;
      RECT 2.105000  2.120000 2.355000 2.290000 ;
      RECT 2.105000  2.290000 4.155000 2.460000 ;
      RECT 2.105000  2.460000 2.355000 2.980000 ;
      RECT 2.180000  0.255000 4.150000 0.425000 ;
      RECT 2.180000  0.425000 2.350000 1.010000 ;
      RECT 2.555000  2.630000 2.805000 3.245000 ;
      RECT 2.960000  0.425000 3.290000 0.710000 ;
      RECT 3.005000  2.460000 3.335000 2.980000 ;
      RECT 3.535000  2.630000 3.705000 3.245000 ;
      RECT 3.820000  0.425000 4.150000 0.710000 ;
      RECT 3.905000  2.460000 4.155000 2.905000 ;
      RECT 3.905000  2.905000 6.035000 3.075000 ;
      RECT 4.830000  0.085000 5.160000 0.840000 ;
      RECT 4.885000  2.290000 5.055000 2.905000 ;
      RECT 5.785000  1.820000 6.035000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
  END
END sky130_fd_sc_hs__a21oi_4
MACRO sky130_fd_sc_hs__a221o_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965000 1.470000 2.295000 1.800000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.375000 1.350000 1.795000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.455000 2.985000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.195000 1.455000 3.715000 1.780000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.865000 0.255000 4.195000 0.670000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.504100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.350000 0.865000 1.130000 ;
        RECT 0.125000 1.130000 0.500000 1.820000 ;
        RECT 0.125000 1.820000 0.900000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.740000  1.300000 1.205000 1.630000 ;
      RECT 1.035000  1.010000 2.860000 1.115000 ;
      RECT 1.035000  1.115000 4.215000 1.180000 ;
      RECT 1.035000  1.180000 1.205000 1.300000 ;
      RECT 1.045000  0.085000 1.965000 0.840000 ;
      RECT 1.100000  1.950000 1.350000 3.245000 ;
      RECT 1.535000  1.950000 1.785000 1.970000 ;
      RECT 1.535000  1.970000 3.285000 2.140000 ;
      RECT 1.535000  2.140000 1.785000 2.980000 ;
      RECT 1.985000  2.310000 2.315000 3.245000 ;
      RECT 2.420000  0.375000 2.860000 1.010000 ;
      RECT 2.465000  1.180000 4.215000 1.285000 ;
      RECT 2.505000  2.310000 2.785000 2.905000 ;
      RECT 2.505000  2.905000 3.685000 3.075000 ;
      RECT 2.955000  1.950000 3.285000 1.970000 ;
      RECT 2.955000  2.140000 3.285000 2.735000 ;
      RECT 3.320000  0.085000 3.690000 0.945000 ;
      RECT 3.485000  1.950000 3.685000 2.905000 ;
      RECT 3.860000  0.840000 4.215000 1.115000 ;
      RECT 3.885000  1.285000 4.215000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__a221o_1
MACRO sky130_fd_sc_hs__a221o_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935000 1.450000 2.275000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.365000 1.260000 1.765000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.455000 1.450000 2.760000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.270000 1.180000 3.695000 1.550000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.865000 1.180000 4.195000 1.550000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 0.960000 0.855000 1.130000 ;
        RECT 0.100000 1.130000 0.335000 1.800000 ;
        RECT 0.100000 1.800000 0.930000 1.970000 ;
        RECT 0.600000 1.970000 0.930000 2.980000 ;
        RECT 0.605000 0.350000 0.855000 0.960000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.150000  2.140000 0.400000 3.245000 ;
      RECT 0.175000  0.085000 0.425000 0.790000 ;
      RECT 0.525000  1.300000 1.195000 1.630000 ;
      RECT 1.025000  0.920000 4.220000 1.010000 ;
      RECT 1.025000  1.010000 3.100000 1.090000 ;
      RECT 1.025000  1.090000 1.195000 1.300000 ;
      RECT 1.035000  0.085000 1.560000 0.750000 ;
      RECT 1.130000  1.950000 1.380000 3.245000 ;
      RECT 1.565000  1.950000 2.730000 2.060000 ;
      RECT 1.565000  2.060000 3.315000 2.120000 ;
      RECT 1.565000  2.120000 1.815000 2.980000 ;
      RECT 2.015000  2.290000 2.345000 3.245000 ;
      RECT 2.020000  0.350000 2.890000 0.840000 ;
      RECT 2.020000  0.840000 4.220000 0.920000 ;
      RECT 2.020000  1.090000 3.100000 1.130000 ;
      RECT 2.535000  2.400000 2.785000 2.905000 ;
      RECT 2.535000  2.905000 3.685000 3.075000 ;
      RECT 2.540000  2.120000 3.315000 2.230000 ;
      RECT 2.930000  1.130000 3.100000 1.720000 ;
      RECT 2.930000  1.720000 4.215000 1.890000 ;
      RECT 2.985000  2.230000 3.315000 2.735000 ;
      RECT 3.350000  0.085000 3.720000 0.670000 ;
      RECT 3.515000  2.060000 3.685000 2.905000 ;
      RECT 3.885000  1.890000 4.215000 2.980000 ;
      RECT 3.890000  0.350000 4.220000 0.840000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__a221o_2
MACRO sky130_fd_sc_hs__a221o_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.600000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435000 0.255000 1.765000 0.565000 ;
        RECT 1.595000 0.565000 1.765000 1.040000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.275000 0.255000 2.755000 0.505000 ;
        RECT 2.525000 0.505000 2.755000 0.670000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.615000 1.300000 9.495000 1.750000 ;
        RECT 9.095000 1.210000 9.495000 1.300000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.470000 0.255000 7.045000 0.505000 ;
        RECT 6.845000 0.505000 7.045000 0.670000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.405000 1.470000 5.735000 2.150000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  1.086400 ;
    ANTENNAPARTIALMETALSIDEAREA  2.205000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.095000 1.180000 0.385000 1.225000 ;
        RECT 0.095000 1.225000 3.265000 1.365000 ;
        RECT 0.095000 1.365000 0.385000 1.410000 ;
        RECT 2.975000 1.180000 3.265000 1.225000 ;
        RECT 2.975000 1.365000 3.265000 1.410000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.600000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.600000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.600000 0.085000 ;
      RECT 0.000000  3.245000 9.600000 3.415000 ;
      RECT 0.125000  1.180000 0.355000 1.920000 ;
      RECT 0.125000  1.920000 4.525000 2.090000 ;
      RECT 0.315000  0.655000 0.565000 0.735000 ;
      RECT 0.315000  0.735000 1.425000 0.905000 ;
      RECT 0.315000  0.905000 0.565000 1.010000 ;
      RECT 0.320000  2.260000 0.650000 3.245000 ;
      RECT 0.745000  1.075000 1.075000 1.580000 ;
      RECT 0.745000  1.580000 4.880000 1.750000 ;
      RECT 0.890000  2.260000 2.565000 2.360000 ;
      RECT 0.890000  2.360000 7.150000 2.430000 ;
      RECT 0.890000  2.430000 1.220000 2.900000 ;
      RECT 1.255000  0.905000 1.425000 1.240000 ;
      RECT 1.255000  1.240000 2.760000 1.410000 ;
      RECT 1.395000  2.600000 2.065000 3.245000 ;
      RECT 1.935000  0.085000 2.105000 0.675000 ;
      RECT 1.935000  0.675000 2.330000 1.070000 ;
      RECT 2.235000  2.430000 7.150000 2.530000 ;
      RECT 2.235000  2.530000 2.565000 2.900000 ;
      RECT 2.510000  0.840000 2.760000 1.240000 ;
      RECT 2.845000  2.700000 3.175000 3.245000 ;
      RECT 2.850000  2.090000 4.525000 2.190000 ;
      RECT 3.000000  0.085000 3.250000 0.840000 ;
      RECT 3.005000  1.010000 4.540000 1.180000 ;
      RECT 3.005000  1.180000 3.235000 1.410000 ;
      RECT 3.430000  0.440000 3.760000 1.010000 ;
      RECT 3.595000  1.350000 4.880000 1.580000 ;
      RECT 3.745000  2.700000 4.075000 3.245000 ;
      RECT 3.940000  0.085000 4.110000 0.840000 ;
      RECT 4.290000  0.480000 4.540000 1.010000 ;
      RECT 4.645000  2.700000 4.975000 3.245000 ;
      RECT 4.710000  1.130000 6.090000 1.300000 ;
      RECT 4.710000  1.300000 4.880000 1.350000 ;
      RECT 4.720000  0.085000 5.440000 0.960000 ;
      RECT 5.470000  2.700000 6.700000 2.905000 ;
      RECT 5.470000  2.905000 8.830000 3.075000 ;
      RECT 5.610000  0.580000 5.940000 1.130000 ;
      RECT 5.920000  1.300000 6.090000 1.600000 ;
      RECT 5.920000  1.600000 8.445000 1.770000 ;
      RECT 5.920000  1.770000 6.250000 2.190000 ;
      RECT 6.130000  0.085000 6.300000 0.675000 ;
      RECT 6.130000  0.675000 6.525000 0.960000 ;
      RECT 6.275000  0.960000 6.525000 1.280000 ;
      RECT 6.705000  0.840000 7.035000 1.260000 ;
      RECT 6.705000  1.260000 7.935000 1.430000 ;
      RECT 6.820000  1.940000 8.380000 2.110000 ;
      RECT 6.820000  2.110000 7.150000 2.360000 ;
      RECT 6.870000  2.530000 7.150000 2.735000 ;
      RECT 7.215000  0.085000 7.465000 1.090000 ;
      RECT 7.425000  2.280000 7.755000 2.905000 ;
      RECT 7.685000  0.255000 8.925000 0.425000 ;
      RECT 7.685000  0.425000 7.935000 1.260000 ;
      RECT 8.010000  2.110000 8.380000 2.735000 ;
      RECT 8.115000  0.595000 8.445000 1.600000 ;
      RECT 8.580000  1.940000 8.830000 2.905000 ;
      RECT 8.625000  0.425000 8.925000 1.040000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  1.210000 0.325000 1.380000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  1.210000 3.205000 1.380000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
  END
END sky130_fd_sc_hs__a221o_4
MACRO sky130_fd_sc_hs__a221oi_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505000 1.350000 2.835000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.180000 3.715000 1.550000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965000 1.350000 2.295000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.350000 1.795000 1.780000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 1.350000 0.875000 1.780000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.177500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.350000 1.090000 1.010000 ;
        RECT 0.125000 1.010000 2.575000 1.180000 ;
        RECT 0.125000 1.180000 0.375000 2.980000 ;
        RECT 2.160000 0.350000 2.575000 1.010000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.575000  1.950000 0.905000 2.905000 ;
      RECT 0.575000  2.905000 2.055000 3.075000 ;
      RECT 1.260000  0.085000 1.630000 0.825000 ;
      RECT 1.275000  1.950000 3.525000 2.120000 ;
      RECT 1.275000  2.120000 1.545000 2.735000 ;
      RECT 1.725000  2.290000 2.055000 2.905000 ;
      RECT 2.255000  2.120000 2.505000 2.980000 ;
      RECT 2.675000  2.290000 3.025000 3.245000 ;
      RECT 3.170000  0.085000 3.500000 1.010000 ;
      RECT 3.195000  1.820000 3.525000 1.950000 ;
      RECT 3.195000  2.120000 3.525000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__a221oi_1
MACRO sky130_fd_sc_hs__a221oi_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405000 1.430000 3.735000 1.950000 ;
        RECT 3.405000 1.950000 5.065000 2.120000 ;
        RECT 4.895000 1.430000 5.635000 1.780000 ;
        RECT 4.895000 1.780000 5.065000 1.950000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.430000 4.675000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.245000 1.430000 1.595000 1.680000 ;
        RECT 1.425000 1.680000 1.595000 1.950000 ;
        RECT 1.425000 1.950000 3.235000 2.120000 ;
        RECT 2.525000 1.550000 3.235000 1.950000 ;
        RECT 2.685000 1.430000 3.015000 1.550000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945000 1.430000 2.275000 1.780000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.585000 1.350000 0.915000 1.780000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.172200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.350000 0.380000 1.010000 ;
        RECT 0.125000 1.010000 1.260000 1.090000 ;
        RECT 0.125000 1.090000 5.430000 1.180000 ;
        RECT 0.125000 1.180000 0.380000 1.950000 ;
        RECT 0.125000 1.950000 0.885000 2.120000 ;
        RECT 0.555000 2.120000 0.885000 2.735000 ;
        RECT 1.090000 0.350000 1.260000 1.010000 ;
        RECT 1.090000 1.180000 5.430000 1.260000 ;
        RECT 2.950000 0.350000 3.180000 1.090000 ;
        RECT 5.180000 0.350000 5.430000 1.090000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.105000  2.290000 0.355000 2.905000 ;
      RECT 0.105000  2.905000 3.165000 2.980000 ;
      RECT 0.105000  2.980000 2.265000 3.075000 ;
      RECT 0.560000  0.085000 0.910000 0.840000 ;
      RECT 1.085000  1.850000 1.255000 2.905000 ;
      RECT 1.440000  0.350000 1.770000 0.750000 ;
      RECT 1.440000  0.750000 2.780000 0.920000 ;
      RECT 1.455000  2.290000 5.035000 2.460000 ;
      RECT 1.455000  2.460000 1.815000 2.735000 ;
      RECT 1.940000  0.085000 2.280000 0.580000 ;
      RECT 2.015000  2.630000 3.165000 2.905000 ;
      RECT 2.450000  0.330000 2.780000 0.750000 ;
      RECT 3.350000  0.330000 4.030000 0.750000 ;
      RECT 3.350000  0.750000 5.000000 0.920000 ;
      RECT 3.355000  2.630000 3.605000 3.245000 ;
      RECT 3.805000  2.460000 4.135000 2.980000 ;
      RECT 4.200000  0.085000 4.530000 0.580000 ;
      RECT 4.335000  2.630000 4.505000 3.245000 ;
      RECT 4.700000  0.330000 5.000000 0.750000 ;
      RECT 4.705000  2.460000 5.035000 2.980000 ;
      RECT 5.235000  1.950000 5.485000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_hs__a221oi_2
MACRO sky130_fd_sc_hs__a221oi_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.56000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.430000 6.115000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.430000 4.265000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365000 1.430000 8.095000 1.780000 ;
        RECT 6.730000 1.350000 8.095000 1.430000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.285000 1.350000 9.955000 1.780000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525000 1.350000 1.875000 1.780000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  2.380200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.350000 0.495000 1.010000 ;
        RECT 0.105000 1.010000 2.295000 1.090000 ;
        RECT 0.105000 1.090000 8.210000 1.180000 ;
        RECT 0.105000 1.180000 0.355000 2.905000 ;
        RECT 0.105000 2.905000 2.235000 3.075000 ;
        RECT 1.005000 2.290000 1.335000 2.905000 ;
        RECT 1.185000 0.350000 1.355000 1.010000 ;
        RECT 1.905000 2.290000 2.235000 2.905000 ;
        RECT 2.045000 0.350000 2.295000 1.010000 ;
        RECT 2.045000 1.180000 6.530000 1.260000 ;
        RECT 4.850000 0.640000 5.040000 1.090000 ;
        RECT 5.710000 0.640000 5.900000 1.090000 ;
        RECT 6.360000 0.850000 8.210000 1.090000 ;
        RECT 7.915000 0.770000 8.210000 0.850000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.560000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.560000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 10.560000 0.085000 ;
      RECT  0.000000  3.245000 10.560000 3.415000 ;
      RECT  0.555000  1.950000  9.925000 2.120000 ;
      RECT  0.555000  2.120000  0.835000 2.735000 ;
      RECT  0.675000  0.085000  1.005000 0.840000 ;
      RECT  1.505000  2.120000  1.735000 2.735000 ;
      RECT  1.535000  0.085000  1.865000 0.840000 ;
      RECT  2.615000  2.290000  6.725000 2.460000 ;
      RECT  2.615000  2.460000  2.945000 2.980000 ;
      RECT  2.630000  0.350000  2.880000 0.750000 ;
      RECT  2.630000  0.750000  4.680000 0.920000 ;
      RECT  3.060000  0.085000  3.390000 0.580000 ;
      RECT  3.145000  2.630000  3.315000 3.245000 ;
      RECT  3.515000  2.460000  3.845000 2.980000 ;
      RECT  3.570000  0.350000  3.740000 0.750000 ;
      RECT  3.920000  0.085000  4.250000 0.580000 ;
      RECT  4.045000  2.630000  4.215000 3.245000 ;
      RECT  4.415000  2.460000  4.745000 2.980000 ;
      RECT  4.430000  0.300000  6.400000 0.470000 ;
      RECT  4.430000  0.470000  4.680000 0.750000 ;
      RECT  4.945000  2.630000  5.115000 3.245000 ;
      RECT  5.210000  0.470000  5.540000 0.920000 ;
      RECT  5.315000  2.460000  5.645000 2.980000 ;
      RECT  5.815000  2.630000  6.275000 3.245000 ;
      RECT  6.070000  0.470000  6.400000 0.680000 ;
      RECT  6.445000  2.460000  6.725000 2.905000 ;
      RECT  6.445000  2.905000 10.375000 3.075000 ;
      RECT  6.590000  0.350000  8.560000 0.600000 ;
      RECT  6.590000  0.600000  6.920000 0.680000 ;
      RECT  6.895000  2.120000  7.225000 2.735000 ;
      RECT  7.395000  2.290000  7.625000 2.905000 ;
      RECT  7.450000  0.600000  7.745000 0.680000 ;
      RECT  7.795000  2.120000  8.125000 2.735000 ;
      RECT  8.295000  2.290000  8.525000 2.905000 ;
      RECT  8.390000  0.600000  8.560000 1.010000 ;
      RECT  8.390000  1.010000 10.360000 1.180000 ;
      RECT  8.695000  2.120000  9.025000 2.735000 ;
      RECT  8.740000  0.085000  9.070000 0.840000 ;
      RECT  9.195000  2.290000  9.425000 2.905000 ;
      RECT  9.250000  0.350000  9.420000 1.010000 ;
      RECT  9.595000  2.120000  9.925000 2.735000 ;
      RECT  9.600000  0.085000  9.930000 0.840000 ;
      RECT 10.110000  0.350000 10.360000 1.010000 ;
      RECT 10.125000  1.820000 10.375000 2.905000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
  END
END sky130_fd_sc_hs__a221oi_4
MACRO sky130_fd_sc_hs__a222o_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925000 1.120000 3.255000 1.520000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.120000 3.825000 1.545000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.220000 1.120000 2.755000 1.790000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.180000 1.930000 1.760000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.120000 0.550000 1.790000 ;
    END
  END C1
  PIN C2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.060000 1.120000 1.390000 1.760000 ;
    END
  END C2
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.355000 0.350000 4.710000 1.130000 ;
        RECT 4.355000 1.820000 4.710000 2.980000 ;
        RECT 4.540000 1.130000 4.710000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.115000  1.960000 0.445000 2.905000 ;
      RECT 0.115000  2.905000 2.590000 3.075000 ;
      RECT 0.140000  0.350000 0.470000 0.780000 ;
      RECT 0.140000  0.780000 4.185000 0.950000 ;
      RECT 0.720000  0.950000 0.890000 1.930000 ;
      RECT 0.720000  1.930000 1.050000 2.735000 ;
      RECT 0.960000  0.085000 1.805000 0.600000 ;
      RECT 1.220000  1.930000 1.550000 2.905000 ;
      RECT 1.720000  1.930000 2.050000 1.960000 ;
      RECT 1.720000  1.960000 3.650000 2.130000 ;
      RECT 1.720000  2.130000 2.050000 2.735000 ;
      RECT 2.260000  2.300000 2.590000 2.905000 ;
      RECT 2.295000  0.330000 3.130000 0.780000 ;
      RECT 2.820000  2.300000 3.150000 3.245000 ;
      RECT 3.320000  1.895000 3.650000 1.960000 ;
      RECT 3.320000  2.130000 3.650000 2.935000 ;
      RECT 3.620000  0.085000 4.185000 0.610000 ;
      RECT 3.855000  1.895000 4.185000 3.245000 ;
      RECT 4.015000  0.950000 4.185000 1.300000 ;
      RECT 4.015000  1.300000 4.370000 1.630000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_hs__a222o_1
MACRO sky130_fd_sc_hs__a222o_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925000 1.350000 3.255000 2.150000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.685000 1.350000 5.155000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.465000 1.350000 3.795000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.350000 4.445000 1.780000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.300000 0.435000 1.780000 ;
    END
  END C1
  PIN C2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.260000 1.140000 1.780000 ;
    END
  END C2
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695000 0.920000 2.025000 1.820000 ;
        RECT 1.695000 1.820000 2.440000 2.200000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.280000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.245000 5.280000 3.415000 ;
      RECT 0.115000  0.390000 0.365000 0.920000 ;
      RECT 0.115000  0.920000 1.525000 1.090000 ;
      RECT 0.115000  1.950000 1.525000 2.200000 ;
      RECT 0.115000  2.200000 0.365000 2.980000 ;
      RECT 0.565000  2.370000 4.165000 2.540000 ;
      RECT 0.565000  2.540000 0.895000 2.980000 ;
      RECT 0.935000  0.085000 1.185000 0.750000 ;
      RECT 1.355000  0.580000 2.400000 0.750000 ;
      RECT 1.355000  0.750000 1.525000 0.920000 ;
      RECT 1.355000  1.090000 1.525000 1.950000 ;
      RECT 1.575000  2.710000 1.905000 3.245000 ;
      RECT 2.205000  0.085000 2.535000 0.410000 ;
      RECT 2.230000  0.750000 2.400000 1.010000 ;
      RECT 2.230000  1.010000 3.750000 1.180000 ;
      RECT 2.230000  1.180000 2.560000 1.590000 ;
      RECT 2.645000  2.710000 2.975000 3.245000 ;
      RECT 2.765000  0.350000 4.090000 0.520000 ;
      RECT 2.765000  0.520000 3.095000 0.840000 ;
      RECT 3.265000  0.700000 3.750000 1.010000 ;
      RECT 3.265000  2.710000 3.630000 2.905000 ;
      RECT 3.265000  2.905000 4.665000 3.075000 ;
      RECT 3.835000  1.950000 4.165000 2.370000 ;
      RECT 3.835000  2.540000 4.165000 2.735000 ;
      RECT 3.920000  0.520000 4.090000 1.010000 ;
      RECT 3.920000  1.010000 5.140000 1.180000 ;
      RECT 4.260000  0.085000 4.590000 0.840000 ;
      RECT 4.335000  1.950000 4.665000 2.905000 ;
      RECT 4.810000  0.350000 5.140000 1.010000 ;
      RECT 4.835000  1.950000 5.165000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
  END
END sky130_fd_sc_hs__a222o_2
MACRO sky130_fd_sc_hs__a222oi_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.155000 1.120000 3.715000 1.790000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.885000 1.180000 4.215000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.120000 2.875000 1.790000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975000 1.120000 2.305000 1.790000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.120000 0.595000 1.790000 ;
    END
  END C1
  PIN C2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985000 1.120000 1.315000 1.790000 ;
    END
  END C2
  PIN Y
    ANTENNADIFFAREA  1.232000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 1.960000 1.655000 2.130000 ;
        RECT 0.115000 2.130000 0.445000 2.980000 ;
        RECT 0.140000 0.350000 0.470000 0.780000 ;
        RECT 0.140000 0.780000 3.360000 0.950000 ;
        RECT 1.115000 2.130000 1.655000 2.735000 ;
        RECT 1.485000 0.950000 1.795000 1.780000 ;
        RECT 1.485000 1.780000 1.655000 1.960000 ;
        RECT 2.525000 0.330000 3.360000 0.780000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.615000  2.300000 0.945000 2.905000 ;
      RECT 0.615000  2.905000 2.655000 3.075000 ;
      RECT 0.960000  0.085000 2.180000 0.600000 ;
      RECT 1.825000  1.960000 4.205000 2.130000 ;
      RECT 1.825000  2.130000 2.155000 2.735000 ;
      RECT 2.325000  2.300000 2.655000 2.905000 ;
      RECT 2.825000  2.130000 3.155000 2.980000 ;
      RECT 3.325000  2.300000 3.655000 3.245000 ;
      RECT 3.850000  0.085000 4.180000 0.950000 ;
      RECT 3.875000  2.130000 4.205000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__a222oi_1
MACRO sky130_fd_sc_hs__a222oi_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.685000 1.450000 5.115000 1.780000 ;
        RECT 4.945000 1.780000 5.115000 1.950000 ;
        RECT 4.945000 1.950000 6.055000 2.120000 ;
        RECT 5.885000 1.450000 6.455000 1.780000 ;
        RECT 5.885000 1.780000 6.055000 1.950000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.305000 1.450000 5.635000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.675000 1.470000 3.235000 1.800000 ;
        RECT 3.065000 1.800000 3.235000 1.950000 ;
        RECT 3.065000 1.950000 4.275000 2.120000 ;
        RECT 4.105000 1.450000 4.475000 1.780000 ;
        RECT 4.105000 1.780000 4.275000 1.950000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405000 1.260000 3.735000 1.780000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.165000 1.335000 1.495000 ;
    END
  END C1
  PIN C2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.165000 0.835000 1.495000 ;
        RECT 0.605000 1.495000 0.835000 1.665000 ;
        RECT 0.605000 1.665000 2.125000 1.835000 ;
        RECT 1.795000 1.130000 2.125000 1.665000 ;
    END
  END C2
  PIN Y
    ANTENNADIFFAREA  1.693200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.825000 1.420000 0.995000 ;
        RECT 0.085000 0.995000 0.255000 1.920000 ;
        RECT 0.085000 1.920000 0.365000 2.005000 ;
        RECT 0.085000 2.005000 2.465000 2.175000 ;
        RECT 0.085000 2.175000 0.365000 2.980000 ;
        RECT 1.065000 2.175000 1.325000 2.735000 ;
        RECT 1.090000 0.780000 1.420000 0.825000 ;
        RECT 1.995000 2.175000 2.465000 2.735000 ;
        RECT 2.295000 1.130000 2.840000 1.300000 ;
        RECT 2.295000 1.300000 2.465000 2.005000 ;
        RECT 2.510000 0.350000 2.840000 0.920000 ;
        RECT 2.510000 0.920000 4.715000 1.090000 ;
        RECT 2.510000 1.090000 2.840000 1.130000 ;
        RECT 4.450000 0.350000 4.715000 0.920000 ;
        RECT 4.450000 1.090000 4.715000 1.110000 ;
        RECT 4.450000 1.110000 6.580000 1.280000 ;
        RECT 6.320000 0.350000 6.580000 1.110000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.720000 0.085000 ;
      RECT 0.000000  3.245000 6.720000 3.415000 ;
      RECT 0.115000  0.085000 0.480000 0.655000 ;
      RECT 0.565000  2.345000 0.895000 2.905000 ;
      RECT 0.565000  2.905000 4.325000 2.980000 ;
      RECT 0.565000  2.980000 3.335000 3.075000 ;
      RECT 0.660000  0.350000 1.780000 0.610000 ;
      RECT 1.495000  2.345000 1.825000 2.905000 ;
      RECT 1.590000  0.610000 1.780000 0.885000 ;
      RECT 1.950000  0.085000 2.280000 0.940000 ;
      RECT 2.635000  1.970000 2.805000 2.290000 ;
      RECT 2.635000  2.290000 6.605000 2.460000 ;
      RECT 2.635000  2.460000 2.805000 2.735000 ;
      RECT 3.005000  2.630000 3.335000 2.650000 ;
      RECT 3.005000  2.650000 4.325000 2.905000 ;
      RECT 3.020000  0.350000 3.270000 0.580000 ;
      RECT 3.020000  0.580000 4.270000 0.750000 ;
      RECT 3.450000  0.085000 3.840000 0.410000 ;
      RECT 4.020000  0.350000 4.270000 0.580000 ;
      RECT 4.445000  1.950000 4.775000 2.290000 ;
      RECT 4.500000  2.460000 6.605000 2.480000 ;
      RECT 4.500000  2.480000 4.715000 2.980000 ;
      RECT 4.885000  0.350000 5.215000 0.770000 ;
      RECT 4.885000  0.770000 6.150000 0.940000 ;
      RECT 4.895000  2.650000 5.255000 3.245000 ;
      RECT 5.385000  0.085000 5.715000 0.600000 ;
      RECT 5.425000  2.480000 5.655000 2.980000 ;
      RECT 5.825000  2.650000 6.155000 3.245000 ;
      RECT 5.900000  0.330000 6.150000 0.770000 ;
      RECT 6.275000  1.950000 6.605000 2.290000 ;
      RECT 6.335000  2.480000 6.605000 3.000000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
  END
END sky130_fd_sc_hs__a222oi_2
MACRO sky130_fd_sc_hs__a22o_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965000 1.350000 2.295000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.255000 0.560000 0.505000 ;
        RECT 0.125000 0.505000 0.355000 0.670000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.425000 1.470000 1.795000 1.800000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.470000 1.215000 1.800000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.504100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925000 0.350000 3.255000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.195000  1.970000 0.445000 3.245000 ;
      RECT 0.220000  0.840000 0.550000 1.130000 ;
      RECT 0.220000  1.130000 1.285000 1.300000 ;
      RECT 0.645000  1.970000 0.895000 2.905000 ;
      RECT 0.645000  2.905000 1.995000 3.075000 ;
      RECT 0.730000  0.085000 0.945000 0.960000 ;
      RECT 1.095000  1.970000 2.755000 2.140000 ;
      RECT 1.095000  2.140000 1.425000 2.735000 ;
      RECT 1.115000  0.375000 2.245000 0.625000 ;
      RECT 1.115000  0.625000 1.285000 1.130000 ;
      RECT 1.485000  0.795000 1.815000 1.010000 ;
      RECT 1.485000  1.010000 2.755000 1.180000 ;
      RECT 1.595000  2.310000 1.995000 2.905000 ;
      RECT 2.165000  2.310000 2.725000 3.245000 ;
      RECT 2.495000  0.085000 2.745000 0.840000 ;
      RECT 2.505000  1.180000 2.755000 1.970000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__a22o_1
MACRO sky130_fd_sc_hs__a22o_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.585000 1.350000 1.905000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405000 1.350000 3.735000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.075000 1.350000 2.495000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.705000 1.350000 3.235000 1.780000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.530000 0.350000 0.860000 1.720000 ;
        RECT 0.530000 1.720000 1.075000 1.890000 ;
        RECT 0.905000 1.890000 1.075000 2.290000 ;
        RECT 0.905000 2.290000 1.185000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.100000  0.085000 0.350000 1.130000 ;
      RECT 0.485000  2.060000 0.735000 3.245000 ;
      RECT 1.040000  0.085000 1.290000 0.840000 ;
      RECT 1.085000  1.010000 2.330000 1.180000 ;
      RECT 1.085000  1.180000 1.415000 1.550000 ;
      RECT 1.245000  1.550000 1.415000 1.950000 ;
      RECT 1.245000  1.950000 2.705000 2.120000 ;
      RECT 1.385000  2.290000 1.715000 3.245000 ;
      RECT 1.500000  0.255000 2.670000 0.425000 ;
      RECT 1.500000  0.425000 1.830000 0.840000 ;
      RECT 1.925000  2.290000 2.255000 2.905000 ;
      RECT 1.925000  2.905000 3.225000 3.075000 ;
      RECT 2.000000  0.595000 2.330000 1.010000 ;
      RECT 2.455000  2.120000 2.705000 2.735000 ;
      RECT 2.500000  0.425000 2.670000 1.010000 ;
      RECT 2.500000  1.010000 3.700000 1.180000 ;
      RECT 2.870000  0.085000 3.200000 0.840000 ;
      RECT 2.875000  1.950000 3.225000 2.905000 ;
      RECT 3.370000  0.350000 3.700000 1.010000 ;
      RECT 3.395000  1.950000 3.725000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__a22o_2
MACRO sky130_fd_sc_hs__a22o_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.405000 1.450000 6.115000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.955000 0.255000 5.320000 0.505000 ;
        RECT 4.955000 0.505000 5.125000 0.670000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.495000 1.435000 3.825000 1.765000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.025000 1.435000 3.325000 1.765000 ;
        RECT 3.155000 1.765000 3.325000 1.935000 ;
        RECT 3.155000 1.935000 4.195000 2.150000 ;
        RECT 4.025000 1.440000 4.655000 1.770000 ;
        RECT 4.025000 1.770000 4.195000 1.935000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.140000 2.515000 1.180000 ;
        RECT 0.125000 1.180000 1.855000 1.410000 ;
        RECT 0.705000 1.410000 1.855000 1.650000 ;
        RECT 0.705000 1.650000 0.875000 2.980000 ;
        RECT 1.405000 0.480000 1.655000 1.010000 ;
        RECT 1.405000 1.010000 2.515000 1.140000 ;
        RECT 1.525000 1.650000 1.855000 2.980000 ;
        RECT 2.265000 0.480000 2.515000 1.010000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.200000 0.085000 ;
      RECT 0.000000  3.245000 7.200000 3.415000 ;
      RECT 0.175000  1.900000 0.505000 3.245000 ;
      RECT 0.975000  0.085000 1.225000 0.970000 ;
      RECT 1.075000  1.820000 1.325000 3.245000 ;
      RECT 1.835000  0.085000 2.085000 0.840000 ;
      RECT 2.025000  1.350000 2.855000 1.680000 ;
      RECT 2.055000  1.850000 2.305000 3.245000 ;
      RECT 2.475000  1.680000 2.645000 2.905000 ;
      RECT 2.475000  2.905000 4.415000 2.980000 ;
      RECT 2.475000  2.980000 3.515000 3.075000 ;
      RECT 2.685000  1.095000 6.055000 1.265000 ;
      RECT 2.685000  1.265000 2.855000 1.350000 ;
      RECT 2.695000  0.085000 3.025000 0.925000 ;
      RECT 2.815000  1.940000 2.985000 2.320000 ;
      RECT 2.815000  2.320000 4.865000 2.490000 ;
      RECT 2.815000  2.490000 2.985000 2.735000 ;
      RECT 3.185000  2.660000 4.415000 2.905000 ;
      RECT 3.200000  0.580000 4.355000 0.830000 ;
      RECT 3.630000  1.000000 3.960000 1.095000 ;
      RECT 4.140000  0.830000 4.355000 0.925000 ;
      RECT 4.535000  0.085000 4.785000 0.925000 ;
      RECT 4.615000  1.940000 4.865000 1.950000 ;
      RECT 4.615000  1.950000 6.910000 2.120000 ;
      RECT 4.615000  2.120000 4.865000 2.320000 ;
      RECT 4.615000  2.490000 4.865000 2.980000 ;
      RECT 5.035000  2.290000 5.510000 3.245000 ;
      RECT 5.295000  0.675000 6.405000 0.845000 ;
      RECT 5.680000  2.120000 5.930000 2.980000 ;
      RECT 5.725000  1.015000 6.055000 1.095000 ;
      RECT 5.725000  1.265000 6.055000 1.275000 ;
      RECT 6.130000  2.290000 6.460000 3.245000 ;
      RECT 6.235000  0.595000 6.405000 0.675000 ;
      RECT 6.235000  0.845000 6.405000 1.275000 ;
      RECT 6.585000  0.085000 6.915000 1.275000 ;
      RECT 6.660000  1.940000 6.910000 1.950000 ;
      RECT 6.660000  2.120000 6.910000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
  END
END sky130_fd_sc_hs__a22o_4
MACRO sky130_fd_sc_hs__a22oi_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.880000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.545000 1.350000 1.875000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.350000 2.755000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.350000 1.335000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.435000 1.780000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.624600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.010000 1.570000 1.180000 ;
        RECT 0.605000 1.180000 0.835000 1.950000 ;
        RECT 0.605000 1.950000 1.015000 2.120000 ;
        RECT 0.845000 2.120000 1.015000 2.735000 ;
        RECT 1.130000 0.350000 1.570000 1.010000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.880000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.880000 0.085000 ;
      RECT 0.000000  3.245000 2.880000 3.415000 ;
      RECT 0.315000  2.290000 0.645000 2.905000 ;
      RECT 0.315000  2.905000 1.545000 3.075000 ;
      RECT 0.340000  0.085000 0.670000 0.840000 ;
      RECT 1.215000  1.950000 2.565000 2.120000 ;
      RECT 1.215000  2.120000 1.545000 2.905000 ;
      RECT 1.715000  2.290000 2.065000 3.245000 ;
      RECT 2.210000  0.085000 2.540000 1.130000 ;
      RECT 2.235000  2.120000 2.565000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
  END
END sky130_fd_sc_hs__a22oi_1
MACRO sky130_fd_sc_hs__a22oi_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.430000 0.880000 1.780000 ;
        RECT 0.710000 1.780000 0.880000 1.950000 ;
        RECT 0.710000 1.950000 2.210000 2.120000 ;
        RECT 1.880000 1.430000 2.210000 1.950000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.050000 1.430000 1.420000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.720000 1.090000 4.075000 1.260000 ;
        RECT 2.720000 1.260000 3.235000 1.550000 ;
        RECT 3.905000 1.260000 4.075000 1.300000 ;
        RECT 3.905000 1.300000 4.370000 1.630000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405000 1.430000 3.735000 1.780000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.497400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.285000 0.350000 0.535000 1.090000 ;
        RECT 0.285000 1.090000 2.550000 1.260000 ;
        RECT 2.040000 0.810000 2.550000 1.090000 ;
        RECT 2.145000 0.350000 2.550000 0.810000 ;
        RECT 2.380000 1.260000 2.550000 1.720000 ;
        RECT 2.380000 1.720000 3.130000 1.890000 ;
        RECT 2.930000 1.890000 3.130000 1.950000 ;
        RECT 2.930000 1.950000 4.710000 2.120000 ;
        RECT 2.930000 2.120000 3.130000 2.735000 ;
        RECT 3.860000 2.120000 4.030000 2.735000 ;
        RECT 4.245000 0.350000 4.710000 1.130000 ;
        RECT 4.540000 1.130000 4.710000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.290000  1.950000 0.540000 2.290000 ;
      RECT 0.290000  2.290000 2.730000 2.460000 ;
      RECT 0.290000  2.460000 0.540000 2.980000 ;
      RECT 0.715000  0.330000 0.965000 0.750000 ;
      RECT 0.715000  0.750000 1.815000 0.920000 ;
      RECT 0.740000  2.630000 0.990000 3.245000 ;
      RECT 1.145000  0.085000 1.475000 0.580000 ;
      RECT 1.190000  2.460000 1.520000 2.980000 ;
      RECT 1.645000  0.350000 1.975000 0.640000 ;
      RECT 1.645000  0.640000 1.815000 0.750000 ;
      RECT 1.690000  2.630000 2.230000 3.245000 ;
      RECT 2.400000  2.060000 2.730000 2.290000 ;
      RECT 2.400000  2.460000 2.730000 2.905000 ;
      RECT 2.400000  2.905000 4.560000 3.075000 ;
      RECT 2.835000  0.330000 3.135000 0.750000 ;
      RECT 2.835000  0.750000 4.065000 0.920000 ;
      RECT 3.305000  0.085000 3.635000 0.580000 ;
      RECT 3.330000  2.290000 3.660000 2.905000 ;
      RECT 3.815000  0.330000 4.065000 0.750000 ;
      RECT 4.230000  2.290000 4.560000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_hs__a22oi_2
MACRO sky130_fd_sc_hs__a22oi_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.350000 5.635000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885000 1.350000 7.465000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.265000 1.350000 3.275000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.350000 1.955000 1.780000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  2.172800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.635000 1.950000 3.615000 2.120000 ;
        RECT 0.635000 2.120000 0.885000 2.735000 ;
        RECT 1.615000 2.120000 1.785000 2.735000 ;
        RECT 2.350000 0.595000 2.680000 1.010000 ;
        RECT 2.350000 1.010000 5.780000 1.130000 ;
        RECT 2.350000 1.130000 4.195000 1.180000 ;
        RECT 2.515000 2.120000 2.685000 2.735000 ;
        RECT 3.210000 0.770000 3.990000 0.850000 ;
        RECT 3.210000 0.850000 5.780000 1.010000 ;
        RECT 3.415000 2.120000 3.615000 2.735000 ;
        RECT 3.445000 1.180000 4.195000 1.520000 ;
        RECT 3.445000 1.520000 3.615000 1.950000 ;
        RECT 5.450000 0.770000 5.780000 0.850000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.185000  1.820000 0.435000 2.905000 ;
      RECT 0.185000  2.905000 4.035000 3.075000 ;
      RECT 0.200000  0.350000 0.450000 1.010000 ;
      RECT 0.200000  1.010000 2.170000 1.180000 ;
      RECT 0.630000  0.085000 0.880000 0.840000 ;
      RECT 1.060000  0.350000 1.310000 1.010000 ;
      RECT 1.085000  2.290000 1.415000 2.905000 ;
      RECT 1.490000  0.085000 1.820000 0.840000 ;
      RECT 1.985000  2.290000 2.315000 2.905000 ;
      RECT 2.000000  0.255000 3.970000 0.425000 ;
      RECT 2.000000  0.425000 2.170000 1.010000 ;
      RECT 2.860000  0.425000 3.970000 0.600000 ;
      RECT 2.860000  0.600000 3.030000 0.840000 ;
      RECT 2.885000  2.290000 3.215000 2.905000 ;
      RECT 3.785000  1.820000 4.035000 1.950000 ;
      RECT 3.785000  1.950000 7.945000 2.120000 ;
      RECT 3.785000  2.120000 4.035000 2.905000 ;
      RECT 4.160000  0.350000 6.130000 0.600000 ;
      RECT 4.160000  0.600000 4.490000 0.680000 ;
      RECT 4.235000  2.290000 4.565000 3.245000 ;
      RECT 4.765000  2.120000 5.015000 2.980000 ;
      RECT 5.185000  2.290000 5.645000 3.245000 ;
      RECT 5.815000  2.120000 6.065000 2.980000 ;
      RECT 5.960000  0.600000 6.130000 1.010000 ;
      RECT 5.960000  1.010000 7.930000 1.180000 ;
      RECT 6.265000  2.290000 6.595000 3.245000 ;
      RECT 6.310000  0.085000 6.560000 0.840000 ;
      RECT 6.740000  0.350000 6.990000 1.010000 ;
      RECT 6.795000  2.120000 6.965000 2.980000 ;
      RECT 7.165000  2.290000 7.495000 3.245000 ;
      RECT 7.170000  0.085000 7.420000 0.840000 ;
      RECT 7.600000  0.350000 7.930000 1.010000 ;
      RECT 7.695000  1.820000 7.945000 1.950000 ;
      RECT 7.695000  2.120000 7.945000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_hs__a22oi_4
MACRO sky130_fd_sc_hs__a2bb2o_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  0.233000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.070000 1.180000 1.335000 1.620000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.233000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.545000 1.180000 1.850000 1.620000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 0.255000 4.195000 0.670000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.875000 1.450000 3.235000 1.780000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.504100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.420000 0.590000 1.150000 ;
        RECT 0.125000 1.150000 0.295000 1.820000 ;
        RECT 0.125000 1.820000 0.560000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.465000  1.320000 0.900000 1.650000 ;
      RECT 0.730000  1.650000 0.900000 1.790000 ;
      RECT 0.730000  1.790000 2.190000 1.960000 ;
      RECT 0.760000  2.130000 1.090000 3.245000 ;
      RECT 0.770000  0.085000 1.100000 1.010000 ;
      RECT 1.285000  0.255000 2.595000 0.520000 ;
      RECT 1.285000  0.520000 1.590000 1.010000 ;
      RECT 1.325000  1.960000 1.495000 2.905000 ;
      RECT 1.325000  2.905000 2.515000 3.075000 ;
      RECT 1.665000  2.130000 2.530000 2.300000 ;
      RECT 1.665000  2.300000 1.995000 2.735000 ;
      RECT 1.760000  0.690000 2.935000 0.860000 ;
      RECT 2.020000  1.030000 2.900000 1.210000 ;
      RECT 2.020000  1.210000 2.190000 1.790000 ;
      RECT 2.185000  2.470000 2.515000 2.905000 ;
      RECT 2.360000  1.450000 2.665000 1.780000 ;
      RECT 2.360000  1.780000 2.530000 2.130000 ;
      RECT 2.715000  1.950000 3.895000 2.120000 ;
      RECT 2.715000  2.120000 2.885000 2.980000 ;
      RECT 2.765000  0.085000 2.935000 0.690000 ;
      RECT 3.085000  2.290000 3.445000 3.245000 ;
      RECT 3.145000  0.085000 3.315000 0.840000 ;
      RECT 3.145000  0.840000 3.870000 1.010000 ;
      RECT 3.540000  1.010000 3.870000 1.290000 ;
      RECT 3.645000  1.940000 3.895000 1.950000 ;
      RECT 3.645000  2.120000 3.895000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__a2bb2o_1
MACRO sky130_fd_sc_hs__a2bb2o_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  0.233000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925000 1.180000 3.255000 2.150000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.233000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.385000 1.180000 2.755000 1.510000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.435000 1.550000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.180000 1.315000 1.550000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 0.350000 3.920000 2.150000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.265000  1.720000 1.415000 1.890000 ;
      RECT 0.265000  1.890000 0.515000 2.980000 ;
      RECT 0.290000  0.085000 0.620000 1.010000 ;
      RECT 0.715000  2.060000 1.045000 3.245000 ;
      RECT 1.080000  0.350000 1.480000 0.840000 ;
      RECT 1.080000  0.840000 1.655000 1.010000 ;
      RECT 1.245000  1.890000 1.415000 2.980000 ;
      RECT 1.485000  1.010000 1.655000 1.380000 ;
      RECT 1.485000  1.380000 1.755000 1.550000 ;
      RECT 1.585000  1.550000 1.755000 2.020000 ;
      RECT 1.585000  2.020000 1.945000 2.810000 ;
      RECT 1.585000  2.810000 2.920000 2.980000 ;
      RECT 1.650000  0.085000 2.520000 0.670000 ;
      RECT 1.925000  0.840000 2.870000 1.010000 ;
      RECT 1.925000  1.010000 2.175000 1.680000 ;
      RECT 1.925000  1.680000 2.580000 1.850000 ;
      RECT 2.265000  1.850000 2.580000 2.640000 ;
      RECT 2.690000  0.350000 2.870000 0.840000 ;
      RECT 2.750000  2.320000 4.470000 2.490000 ;
      RECT 2.750000  2.490000 2.920000 2.810000 ;
      RECT 3.050000  0.085000 3.315000 0.940000 ;
      RECT 3.105000  2.660000 3.495000 3.245000 ;
      RECT 4.065000  2.660000 4.395000 3.245000 ;
      RECT 4.090000  1.350000 4.470000 2.320000 ;
      RECT 4.100000  0.085000 4.350000 1.130000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_hs__a2bb2o_2
MACRO sky130_fd_sc_hs__a2bb2o_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  0.264000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555000 1.350000 2.850000 1.780000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.264000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.360000 1.350000 3.685000 1.780000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365000 1.260000 7.075000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.405000 1.260000 6.115000 1.780000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.960000 2.045000 1.130000 ;
        RECT 0.125000 1.130000 0.835000 1.780000 ;
        RECT 0.665000 1.780000 0.835000 1.800000 ;
        RECT 0.665000 1.800000 2.240000 1.970000 ;
        RECT 0.935000 0.350000 1.185000 0.960000 ;
        RECT 1.010000 1.970000 1.340000 2.980000 ;
        RECT 1.795000 0.350000 2.045000 0.960000 ;
        RECT 1.910000 1.970000 2.240000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.200000 0.085000 ;
      RECT 0.000000  3.245000 7.200000 3.415000 ;
      RECT 0.505000  0.085000 0.755000 0.790000 ;
      RECT 0.560000  2.140000 0.810000 3.245000 ;
      RECT 1.035000  1.300000 2.385000 1.630000 ;
      RECT 1.365000  0.085000 1.615000 0.790000 ;
      RECT 1.540000  2.140000 1.710000 3.245000 ;
      RECT 2.215000  1.010000 2.815000 1.180000 ;
      RECT 2.215000  1.180000 2.385000 1.300000 ;
      RECT 2.225000  0.085000 2.475000 0.840000 ;
      RECT 2.410000  1.950000 2.780000 3.245000 ;
      RECT 2.645000  0.255000 3.530000 0.425000 ;
      RECT 2.645000  0.425000 2.815000 1.010000 ;
      RECT 2.985000  0.595000 3.190000 1.130000 ;
      RECT 3.020000  1.130000 3.190000 1.950000 ;
      RECT 3.020000  1.950000 4.150000 2.120000 ;
      RECT 3.290000  2.120000 3.620000 2.980000 ;
      RECT 3.360000  0.425000 3.530000 1.010000 ;
      RECT 3.360000  1.010000 4.815000 1.180000 ;
      RECT 3.700000  0.085000 4.385000 0.840000 ;
      RECT 3.855000  1.470000 4.150000 1.950000 ;
      RECT 4.060000  2.290000 4.390000 2.905000 ;
      RECT 4.060000  2.905000 5.210000 3.075000 ;
      RECT 4.565000  0.350000 5.765000 0.600000 ;
      RECT 4.565000  0.600000 4.815000 1.010000 ;
      RECT 4.565000  1.180000 4.760000 2.735000 ;
      RECT 4.960000  1.950000 7.090000 2.120000 ;
      RECT 4.960000  2.120000 5.210000 2.905000 ;
      RECT 5.005000  0.770000 6.115000 0.920000 ;
      RECT 5.005000  0.920000 7.095000 1.090000 ;
      RECT 5.410000  2.290000 5.660000 3.245000 ;
      RECT 5.860000  2.120000 6.190000 2.980000 ;
      RECT 5.945000  0.350000 6.115000 0.770000 ;
      RECT 6.295000  0.350000 6.665000 0.750000 ;
      RECT 6.390000  2.290000 6.560000 3.245000 ;
      RECT 6.495000  0.085000 6.665000 0.350000 ;
      RECT 6.760000  2.120000 7.090000 2.980000 ;
      RECT 6.845000  0.350000 7.095000 0.920000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
  END
END sky130_fd_sc_hs__a2bb2o_4
MACRO sky130_fd_sc_hs__a2bb2oi_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  0.233000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.260000 0.435000 1.780000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.233000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.450000 1.100000 1.780000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925000 1.180000 3.255000 1.550000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.220000 1.220000 2.755000 1.540000 ;
        RECT 2.525000 1.540000 2.755000 2.150000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.515200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.530000 2.290000 1.780000 2.980000 ;
        RECT 1.610000 1.750000 2.050000 1.920000 ;
        RECT 1.610000 1.920000 2.275000 2.220000 ;
        RECT 1.610000 2.220000 1.780000 2.290000 ;
        RECT 1.880000 0.880000 2.315000 1.050000 ;
        RECT 1.880000 1.050000 2.050000 1.750000 ;
        RECT 2.055000 0.350000 2.315000 0.880000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.120000  1.950000 0.450000 3.245000 ;
      RECT 0.175000  0.085000 0.425000 1.090000 ;
      RECT 0.605000  0.540000 0.935000 0.960000 ;
      RECT 0.605000  0.960000 1.440000 1.130000 ;
      RECT 0.960000  1.950000 1.440000 2.120000 ;
      RECT 0.960000  2.120000 1.290000 2.980000 ;
      RECT 1.105000  0.085000 1.885000 0.710000 ;
      RECT 1.105000  0.710000 1.710000 0.790000 ;
      RECT 1.270000  1.130000 1.440000 1.220000 ;
      RECT 1.270000  1.220000 1.710000 1.550000 ;
      RECT 1.270000  1.550000 1.440000 1.950000 ;
      RECT 1.980000  2.390000 3.240000 2.560000 ;
      RECT 1.980000  2.560000 2.230000 2.980000 ;
      RECT 2.430000  2.730000 2.790000 2.980000 ;
      RECT 2.430000  2.980000 2.600000 3.245000 ;
      RECT 2.885000  0.085000 3.215000 1.010000 ;
      RECT 2.990000  1.820000 3.240000 2.390000 ;
      RECT 2.990000  2.560000 3.240000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__a2bb2oi_1
MACRO sky130_fd_sc_hs__a2bb2oi_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.285000 0.435000 0.670000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.450000 1.570000 1.780000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.350000 4.675000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405000 1.320000 3.735000 1.780000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.750400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.080000 0.390000 2.250000 0.980000 ;
        RECT 2.080000 0.980000 3.795000 1.150000 ;
        RECT 2.525000 1.150000 3.235000 1.410000 ;
        RECT 2.525000 1.410000 2.780000 2.735000 ;
        RECT 3.465000 0.770000 3.795000 0.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.280000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.245000 5.280000 3.415000 ;
      RECT 0.580000  1.940000 0.910000 3.245000 ;
      RECT 0.605000  0.085000 0.855000 1.170000 ;
      RECT 1.035000  0.490000 1.330000 1.110000 ;
      RECT 1.035000  1.110000 1.910000 1.280000 ;
      RECT 1.420000  1.950000 1.910000 2.980000 ;
      RECT 1.570000  0.085000 1.900000 0.940000 ;
      RECT 1.740000  1.280000 1.910000 1.320000 ;
      RECT 1.740000  1.320000 2.205000 1.650000 ;
      RECT 1.740000  1.650000 1.910000 1.950000 ;
      RECT 2.080000  1.820000 2.330000 2.905000 ;
      RECT 2.080000  2.905000 3.230000 3.075000 ;
      RECT 2.430000  0.085000 2.760000 0.810000 ;
      RECT 2.980000  1.820000 3.230000 1.950000 ;
      RECT 2.980000  1.950000 5.110000 2.120000 ;
      RECT 2.980000  2.120000 3.230000 2.905000 ;
      RECT 3.035000  0.350000 4.145000 0.600000 ;
      RECT 3.430000  2.290000 3.760000 3.245000 ;
      RECT 3.960000  2.120000 4.130000 2.980000 ;
      RECT 3.975000  0.600000 4.145000 1.010000 ;
      RECT 3.975000  1.010000 5.085000 1.180000 ;
      RECT 4.325000  0.085000 4.575000 0.840000 ;
      RECT 4.330000  2.290000 4.660000 3.245000 ;
      RECT 4.755000  0.350000 5.085000 1.010000 ;
      RECT 4.860000  1.820000 5.110000 1.950000 ;
      RECT 4.860000  2.120000 5.110000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
  END
END sky130_fd_sc_hs__a2bb2oi_2
MACRO sky130_fd_sc_hs__a2bb2oi_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.470000 2.275000 1.800000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.420000 0.455000 1.770000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.735000 1.350000 8.515000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.350000 6.115000 1.780000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.500800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.270000 0.350000 2.520000 0.790000 ;
        RECT 2.270000 0.790000 6.150000 0.960000 ;
        RECT 3.185000 1.720000 4.255000 1.890000 ;
        RECT 3.185000 1.890000 3.355000 2.735000 ;
        RECT 3.210000 0.350000 3.380000 0.790000 ;
        RECT 3.965000 0.960000 6.150000 1.130000 ;
        RECT 3.965000 1.130000 4.255000 1.720000 ;
        RECT 4.085000 1.890000 4.255000 2.735000 ;
        RECT 4.960000 0.770000 6.150000 0.790000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
      RECT 0.000000  3.245000 8.640000 3.415000 ;
      RECT 0.105000  1.940000 0.435000 2.905000 ;
      RECT 0.105000  2.905000 1.255000 3.075000 ;
      RECT 0.635000  1.130000 3.585000 1.300000 ;
      RECT 0.635000  1.300000 0.885000 2.735000 ;
      RECT 0.940000  0.085000 1.270000 0.960000 ;
      RECT 1.085000  1.940000 1.255000 1.970000 ;
      RECT 1.085000  1.970000 2.235000 2.140000 ;
      RECT 1.085000  2.140000 1.255000 2.905000 ;
      RECT 1.450000  0.350000 1.620000 1.130000 ;
      RECT 1.455000  2.310000 1.705000 3.245000 ;
      RECT 1.800000  0.085000 2.090000 0.885000 ;
      RECT 1.905000  2.140000 2.235000 2.980000 ;
      RECT 2.575000  1.300000 3.585000 1.550000 ;
      RECT 2.655000  1.820000 2.985000 2.905000 ;
      RECT 2.655000  2.905000 4.785000 3.075000 ;
      RECT 2.700000  0.085000 3.030000 0.620000 ;
      RECT 3.555000  2.060000 3.885000 2.905000 ;
      RECT 3.560000  0.085000 3.890000 0.620000 ;
      RECT 4.455000  1.950000 8.385000 2.120000 ;
      RECT 4.455000  2.120000 4.785000 2.905000 ;
      RECT 4.530000  0.350000 6.500000 0.600000 ;
      RECT 4.985000  2.290000 5.155000 3.245000 ;
      RECT 5.355000  2.120000 5.685000 2.980000 ;
      RECT 5.885000  2.290000 6.135000 3.245000 ;
      RECT 6.330000  0.600000 6.500000 1.010000 ;
      RECT 6.330000  1.010000 8.300000 1.180000 ;
      RECT 6.335000  1.820000 6.505000 1.950000 ;
      RECT 6.335000  2.120000 6.505000 2.980000 ;
      RECT 6.680000  0.085000 6.930000 0.840000 ;
      RECT 6.705000  2.290000 6.955000 3.245000 ;
      RECT 7.110000  0.350000 7.360000 1.010000 ;
      RECT 7.155000  2.120000 7.485000 2.980000 ;
      RECT 7.540000  0.085000 7.790000 0.840000 ;
      RECT 7.685000  2.290000 7.855000 3.245000 ;
      RECT 7.970000  0.350000 8.300000 1.010000 ;
      RECT 8.055000  2.120000 8.385000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
  END
END sky130_fd_sc_hs__a2bb2oi_4
MACRO sky130_fd_sc_hs__a311o_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 0.440000 2.335000 0.670000 ;
        RECT 2.005000 0.255000 2.335000 0.440000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.450000 1.905000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.115000 1.450000 1.365000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 0.255000 2.875000 0.505000 ;
        RECT 2.525000 0.505000 2.725000 0.670000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.385000 0.255000 3.715000 0.670000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.504100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.010000 0.605000 1.180000 ;
        RECT 0.125000 1.180000 0.295000 1.850000 ;
        RECT 0.125000 1.850000 0.475000 2.980000 ;
        RECT 0.355000 0.480000 0.605000 1.010000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.480000  1.350000 0.945000 1.680000 ;
      RECT 0.645000  1.950000 1.105000 3.245000 ;
      RECT 0.775000  1.110000 2.570000 1.280000 ;
      RECT 0.775000  1.280000 0.945000 1.350000 ;
      RECT 0.785000  0.085000 1.115000 0.940000 ;
      RECT 1.275000  1.950000 2.595000 2.120000 ;
      RECT 1.275000  2.120000 1.605000 2.980000 ;
      RECT 1.805000  2.290000 2.095000 3.245000 ;
      RECT 2.240000  0.840000 2.570000 1.110000 ;
      RECT 2.240000  1.280000 2.570000 1.445000 ;
      RECT 2.240000  1.445000 3.575000 1.615000 ;
      RECT 2.265000  1.940000 2.595000 1.950000 ;
      RECT 2.265000  2.120000 2.595000 2.980000 ;
      RECT 2.750000  0.855000 3.075000 1.185000 ;
      RECT 2.895000  0.675000 3.215000 0.845000 ;
      RECT 2.895000  0.845000 3.075000 0.855000 ;
      RECT 3.045000  0.085000 3.215000 0.675000 ;
      RECT 3.105000  1.940000 3.575000 2.980000 ;
      RECT 3.245000  1.015000 3.575000 1.445000 ;
      RECT 3.245000  1.615000 3.575000 1.940000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__a311o_1
MACRO sky130_fd_sc_hs__a311o_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505000 1.450000 2.835000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965000 1.450000 2.295000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505000 1.260000 1.795000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.260000 3.715000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.885000 1.440000 4.215000 1.780000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.550000 0.995000 2.060000 ;
        RECT 0.730000 0.350000 1.060000 0.750000 ;
        RECT 0.730000 0.750000 0.995000 1.550000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.105000  1.350000 0.435000 2.230000 ;
      RECT 0.105000  2.230000 1.335000 2.400000 ;
      RECT 0.215000  2.570000 0.545000 3.245000 ;
      RECT 0.300000  0.085000 0.550000 1.130000 ;
      RECT 1.115000  2.570000 1.445000 3.245000 ;
      RECT 1.165000  0.920000 4.040000 1.090000 ;
      RECT 1.165000  1.090000 1.335000 1.950000 ;
      RECT 1.165000  1.950000 4.035000 2.120000 ;
      RECT 1.165000  2.120000 1.335000 2.230000 ;
      RECT 1.230000  0.085000 1.630000 0.750000 ;
      RECT 1.635000  2.290000 3.165000 2.570000 ;
      RECT 1.635000  2.570000 1.965000 2.980000 ;
      RECT 2.135000  2.740000 2.665000 3.245000 ;
      RECT 2.630000  0.350000 3.000000 0.920000 ;
      RECT 2.835000  2.570000 3.165000 2.980000 ;
      RECT 3.170000  0.085000 3.540000 0.750000 ;
      RECT 3.705000  2.120000 4.035000 2.980000 ;
      RECT 3.710000  0.350000 4.040000 0.920000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__a311o_2
MACRO sky130_fd_sc_hs__a311o_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885000 1.450000 7.075000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.245000 1.450000 7.575000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925000 1.420000 5.295000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.535000 1.470000 1.865000 1.800000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.495000 1.470000 0.825000 1.800000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  1.086400 ;
    ANTENNAPARTIALMETALSIDEAREA  1.869000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.095000 0.810000 0.385000 0.855000 ;
        RECT 0.095000 0.855000 2.785000 0.995000 ;
        RECT 0.095000 0.995000 0.385000 1.040000 ;
        RECT 2.495000 0.810000 2.785000 0.855000 ;
        RECT 2.495000 0.995000 2.785000 1.040000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.680000 0.085000 ;
      RECT 0.000000  3.245000 7.680000 3.415000 ;
      RECT 0.125000  0.810000 0.355000 1.040000 ;
      RECT 0.125000  1.040000 0.295000 2.360000 ;
      RECT 0.125000  2.360000 1.505000 2.530000 ;
      RECT 0.305000  2.700000 1.535000 2.905000 ;
      RECT 0.305000  2.905000 2.435000 2.980000 ;
      RECT 0.395000  0.085000 0.725000 0.640000 ;
      RECT 0.755000  2.020000 1.165000 2.190000 ;
      RECT 0.905000  0.390000 1.085000 1.130000 ;
      RECT 0.905000  1.130000 2.325000 1.300000 ;
      RECT 0.995000  1.300000 1.165000 2.020000 ;
      RECT 1.205000  2.980000 2.435000 3.075000 ;
      RECT 1.255000  0.085000 1.585000 0.960000 ;
      RECT 1.335000  1.970000 4.305000 2.140000 ;
      RECT 1.335000  2.140000 1.505000 2.360000 ;
      RECT 1.735000  2.310000 1.905000 2.320000 ;
      RECT 1.735000  2.320000 6.090000 2.460000 ;
      RECT 1.735000  2.460000 5.270000 2.490000 ;
      RECT 1.735000  2.490000 1.905000 2.735000 ;
      RECT 1.755000  0.390000 1.935000 1.130000 ;
      RECT 2.055000  1.300000 2.325000 1.320000 ;
      RECT 2.055000  1.320000 3.905000 1.480000 ;
      RECT 2.055000  1.480000 4.645000 1.650000 ;
      RECT 2.105000  2.660000 2.435000 2.905000 ;
      RECT 2.115000  0.085000 2.365000 0.960000 ;
      RECT 2.525000  1.820000 4.305000 1.970000 ;
      RECT 2.525000  2.140000 4.305000 2.150000 ;
      RECT 2.535000  0.390000 2.920000 0.980000 ;
      RECT 2.535000  0.980000 3.745000 1.150000 ;
      RECT 2.625000  2.660000 2.955000 3.245000 ;
      RECT 3.100000  0.085000 3.315000 0.810000 ;
      RECT 3.495000  0.405000 3.745000 0.980000 ;
      RECT 3.525000  2.660000 3.855000 3.245000 ;
      RECT 3.925000  0.085000 4.175000 0.935000 ;
      RECT 3.925000  0.935000 5.175000 1.150000 ;
      RECT 4.175000  1.150000 5.175000 1.185000 ;
      RECT 4.415000  0.505000 4.745000 0.595000 ;
      RECT 4.415000  0.595000 7.105000 0.765000 ;
      RECT 4.425000  2.660000 4.755000 3.245000 ;
      RECT 4.475000  1.650000 4.645000 1.950000 ;
      RECT 4.475000  1.950000 5.715000 2.120000 ;
      RECT 4.940000  2.290000 6.090000 2.320000 ;
      RECT 4.940000  2.490000 5.270000 2.980000 ;
      RECT 5.365000  0.255000 7.535000 0.425000 ;
      RECT 5.470000  2.630000 5.720000 3.245000 ;
      RECT 5.545000  0.935000 6.105000 1.265000 ;
      RECT 5.545000  1.265000 5.715000 1.950000 ;
      RECT 5.920000  1.950000 7.020000 2.120000 ;
      RECT 5.920000  2.120000 6.090000 2.290000 ;
      RECT 5.920000  2.460000 6.090000 2.980000 ;
      RECT 6.285000  0.985000 7.535000 1.245000 ;
      RECT 6.290000  2.290000 6.650000 3.245000 ;
      RECT 6.775000  0.765000 7.105000 0.815000 ;
      RECT 6.850000  2.120000 7.020000 2.980000 ;
      RECT 7.220000  1.950000 7.550000 3.245000 ;
      RECT 7.285000  0.425000 7.535000 0.985000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  0.840000 0.325000 1.010000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  0.840000 2.725000 1.010000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
  END
END sky130_fd_sc_hs__a311o_4
MACRO sky130_fd_sc_hs__a311oi_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.545000 1.350000 1.875000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.350000 1.335000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 0.495000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.350000 2.755000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925000 1.350000 3.255000 1.780000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.792700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.665000 1.010000 3.080000 1.180000 ;
        RECT 0.665000 1.180000 0.835000 1.950000 ;
        RECT 0.665000 1.950000 3.105000 2.120000 ;
        RECT 1.085000 0.350000 2.040000 1.010000 ;
        RECT 2.750000 0.350000 3.080000 1.010000 ;
        RECT 2.775000 2.120000 3.105000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.315000  2.290000 0.565000 3.245000 ;
      RECT 0.340000  0.085000 0.670000 0.840000 ;
      RECT 0.765000  2.290000 2.175000 2.460000 ;
      RECT 0.765000  2.460000 1.095000 2.980000 ;
      RECT 1.265000  2.630000 1.675000 3.245000 ;
      RECT 1.845000  2.460000 2.175000 2.980000 ;
      RECT 2.210000  0.085000 2.580000 0.840000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__a311oi_1
MACRO sky130_fd_sc_hs__a311oi_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.300000 1.350000 3.235000 1.550000 ;
        RECT 2.870000 1.550000 3.235000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.180000 1.315000 1.220000 ;
        RECT 1.085000 1.220000 2.090000 1.550000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.470000 1.220000 0.835000 1.550000 ;
        RECT 0.605000 1.180000 0.835000 1.220000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.350000 4.675000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.845000 1.350000 5.175000 1.780000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.935400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555000 0.850000 3.745000 1.010000 ;
        RECT 2.555000 1.010000 5.635000 1.180000 ;
        RECT 3.495000 0.350000 3.745000 0.850000 ;
        RECT 4.685000 0.350000 5.635000 1.010000 ;
        RECT 4.850000 1.950000 5.635000 2.120000 ;
        RECT 4.850000 2.120000 5.020000 2.735000 ;
        RECT 5.405000 1.180000 5.635000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.170000  1.820000 0.420000 3.245000 ;
      RECT 0.185000  0.350000 0.435000 0.840000 ;
      RECT 0.185000  0.840000 2.235000 1.010000 ;
      RECT 0.185000  1.010000 0.435000 1.050000 ;
      RECT 0.615000  0.085000 0.945000 0.670000 ;
      RECT 0.620000  1.720000 2.700000 1.890000 ;
      RECT 0.620000  1.890000 0.950000 2.980000 ;
      RECT 1.125000  0.330000 1.295000 0.770000 ;
      RECT 1.125000  0.770000 2.235000 0.840000 ;
      RECT 1.150000  2.060000 1.320000 3.245000 ;
      RECT 1.475000  0.350000 3.315000 0.600000 ;
      RECT 1.520000  1.890000 1.850000 2.980000 ;
      RECT 1.905000  1.010000 2.235000 1.050000 ;
      RECT 2.050000  2.060000 2.330000 3.245000 ;
      RECT 2.530000  1.890000 2.700000 1.950000 ;
      RECT 2.530000  1.950000 4.120000 2.120000 ;
      RECT 2.530000  2.120000 2.700000 2.980000 ;
      RECT 2.900000  2.290000 3.230000 3.245000 ;
      RECT 2.985000  0.600000 3.315000 0.680000 ;
      RECT 3.420000  2.290000 3.755000 2.905000 ;
      RECT 3.420000  2.905000 5.550000 3.075000 ;
      RECT 3.915000  0.085000 4.515000 0.840000 ;
      RECT 3.925000  2.120000 4.120000 2.735000 ;
      RECT 4.320000  1.950000 4.650000 2.905000 ;
      RECT 5.220000  2.290000 5.550000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_hs__a311oi_2
MACRO sky130_fd_sc_hs__a311oi_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.635000 1.350000 6.115000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.350000 3.715000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525000 1.350000 1.875000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.775000 1.180000 7.555000 1.320000 ;
        RECT 6.775000 1.320000 7.785000 1.650000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.065000 1.220000 9.075000 1.550000 ;
        RECT 8.285000 1.180000 9.075000 1.220000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.700600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.330000 0.770000 4.660000 0.850000 ;
        RECT 4.330000 0.850000 9.425000 1.010000 ;
        RECT 4.330000 1.010000 6.380000 1.130000 ;
        RECT 6.130000 0.350000 6.380000 0.840000 ;
        RECT 6.130000 0.840000 9.425000 0.850000 ;
        RECT 7.760000 0.350000 8.010000 0.840000 ;
        RECT 7.760000 1.010000 8.010000 1.050000 ;
        RECT 8.355000 1.720000 9.425000 1.890000 ;
        RECT 8.355000 1.890000 8.525000 2.735000 ;
        RECT 8.700000 0.350000 9.955000 0.670000 ;
        RECT 8.700000 0.670000 9.425000 0.840000 ;
        RECT 9.255000 1.010000 9.425000 1.720000 ;
        RECT 9.255000 1.890000 9.425000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.105000  1.820000  0.355000 3.245000 ;
      RECT 0.150000  0.350000  0.400000 1.010000 ;
      RECT 0.150000  1.010000  3.920000 1.180000 ;
      RECT 0.555000  1.950000  7.655000 2.120000 ;
      RECT 0.555000  2.120000  0.805000 2.980000 ;
      RECT 0.580000  0.085000  0.830000 0.840000 ;
      RECT 1.005000  2.290000  1.335000 3.245000 ;
      RECT 1.010000  0.350000  1.260000 1.010000 ;
      RECT 1.440000  0.085000  1.770000 0.840000 ;
      RECT 1.535000  2.120000  1.705000 2.980000 ;
      RECT 1.905000  2.290000  2.235000 3.245000 ;
      RECT 1.950000  0.350000  2.120000 0.975000 ;
      RECT 1.950000  0.975000  3.920000 1.010000 ;
      RECT 2.300000  0.350000  5.950000 0.600000 ;
      RECT 2.300000  0.600000  2.560000 0.680000 ;
      RECT 2.435000  2.120000  2.605000 2.980000 ;
      RECT 2.730000  0.770000  3.060000 0.975000 ;
      RECT 2.805000  2.290000  3.135000 3.245000 ;
      RECT 3.230000  0.600000  3.420000 0.680000 ;
      RECT 3.335000  2.120000  3.505000 2.980000 ;
      RECT 3.590000  0.770000  3.920000 0.975000 ;
      RECT 3.705000  2.290000  4.035000 3.245000 ;
      RECT 4.235000  1.820000  4.405000 1.950000 ;
      RECT 4.235000  2.120000  4.405000 2.980000 ;
      RECT 4.605000  2.290000  4.855000 3.245000 ;
      RECT 5.055000  2.120000  5.305000 2.980000 ;
      RECT 5.505000  2.290000  5.835000 3.245000 ;
      RECT 5.620000  0.600000  5.950000 0.680000 ;
      RECT 6.025000  2.320000  6.355000 2.905000 ;
      RECT 6.025000  2.905000  9.955000 3.075000 ;
      RECT 6.475000  1.820000  7.655000 1.950000 ;
      RECT 6.475000  2.120000  7.655000 2.150000 ;
      RECT 6.525000  2.150000  6.755000 2.735000 ;
      RECT 6.550000  0.085000  7.590000 0.670000 ;
      RECT 6.925000  2.320000  7.255000 2.905000 ;
      RECT 7.425000  2.150000  7.655000 2.735000 ;
      RECT 7.825000  1.820000  8.155000 2.905000 ;
      RECT 8.190000  0.085000  8.520000 0.670000 ;
      RECT 8.725000  2.060000  9.055000 2.905000 ;
      RECT 9.625000  1.820000  9.955000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
  END
END sky130_fd_sc_hs__a311oi_4
MACRO sky130_fd_sc_hs__a31o_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.490000 2.405000 1.800000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.535000 1.490000 1.865000 1.800000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.995000 1.490000 1.325000 1.800000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 0.255000 2.815000 0.640000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.504100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.480000 0.450000 1.180000 ;
        RECT 0.085000 1.180000 0.255000 1.850000 ;
        RECT 0.085000 1.850000 0.435000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.425000  1.350000 0.825000 1.680000 ;
      RECT 0.605000  1.970000 1.065000 3.245000 ;
      RECT 0.620000  0.085000 1.200000 0.980000 ;
      RECT 0.620000  1.150000 3.095000 1.320000 ;
      RECT 0.620000  1.320000 0.825000 1.350000 ;
      RECT 1.235000  1.970000 2.645000 2.140000 ;
      RECT 1.235000  2.140000 1.565000 2.980000 ;
      RECT 1.735000  2.310000 2.145000 3.245000 ;
      RECT 2.280000  0.810000 2.610000 1.150000 ;
      RECT 2.315000  2.140000 2.645000 2.980000 ;
      RECT 2.790000  0.810000 3.155000 0.980000 ;
      RECT 2.845000  1.320000 3.095000 2.980000 ;
      RECT 2.985000  0.085000 3.155000 0.810000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__a31o_1
MACRO sky130_fd_sc_hs__a31o_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.665000 1.180000 3.235000 1.550000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.180000 2.425000 1.550000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 1.180000 1.855000 1.550000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405000 1.180000 3.735000 1.550000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.820000 0.920000 2.980000 ;
        RECT 0.615000 0.350000 0.890000 1.130000 ;
        RECT 0.615000 1.130000 0.785000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 1.130000 ;
      RECT 0.185000  1.820000 0.435000 3.245000 ;
      RECT 0.955000  1.300000 1.305000 1.630000 ;
      RECT 1.060000  0.085000 1.730000 0.600000 ;
      RECT 1.090000  2.060000 1.625000 3.245000 ;
      RECT 1.135000  0.840000 3.180000 1.010000 ;
      RECT 1.135000  1.010000 1.305000 1.300000 ;
      RECT 1.135000  1.630000 1.305000 1.720000 ;
      RECT 1.135000  1.720000 3.725000 1.890000 ;
      RECT 1.795000  2.060000 3.215000 2.230000 ;
      RECT 1.795000  2.230000 2.125000 2.860000 ;
      RECT 2.350000  2.400000 2.680000 3.245000 ;
      RECT 2.850000  0.350000 3.180000 0.840000 ;
      RECT 2.885000  2.230000 3.215000 2.860000 ;
      RECT 3.360000  0.085000 3.690000 1.010000 ;
      RECT 3.385000  1.890000 3.725000 2.860000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__a31o_2
MACRO sky130_fd_sc_hs__a31o_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.450000 4.675000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925000 1.450000 5.865000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.115000 1.450000 7.075000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.565000 1.470000 3.235000 1.800000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  1.138200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565000 1.550000 0.895000 1.720000 ;
        RECT 0.565000 1.720000 1.895000 1.890000 ;
        RECT 0.565000 1.890000 0.895000 2.980000 ;
        RECT 0.615000 0.350000 0.865000 0.830000 ;
        RECT 0.615000 0.830000 1.725000 1.000000 ;
        RECT 0.615000 1.000000 0.865000 1.550000 ;
        RECT 1.555000 0.330000 1.725000 0.830000 ;
        RECT 1.565000 1.890000 1.895000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.200000 0.085000 ;
      RECT 0.000000  3.245000 7.200000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 1.130000 ;
      RECT 0.115000  1.820000 0.365000 3.245000 ;
      RECT 1.045000  0.085000 1.375000 0.660000 ;
      RECT 1.065000  1.220000 4.750000 1.280000 ;
      RECT 1.065000  1.280000 3.590000 1.300000 ;
      RECT 1.065000  1.300000 2.335000 1.550000 ;
      RECT 1.065000  2.060000 1.395000 3.245000 ;
      RECT 1.895000  1.130000 4.750000 1.220000 ;
      RECT 1.930000  0.085000 2.260000 0.960000 ;
      RECT 2.065000  1.820000 2.395000 3.245000 ;
      RECT 2.490000  0.350000 2.740000 1.130000 ;
      RECT 2.625000  1.970000 2.955000 2.810000 ;
      RECT 2.625000  2.810000 4.075000 2.980000 ;
      RECT 2.920000  0.085000 3.250000 0.960000 ;
      RECT 3.125000  1.970000 3.575000 2.640000 ;
      RECT 3.405000  1.300000 3.575000 1.970000 ;
      RECT 3.420000  0.350000 3.750000 1.110000 ;
      RECT 3.420000  1.110000 4.750000 1.130000 ;
      RECT 3.745000  1.950000 7.085000 2.120000 ;
      RECT 3.745000  2.120000 4.075000 2.810000 ;
      RECT 3.920000  0.255000 5.740000 0.425000 ;
      RECT 3.920000  0.425000 4.250000 0.940000 ;
      RECT 4.245000  2.290000 4.575000 3.245000 ;
      RECT 4.420000  0.595000 4.750000 1.110000 ;
      RECT 4.745000  2.120000 5.075000 2.980000 ;
      RECT 4.980000  0.595000 5.230000 1.110000 ;
      RECT 4.980000  1.110000 7.030000 1.280000 ;
      RECT 5.245000  2.290000 5.575000 3.245000 ;
      RECT 5.410000  0.425000 5.740000 0.940000 ;
      RECT 5.755000  2.120000 6.085000 2.980000 ;
      RECT 5.920000  0.350000 6.090000 1.110000 ;
      RECT 6.255000  2.290000 6.585000 3.245000 ;
      RECT 6.270000  0.085000 6.600000 0.940000 ;
      RECT 6.755000  2.120000 7.085000 2.980000 ;
      RECT 6.780000  0.350000 7.030000 1.110000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
  END
END sky130_fd_sc_hs__a31o_4
MACRO sky130_fd_sc_hs__a31oi_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.880000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.535000 1.180000 1.865000 1.550000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965000 0.810000 1.315000 1.550000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 0.455000 1.550000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.180000 2.775000 1.550000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.641200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.625000 0.350000 2.060000 0.520000 ;
        RECT 0.625000 0.520000 0.795000 1.720000 ;
        RECT 0.625000 1.720000 2.755000 1.890000 ;
        RECT 1.730000 0.520000 2.060000 1.010000 ;
        RECT 2.255000 1.890000 2.755000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.880000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.880000 0.085000 ;
      RECT 0.000000  3.245000 2.880000 3.415000 ;
      RECT 0.125000  0.085000 0.455000 1.010000 ;
      RECT 0.125000  1.820000 0.455000 3.245000 ;
      RECT 0.665000  2.060000 2.085000 2.230000 ;
      RECT 0.665000  2.230000 0.995000 2.980000 ;
      RECT 1.205000  2.400000 1.535000 3.245000 ;
      RECT 1.755000  2.230000 2.085000 2.980000 ;
      RECT 2.230000  0.085000 2.560000 1.010000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
  END
END sky130_fd_sc_hs__a31oi_1
MACRO sky130_fd_sc_hs__a31oi_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.505000 1.430000 4.195000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.430000 1.545000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.090000 2.115000 1.260000 ;
        RECT 0.105000 1.260000 0.435000 1.550000 ;
        RECT 1.785000 1.260000 2.115000 1.550000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.325000 1.180000 2.995000 1.550000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.090800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.475000 1.720000 3.335000 1.890000 ;
        RECT 2.475000 1.890000 2.805000 2.735000 ;
        RECT 2.545000 0.255000 4.205000 0.425000 ;
        RECT 2.545000 0.425000 3.260000 0.580000 ;
        RECT 3.165000 1.090000 4.205000 1.260000 ;
        RECT 3.165000 1.260000 3.335000 1.720000 ;
        RECT 3.875000 0.425000 4.205000 1.090000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  0.085000 0.365000 0.920000 ;
      RECT 0.115000  1.820000 0.365000 1.950000 ;
      RECT 0.115000  1.950000 2.275000 2.120000 ;
      RECT 0.115000  2.120000 0.365000 2.980000 ;
      RECT 0.545000  0.255000 1.875000 0.425000 ;
      RECT 0.545000  0.425000 0.875000 0.920000 ;
      RECT 0.565000  2.290000 0.895000 3.245000 ;
      RECT 1.045000  0.595000 1.375000 0.750000 ;
      RECT 1.045000  0.750000 3.705000 0.920000 ;
      RECT 1.065000  2.120000 1.395000 2.980000 ;
      RECT 1.545000  0.425000 1.875000 0.580000 ;
      RECT 1.595000  2.290000 1.845000 3.245000 ;
      RECT 2.015000  2.120000 2.275000 2.905000 ;
      RECT 2.015000  2.905000 3.255000 3.075000 ;
      RECT 2.045000  0.085000 2.375000 0.580000 ;
      RECT 2.975000  2.060000 4.205000 2.230000 ;
      RECT 2.975000  2.230000 3.255000 2.905000 ;
      RECT 3.425000  2.400000 3.755000 3.245000 ;
      RECT 3.430000  0.670000 3.705000 0.750000 ;
      RECT 3.875000  1.950000 4.205000 2.060000 ;
      RECT 3.925000  2.230000 4.205000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__a31oi_2
MACRO sky130_fd_sc_hs__a31oi_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925000 1.350000 6.115000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.415000 1.350000 4.195000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.745000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365000 1.350000 8.515000 1.780000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.621350 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.350000 0.770000 4.685000 0.965000 ;
        RECT 4.350000 0.965000 5.840000 1.010000 ;
        RECT 4.350000 1.010000 8.525000 1.130000 ;
        RECT 4.445000 1.130000 8.525000 1.180000 ;
        RECT 4.445000 1.180000 4.690000 1.950000 ;
        RECT 4.445000 1.950000 8.075000 2.120000 ;
        RECT 5.510000 0.595000 5.840000 0.965000 ;
        RECT 6.510000 0.350000 6.840000 1.010000 ;
        RECT 6.845000 2.120000 7.175000 2.735000 ;
        RECT 7.745000 2.120000 8.075000 2.735000 ;
        RECT 8.195000 0.350000 8.525000 1.010000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
      RECT 0.000000  3.245000 8.640000 3.415000 ;
      RECT 0.115000  1.950000 4.195000 2.120000 ;
      RECT 0.115000  2.120000 0.395000 2.980000 ;
      RECT 0.130000  0.350000 0.380000 1.010000 ;
      RECT 0.130000  1.010000 4.120000 1.180000 ;
      RECT 0.560000  0.085000 0.890000 0.840000 ;
      RECT 0.565000  2.290000 0.895000 3.245000 ;
      RECT 1.065000  2.120000 1.295000 2.935000 ;
      RECT 1.070000  0.350000 1.240000 1.010000 ;
      RECT 1.420000  0.085000 1.750000 0.840000 ;
      RECT 1.465000  2.290000 1.795000 3.245000 ;
      RECT 1.915000  1.820000 2.245000 1.950000 ;
      RECT 1.920000  0.330000 2.170000 1.010000 ;
      RECT 1.965000  2.120000 3.195000 2.150000 ;
      RECT 1.965000  2.150000 2.195000 2.950000 ;
      RECT 2.350000  0.255000 6.340000 0.425000 ;
      RECT 2.350000  0.425000 2.655000 0.840000 ;
      RECT 2.365000  2.320000 2.695000 3.245000 ;
      RECT 2.825000  0.595000 3.120000 1.010000 ;
      RECT 2.865000  2.150000 3.195000 2.980000 ;
      RECT 3.290000  0.425000 3.620000 0.840000 ;
      RECT 3.365000  2.290000 3.695000 3.245000 ;
      RECT 3.790000  0.595000 4.120000 1.010000 ;
      RECT 3.865000  2.120000 4.195000 2.290000 ;
      RECT 3.865000  2.290000 6.675000 2.460000 ;
      RECT 3.865000  2.460000 4.195000 2.980000 ;
      RECT 4.365000  2.630000 4.695000 3.245000 ;
      RECT 4.865000  2.460000 5.675000 2.930000 ;
      RECT 4.935000  0.425000 5.265000 0.795000 ;
      RECT 5.845000  2.630000 6.175000 3.245000 ;
      RECT 6.010000  0.425000 6.340000 0.840000 ;
      RECT 6.345000  2.460000 6.675000 2.905000 ;
      RECT 6.345000  2.905000 8.525000 3.075000 ;
      RECT 7.010000  0.085000 8.025000 0.840000 ;
      RECT 7.375000  2.290000 7.575000 2.905000 ;
      RECT 8.255000  1.950000 8.525000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
  END
END sky130_fd_sc_hs__a31oi_4
MACRO sky130_fd_sc_hs__a32o_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.190000 2.375000 1.550000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505000 1.190000 1.835000 1.550000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965000 1.190000 1.315000 1.550000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.545000 1.190000 3.005000 1.550000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.290000 1.210000 3.715000 1.550000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.350000 0.445000 1.130000 ;
        RECT 0.085000 1.130000 0.255000 1.820000 ;
        RECT 0.085000 1.820000 0.455000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.425000  1.300000 0.795000 1.630000 ;
      RECT 0.625000  0.850000 2.880000 1.020000 ;
      RECT 0.625000  1.020000 0.795000 1.300000 ;
      RECT 0.625000  1.630000 0.795000 1.720000 ;
      RECT 0.625000  1.720000 3.225000 1.890000 ;
      RECT 0.625000  2.060000 1.015000 3.245000 ;
      RECT 0.650000  0.085000 1.050000 0.680000 ;
      RECT 1.205000  2.060000 2.725000 2.230000 ;
      RECT 1.205000  2.230000 1.535000 2.860000 ;
      RECT 1.800000  2.400000 2.130000 3.245000 ;
      RECT 2.200000  0.430000 2.880000 0.850000 ;
      RECT 2.395000  2.230000 2.725000 2.905000 ;
      RECT 2.395000  2.905000 3.725000 3.075000 ;
      RECT 2.895000  1.890000 3.225000 2.735000 ;
      RECT 3.370000  0.085000 3.700000 1.040000 ;
      RECT 3.395000  1.820000 3.725000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__a32o_1
MACRO sky130_fd_sc_hs__a32o_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.350000 2.915000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.015000 1.350000 2.345000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.445000 1.350000 1.775000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.155000 1.350000 3.715000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.885000 1.300000 4.215000 1.780000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.550600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565000 1.820000 0.935000 2.150000 ;
        RECT 0.615000 0.330000 0.935000 1.150000 ;
        RECT 0.725000 1.150000 0.935000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 1.130000 ;
      RECT 0.115000  2.660000 0.445000 3.245000 ;
      RECT 0.225000  1.320000 0.555000 1.650000 ;
      RECT 0.225000  1.650000 0.395000 2.320000 ;
      RECT 0.225000  2.320000 1.275000 2.490000 ;
      RECT 1.100000  2.660000 1.510000 3.245000 ;
      RECT 1.105000  1.010000 3.105000 1.180000 ;
      RECT 1.105000  1.180000 1.275000 1.950000 ;
      RECT 1.105000  1.950000 3.705000 2.120000 ;
      RECT 1.105000  2.120000 1.275000 2.320000 ;
      RECT 1.185000  0.085000 1.515000 0.840000 ;
      RECT 1.715000  2.290000 3.205000 2.460000 ;
      RECT 1.715000  2.460000 2.045000 2.860000 ;
      RECT 2.265000  2.630000 2.645000 3.245000 ;
      RECT 2.775000  0.350000 3.105000 1.010000 ;
      RECT 2.875000  2.460000 3.205000 2.905000 ;
      RECT 2.875000  2.905000 4.205000 3.075000 ;
      RECT 3.375000  2.120000 3.705000 2.735000 ;
      RECT 3.850000  0.085000 4.180000 1.130000 ;
      RECT 3.875000  1.950000 4.205000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__a32o_2
MACRO sky130_fd_sc_hs__a32o_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.635000 1.450000 6.115000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.440000 1.470000 5.350000 1.790000 ;
        RECT 5.180000 1.790000 5.350000 1.950000 ;
        RECT 5.180000 1.950000 6.595000 2.120000 ;
        RECT 6.425000 1.440000 6.825000 1.770000 ;
        RECT 6.425000 1.770000 6.595000 1.950000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.065000 1.450000 8.035000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.450000 3.715000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505000 1.450000 2.835000 1.780000 ;
        RECT 2.570000 0.255000 4.415000 0.425000 ;
        RECT 2.570000 0.425000 2.740000 1.450000 ;
        RECT 4.085000 0.425000 4.415000 0.585000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  1.097500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.930000 1.900000 1.180000 ;
        RECT 0.125000 1.180000 0.355000 1.480000 ;
        RECT 0.125000 1.480000 0.815000 1.650000 ;
        RECT 0.565000 1.650000 0.815000 1.850000 ;
        RECT 0.565000 1.850000 1.795000 2.020000 ;
        RECT 0.565000 2.020000 0.815000 2.980000 ;
        RECT 0.615000 0.410000 0.820000 0.930000 ;
        RECT 1.515000 2.020000 1.795000 3.000000 ;
        RECT 1.570000 0.430000 1.900000 0.930000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 0.760000 ;
      RECT 0.115000  1.820000 0.365000 3.245000 ;
      RECT 0.985000  1.350000 2.185000 1.680000 ;
      RECT 0.990000  0.085000 1.400000 0.760000 ;
      RECT 1.015000  2.190000 1.345000 3.245000 ;
      RECT 1.965000  2.290000 2.295000 3.245000 ;
      RECT 2.015000  1.680000 2.185000 1.950000 ;
      RECT 2.015000  1.950000 4.355000 2.120000 ;
      RECT 2.070000  0.085000 2.400000 1.180000 ;
      RECT 2.525000  2.290000 2.855000 2.905000 ;
      RECT 2.525000  2.905000 4.925000 3.075000 ;
      RECT 2.910000  0.595000 3.240000 0.755000 ;
      RECT 2.910000  0.755000 4.180000 0.925000 ;
      RECT 2.910000  0.925000 3.240000 1.210000 ;
      RECT 3.025000  2.120000 3.355000 2.735000 ;
      RECT 3.420000  1.095000 3.750000 1.110000 ;
      RECT 3.420000  1.110000 6.130000 1.280000 ;
      RECT 3.525000  2.290000 3.855000 2.905000 ;
      RECT 3.885000  1.280000 4.055000 1.950000 ;
      RECT 4.025000  2.120000 4.355000 2.735000 ;
      RECT 4.350000  0.755000 4.755000 0.940000 ;
      RECT 4.585000  0.085000 4.755000 0.755000 ;
      RECT 4.595000  1.960000 4.925000 2.290000 ;
      RECT 4.595000  2.290000 7.095000 2.460000 ;
      RECT 4.595000  2.460000 4.925000 2.905000 ;
      RECT 4.940000  0.255000 6.990000 0.425000 ;
      RECT 4.940000  0.425000 5.190000 0.940000 ;
      RECT 5.210000  2.630000 5.615000 3.245000 ;
      RECT 5.370000  0.595000 6.560000 0.765000 ;
      RECT 5.370000  0.765000 5.620000 0.940000 ;
      RECT 5.785000  2.460000 6.115000 2.900000 ;
      RECT 5.800000  0.935000 6.130000 1.110000 ;
      RECT 6.285000  2.630000 6.645000 3.245000 ;
      RECT 6.310000  0.765000 6.560000 1.270000 ;
      RECT 6.740000  0.425000 6.990000 1.100000 ;
      RECT 6.740000  1.100000 8.045000 1.270000 ;
      RECT 6.765000  1.950000 8.045000 2.120000 ;
      RECT 6.765000  2.120000 7.095000 2.290000 ;
      RECT 6.815000  2.460000 7.095000 3.000000 ;
      RECT 7.190000  0.085000 7.545000 0.920000 ;
      RECT 7.265000  2.290000 7.545000 3.245000 ;
      RECT 7.715000  0.590000 8.045000 1.100000 ;
      RECT 7.715000  2.120000 8.045000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_hs__a32o_4
MACRO sky130_fd_sc_hs__a32oi_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 1.180000 1.855000 1.550000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 0.440000 2.525000 1.550000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.765000 1.180000 3.235000 1.550000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955000 1.180000 1.315000 1.550000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 1.180000 0.445000 1.550000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.998800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.615000 0.350000 1.830000 1.010000 ;
        RECT 0.615000 1.010000 0.785000 1.720000 ;
        RECT 0.615000 1.720000 2.275000 1.890000 ;
        RECT 0.615000 1.890000 0.945000 2.735000 ;
        RECT 1.590000 1.890000 2.275000 2.150000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 1.010000 ;
      RECT 0.115000  1.820000 0.445000 2.905000 ;
      RECT 0.115000  2.905000 1.445000 3.075000 ;
      RECT 1.115000  2.060000 1.420000 2.320000 ;
      RECT 1.115000  2.320000 2.795000 2.490000 ;
      RECT 1.115000  2.490000 1.445000 2.905000 ;
      RECT 1.675000  2.660000 2.345000 3.245000 ;
      RECT 2.465000  1.820000 2.795000 2.320000 ;
      RECT 2.515000  2.490000 2.795000 2.980000 ;
      RECT 2.890000  0.085000 3.220000 1.010000 ;
      RECT 2.995000  1.820000 3.245000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__a32oi_1
MACRO sky130_fd_sc_hs__a32oi_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 1.180000 2.775000 1.550000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.350000 4.375000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.785000 1.180000 6.115000 1.550000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505000 1.180000 2.275000 1.550000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 1.090000 1.630000 ;
        RECT 0.125000 1.630000 0.355000 1.780000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.192800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.615000 1.800000 3.235000 1.890000 ;
        RECT 0.615000 1.890000 1.945000 1.970000 ;
        RECT 0.615000 1.970000 0.945000 2.735000 ;
        RECT 1.455000 0.595000 1.785000 0.840000 ;
        RECT 1.455000 0.840000 3.205000 1.010000 ;
        RECT 1.615000 1.720000 3.235000 1.800000 ;
        RECT 1.615000 1.970000 1.945000 2.735000 ;
        RECT 3.005000 1.010000 3.205000 1.235000 ;
        RECT 3.005000 1.235000 3.235000 1.720000 ;
        RECT 3.015000 0.595000 3.205000 0.840000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.240000 0.085000 ;
      RECT 0.000000  3.245000 6.240000 3.415000 ;
      RECT 0.115000  0.350000 0.365000 0.960000 ;
      RECT 0.115000  0.960000 1.275000 1.130000 ;
      RECT 0.115000  1.950000 0.445000 2.905000 ;
      RECT 0.115000  2.905000 2.400000 3.075000 ;
      RECT 0.545000  0.085000 0.875000 0.790000 ;
      RECT 1.105000  0.255000 2.285000 0.425000 ;
      RECT 1.105000  0.425000 1.275000 0.960000 ;
      RECT 1.115000  2.140000 1.445000 2.905000 ;
      RECT 1.955000  0.425000 2.285000 0.670000 ;
      RECT 2.115000  2.060000 4.875000 2.120000 ;
      RECT 2.115000  2.120000 3.735000 2.230000 ;
      RECT 2.115000  2.230000 2.400000 2.905000 ;
      RECT 2.515000  0.255000 4.705000 0.425000 ;
      RECT 2.515000  0.425000 2.845000 0.670000 ;
      RECT 2.570000  2.400000 3.280000 3.245000 ;
      RECT 3.375000  0.425000 3.705000 1.130000 ;
      RECT 3.405000  1.950000 4.875000 2.060000 ;
      RECT 3.450000  2.230000 3.735000 2.980000 ;
      RECT 3.875000  0.595000 4.205000 1.010000 ;
      RECT 3.875000  1.010000 5.615000 1.180000 ;
      RECT 3.905000  2.290000 4.250000 3.245000 ;
      RECT 4.375000  0.425000 4.705000 0.840000 ;
      RECT 4.420000  2.120000 4.875000 2.980000 ;
      RECT 4.545000  1.720000 5.875000 1.890000 ;
      RECT 4.545000  1.890000 4.875000 1.950000 ;
      RECT 4.935000  0.085000 5.185000 0.840000 ;
      RECT 5.045000  2.060000 5.375000 3.245000 ;
      RECT 5.365000  0.350000 5.615000 1.010000 ;
      RECT 5.545000  1.890000 5.875000 2.980000 ;
      RECT 5.795000  0.085000 6.125000 1.010000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
  END
END sky130_fd_sc_hs__a32oi_2
MACRO sky130_fd_sc_hs__a32oi_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.56000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.350000 5.805000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.735000 1.350000 8.515000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.765000 1.350000 10.435000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.350000 4.195000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.795000 1.780000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  2.387000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.615000 1.950000 6.350000 2.120000 ;
        RECT 0.615000 2.120000 0.945000 2.735000 ;
        RECT 1.515000 2.120000 1.845000 2.735000 ;
        RECT 2.400000 0.595000 2.730000 0.880000 ;
        RECT 2.400000 0.880000 3.660000 1.010000 ;
        RECT 2.400000 1.010000 6.350000 1.130000 ;
        RECT 2.400000 1.130000 5.150000 1.180000 ;
        RECT 2.515000 2.120000 2.845000 2.735000 ;
        RECT 3.515000 2.120000 3.845000 2.735000 ;
        RECT 4.820000 0.770000 6.350000 1.010000 ;
        RECT 6.180000 1.130000 6.350000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.560000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.560000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 10.560000 0.085000 ;
      RECT  0.000000  3.245000 10.560000 3.415000 ;
      RECT  0.115000  0.350000  0.445000 1.010000 ;
      RECT  0.115000  1.010000  2.220000 1.180000 ;
      RECT  0.115000  1.950000  0.445000 2.905000 ;
      RECT  0.115000  2.905000  4.345000 3.075000 ;
      RECT  0.615000  0.085000  0.945000 0.840000 ;
      RECT  1.125000  0.350000  1.295000 1.010000 ;
      RECT  1.145000  2.290000  1.315000 2.905000 ;
      RECT  1.475000  0.085000  1.805000 0.840000 ;
      RECT  2.015000  2.290000  2.345000 2.905000 ;
      RECT  2.050000  0.255000  4.090000 0.425000 ;
      RECT  2.050000  0.425000  2.220000 1.010000 ;
      RECT  2.900000  0.425000  3.230000 0.710000 ;
      RECT  3.015000  2.290000  3.345000 2.905000 ;
      RECT  3.760000  0.425000  4.090000 0.710000 ;
      RECT  4.015000  2.290000  7.435000 2.460000 ;
      RECT  4.015000  2.460000  4.345000 2.905000 ;
      RECT  4.320000  0.350000  8.165000 0.600000 ;
      RECT  4.320000  0.600000  4.650000 0.840000 ;
      RECT  4.605000  2.630000  4.935000 3.245000 ;
      RECT  5.105000  2.460000  5.435000 2.980000 ;
      RECT  5.605000  2.630000  5.935000 3.245000 ;
      RECT  6.105000  2.460000  6.435000 2.980000 ;
      RECT  6.540000  0.770000  6.870000 0.850000 ;
      RECT  6.540000  0.850000  7.735000 1.010000 ;
      RECT  6.540000  1.010000  9.935000 1.180000 ;
      RECT  6.605000  2.630000  6.935000 3.245000 ;
      RECT  7.105000  1.950000 10.440000 2.120000 ;
      RECT  7.105000  2.120000  7.435000 2.290000 ;
      RECT  7.105000  2.460000  7.435000 2.980000 ;
      RECT  7.605000  2.290000  7.935000 3.245000 ;
      RECT  7.835000  0.600000  8.165000 0.680000 ;
      RECT  8.105000  2.120000  8.435000 2.980000 ;
      RECT  8.395000  0.085000  8.725000 0.840000 ;
      RECT  8.605000  2.290000  8.935000 3.245000 ;
      RECT  8.905000  0.350000  9.075000 1.010000 ;
      RECT  9.105000  2.120000  9.435000 2.980000 ;
      RECT  9.255000  0.085000  9.585000 0.840000 ;
      RECT  9.605000  2.290000  9.935000 3.245000 ;
      RECT  9.765000  0.350000  9.935000 1.010000 ;
      RECT 10.110000  2.120000 10.440000 2.980000 ;
      RECT 10.115000  0.085000 10.445000 1.130000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
  END
END sky130_fd_sc_hs__a32oi_4
MACRO sky130_fd_sc_hs__a41o_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.025000 1.450000 2.355000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 0.440000 2.895000 1.550000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.135000 1.180000 3.715000 1.550000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.885000 1.180000 4.215000 1.550000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 1.450000 1.815000 1.780000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  1.040800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.290000 1.120000 0.940000 ;
        RECT 0.115000 0.940000 0.355000 1.820000 ;
        RECT 0.115000 1.820000 0.445000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.575000  1.110000 2.120000 1.280000 ;
      RECT 0.575000  1.280000 1.315000 1.550000 ;
      RECT 0.645000  1.820000 0.895000 3.245000 ;
      RECT 1.145000  1.550000 1.315000 1.950000 ;
      RECT 1.145000  1.950000 1.635000 2.980000 ;
      RECT 1.290000  0.085000 1.620000 0.940000 ;
      RECT 1.790000  0.350000 2.120000 1.110000 ;
      RECT 1.805000  1.950000 3.165000 2.120000 ;
      RECT 1.805000  2.120000 2.135000 2.980000 ;
      RECT 2.305000  2.290000 2.635000 3.245000 ;
      RECT 2.835000  1.720000 4.185000 1.890000 ;
      RECT 2.835000  1.890000 3.165000 1.950000 ;
      RECT 2.835000  2.120000 3.165000 2.980000 ;
      RECT 3.335000  2.060000 3.665000 3.245000 ;
      RECT 3.830000  0.085000 4.160000 1.010000 ;
      RECT 3.855000  1.890000 4.185000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__a41o_1
MACRO sky130_fd_sc_hs__a41o_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.025000 1.450000 2.355000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 0.440000 1.815000 1.550000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.845000 0.440000 1.315000 1.550000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 0.455000 1.550000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.450000 2.925000 1.780000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.639400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.385000 0.350000 3.715000 0.770000 ;
        RECT 3.385000 0.770000 4.185000 0.940000 ;
        RECT 3.855000 1.820000 4.185000 2.980000 ;
        RECT 4.015000 0.940000 4.185000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.115000  1.720000 1.445000 1.890000 ;
      RECT 0.115000  1.890000 0.445000 2.980000 ;
      RECT 0.150000  0.085000 0.480000 1.010000 ;
      RECT 0.615000  2.060000 0.945000 3.245000 ;
      RECT 1.115000  1.890000 1.445000 1.950000 ;
      RECT 1.115000  1.950000 2.625000 2.120000 ;
      RECT 1.115000  2.120000 1.445000 2.980000 ;
      RECT 1.615000  2.290000 2.125000 3.245000 ;
      RECT 2.230000  0.350000 2.560000 1.110000 ;
      RECT 2.230000  1.110000 3.845000 1.280000 ;
      RECT 2.295000  2.120000 2.625000 2.980000 ;
      RECT 2.790000  0.085000 3.120000 0.940000 ;
      RECT 2.795000  1.950000 3.265000 2.120000 ;
      RECT 2.795000  2.120000 3.125000 2.980000 ;
      RECT 3.095000  1.280000 3.845000 1.550000 ;
      RECT 3.095000  1.550000 3.265000 1.950000 ;
      RECT 3.355000  2.270000 3.685000 3.245000 ;
      RECT 3.885000  0.085000 4.685000 0.600000 ;
      RECT 4.355000  1.820000 4.685000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_hs__a41o_2
MACRO sky130_fd_sc_hs__a41o_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.522000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.450000 4.195000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.522000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.900000 1.450000 5.635000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.522000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885000 1.450000 7.075000 1.780000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.522000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.325000 1.450000 8.035000 1.780000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.522000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.450000 0.550000 1.780000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.550000 1.000000 3.305000 1.170000 ;
        RECT 2.075000 1.840000 3.305000 2.120000 ;
        RECT 2.555000 1.170000 3.305000 1.840000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.110000  0.085000 0.360000 1.250000 ;
      RECT 0.115000  1.950000 0.445000 2.905000 ;
      RECT 0.115000  2.905000 1.395000 3.075000 ;
      RECT 0.540000  0.470000 0.870000 0.660000 ;
      RECT 0.540000  0.660000 3.645000 0.830000 ;
      RECT 0.540000  0.830000 1.225000 1.250000 ;
      RECT 0.615000  1.950000 0.890000 2.735000 ;
      RECT 0.720000  1.250000 1.225000 1.340000 ;
      RECT 0.720000  1.340000 2.385000 1.670000 ;
      RECT 0.720000  1.670000 0.890000 1.950000 ;
      RECT 1.045000  0.085000 1.375000 0.490000 ;
      RECT 1.065000  1.940000 1.395000 2.290000 ;
      RECT 1.065000  2.290000 4.375000 2.460000 ;
      RECT 1.065000  2.460000 1.395000 2.905000 ;
      RECT 1.625000  2.630000 1.955000 3.245000 ;
      RECT 2.055000  0.085000 2.385000 0.490000 ;
      RECT 2.525000  2.630000 2.855000 3.245000 ;
      RECT 3.055000  0.085000 3.305000 0.490000 ;
      RECT 3.425000  2.650000 3.775000 3.245000 ;
      RECT 3.475000  0.255000 4.495000 0.425000 ;
      RECT 3.475000  0.425000 3.645000 0.660000 ;
      RECT 3.815000  0.700000 3.985000 0.770000 ;
      RECT 3.815000  0.770000 4.845000 1.150000 ;
      RECT 4.045000  1.950000 7.595000 2.120000 ;
      RECT 4.045000  2.120000 4.375000 2.290000 ;
      RECT 4.045000  2.460000 4.375000 2.980000 ;
      RECT 4.165000  0.425000 4.495000 0.600000 ;
      RECT 4.635000  2.290000 5.095000 3.245000 ;
      RECT 4.675000  0.330000 5.785000 0.600000 ;
      RECT 4.675000  0.600000 4.845000 0.770000 ;
      RECT 5.025000  0.770000 5.285000 1.110000 ;
      RECT 5.025000  1.110000 6.680000 1.280000 ;
      RECT 5.265000  2.120000 5.595000 2.980000 ;
      RECT 5.455000  0.600000 5.785000 0.940000 ;
      RECT 5.765000  2.290000 6.095000 3.245000 ;
      RECT 6.000000  0.255000 7.110000 0.425000 ;
      RECT 6.000000  0.425000 6.330000 0.940000 ;
      RECT 6.265000  2.120000 6.595000 2.980000 ;
      RECT 6.510000  0.595000 6.680000 1.110000 ;
      RECT 6.765000  2.290000 7.095000 3.245000 ;
      RECT 6.860000  0.425000 7.110000 1.110000 ;
      RECT 6.860000  1.110000 8.050000 1.280000 ;
      RECT 7.265000  2.120000 7.595000 2.980000 ;
      RECT 7.290000  0.085000 7.620000 0.940000 ;
      RECT 7.790000  0.350000 8.050000 1.110000 ;
      RECT 7.795000  1.950000 8.045000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_hs__a41o_4
MACRO sky130_fd_sc_hs__a41oi_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925000 1.300000 3.255000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.195000 1.350000 2.755000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.350000 1.955000 1.780000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.350000 1.335000 1.780000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.300000 0.435000 1.780000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.752200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.350000 0.445000 0.960000 ;
        RECT 0.115000 0.960000 3.220000 1.130000 ;
        RECT 0.115000 1.950000 0.835000 2.120000 ;
        RECT 0.115000 2.120000 0.445000 2.980000 ;
        RECT 0.605000 1.130000 0.835000 1.950000 ;
        RECT 2.890000 0.350000 3.220000 0.960000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.615000  0.085000 1.260000 0.680000 ;
      RECT 0.615000  2.290000 1.275000 2.460000 ;
      RECT 0.615000  2.460000 0.945000 2.980000 ;
      RECT 1.105000  1.950000 3.245000 2.290000 ;
      RECT 1.115000  2.630000 1.785000 3.245000 ;
      RECT 1.445000  2.460000 1.785000 2.630000 ;
      RECT 2.405000  2.460000 2.745000 3.245000 ;
      RECT 2.915000  2.290000 3.245000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__a41oi_1
MACRO sky130_fd_sc_hs__a41oi_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415000 1.430000 1.795000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.665000 1.300000 3.715000 1.630000 ;
        RECT 3.005000 1.630000 3.715000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.350000 4.675000 1.780000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925000 1.350000 5.635000 1.780000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.085000 1.780000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.810100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.615000 0.400000 0.945000 1.010000 ;
        RECT 0.615000 1.010000 1.935000 1.090000 ;
        RECT 0.615000 1.090000 2.275000 1.180000 ;
        RECT 0.615000 1.950000 2.135000 2.120000 ;
        RECT 0.615000 2.120000 0.945000 2.735000 ;
        RECT 1.685000 0.595000 1.935000 1.010000 ;
        RECT 1.685000 1.180000 2.275000 1.260000 ;
        RECT 1.965000 1.260000 2.275000 1.650000 ;
        RECT 1.965000 1.650000 2.135000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 1.180000 ;
      RECT 0.115000  1.950000 0.445000 2.905000 ;
      RECT 0.115000  2.905000 1.445000 3.075000 ;
      RECT 1.115000  2.290000 2.635000 2.460000 ;
      RECT 1.115000  2.460000 1.445000 2.905000 ;
      RECT 1.175000  0.255000 2.355000 0.425000 ;
      RECT 1.175000  0.425000 1.505000 0.840000 ;
      RECT 1.615000  2.650000 2.135000 3.245000 ;
      RECT 2.105000  0.425000 2.355000 0.750000 ;
      RECT 2.105000  0.750000 3.295000 0.920000 ;
      RECT 2.305000  1.820000 2.635000 1.950000 ;
      RECT 2.305000  1.950000 5.645000 2.120000 ;
      RECT 2.305000  2.120000 2.635000 2.290000 ;
      RECT 2.305000  2.460000 2.635000 2.980000 ;
      RECT 2.535000  0.330000 4.285000 0.580000 ;
      RECT 2.805000  2.290000 3.135000 3.245000 ;
      RECT 2.965000  0.920000 3.295000 1.080000 ;
      RECT 3.305000  2.120000 3.635000 2.980000 ;
      RECT 3.525000  0.850000 4.635000 1.010000 ;
      RECT 3.525000  1.010000 5.645000 1.130000 ;
      RECT 3.805000  2.290000 4.135000 3.245000 ;
      RECT 3.955000  0.580000 4.285000 0.680000 ;
      RECT 4.305000  2.120000 4.670000 3.000000 ;
      RECT 4.465000  0.350000 4.635000 0.850000 ;
      RECT 4.465000  1.130000 5.645000 1.180000 ;
      RECT 4.815000  0.085000 5.145000 0.840000 ;
      RECT 4.840000  2.290000 5.170000 3.245000 ;
      RECT 5.315000  0.350000 5.645000 1.010000 ;
      RECT 5.340000  2.120000 5.645000 3.000000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_hs__a41oi_2
MACRO sky130_fd_sc_hs__a41oi_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.285000 1.350000 3.295000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.320000 5.620000 1.650000 ;
        RECT 3.965000 1.650000 4.675000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885000 1.350000 8.035000 1.780000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.285000 1.350000 9.955000 1.780000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.430000 1.780000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.447600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.350000 0.875000 1.010000 ;
        RECT 0.545000 1.010000 2.435000 1.180000 ;
        RECT 0.615000 1.950000 3.715000 2.120000 ;
        RECT 0.615000 2.120000 0.945000 2.735000 ;
        RECT 1.645000 1.820000 2.105000 1.950000 ;
        RECT 1.645000 2.120000 1.815000 2.735000 ;
        RECT 1.815000 1.180000 2.105000 1.820000 ;
        RECT 2.105000 0.595000 2.435000 1.010000 ;
        RECT 3.305000 0.595000 3.635000 1.000000 ;
        RECT 3.465000 1.000000 3.635000 1.550000 ;
        RECT 3.465000 1.550000 3.715000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.115000  0.085000  0.365000 1.130000 ;
      RECT 0.115000  1.950000  0.445000 2.905000 ;
      RECT 0.115000  2.905000  2.345000 3.075000 ;
      RECT 1.045000  0.085000  1.375000 0.840000 ;
      RECT 1.115000  2.290000  1.445000 2.905000 ;
      RECT 1.605000  0.255000  5.925000 0.425000 ;
      RECT 1.605000  0.425000  1.935000 0.840000 ;
      RECT 2.015000  2.290000  4.300000 2.460000 ;
      RECT 2.015000  2.460000  2.345000 2.905000 ;
      RECT 2.515000  2.630000  2.845000 3.245000 ;
      RECT 2.605000  0.425000  3.135000 1.130000 ;
      RECT 3.015000  2.460000  3.345000 2.980000 ;
      RECT 3.545000  2.630000  3.795000 3.245000 ;
      RECT 3.805000  0.425000  5.925000 0.620000 ;
      RECT 3.805000  0.620000  4.135000 1.130000 ;
      RECT 3.970000  1.950000  9.960000 2.120000 ;
      RECT 3.970000  2.120000  4.300000 2.290000 ;
      RECT 3.970000  2.460000  4.300000 2.980000 ;
      RECT 4.305000  0.790000  7.775000 1.130000 ;
      RECT 4.500000  2.290000  4.750000 3.245000 ;
      RECT 4.930000  1.820000  5.260000 1.950000 ;
      RECT 4.930000  2.120000  5.260000 2.980000 ;
      RECT 5.460000  2.290000  5.710000 3.245000 ;
      RECT 5.880000  2.120000  6.210000 2.980000 ;
      RECT 6.155000  0.350000  8.125000 0.600000 ;
      RECT 6.155000  0.600000  6.485000 0.620000 ;
      RECT 6.410000  2.290000  6.660000 3.245000 ;
      RECT 6.830000  2.120000  7.160000 2.980000 ;
      RECT 7.360000  2.290000  7.610000 3.245000 ;
      RECT 7.445000  0.770000  7.775000 0.790000 ;
      RECT 7.780000  2.120000  8.110000 2.980000 ;
      RECT 7.955000  0.600000  8.125000 1.010000 ;
      RECT 7.955000  1.010000  9.965000 1.180000 ;
      RECT 8.280000  2.290000  8.530000 3.245000 ;
      RECT 8.305000  0.085000  8.635000 0.840000 ;
      RECT 8.730000  2.120000  9.060000 2.980000 ;
      RECT 8.815000  0.350000  8.985000 1.010000 ;
      RECT 9.165000  0.085000  9.495000 0.840000 ;
      RECT 9.260000  2.290000  9.430000 3.245000 ;
      RECT 9.630000  2.120000  9.960000 2.980000 ;
      RECT 9.715000  0.350000  9.965000 1.010000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
  END
END sky130_fd_sc_hs__a41oi_4
MACRO sky130_fd_sc_hs__and2_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.400000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.255000 0.835000 0.670000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.075000 1.180000 1.405000 1.680000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.840000 0.470000 2.315000 1.180000 ;
        RECT 1.920000 1.850000 2.315000 2.980000 ;
        RECT 2.145000 1.180000 2.315000 1.850000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.400000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.400000 0.085000 ;
      RECT 0.000000  3.245000 2.400000 3.415000 ;
      RECT 0.260000  0.840000 0.590000 1.850000 ;
      RECT 0.260000  1.850000 1.750000 2.020000 ;
      RECT 0.350000  2.190000 0.685000 3.245000 ;
      RECT 0.855000  2.020000 1.185000 3.000000 ;
      RECT 1.340000  0.085000 1.670000 1.010000 ;
      RECT 1.390000  2.190000 1.720000 3.245000 ;
      RECT 1.580000  1.350000 1.975000 1.680000 ;
      RECT 1.580000  1.680000 1.750000 1.850000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
  END
END sky130_fd_sc_hs__and2_1
MACRO sky130_fd_sc_hs__and2_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.400000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.300000 0.435000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.300000 1.085000 1.780000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 0.350000 1.795000 0.790000 ;
        RECT 1.595000 1.720000 2.010000 1.890000 ;
        RECT 1.595000 1.890000 1.845000 2.980000 ;
        RECT 1.625000 0.790000 1.795000 0.850000 ;
        RECT 1.625000 0.850000 2.010000 1.020000 ;
        RECT 1.840000 1.020000 2.010000 1.720000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.400000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.400000 0.085000 ;
      RECT 0.000000  3.245000 2.400000 3.415000 ;
      RECT 0.110000  1.950000 0.440000 3.245000 ;
      RECT 0.135000  0.350000 0.465000 0.960000 ;
      RECT 0.135000  0.960000 1.425000 1.130000 ;
      RECT 0.640000  1.950000 1.425000 2.120000 ;
      RECT 0.640000  2.120000 0.890000 2.980000 ;
      RECT 0.955000  0.085000 1.285000 0.790000 ;
      RECT 1.060000  2.290000 1.390000 3.245000 ;
      RECT 1.255000  1.130000 1.425000 1.220000 ;
      RECT 1.255000  1.220000 1.670000 1.550000 ;
      RECT 1.255000  1.550000 1.425000 1.950000 ;
      RECT 1.975000  0.085000 2.285000 0.680000 ;
      RECT 2.045000  2.060000 2.295000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
  END
END sky130_fd_sc_hs__and2_2
MACRO sky130_fd_sc_hs__and2_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.444000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925000 1.450000 3.255000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.444000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.255000 1.345000 2.755000 1.780000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  1.219800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.475000 0.795000 1.005000 ;
        RECT 0.545000 1.005000 1.725000 1.175000 ;
        RECT 0.545000 1.175000 0.795000 1.550000 ;
        RECT 0.545000 1.550000 0.835000 1.845000 ;
        RECT 0.545000 1.845000 1.715000 2.015000 ;
        RECT 0.545000 2.015000 0.815000 2.980000 ;
        RECT 1.465000 2.015000 1.715000 2.980000 ;
        RECT 1.475000 0.475000 1.725000 1.005000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  0.085000 0.365000 1.255000 ;
      RECT 0.115000  1.820000 0.365000 3.245000 ;
      RECT 0.975000  0.085000 1.305000 0.835000 ;
      RECT 1.005000  1.345000 2.055000 1.675000 ;
      RECT 1.015000  2.185000 1.265000 3.245000 ;
      RECT 1.885000  1.675000 2.055000 1.950000 ;
      RECT 1.885000  1.950000 3.670000 2.120000 ;
      RECT 1.935000  2.290000 2.265000 3.245000 ;
      RECT 1.985000  0.085000 2.315000 1.175000 ;
      RECT 2.470000  2.120000 2.800000 2.905000 ;
      RECT 2.495000  0.255000 3.675000 0.425000 ;
      RECT 2.495000  0.425000 2.825000 1.175000 ;
      RECT 2.970000  2.290000 3.300000 3.245000 ;
      RECT 2.995000  0.595000 3.325000 1.110000 ;
      RECT 2.995000  1.110000 3.670000 1.280000 ;
      RECT 3.500000  1.280000 3.670000 1.950000 ;
      RECT 3.500000  2.120000 3.670000 2.905000 ;
      RECT 3.505000  0.425000 3.675000 0.940000 ;
      RECT 3.870000  2.025000 4.200000 3.245000 ;
      RECT 3.875000  0.085000 4.205000 1.255000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__and2_4
MACRO sky130_fd_sc_hs__and2b_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 0.550000 2.150000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.350000 2.375000 1.780000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.770000 1.820000 3.255000 2.980000 ;
        RECT 2.915000 0.370000 3.255000 1.150000 ;
        RECT 3.085000 1.150000 3.255000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.115000  0.350000 0.445000 1.010000 ;
      RECT 0.115000  1.010000 1.140000 1.180000 ;
      RECT 0.115000  2.320000 1.165000 2.650000 ;
      RECT 0.615000  0.085000 0.945000 0.840000 ;
      RECT 0.810000  1.180000 1.140000 2.320000 ;
      RECT 1.310000  0.470000 1.640000 0.980000 ;
      RECT 1.310000  0.980000 2.745000 1.150000 ;
      RECT 1.365000  1.820000 1.535000 3.245000 ;
      RECT 1.705000  1.150000 1.875000 1.950000 ;
      RECT 1.705000  1.950000 2.065000 2.700000 ;
      RECT 2.130000  0.085000 2.745000 0.810000 ;
      RECT 2.270000  1.950000 2.600000 3.245000 ;
      RECT 2.575000  1.150000 2.745000 1.320000 ;
      RECT 2.575000  1.320000 2.915000 1.650000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__and2b_1
MACRO sky130_fd_sc_hs__and2b_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 0.550000 1.780000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.180000 2.525000 1.550000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.820000 1.515000 2.150000 ;
        RECT 1.115000 0.350000 1.445000 1.130000 ;
        RECT 1.115000 1.130000 1.285000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.115000  0.350000 0.445000 1.010000 ;
      RECT 0.115000  1.010000 0.890000 1.180000 ;
      RECT 0.115000  1.950000 0.890000 2.320000 ;
      RECT 0.115000  2.320000 3.135000 2.490000 ;
      RECT 0.115000  2.490000 0.445000 2.700000 ;
      RECT 0.615000  0.085000 0.945000 0.840000 ;
      RECT 0.650000  2.660000 0.980000 3.245000 ;
      RECT 0.720000  1.180000 0.890000 1.950000 ;
      RECT 1.455000  1.300000 1.855000 1.630000 ;
      RECT 1.615000  0.085000 2.400000 0.600000 ;
      RECT 1.635000  2.660000 2.260000 3.245000 ;
      RECT 1.685000  0.840000 3.220000 1.010000 ;
      RECT 1.685000  1.010000 1.855000 1.300000 ;
      RECT 1.685000  1.630000 1.855000 1.870000 ;
      RECT 1.685000  1.870000 2.795000 2.150000 ;
      RECT 2.765000  1.300000 3.135000 1.630000 ;
      RECT 2.890000  0.350000 3.220000 0.840000 ;
      RECT 2.890000  1.010000 3.220000 1.130000 ;
      RECT 2.915000  2.660000 3.245000 3.245000 ;
      RECT 2.965000  1.630000 3.135000 2.320000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__and2b_2
MACRO sky130_fd_sc_hs__and2b_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.450000 0.805000 1.780000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.444000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.975000 1.435000 1.305000 1.620000 ;
        RECT 0.975000 1.620000 2.585000 1.790000 ;
        RECT 2.045000 1.180000 2.585000 1.620000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  1.093800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.095000 0.350000 3.265000 0.980000 ;
        RECT 3.095000 0.980000 4.675000 1.150000 ;
        RECT 3.095000 1.820000 4.165000 1.990000 ;
        RECT 3.095000 1.990000 3.265000 2.980000 ;
        RECT 3.910000 0.350000 4.160000 0.980000 ;
        RECT 3.995000 1.480000 4.675000 1.650000 ;
        RECT 3.995000 1.650000 4.165000 1.820000 ;
        RECT 3.995000 1.990000 4.165000 2.980000 ;
        RECT 4.445000 1.150000 4.675000 1.480000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.085000  0.350000 0.540000 1.095000 ;
      RECT 0.085000  1.095000 1.845000 1.265000 ;
      RECT 0.085000  1.265000 0.255000 1.950000 ;
      RECT 0.085000  1.950000 0.355000 2.980000 ;
      RECT 0.555000  2.100000 0.885000 3.245000 ;
      RECT 0.710000  0.085000 1.040000 0.925000 ;
      RECT 1.075000  1.960000 2.925000 2.130000 ;
      RECT 1.075000  2.130000 1.405000 2.980000 ;
      RECT 1.210000  0.335000 2.400000 0.585000 ;
      RECT 1.210000  0.585000 1.470000 0.925000 ;
      RECT 1.515000  1.265000 1.845000 1.450000 ;
      RECT 1.605000  2.300000 1.855000 3.245000 ;
      RECT 1.640000  0.755000 2.925000 0.925000 ;
      RECT 2.045000  2.130000 2.375000 2.980000 ;
      RECT 2.565000  2.300000 2.895000 3.245000 ;
      RECT 2.570000  0.085000 2.900000 0.585000 ;
      RECT 2.755000  0.925000 2.925000 1.320000 ;
      RECT 2.755000  1.320000 3.825000 1.650000 ;
      RECT 2.755000  1.650000 2.925000 1.960000 ;
      RECT 3.445000  0.085000 3.695000 0.810000 ;
      RECT 3.465000  2.160000 3.795000 3.245000 ;
      RECT 4.340000  0.085000 4.670000 0.810000 ;
      RECT 4.365000  1.820000 4.695000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_hs__and2b_4
MACRO sky130_fd_sc_hs__and3_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.880000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.255000 1.315000 0.570000 ;
        RECT 1.085000 0.570000 1.315000 0.670000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.845000 1.180000 1.315000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 1.450000 1.815000 1.780000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.195000 0.480000 2.525000 1.010000 ;
        RECT 2.195000 1.010000 2.765000 1.180000 ;
        RECT 2.480000 1.850000 2.765000 2.980000 ;
        RECT 2.595000 1.180000 2.765000 1.850000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.880000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.880000 0.085000 ;
      RECT 0.000000  3.245000 2.880000 3.415000 ;
      RECT 0.115000  0.740000 0.480000 1.950000 ;
      RECT 0.115000  1.950000 2.240000 2.120000 ;
      RECT 0.115000  2.120000 0.445000 2.850000 ;
      RECT 0.615000  2.290000 0.945000 3.245000 ;
      RECT 1.115000  2.120000 1.400000 2.850000 ;
      RECT 1.570000  2.290000 2.310000 3.245000 ;
      RECT 1.695000  0.085000 2.025000 1.180000 ;
      RECT 2.070000  1.350000 2.400000 1.680000 ;
      RECT 2.070000  1.680000 2.240000 1.950000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
  END
END sky130_fd_sc_hs__and3_1
MACRO sky130_fd_sc_hs__and3_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.255000 1.315000 0.670000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.905000 1.180000 1.315000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 1.430000 1.815000 1.780000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.572800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.180000 0.390000 2.510000 0.810000 ;
        RECT 2.180000 0.810000 2.755000 1.170000 ;
        RECT 2.375000 1.840000 2.725000 2.980000 ;
        RECT 2.555000 1.170000 2.725000 1.840000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.185000  0.840000 0.540000 1.340000 ;
      RECT 0.185000  1.340000 0.515000 1.950000 ;
      RECT 0.185000  1.950000 2.205000 2.120000 ;
      RECT 0.185000  2.120000 0.515000 2.780000 ;
      RECT 0.685000  2.290000 1.015000 3.245000 ;
      RECT 1.205000  2.120000 1.535000 2.780000 ;
      RECT 1.680000  0.085000 2.010000 1.170000 ;
      RECT 1.875000  2.290000 2.205000 3.245000 ;
      RECT 2.035000  1.340000 2.385000 1.670000 ;
      RECT 2.035000  1.670000 2.205000 1.950000 ;
      RECT 2.680000  0.085000 3.245000 0.640000 ;
      RECT 2.895000  1.820000 3.225000 3.245000 ;
      RECT 2.925000  0.640000 3.245000 1.170000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__and3_2
MACRO sky130_fd_sc_hs__and3_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.444000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.615000 1.450000 5.285000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.444000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.325000 4.335000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.444000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.450000 3.230000 1.780000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.560000 0.350000 0.890000 0.960000 ;
        RECT 0.560000 0.960000 1.740000 1.130000 ;
        RECT 0.560000 1.130000 0.835000 1.800000 ;
        RECT 0.560000 1.800000 1.895000 1.970000 ;
        RECT 0.560000 1.970000 0.895000 2.980000 ;
        RECT 1.490000 0.350000 1.740000 0.960000 ;
        RECT 1.565000 1.970000 1.895000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.115000  1.820000 0.365000 3.245000 ;
      RECT 0.130000  0.085000 0.380000 1.130000 ;
      RECT 1.035000  1.300000 2.235000 1.630000 ;
      RECT 1.065000  2.140000 1.395000 3.245000 ;
      RECT 1.070000  0.085000 1.320000 0.790000 ;
      RECT 1.920000  0.085000 2.250000 1.030000 ;
      RECT 2.065000  1.630000 2.235000 1.950000 ;
      RECT 2.065000  1.950000 5.625000 2.120000 ;
      RECT 2.065000  2.290000 2.395000 3.245000 ;
      RECT 2.420000  0.350000 2.670000 0.985000 ;
      RECT 2.420000  0.985000 4.090000 1.155000 ;
      RECT 2.565000  2.120000 2.895000 2.980000 ;
      RECT 2.850000  0.085000 3.180000 0.815000 ;
      RECT 3.065000  2.290000 3.645000 3.245000 ;
      RECT 3.410000  0.255000 5.640000 0.425000 ;
      RECT 3.410000  0.425000 3.740000 0.815000 ;
      RECT 3.815000  2.120000 4.145000 2.980000 ;
      RECT 3.920000  0.595000 4.090000 0.985000 ;
      RECT 4.310000  0.425000 4.640000 1.030000 ;
      RECT 4.315000  2.290000 4.645000 3.245000 ;
      RECT 4.810000  0.595000 5.140000 1.110000 ;
      RECT 4.810000  1.110000 5.625000 1.280000 ;
      RECT 4.815000  2.120000 5.145000 2.980000 ;
      RECT 5.310000  0.425000 5.640000 0.940000 ;
      RECT 5.315000  2.290000 5.645000 3.245000 ;
      RECT 5.455000  1.280000 5.625000 1.950000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_hs__and3_4
MACRO sky130_fd_sc_hs__and3b_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.110000 0.570000 1.780000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.005000 1.390000 2.335000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.390000 2.875000 1.780000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.345000 1.820000 3.755000 2.980000 ;
        RECT 3.385000 0.350000 3.755000 1.130000 ;
        RECT 3.585000 1.130000 3.755000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 0.940000 ;
      RECT 0.115000  2.100000 0.445000 3.245000 ;
      RECT 0.615000  0.350000 0.945000 0.940000 ;
      RECT 0.615000  2.100000 0.945000 2.980000 ;
      RECT 0.775000  0.940000 0.945000 1.030000 ;
      RECT 0.775000  1.030000 1.140000 1.700000 ;
      RECT 0.775000  1.700000 0.945000 2.100000 ;
      RECT 1.310000  0.450000 1.640000 1.050000 ;
      RECT 1.310000  1.050000 3.215000 1.220000 ;
      RECT 1.310000  1.220000 1.640000 1.950000 ;
      RECT 1.310000  1.950000 2.640000 2.120000 ;
      RECT 1.310000  2.120000 1.640000 2.700000 ;
      RECT 1.810000  2.290000 2.140000 3.245000 ;
      RECT 2.310000  2.120000 2.640000 2.700000 ;
      RECT 2.625000  0.085000 3.215000 0.880000 ;
      RECT 2.845000  1.950000 3.175000 3.245000 ;
      RECT 3.045000  1.220000 3.215000 1.300000 ;
      RECT 3.045000  1.300000 3.415000 1.630000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__and3b_1
MACRO sky130_fd_sc_hs__and3b_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.260000 0.550000 1.930000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 0.440000 2.450000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.690000 1.350000 3.235000 1.780000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.560000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.385000 0.350000 3.715000 1.130000 ;
        RECT 3.410000 1.130000 3.715000 1.820000 ;
        RECT 3.410000 1.820000 3.755000 2.070000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  0.420000 0.375000 0.920000 ;
      RECT 0.115000  0.920000 1.230000 1.090000 ;
      RECT 0.115000  2.100000 1.070000 2.270000 ;
      RECT 0.115000  2.270000 0.400000 2.980000 ;
      RECT 0.545000  0.085000 0.875000 0.750000 ;
      RECT 0.570000  2.440000 0.900000 3.245000 ;
      RECT 0.900000  1.090000 1.230000 1.855000 ;
      RECT 0.900000  1.855000 1.070000 2.100000 ;
      RECT 1.400000  0.350000 1.755000 1.950000 ;
      RECT 1.400000  1.950000 2.750000 2.120000 ;
      RECT 1.400000  2.120000 1.730000 2.860000 ;
      RECT 1.900000  2.290000 2.230000 3.245000 ;
      RECT 2.420000  2.120000 2.750000 2.240000 ;
      RECT 2.420000  2.240000 4.215000 2.410000 ;
      RECT 2.420000  2.410000 2.750000 2.860000 ;
      RECT 2.815000  0.085000 3.145000 1.130000 ;
      RECT 2.960000  2.580000 3.290000 3.245000 ;
      RECT 3.875000  2.580000 4.205000 3.245000 ;
      RECT 3.885000  1.300000 4.215000 1.630000 ;
      RECT 3.895000  0.085000 4.145000 1.130000 ;
      RECT 4.045000  1.630000 4.215000 2.240000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__and3b_2
MACRO sky130_fd_sc_hs__and3b_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.505000 1.180000 0.835000 1.510000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.350000 2.755000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.350000 3.560000 1.780000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  1.138200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.570000 1.800000 6.595000 1.970000 ;
        RECT 4.570000 1.970000 4.900000 2.980000 ;
        RECT 4.965000 0.350000 5.215000 0.960000 ;
        RECT 4.965000 0.960000 6.105000 1.130000 ;
        RECT 5.570000 1.970000 5.900000 2.980000 ;
        RECT 5.925000 0.350000 6.105000 0.960000 ;
        RECT 5.935000 1.130000 6.105000 1.800000 ;
        RECT 6.365000 1.550000 6.595000 1.800000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.720000 0.085000 ;
      RECT 0.000000  3.245000 6.720000 3.415000 ;
      RECT 0.115000  0.350000 0.445000 1.010000 ;
      RECT 0.115000  1.010000 0.285000 1.680000 ;
      RECT 0.115000  1.680000 1.305000 1.850000 ;
      RECT 0.475000  1.850000 0.805000 2.860000 ;
      RECT 0.615000  0.085000 0.875000 1.010000 ;
      RECT 0.975000  2.020000 1.305000 3.245000 ;
      RECT 1.135000  1.320000 1.525000 1.650000 ;
      RECT 1.135000  1.650000 1.305000 1.680000 ;
      RECT 1.175000  0.255000 2.365000 0.425000 ;
      RECT 1.175000  0.425000 1.505000 1.150000 ;
      RECT 1.475000  1.820000 1.865000 1.950000 ;
      RECT 1.475000  1.950000 3.900000 2.120000 ;
      RECT 1.475000  2.120000 1.805000 2.860000 ;
      RECT 1.685000  0.595000 1.865000 1.150000 ;
      RECT 1.695000  1.150000 1.865000 1.820000 ;
      RECT 1.975000  2.290000 2.305000 3.245000 ;
      RECT 2.035000  0.425000 2.365000 0.470000 ;
      RECT 2.035000  0.470000 3.295000 0.720000 ;
      RECT 2.035000  0.720000 2.365000 1.150000 ;
      RECT 2.475000  2.120000 2.805000 2.860000 ;
      RECT 2.535000  0.890000 2.865000 1.010000 ;
      RECT 2.535000  1.010000 4.285000 1.180000 ;
      RECT 2.975000  2.290000 3.305000 3.245000 ;
      RECT 3.525000  0.085000 3.855000 0.840000 ;
      RECT 3.535000  2.120000 3.900000 2.860000 ;
      RECT 3.730000  1.460000 5.765000 1.630000 ;
      RECT 3.730000  1.630000 3.900000 1.950000 ;
      RECT 4.035000  0.450000 4.285000 1.010000 ;
      RECT 4.070000  1.820000 4.400000 3.245000 ;
      RECT 4.465000  0.085000 4.795000 1.130000 ;
      RECT 4.755000  1.300000 5.765000 1.460000 ;
      RECT 5.070000  2.140000 5.400000 3.245000 ;
      RECT 5.395000  0.085000 5.725000 0.790000 ;
      RECT 6.070000  2.140000 6.400000 3.245000 ;
      RECT 6.275000  0.085000 6.605000 1.130000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
  END
END sky130_fd_sc_hs__and3b_4
MACRO sky130_fd_sc_hs__and4_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.120000 0.815000 1.790000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985000 0.440000 1.315000 1.805000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 0.440000 1.855000 1.790000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.350000 2.395000 1.780000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.730000 0.350000 3.275000 1.130000 ;
        RECT 2.910000 1.820000 3.275000 2.980000 ;
        RECT 3.105000 1.130000 3.275000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.085000  0.355000 0.770000 0.950000 ;
      RECT 0.085000  0.950000 0.255000 1.975000 ;
      RECT 0.085000  1.975000 2.740000 2.130000 ;
      RECT 0.085000  2.130000 2.205000 2.145000 ;
      RECT 0.115000  2.315000 0.445000 3.245000 ;
      RECT 0.615000  2.145000 0.945000 2.980000 ;
      RECT 1.115000  2.315000 1.705000 3.245000 ;
      RECT 1.875000  1.960000 2.740000 1.975000 ;
      RECT 1.875000  2.145000 2.205000 2.980000 ;
      RECT 2.220000  0.085000 2.550000 1.030000 ;
      RECT 2.410000  2.300000 2.740000 3.245000 ;
      RECT 2.570000  1.320000 2.935000 1.650000 ;
      RECT 2.570000  1.650000 2.740000 1.960000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__and4_1
MACRO sky130_fd_sc_hs__and4_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 1.300000 0.445000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955000 0.440000 1.315000 1.550000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 0.440000 1.855000 1.550000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.180000 2.425000 1.550000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.790000 0.770000 3.235000 1.130000 ;
        RECT 2.835000 1.130000 3.235000 2.150000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.115000  1.950000 0.445000 3.245000 ;
      RECT 0.260000  0.350000 0.590000 0.960000 ;
      RECT 0.260000  0.960000 0.785000 1.130000 ;
      RECT 0.615000  1.130000 0.785000 1.720000 ;
      RECT 0.615000  1.720000 2.095000 1.890000 ;
      RECT 0.615000  1.890000 0.985000 2.980000 ;
      RECT 1.215000  2.060000 1.545000 3.245000 ;
      RECT 1.765000  1.890000 2.095000 2.320000 ;
      RECT 1.765000  2.320000 3.735000 2.490000 ;
      RECT 1.765000  2.490000 2.095000 2.980000 ;
      RECT 2.265000  0.085000 2.595000 1.010000 ;
      RECT 2.300000  2.660000 2.630000 3.245000 ;
      RECT 3.220000  0.085000 3.655000 0.600000 ;
      RECT 3.370000  2.660000 3.725000 3.245000 ;
      RECT 3.405000  0.600000 3.655000 1.080000 ;
      RECT 3.405000  1.300000 3.735000 2.320000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__and4_2
MACRO sky130_fd_sc_hs__and4_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.060000 1.450000 1.390000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.450000 0.550000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.980000 1.345000 4.365000 1.780000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.930000 1.470000 3.260000 1.800000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  1.164600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.830000 0.350000 5.080000 0.960000 ;
        RECT 4.830000 0.960000 6.595000 1.130000 ;
        RECT 4.875000 1.800000 6.105000 1.970000 ;
        RECT 4.875000 1.970000 5.205000 2.980000 ;
        RECT 5.760000 0.350000 6.090000 0.960000 ;
        RECT 5.855000 1.480000 6.595000 1.650000 ;
        RECT 5.855000 1.650000 6.105000 1.800000 ;
        RECT 5.855000 1.970000 6.105000 2.980000 ;
        RECT 6.365000 1.130000 6.595000 1.480000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.720000 0.085000 ;
      RECT 0.000000  3.245000 6.720000 3.415000 ;
      RECT 0.115000  1.950000 0.395000 3.245000 ;
      RECT 0.140000  0.315000 2.110000 0.485000 ;
      RECT 0.140000  0.485000 0.390000 1.255000 ;
      RECT 0.565000  1.950000 1.730000 2.240000 ;
      RECT 0.570000  0.655000 1.760000 0.835000 ;
      RECT 0.720000  1.005000 1.330000 1.255000 ;
      RECT 0.720000  1.255000 0.890000 1.950000 ;
      RECT 1.015000  2.410000 1.345000 3.245000 ;
      RECT 1.560000  1.600000 2.760000 1.770000 ;
      RECT 1.560000  1.770000 1.730000 1.950000 ;
      RECT 1.560000  2.240000 1.730000 2.980000 ;
      RECT 1.930000  1.940000 2.260000 3.245000 ;
      RECT 1.940000  0.485000 2.110000 1.130000 ;
      RECT 1.940000  1.130000 4.070000 1.175000 ;
      RECT 1.940000  1.175000 3.810000 1.300000 ;
      RECT 2.290000  0.575000 2.620000 0.790000 ;
      RECT 2.290000  0.790000 3.640000 0.825000 ;
      RECT 2.290000  0.825000 3.470000 0.960000 ;
      RECT 2.430000  1.770000 2.760000 1.970000 ;
      RECT 2.430000  1.970000 4.705000 2.120000 ;
      RECT 2.430000  2.120000 4.145000 2.140000 ;
      RECT 2.430000  2.140000 2.760000 2.980000 ;
      RECT 2.800000  0.085000 3.130000 0.620000 ;
      RECT 2.930000  2.310000 3.645000 3.245000 ;
      RECT 3.300000  0.575000 3.640000 0.790000 ;
      RECT 3.640000  0.995000 4.070000 1.130000 ;
      RECT 3.815000  1.950000 4.705000 1.970000 ;
      RECT 3.815000  2.140000 4.145000 2.980000 ;
      RECT 4.315000  2.290000 4.645000 3.245000 ;
      RECT 4.330000  0.085000 4.660000 1.130000 ;
      RECT 4.535000  1.300000 5.685000 1.630000 ;
      RECT 4.535000  1.630000 4.705000 1.950000 ;
      RECT 5.260000  0.085000 5.590000 0.790000 ;
      RECT 5.405000  2.140000 5.655000 3.245000 ;
      RECT 6.260000  0.085000 6.520000 0.680000 ;
      RECT 6.275000  1.820000 6.605000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
  END
END sky130_fd_sc_hs__and4_4
MACRO sky130_fd_sc_hs__and4b_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.190000 0.595000 1.860000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.550000 2.275000 1.960000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 0.255000 2.810000 0.670000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.985000 1.550000 3.315000 1.880000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.875000 0.480000 4.230000 1.180000 ;
        RECT 3.875000 1.850000 4.230000 2.980000 ;
        RECT 4.060000 1.180000 4.230000 1.850000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  0.350000 0.405000 0.850000 ;
      RECT 0.115000  0.850000 0.945000 1.020000 ;
      RECT 0.115000  2.030000 0.945000 2.200000 ;
      RECT 0.115000  2.200000 0.445000 2.980000 ;
      RECT 0.575000  0.085000 0.875000 0.680000 ;
      RECT 0.615000  2.370000 0.945000 3.245000 ;
      RECT 0.775000  1.020000 0.945000 1.550000 ;
      RECT 0.775000  1.550000 1.255000 1.880000 ;
      RECT 0.775000  1.880000 0.945000 2.030000 ;
      RECT 1.115000  2.130000 3.095000 2.350000 ;
      RECT 1.115000  2.350000 1.460000 2.460000 ;
      RECT 1.310000  0.600000 1.640000 1.210000 ;
      RECT 1.310000  1.210000 3.705000 1.350000 ;
      RECT 1.310000  1.350000 3.890000 1.380000 ;
      RECT 1.645000  2.535000 2.595000 3.245000 ;
      RECT 2.595000  1.380000 2.765000 2.100000 ;
      RECT 2.595000  2.100000 3.095000 2.130000 ;
      RECT 2.765000  2.350000 3.095000 2.980000 ;
      RECT 3.335000  2.100000 3.665000 3.245000 ;
      RECT 3.375000  0.085000 3.705000 1.040000 ;
      RECT 3.535000  1.380000 3.890000 1.680000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__and4b_1
MACRO sky130_fd_sc_hs__and4b_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.455000 1.780000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.350000 3.405000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505000 1.350000 2.835000 1.780000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965000 1.350000 2.295000 1.780000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055000 0.350000 1.385000 1.130000 ;
        RECT 1.055000 1.130000 1.225000 1.820000 ;
        RECT 1.055000 1.820000 1.440000 2.200000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  0.540000 0.445000 0.960000 ;
      RECT 0.115000  0.960000 0.795000 1.130000 ;
      RECT 0.115000  1.950000 0.795000 2.370000 ;
      RECT 0.115000  2.370000 3.985000 2.540000 ;
      RECT 0.115000  2.540000 0.445000 2.700000 ;
      RECT 0.625000  0.085000 0.875000 0.790000 ;
      RECT 0.625000  1.130000 0.795000 1.950000 ;
      RECT 0.650000  2.710000 0.980000 3.245000 ;
      RECT 1.395000  1.300000 1.780000 1.630000 ;
      RECT 1.555000  0.085000 2.165000 0.790000 ;
      RECT 1.610000  0.960000 4.070000 1.130000 ;
      RECT 1.610000  1.130000 1.780000 1.300000 ;
      RECT 1.610000  1.630000 1.780000 1.950000 ;
      RECT 1.610000  1.950000 3.645000 2.200000 ;
      RECT 1.645000  2.710000 1.975000 3.245000 ;
      RECT 2.740000  2.710000 3.070000 3.245000 ;
      RECT 3.615000  1.350000 3.985000 1.680000 ;
      RECT 3.740000  0.350000 4.070000 0.960000 ;
      RECT 3.815000  1.680000 3.985000 2.370000 ;
      RECT 3.850000  2.710000 4.205000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__and4b_2
MACRO sky130_fd_sc_hs__and4b_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.190000 0.835000 1.550000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.845000 1.470000 7.180000 1.800000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.915000 1.350000 3.245000 1.780000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.470000 5.155000 1.800000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  1.209600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 0.350000 1.470000 0.980000 ;
        RECT 1.085000 0.980000 2.540000 1.150000 ;
        RECT 1.085000 1.150000 1.315000 1.820000 ;
        RECT 1.085000 1.820000 2.405000 2.220000 ;
        RECT 2.210000 0.350000 2.540000 0.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.680000 0.085000 ;
      RECT 0.000000  3.245000 7.680000 3.415000 ;
      RECT 0.085000  0.450000 0.405000 1.020000 ;
      RECT 0.085000  1.020000 0.255000 1.820000 ;
      RECT 0.085000  1.820000 0.445000 2.390000 ;
      RECT 0.085000  2.390000 7.520000 2.560000 ;
      RECT 0.085000  2.560000 0.445000 2.860000 ;
      RECT 0.585000  0.085000 0.915000 1.020000 ;
      RECT 0.650000  2.730000 1.025000 3.245000 ;
      RECT 1.485000  1.320000 2.745000 1.650000 ;
      RECT 1.595000  2.730000 1.955000 3.245000 ;
      RECT 1.670000  0.085000 2.000000 0.810000 ;
      RECT 2.575000  1.650000 2.745000 1.950000 ;
      RECT 2.575000  1.950000 3.515000 1.970000 ;
      RECT 2.575000  1.970000 6.880000 2.220000 ;
      RECT 2.635000  2.730000 2.980000 3.245000 ;
      RECT 2.710000  0.085000 3.040000 1.130000 ;
      RECT 3.300000  0.605000 3.630000 1.130000 ;
      RECT 3.300000  1.130000 5.475000 1.180000 ;
      RECT 3.460000  1.180000 5.475000 1.300000 ;
      RECT 3.720000  2.730000 4.050000 3.245000 ;
      RECT 3.810000  0.630000 4.105000 0.790000 ;
      RECT 3.810000  0.790000 5.125000 0.960000 ;
      RECT 4.285000  0.085000 4.615000 0.620000 ;
      RECT 4.795000  0.605000 5.125000 0.790000 ;
      RECT 5.180000  2.730000 5.530000 3.245000 ;
      RECT 5.305000  0.255000 7.495000 0.425000 ;
      RECT 5.305000  0.425000 5.475000 1.130000 ;
      RECT 5.650000  1.940000 6.080000 1.970000 ;
      RECT 5.655000  0.595000 6.955000 0.765000 ;
      RECT 5.655000  0.765000 5.905000 0.960000 ;
      RECT 5.910000  1.130000 6.335000 1.300000 ;
      RECT 5.910000  1.300000 6.080000 1.940000 ;
      RECT 6.080000  0.935000 6.335000 1.130000 ;
      RECT 6.100000  2.730000 6.430000 3.245000 ;
      RECT 6.250000  1.470000 6.675000 1.800000 ;
      RECT 6.505000  1.130000 7.520000 1.300000 ;
      RECT 6.505000  1.300000 6.675000 1.470000 ;
      RECT 6.625000  0.765000 6.955000 0.935000 ;
      RECT 7.000000  2.730000 7.565000 3.245000 ;
      RECT 7.165000  0.425000 7.495000 0.960000 ;
      RECT 7.350000  1.300000 7.520000 2.390000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
  END
END sky130_fd_sc_hs__and4b_4
MACRO sky130_fd_sc_hs__and4bb_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.300000 0.400000 1.780000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.400000 1.300000 4.695000 1.780000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.015000 1.190000 3.345000 1.860000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.515000 1.190000 3.890000 1.860000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.692500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.910000 0.960000 1.270000 1.130000 ;
        RECT 0.910000 1.130000 1.080000 1.820000 ;
        RECT 0.910000 1.820000 1.565000 2.150000 ;
        RECT 1.080000 0.350000 1.270000 0.960000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.115000  0.350000 0.365000 0.960000 ;
      RECT 0.115000  0.960000 0.740000 1.130000 ;
      RECT 0.115000  1.950000 0.740000 2.320000 ;
      RECT 0.115000  2.320000 2.045000 2.490000 ;
      RECT 0.115000  2.490000 0.445000 2.700000 ;
      RECT 0.545000  0.085000 0.875000 0.790000 ;
      RECT 0.570000  1.130000 0.740000 1.950000 ;
      RECT 0.650000  2.660000 0.980000 3.245000 ;
      RECT 1.250000  1.300000 1.610000 1.630000 ;
      RECT 1.440000  0.860000 2.385000 1.030000 ;
      RECT 1.440000  1.030000 1.610000 1.300000 ;
      RECT 1.780000  1.290000 2.045000 2.320000 ;
      RECT 1.795000  2.660000 2.125000 3.245000 ;
      RECT 1.820000  0.350000 2.385000 0.860000 ;
      RECT 2.215000  1.030000 2.385000 2.030000 ;
      RECT 2.215000  2.030000 3.625000 2.200000 ;
      RECT 2.295000  2.200000 2.625000 2.980000 ;
      RECT 2.555000  0.850000 4.685000 1.020000 ;
      RECT 2.555000  1.020000 2.845000 1.790000 ;
      RECT 2.795000  2.370000 3.125000 3.245000 ;
      RECT 3.295000  2.200000 3.625000 2.980000 ;
      RECT 3.720000  0.085000 4.110000 0.680000 ;
      RECT 3.815000  2.290000 4.145000 3.245000 ;
      RECT 4.060000  1.020000 4.685000 1.030000 ;
      RECT 4.060000  1.030000 4.230000 1.950000 ;
      RECT 4.060000  1.950000 4.645000 2.120000 ;
      RECT 4.315000  2.120000 4.645000 2.980000 ;
      RECT 4.355000  0.440000 4.685000 0.850000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_hs__and4bb_1
MACRO sky130_fd_sc_hs__and4bb_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.450000 0.550000 1.780000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.825000 1.180000 5.155000 1.590000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.310000 1.420000 2.755000 1.780000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925000 1.420000 3.255000 1.780000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.815000 0.920000 4.195000 1.170000 ;
        RECT 3.835000 1.840000 4.195000 2.980000 ;
        RECT 4.025000 1.170000 4.195000 1.840000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.280000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.245000 5.280000 3.415000 ;
      RECT 0.115000  0.350000 0.365000 1.110000 ;
      RECT 0.115000  1.110000 0.935000 1.280000 ;
      RECT 0.210000  1.950000 0.935000 2.120000 ;
      RECT 0.210000  2.120000 0.540000 2.820000 ;
      RECT 0.545000  0.085000 0.875000 0.940000 ;
      RECT 0.765000  1.280000 0.935000 1.340000 ;
      RECT 0.765000  1.340000 1.260000 1.670000 ;
      RECT 0.765000  1.670000 0.935000 1.950000 ;
      RECT 0.780000  2.290000 1.110000 3.245000 ;
      RECT 1.105000  0.390000 1.600000 1.170000 ;
      RECT 1.430000  1.170000 1.600000 1.940000 ;
      RECT 1.430000  1.940000 1.760000 1.950000 ;
      RECT 1.430000  1.950000 3.665000 2.120000 ;
      RECT 1.430000  2.120000 1.760000 2.980000 ;
      RECT 1.770000  1.000000 3.645000 1.170000 ;
      RECT 1.770000  1.170000 2.100000 1.590000 ;
      RECT 2.065000  2.290000 2.395000 3.245000 ;
      RECT 2.610000  2.120000 2.940000 2.980000 ;
      RECT 2.975000  0.085000 3.305000 0.830000 ;
      RECT 3.200000  2.290000 3.530000 3.245000 ;
      RECT 3.475000  0.580000 5.165000 0.750000 ;
      RECT 3.475000  0.750000 3.645000 1.000000 ;
      RECT 3.495000  1.340000 3.855000 1.670000 ;
      RECT 3.495000  1.670000 3.665000 1.950000 ;
      RECT 4.325000  0.085000 4.655000 0.410000 ;
      RECT 4.365000  0.750000 4.535000 1.760000 ;
      RECT 4.365000  1.760000 5.165000 1.930000 ;
      RECT 4.365000  2.100000 4.615000 3.245000 ;
      RECT 4.820000  1.930000 5.165000 2.700000 ;
      RECT 4.835000  0.750000 5.165000 1.010000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
  END
END sky130_fd_sc_hs__and4bb_2
MACRO sky130_fd_sc_hs__and4bb_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.450000 1.335000 1.780000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.450000 0.835000 1.780000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.965000 1.450000 6.115000 1.780000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365000 1.350000 6.875000 1.780000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  1.116000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.240000 0.350000 7.570000 0.980000 ;
        RECT 7.240000 0.980000 8.995000 1.150000 ;
        RECT 7.405000 1.820000 8.995000 2.150000 ;
        RECT 7.405000 2.150000 7.575000 2.980000 ;
        RECT 8.240000 0.770000 8.995000 0.980000 ;
        RECT 8.765000 1.150000 8.995000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.120000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.120000 0.085000 ;
      RECT 0.000000  3.245000 9.120000 3.415000 ;
      RECT 0.115000  0.350000 0.365000 1.110000 ;
      RECT 0.115000  1.110000 1.870000 1.280000 ;
      RECT 0.115000  1.950000 1.675000 2.120000 ;
      RECT 0.115000  2.120000 0.445000 2.980000 ;
      RECT 0.545000  0.085000 0.875000 0.940000 ;
      RECT 0.615000  2.290000 0.945000 3.245000 ;
      RECT 1.045000  0.255000 1.690000 0.585000 ;
      RECT 1.045000  0.585000 1.530000 0.940000 ;
      RECT 1.115000  2.290000 2.260000 2.460000 ;
      RECT 1.115000  2.460000 1.445000 2.980000 ;
      RECT 1.505000  1.280000 1.675000 1.950000 ;
      RECT 1.700000  0.755000 2.030000 0.925000 ;
      RECT 1.700000  0.925000 1.870000 1.110000 ;
      RECT 1.860000  0.255000 3.605000 0.585000 ;
      RECT 1.860000  0.585000 2.030000 0.755000 ;
      RECT 1.890000  2.630000 2.225000 3.245000 ;
      RECT 1.930000  1.450000 2.260000 2.290000 ;
      RECT 2.040000  1.095000 2.370000 1.280000 ;
      RECT 2.200000  0.755000 3.220000 0.925000 ;
      RECT 2.200000  0.925000 2.370000 1.095000 ;
      RECT 2.430000  1.595000 4.795000 1.765000 ;
      RECT 2.430000  1.765000 2.760000 2.960000 ;
      RECT 2.540000  1.095000 2.870000 1.360000 ;
      RECT 2.540000  1.360000 2.760000 1.595000 ;
      RECT 2.965000  1.935000 3.295000 3.245000 ;
      RECT 3.050000  0.925000 3.220000 1.255000 ;
      RECT 3.050000  1.255000 4.160000 1.425000 ;
      RECT 3.400000  0.755000 5.220000 0.925000 ;
      RECT 3.400000  0.925000 3.650000 1.085000 ;
      RECT 3.465000  1.765000 3.795000 2.960000 ;
      RECT 3.830000  1.095000 4.160000 1.255000 ;
      RECT 3.965000  1.935000 4.295000 3.245000 ;
      RECT 4.390000  1.095000 4.720000 1.110000 ;
      RECT 4.390000  1.110000 6.560000 1.180000 ;
      RECT 4.390000  1.180000 5.650000 1.280000 ;
      RECT 4.390000  1.280000 4.720000 1.345000 ;
      RECT 4.465000  1.765000 4.795000 1.950000 ;
      RECT 4.465000  1.950000 7.235000 2.120000 ;
      RECT 4.465000  2.120000 4.795000 2.960000 ;
      RECT 4.890000  0.665000 5.220000 0.755000 ;
      RECT 4.890000  0.925000 5.220000 0.940000 ;
      RECT 4.965000  2.290000 6.165000 3.245000 ;
      RECT 5.400000  0.665000 5.650000 1.010000 ;
      RECT 5.400000  1.010000 6.560000 1.110000 ;
      RECT 5.880000  0.085000 6.130000 0.840000 ;
      RECT 6.310000  0.450000 6.560000 1.010000 ;
      RECT 6.335000  2.120000 6.665000 2.860000 ;
      RECT 6.740000  0.085000 7.070000 1.130000 ;
      RECT 6.875000  2.290000 7.205000 3.245000 ;
      RECT 7.065000  1.320000 8.565000 1.650000 ;
      RECT 7.065000  1.650000 7.235000 1.950000 ;
      RECT 7.740000  0.085000 8.070000 0.810000 ;
      RECT 7.775000  2.320000 8.105000 3.245000 ;
      RECT 8.670000  0.085000 9.005000 0.600000 ;
      RECT 8.675000  2.320000 9.005000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
  END
END sky130_fd_sc_hs__and4bb_4
MACRO sky130_fd_sc_hs__buf_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.920000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.450000 0.910000 1.780000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.470000 1.820000 1.830000 2.980000 ;
        RECT 1.475000 0.350000 1.830000 1.130000 ;
        RECT 1.660000 1.130000 1.830000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 1.920000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 1.920000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.920000 0.085000 ;
      RECT 0.000000  3.245000 1.920000 3.415000 ;
      RECT 0.115000  0.800000 0.795000 1.110000 ;
      RECT 0.115000  1.110000 1.300000 1.280000 ;
      RECT 0.470000  1.950000 1.300000 2.120000 ;
      RECT 0.470000  2.120000 0.800000 2.980000 ;
      RECT 0.970000  2.290000 1.300000 3.245000 ;
      RECT 0.975000  0.085000 1.305000 0.940000 ;
      RECT 1.130000  1.280000 1.300000 1.300000 ;
      RECT 1.130000  1.300000 1.490000 1.630000 ;
      RECT 1.130000  1.630000 1.300000 1.950000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
  END
END sky130_fd_sc_hs__buf_1
MACRO sky130_fd_sc_hs__buf_16
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.56000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.674000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.775000 1.350000 10.435000 1.780000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  4.345600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.575000 1.920000 7.255000 2.150000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.560000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.560000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 10.560000 0.085000 ;
      RECT  0.000000  3.245000 10.560000 3.415000 ;
      RECT  0.115000  1.820000  0.365000 3.245000 ;
      RECT  0.130000  0.085000  0.380000 1.130000 ;
      RECT  0.560000  0.350000  0.815000 2.980000 ;
      RECT  0.985000  1.300000  1.295000 1.780000 ;
      RECT  0.990000  0.085000  1.285000 1.130000 ;
      RECT  1.095000  1.965000  1.265000 3.245000 ;
      RECT  1.465000  0.350000  1.720000 2.980000 ;
      RECT  1.890000  1.300000  2.175000 1.780000 ;
      RECT  1.895000  0.085000  2.100000 1.130000 ;
      RECT  1.965000  1.965000  2.215000 3.245000 ;
      RECT  2.345000  0.350000  2.610000 1.185000 ;
      RECT  2.345000  1.185000  2.675000 1.355000 ;
      RECT  2.415000  1.355000  2.675000 2.980000 ;
      RECT  2.790000  0.085000  2.960000 1.015000 ;
      RECT  2.845000  1.300000  3.140000 1.780000 ;
      RECT  2.945000  1.965000  3.115000 3.245000 ;
      RECT  3.220000  0.350000  3.480000 1.130000 ;
      RECT  3.310000  1.130000  3.480000 1.820000 ;
      RECT  3.310000  1.820000  3.565000 2.980000 ;
      RECT  3.650000  0.085000  3.820000 1.130000 ;
      RECT  3.655000  1.300000  4.045000 1.655000 ;
      RECT  3.735000  1.655000  4.045000 1.780000 ;
      RECT  3.845000  1.965000  4.015000 3.245000 ;
      RECT  4.000000  0.350000  4.385000 1.130000 ;
      RECT  4.215000  1.130000  4.385000 1.900000 ;
      RECT  4.215000  1.900000  4.545000 2.980000 ;
      RECT  4.555000  0.085000  4.830000 1.130000 ;
      RECT  4.555000  1.300000  4.865000 1.730000 ;
      RECT  4.675000  1.730000  4.865000 1.780000 ;
      RECT  4.745000  1.965000  4.915000 3.245000 ;
      RECT  5.035000  0.350000  5.330000 1.205000 ;
      RECT  5.035000  1.205000  5.410000 1.375000 ;
      RECT  5.115000  1.375000  5.410000 2.980000 ;
      RECT  5.500000  0.085000  5.830000 1.035000 ;
      RECT  5.580000  1.300000  5.890000 1.780000 ;
      RECT  5.645000  1.965000  5.815000 3.245000 ;
      RECT  6.000000  0.350000  6.330000 1.130000 ;
      RECT  6.060000  1.130000  6.330000 2.980000 ;
      RECT  6.500000  0.085000  6.830000 1.130000 ;
      RECT  6.500000  1.300000  6.810000 1.780000 ;
      RECT  6.545000  1.965000  6.715000 3.245000 ;
      RECT  6.980000  1.250000  7.245000 2.980000 ;
      RECT  7.000000  0.350000  7.250000 1.250000 ;
      RECT  7.420000  1.010000  9.945000 1.180000 ;
      RECT  7.420000  1.180000  7.590000 1.950000 ;
      RECT  7.420000  1.950000  9.995000 2.120000 ;
      RECT  7.430000  0.085000  7.760000 0.840000 ;
      RECT  7.445000  2.290000  7.695000 3.245000 ;
      RECT  7.865000  2.120000  8.195000 2.980000 ;
      RECT  7.940000  0.350000  8.110000 1.010000 ;
      RECT  8.290000  0.085000  8.620000 0.840000 ;
      RECT  8.395000  2.290000  8.565000 3.245000 ;
      RECT  8.765000  2.120000  9.095000 2.980000 ;
      RECT  8.800000  0.350000  8.970000 1.010000 ;
      RECT  9.150000  0.085000  9.480000 0.840000 ;
      RECT  9.295000  2.290000  9.465000 3.245000 ;
      RECT  9.665000  2.120000  9.995000 2.980000 ;
      RECT  9.695000  0.350000  9.945000 1.010000 ;
      RECT 10.115000  0.085000 10.445000 1.130000 ;
      RECT 10.195000  1.950000 10.445000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  1.950000  0.805000 2.120000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.055000  1.580000  1.225000 1.750000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.515000  1.950000  1.685000 2.120000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  1.950000  1.580000  2.120000 1.750000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.470000  1.950000  2.640000 2.120000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  2.910000  1.580000  3.080000 1.750000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.360000  1.950000  3.530000 2.120000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.800000  1.580000  3.970000 1.750000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.300000  1.950000  4.470000 2.120000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.680000  1.580000  4.850000 1.750000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.195000  1.950000  5.365000 2.120000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.650000  1.580000  5.820000 1.750000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.095000  1.950000  6.265000 2.120000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.565000  1.580000  6.735000 1.750000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.025000  1.950000  7.195000 2.120000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.420000  1.580000  7.590000 1.750000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
    LAYER met1 ;
      RECT 0.985000 1.550000 7.650000 1.780000 ;
  END
END sky130_fd_sc_hs__buf_16
MACRO sky130_fd_sc_hs__buf_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.400000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.825000 1.350000 2.275000 1.780000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945000 0.350000 1.275000 1.180000 ;
        RECT 0.945000 1.180000 1.315000 2.150000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.400000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.400000 0.085000 ;
      RECT 0.000000  3.245000 2.400000 3.415000 ;
      RECT 0.105000  1.300000 0.775000 1.630000 ;
      RECT 0.115000  1.820000 0.420000 2.735000 ;
      RECT 0.115000  2.735000 0.825000 3.245000 ;
      RECT 0.515000  0.085000 0.765000 1.130000 ;
      RECT 0.605000  1.630000 0.775000 2.320000 ;
      RECT 0.605000  2.320000 2.285000 2.490000 ;
      RECT 1.395000  2.660000 1.725000 3.245000 ;
      RECT 1.445000  0.085000 1.775000 0.840000 ;
      RECT 1.485000  1.010000 2.285000 1.180000 ;
      RECT 1.485000  1.180000 1.655000 2.320000 ;
      RECT 1.930000  1.950000 2.285000 2.320000 ;
      RECT 1.930000  2.490000 2.285000 2.880000 ;
      RECT 1.955000  0.450000 2.285000 1.010000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
  END
END sky130_fd_sc_hs__buf_2
MACRO sky130_fd_sc_hs__buf_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.363000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.350000 2.905000 1.780000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.180000 0.835000 1.410000 ;
        RECT 0.615000 0.350000 0.945000 0.960000 ;
        RECT 0.615000 0.960000 1.945000 1.130000 ;
        RECT 0.615000 1.130000 0.835000 1.180000 ;
        RECT 0.660000 1.410000 0.835000 1.800000 ;
        RECT 0.660000 1.800000 1.730000 1.970000 ;
        RECT 0.660000 1.970000 0.835000 2.980000 ;
        RECT 1.560000 1.970000 1.730000 2.980000 ;
        RECT 1.615000 0.350000 1.945000 0.960000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 1.010000 ;
      RECT 0.130000  1.820000 0.460000 3.245000 ;
      RECT 1.030000  2.140000 1.360000 3.245000 ;
      RECT 1.060000  1.300000 2.285000 1.630000 ;
      RECT 1.115000  0.085000 1.445000 0.790000 ;
      RECT 1.930000  1.820000 2.260000 3.245000 ;
      RECT 2.115000  0.085000 2.745000 0.680000 ;
      RECT 2.115000  0.960000 3.245000 1.130000 ;
      RECT 2.115000  1.130000 2.285000 1.300000 ;
      RECT 2.465000  1.950000 3.245000 2.200000 ;
      RECT 2.915000  0.350000 3.245000 0.960000 ;
      RECT 2.915000  2.370000 3.245000 3.245000 ;
      RECT 3.075000  1.130000 3.245000 1.950000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__buf_4
MACRO sky130_fd_sc_hs__buf_8
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.837000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.430000 1.780000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  2.249300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.960000 0.350000 2.130000 0.960000 ;
        RECT 1.960000 0.960000 5.145000 1.130000 ;
        RECT 1.970000 1.800000 5.155000 1.970000 ;
        RECT 1.970000 1.970000 2.300000 2.980000 ;
        RECT 2.810000 0.350000 3.140000 0.960000 ;
        RECT 2.920000 1.970000 3.250000 2.980000 ;
        RECT 3.810000 0.350000 4.140000 0.960000 ;
        RECT 3.870000 1.970000 4.200000 2.980000 ;
        RECT 4.810000 0.350000 5.145000 0.960000 ;
        RECT 4.820000 1.970000 5.155000 2.980000 ;
        RECT 4.975000 1.130000 5.145000 1.800000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.115000  0.350000 0.365000 1.010000 ;
      RECT 0.115000  1.010000 1.770000 1.180000 ;
      RECT 0.120000  1.950000 1.770000 2.120000 ;
      RECT 0.120000  2.120000 0.450000 2.980000 ;
      RECT 0.545000  0.085000 0.875000 0.840000 ;
      RECT 0.650000  2.290000 0.820000 3.245000 ;
      RECT 1.020000  2.120000 1.350000 2.980000 ;
      RECT 1.100000  0.350000 1.270000 1.010000 ;
      RECT 1.450000  0.085000 1.780000 0.840000 ;
      RECT 1.550000  2.290000 1.800000 3.245000 ;
      RECT 1.600000  1.180000 1.770000 1.300000 ;
      RECT 1.600000  1.300000 4.805000 1.630000 ;
      RECT 1.600000  1.630000 1.770000 1.950000 ;
      RECT 2.310000  0.085000 2.640000 0.790000 ;
      RECT 2.500000  2.140000 2.750000 3.245000 ;
      RECT 3.310000  0.085000 3.640000 0.790000 ;
      RECT 3.450000  2.140000 3.700000 3.245000 ;
      RECT 4.310000  0.085000 4.640000 0.790000 ;
      RECT 4.400000  2.140000 4.650000 3.245000 ;
      RECT 5.315000  0.085000 5.645000 1.130000 ;
      RECT 5.350000  1.820000 5.600000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_hs__buf_8
MACRO sky130_fd_sc_hs__bufbuf_16
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.96000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.505000 1.780000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  4.401600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 5.700000 1.920000 12.380000 2.150000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.960000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 12.960000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.960000 0.085000 ;
      RECT  0.000000  3.245000 12.960000 3.415000 ;
      RECT  0.115000  1.950000  0.845000 2.120000 ;
      RECT  0.115000  2.120000  0.445000 2.980000 ;
      RECT  0.130000  0.350000  0.380000 0.960000 ;
      RECT  0.130000  0.960000  0.845000 1.130000 ;
      RECT  0.560000  0.085000  0.890000 0.790000 ;
      RECT  0.645000  2.290000  0.815000 3.245000 ;
      RECT  0.675000  1.130000  0.845000 1.300000 ;
      RECT  0.675000  1.300000  1.875000 1.630000 ;
      RECT  0.675000  1.630000  0.845000 1.950000 ;
      RECT  1.015000  1.800000  2.245000 1.970000 ;
      RECT  1.015000  1.970000  1.345000 2.980000 ;
      RECT  1.070000  0.350000  1.240000 0.960000 ;
      RECT  1.070000  0.960000  2.215000 1.130000 ;
      RECT  1.420000  0.085000  1.670000 0.790000 ;
      RECT  1.545000  2.140000  1.715000 3.245000 ;
      RECT  1.855000  0.350000  2.215000 0.960000 ;
      RECT  1.915000  1.970000  2.245000 2.980000 ;
      RECT  2.045000  1.130000  2.215000 1.320000 ;
      RECT  2.045000  1.320000  4.480000 1.650000 ;
      RECT  2.045000  1.650000  2.245000 1.800000 ;
      RECT  2.415000  0.085000  2.745000 1.130000 ;
      RECT  2.490000  1.820000  2.740000 3.245000 ;
      RECT  2.915000  0.350000  3.165000 0.980000 ;
      RECT  2.915000  0.980000  5.105000 1.150000 ;
      RECT  2.940000  1.820000  5.080000 1.990000 ;
      RECT  2.940000  1.990000  3.270000 2.980000 ;
      RECT  3.345000  0.085000  3.675000 0.810000 ;
      RECT  3.470000  2.160000  3.640000 3.245000 ;
      RECT  3.840000  1.990000  4.170000 2.980000 ;
      RECT  3.845000  0.350000  4.095000 0.980000 ;
      RECT  4.275000  0.085000  4.605000 0.810000 ;
      RECT  4.370000  2.160000  4.540000 3.245000 ;
      RECT  4.750000  1.990000  5.080000 2.980000 ;
      RECT  4.775000  0.350000  5.025000 0.980000 ;
      RECT  4.845000  1.150000  5.105000 1.320000 ;
      RECT  4.845000  1.320000  5.405000 1.755000 ;
      RECT  4.845000  1.755000  5.080000 1.820000 ;
      RECT  5.275000  0.085000  5.455000 1.130000 ;
      RECT  5.280000  1.925000  5.450000 3.245000 ;
      RECT  5.635000  0.350000  5.885000 1.900000 ;
      RECT  5.660000  1.900000  5.885000 1.920000 ;
      RECT  5.660000  1.920000  5.990000 2.980000 ;
      RECT  6.055000  1.320000  6.365000 1.750000 ;
      RECT  6.065000  0.085000  6.315000 1.130000 ;
      RECT  6.160000  1.925000  6.410000 3.245000 ;
      RECT  6.535000  0.350000  6.780000 1.650000 ;
      RECT  6.610000  1.650000  6.780000 1.920000 ;
      RECT  6.610000  1.920000  6.940000 2.980000 ;
      RECT  6.950000  1.320000  7.215000 1.750000 ;
      RECT  6.960000  0.085000  7.175000 1.130000 ;
      RECT  7.140000  1.925000  7.310000 3.245000 ;
      RECT  7.385000  0.350000  7.680000 1.650000 ;
      RECT  7.510000  1.650000  7.680000 1.920000 ;
      RECT  7.510000  1.920000  7.840000 2.980000 ;
      RECT  7.850000  0.085000  8.115000 1.130000 ;
      RECT  7.850000  1.320000  8.115000 1.750000 ;
      RECT  8.040000  1.925000  8.210000 3.245000 ;
      RECT  8.285000  0.350000  8.580000 1.650000 ;
      RECT  8.410000  1.650000  8.580000 1.920000 ;
      RECT  8.410000  1.920000  8.740000 2.980000 ;
      RECT  8.750000  0.085000  9.045000 1.130000 ;
      RECT  8.750000  1.320000  9.045000 1.750000 ;
      RECT  8.940000  1.925000  9.110000 3.245000 ;
      RECT  9.215000  0.350000  9.480000 1.650000 ;
      RECT  9.310000  1.650000  9.480000 1.920000 ;
      RECT  9.310000  1.920000  9.640000 2.980000 ;
      RECT  9.650000  1.320000  9.975000 1.750000 ;
      RECT  9.665000  0.085000  9.975000 1.130000 ;
      RECT  9.840000  1.925000 10.010000 3.245000 ;
      RECT 10.145000  0.350000 10.395000 1.650000 ;
      RECT 10.210000  1.650000 10.395000 1.920000 ;
      RECT 10.210000  1.920000 10.540000 2.980000 ;
      RECT 10.565000  1.320000 10.940000 1.750000 ;
      RECT 10.575000  0.085000 10.905000 1.130000 ;
      RECT 10.740000  1.925000 10.910000 3.245000 ;
      RECT 11.110000  0.350000 11.325000 1.920000 ;
      RECT 11.110000  1.920000 11.440000 2.980000 ;
      RECT 11.495000  1.320000 11.890000 1.750000 ;
      RECT 11.505000  0.085000 11.835000 1.130000 ;
      RECT 11.640000  1.925000 11.890000 3.245000 ;
      RECT 12.015000  0.350000 12.345000 1.150000 ;
      RECT 12.060000  1.150000 12.345000 2.020000 ;
      RECT 12.060000  2.020000 12.390000 2.980000 ;
      RECT 12.515000  0.085000 12.845000 1.130000 ;
      RECT 12.590000  1.820000 12.840000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.180000  1.580000  5.350000 1.750000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.760000  1.950000  5.930000 2.120000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.125000  1.580000  6.295000 1.750000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.675000  1.950000  6.845000 2.120000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.000000  1.580000  7.170000 1.750000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.595000  1.950000  7.765000 2.120000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  7.900000  1.580000  8.070000 1.750000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.485000  1.950000  8.655000 2.120000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  8.820000  1.580000  8.990000 1.750000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.405000  1.950000  9.575000 2.120000 ;
      RECT  9.730000  1.580000  9.900000 1.750000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.295000  1.950000 10.465000 2.120000 ;
      RECT 10.675000  1.580000 10.845000 1.750000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  1.950000 11.365000 2.120000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.600000  1.580000 11.770000 1.750000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.115000  1.950000 12.285000 2.120000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
    LAYER met1 ;
      RECT 5.110000 1.550000 11.830000 1.780000 ;
  END
END sky130_fd_sc_hs__bufbuf_16
MACRO sky130_fd_sc_hs__bufbuf_8
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 0.570000 1.780000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  2.273200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.475000 0.350000 3.805000 0.880000 ;
        RECT 3.475000 0.880000 6.585000 1.130000 ;
        RECT 3.565000 1.800000 6.555000 1.970000 ;
        RECT 3.565000 1.970000 3.830000 2.980000 ;
        RECT 4.495000 1.970000 4.745000 2.980000 ;
        RECT 5.385000 1.970000 5.655000 2.980000 ;
        RECT 6.255000 0.350000 6.585000 0.880000 ;
        RECT 6.255000 1.130000 6.585000 1.270000 ;
        RECT 6.255000 1.270000 7.075000 1.780000 ;
        RECT 6.255000 1.780000 6.555000 1.800000 ;
        RECT 6.285000 1.970000 6.555000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.200000 0.085000 ;
      RECT 0.000000  3.245000 7.200000 3.415000 ;
      RECT 0.115000  0.540000 0.445000 1.010000 ;
      RECT 0.115000  1.010000 0.920000 1.180000 ;
      RECT 0.115000  1.950000 0.920000 2.200000 ;
      RECT 0.115000  2.200000 0.380000 2.700000 ;
      RECT 0.565000  2.370000 0.920000 3.245000 ;
      RECT 0.625000  0.085000 0.955000 0.840000 ;
      RECT 0.750000  1.180000 0.920000 1.300000 ;
      RECT 0.750000  1.300000 1.140000 1.630000 ;
      RECT 0.750000  1.630000 0.920000 1.950000 ;
      RECT 1.090000  1.820000 1.480000 2.980000 ;
      RECT 1.125000  0.350000 1.480000 1.130000 ;
      RECT 1.310000  1.130000 1.480000 1.300000 ;
      RECT 1.310000  1.300000 2.500000 1.630000 ;
      RECT 1.310000  1.630000 1.480000 1.820000 ;
      RECT 1.650000  1.820000 2.880000 1.990000 ;
      RECT 1.650000  1.990000 1.980000 2.980000 ;
      RECT 1.685000  0.350000 1.935000 0.880000 ;
      RECT 1.685000  0.880000 3.125000 1.130000 ;
      RECT 2.115000  0.085000 2.445000 0.710000 ;
      RECT 2.150000  2.160000 2.380000 3.245000 ;
      RECT 2.550000  1.990000 2.880000 2.980000 ;
      RECT 2.670000  1.130000 3.125000 1.300000 ;
      RECT 2.670000  1.300000 6.020000 1.630000 ;
      RECT 2.670000  1.630000 2.880000 1.820000 ;
      RECT 2.975000  0.085000 3.305000 0.710000 ;
      RECT 3.050000  1.820000 3.380000 3.245000 ;
      RECT 3.975000  0.085000 4.305000 0.710000 ;
      RECT 4.035000  2.140000 4.290000 3.245000 ;
      RECT 4.835000  0.085000 5.165000 0.710000 ;
      RECT 4.930000  2.140000 5.205000 3.245000 ;
      RECT 5.755000  0.085000 6.085000 0.710000 ;
      RECT 5.835000  2.140000 6.105000 3.245000 ;
      RECT 6.735000  1.950000 7.040000 3.245000 ;
      RECT 6.755000  0.085000 7.085000 1.100000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
  END
END sky130_fd_sc_hs__bufbuf_8
MACRO sky130_fd_sc_hs__bufinv_16
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.837000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.430000 1.780000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  4.390400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 4.660000 1.920000 11.400000 2.150000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.000000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 12.000000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.000000 0.085000 ;
      RECT  0.000000  3.245000 12.000000 3.415000 ;
      RECT  0.115000  0.350000  0.365000 1.010000 ;
      RECT  0.115000  1.010000  1.770000 1.180000 ;
      RECT  0.120000  1.950000  1.770000 2.120000 ;
      RECT  0.120000  2.120000  0.450000 2.980000 ;
      RECT  0.545000  0.085000  0.875000 0.840000 ;
      RECT  0.650000  2.290000  0.820000 3.245000 ;
      RECT  1.020000  2.120000  1.350000 2.980000 ;
      RECT  1.115000  0.350000  1.285000 1.010000 ;
      RECT  1.465000  0.085000  1.795000 0.840000 ;
      RECT  1.550000  2.290000  1.720000 3.245000 ;
      RECT  1.600000  1.180000  1.770000 1.300000 ;
      RECT  1.600000  1.300000  3.460000 1.630000 ;
      RECT  1.600000  1.630000  1.770000 1.950000 ;
      RECT  1.940000  1.800000  4.070000 1.970000 ;
      RECT  1.940000  1.970000  2.270000 2.980000 ;
      RECT  1.975000  0.350000  2.145000 0.960000 ;
      RECT  1.975000  0.960000  3.935000 1.130000 ;
      RECT  2.325000  0.085000  2.575000 0.790000 ;
      RECT  2.470000  2.140000  2.640000 3.245000 ;
      RECT  2.755000  0.350000  3.005000 0.960000 ;
      RECT  2.840000  1.970000  3.170000 2.980000 ;
      RECT  3.185000  0.085000  3.515000 0.790000 ;
      RECT  3.370000  2.140000  3.540000 3.245000 ;
      RECT  3.685000  0.350000  3.935000 0.960000 ;
      RECT  3.685000  1.130000  3.935000 1.300000 ;
      RECT  3.740000  1.300000  4.435000 1.750000 ;
      RECT  3.740000  1.750000  4.070000 1.800000 ;
      RECT  3.740000  1.970000  4.070000 2.980000 ;
      RECT  4.115000  0.085000  4.445000 1.130000 ;
      RECT  4.270000  1.920000  4.440000 3.245000 ;
      RECT  4.615000  0.350000  4.865000 1.920000 ;
      RECT  4.615000  1.920000  4.970000 2.020000 ;
      RECT  4.640000  2.020000  4.970000 2.980000 ;
      RECT  5.035000  1.300000  5.305000 1.750000 ;
      RECT  5.045000  0.085000  5.295000 1.105000 ;
      RECT  5.170000  1.920000  5.340000 3.245000 ;
      RECT  5.510000  0.350000  5.725000 1.920000 ;
      RECT  5.510000  1.920000  5.870000 2.020000 ;
      RECT  5.540000  2.020000  5.870000 2.980000 ;
      RECT  5.900000  1.300000  6.230000 1.750000 ;
      RECT  5.905000  0.085000  6.235000 1.105000 ;
      RECT  6.070000  1.920000  6.240000 3.245000 ;
      RECT  6.420000  0.350000  6.655000 1.920000 ;
      RECT  6.420000  1.920000  6.770000 2.020000 ;
      RECT  6.440000  2.020000  6.770000 2.980000 ;
      RECT  6.835000  0.085000  7.165000 1.105000 ;
      RECT  6.840000  1.300000  7.170000 1.750000 ;
      RECT  6.970000  1.920000  7.140000 3.245000 ;
      RECT  7.340000  0.350000  7.585000 1.920000 ;
      RECT  7.340000  1.920000  7.670000 2.980000 ;
      RECT  7.760000  1.300000  8.090000 1.750000 ;
      RECT  7.765000  0.085000  8.095000 1.105000 ;
      RECT  7.870000  1.920000  8.040000 3.245000 ;
      RECT  8.240000  2.020000  8.570000 2.980000 ;
      RECT  8.265000  0.350000  8.515000 1.920000 ;
      RECT  8.265000  1.920000  8.570000 2.020000 ;
      RECT  8.685000  1.300000  9.015000 1.750000 ;
      RECT  8.695000  0.085000  9.025000 1.105000 ;
      RECT  8.770000  1.920000  8.995000 3.245000 ;
      RECT  9.190000  2.020000  9.520000 2.980000 ;
      RECT  9.195000  0.350000  9.445000 1.920000 ;
      RECT  9.195000  1.920000  9.520000 2.020000 ;
      RECT  9.615000  1.300000  9.945000 1.750000 ;
      RECT  9.625000  0.085000  9.955000 1.105000 ;
      RECT  9.720000  1.920000  9.955000 3.245000 ;
      RECT 10.125000  0.350000 10.375000 1.920000 ;
      RECT 10.125000  1.920000 10.470000 2.020000 ;
      RECT 10.140000  2.020000 10.470000 2.980000 ;
      RECT 10.545000  1.300000 10.875000 1.750000 ;
      RECT 10.555000  0.085000 10.885000 1.105000 ;
      RECT 10.670000  1.920000 10.885000 3.245000 ;
      RECT 11.055000  0.350000 11.385000 1.790000 ;
      RECT 11.055000  1.790000 11.420000 2.020000 ;
      RECT 11.090000  2.020000 11.420000 2.980000 ;
      RECT 11.555000  0.085000 11.885000 1.130000 ;
      RECT 11.620000  1.820000 11.870000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.225000  1.580000  4.395000 1.750000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.730000  1.950000  4.900000 2.120000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.090000  1.580000  5.260000 1.750000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.620000  1.950000  5.790000 2.120000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  5.980000  1.580000  6.150000 1.750000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.520000  1.950000  6.690000 2.120000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  6.920000  1.580000  7.090000 1.750000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.420000  1.950000  7.590000 2.120000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  1.580000  8.005000 1.750000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.320000  1.950000  8.490000 2.120000 ;
      RECT  8.765000  1.580000  8.935000 1.750000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.270000  1.950000  9.440000 2.120000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.690000  1.580000  9.860000 1.750000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.220000  1.950000 10.390000 2.120000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.625000  1.580000 10.795000 1.750000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.170000  1.950000 11.340000 2.120000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
    LAYER met1 ;
      RECT 4.155000 1.550000 10.855000 1.780000 ;
  END
END sky130_fd_sc_hs__bufinv_16
MACRO sky130_fd_sc_hs__bufinv_8
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 0.550000 1.780000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  2.385000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.060000 0.350000 1.390000 0.880000 ;
        RECT 1.060000 0.880000 3.250000 0.960000 ;
        RECT 1.060000 0.960000 4.250000 1.130000 ;
        RECT 1.060000 1.130000 1.390000 1.800000 ;
        RECT 1.060000 1.800000 4.225000 2.070000 ;
        RECT 2.060000 0.350000 2.250000 0.880000 ;
        RECT 2.920000 0.350000 3.250000 0.880000 ;
        RECT 3.920000 0.350000 4.250000 0.960000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.240000 0.085000 ;
      RECT 0.000000  3.245000 6.240000 3.415000 ;
      RECT 0.115000  1.950000 0.445000 2.240000 ;
      RECT 0.115000  2.240000 4.565000 2.410000 ;
      RECT 0.115000  2.410000 0.445000 2.980000 ;
      RECT 0.130000  0.350000 0.380000 1.010000 ;
      RECT 0.130000  1.010000 0.890000 1.180000 ;
      RECT 0.560000  0.085000 0.890000 0.840000 ;
      RECT 0.615000  2.580000 0.945000 3.245000 ;
      RECT 0.720000  1.180000 0.890000 2.240000 ;
      RECT 1.515000  2.580000 1.845000 3.245000 ;
      RECT 1.560000  0.085000 1.890000 0.710000 ;
      RECT 1.665000  1.300000 4.820000 1.630000 ;
      RECT 2.415000  2.580000 2.745000 3.245000 ;
      RECT 2.420000  0.085000 2.750000 0.710000 ;
      RECT 3.315000  2.580000 3.645000 3.245000 ;
      RECT 3.420000  0.085000 3.750000 0.790000 ;
      RECT 4.345000  2.580000 4.675000 3.245000 ;
      RECT 4.395000  1.800000 5.605000 1.970000 ;
      RECT 4.395000  1.970000 4.565000 2.240000 ;
      RECT 4.420000  0.085000 4.750000 0.710000 ;
      RECT 4.650000  0.880000 6.125000 1.130000 ;
      RECT 4.650000  1.130000 4.820000 1.300000 ;
      RECT 4.845000  2.140000 6.125000 2.310000 ;
      RECT 4.845000  2.310000 5.175000 2.980000 ;
      RECT 4.920000  0.350000 5.125000 0.880000 ;
      RECT 4.990000  1.320000 5.605000 1.800000 ;
      RECT 5.295000  0.085000 5.625000 0.710000 ;
      RECT 5.345000  2.480000 5.675000 3.245000 ;
      RECT 5.795000  0.350000 6.125000 0.880000 ;
      RECT 5.795000  1.130000 6.125000 2.140000 ;
      RECT 5.845000  2.310000 6.125000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
  END
END sky130_fd_sc_hs__bufinv_8
MACRO sky130_fd_sc_hs__clkbuf_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.920000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.231000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.835000 1.780000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.449400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.345000 1.820000 1.805000 2.980000 ;
        RECT 1.475000 0.350000 1.805000 0.790000 ;
        RECT 1.565000 0.790000 1.805000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 1.920000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 1.920000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.920000 0.085000 ;
      RECT 0.000000  3.245000 1.920000 3.415000 ;
      RECT 0.115000  0.350000 0.445000 0.960000 ;
      RECT 0.115000  0.960000 1.395000 1.130000 ;
      RECT 0.345000  1.950000 1.175000 2.120000 ;
      RECT 0.345000  2.120000 0.675000 2.980000 ;
      RECT 0.615000  0.085000 1.305000 0.680000 ;
      RECT 0.845000  2.290000 1.175000 3.245000 ;
      RECT 1.005000  1.130000 1.395000 1.630000 ;
      RECT 1.005000  1.630000 1.175000 1.950000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
  END
END sky130_fd_sc_hs__clkbuf_1
MACRO sky130_fd_sc_hs__clkbuf_16
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.600000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.924000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.795000 1.780000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  3.628800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2.390000 1.920000 9.090000 2.150000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.600000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.600000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.600000 0.085000 ;
      RECT 0.000000  3.245000 9.600000 3.415000 ;
      RECT 0.115000  0.085000 0.365000 0.810000 ;
      RECT 0.120000  1.950000 0.370000 3.245000 ;
      RECT 0.545000  0.350000 0.795000 0.980000 ;
      RECT 0.545000  0.980000 2.135000 1.150000 ;
      RECT 0.570000  1.950000 2.135000 2.120000 ;
      RECT 0.570000  2.120000 0.900000 2.980000 ;
      RECT 0.975000  0.085000 1.225000 0.810000 ;
      RECT 1.100000  2.290000 1.270000 3.245000 ;
      RECT 1.425000  0.350000 1.675000 0.980000 ;
      RECT 1.470000  2.120000 1.800000 2.980000 ;
      RECT 1.855000  0.085000 2.185000 0.810000 ;
      RECT 1.965000  1.150000 2.135000 1.180000 ;
      RECT 1.965000  1.180000 2.210000 1.410000 ;
      RECT 1.965000  1.410000 2.135000 1.950000 ;
      RECT 2.000000  2.290000 2.250000 3.245000 ;
      RECT 2.390000  0.350000 2.660000 2.120000 ;
      RECT 2.430000  2.120000 2.660000 2.980000 ;
      RECT 2.830000  2.030000 3.160000 3.245000 ;
      RECT 2.835000  1.190000 3.105000 1.520000 ;
      RECT 2.865000  0.085000 3.035000 0.680000 ;
      RECT 3.275000  0.350000 3.500000 1.690000 ;
      RECT 3.275000  1.690000 3.545000 1.860000 ;
      RECT 3.340000  1.860000 3.545000 2.980000 ;
      RECT 3.670000  0.085000 3.895000 0.725000 ;
      RECT 3.670000  1.190000 4.000000 1.520000 ;
      RECT 3.730000  2.030000 4.060000 3.245000 ;
      RECT 4.075000  0.350000 4.340000 0.745000 ;
      RECT 4.170000  0.745000 4.340000 1.690000 ;
      RECT 4.170000  1.690000 4.430000 1.860000 ;
      RECT 4.230000  1.860000 4.430000 2.980000 ;
      RECT 4.510000  0.085000 4.835000 0.740000 ;
      RECT 4.510000  1.190000 4.840000 1.520000 ;
      RECT 4.630000  2.030000 4.960000 3.245000 ;
      RECT 5.025000  0.350000 5.255000 1.690000 ;
      RECT 5.025000  1.690000 5.350000 1.860000 ;
      RECT 5.140000  1.860000 5.350000 2.980000 ;
      RECT 5.425000  1.190000 5.755000 1.520000 ;
      RECT 5.435000  0.085000 5.765000 0.680000 ;
      RECT 5.530000  2.030000 5.860000 3.245000 ;
      RECT 5.935000  0.350000 6.185000 1.690000 ;
      RECT 5.935000  1.690000 6.245000 1.860000 ;
      RECT 6.040000  1.860000 6.245000 2.980000 ;
      RECT 6.365000  0.085000 6.695000 0.680000 ;
      RECT 6.365000  1.190000 6.695000 1.520000 ;
      RECT 6.430000  2.030000 6.760000 3.245000 ;
      RECT 6.865000  0.350000 7.115000 1.690000 ;
      RECT 6.865000  1.690000 7.150000 1.860000 ;
      RECT 6.945000  1.860000 7.150000 2.980000 ;
      RECT 7.295000  0.085000 7.625000 0.680000 ;
      RECT 7.295000  1.190000 7.625000 1.520000 ;
      RECT 7.330000  2.030000 7.660000 3.245000 ;
      RECT 7.795000  0.350000 8.045000 1.690000 ;
      RECT 7.795000  1.690000 8.050000 1.860000 ;
      RECT 7.840000  1.860000 8.050000 2.980000 ;
      RECT 8.225000  0.085000 8.555000 0.680000 ;
      RECT 8.225000  1.190000 8.555000 1.520000 ;
      RECT 8.230000  2.030000 8.560000 3.245000 ;
      RECT 8.725000  0.350000 8.975000 1.830000 ;
      RECT 8.725000  1.830000 8.970000 1.860000 ;
      RECT 8.750000  1.860000 8.970000 2.980000 ;
      RECT 9.150000  2.030000 9.480000 3.245000 ;
      RECT 9.155000  0.085000 9.485000 0.745000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.010000  1.210000 2.180000 1.380000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.460000  1.950000 2.630000 2.120000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 2.890000  1.210000 3.060000 1.380000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.360000  1.950000 3.530000 2.120000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.750000  1.210000 3.920000 1.380000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.245000  1.950000 4.415000 2.120000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.590000  1.210000 4.760000 1.380000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.160000  1.950000 5.330000 2.120000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.505000  1.210000 5.675000 1.380000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.060000  1.950000 6.230000 2.120000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.445000  1.210000 6.615000 1.380000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 6.960000  1.950000 7.130000 2.120000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.375000  1.210000 7.545000 1.380000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 7.860000  1.950000 8.030000 2.120000 ;
      RECT 8.305000  1.210000 8.475000 1.380000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.780000  1.950000 8.950000 2.120000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
    LAYER met1 ;
      RECT 1.940000 1.180000 8.640000 1.410000 ;
  END
END sky130_fd_sc_hs__clkbuf_16
MACRO sky130_fd_sc_hs__clkbuf_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.920000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.231000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.010000 1.495000 2.150000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.453600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.350000 0.885000 0.790000 ;
        RECT 0.555000 1.820000 0.885000 2.150000 ;
        RECT 0.715000 0.790000 0.885000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 1.920000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 1.920000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.920000 0.085000 ;
      RECT 0.000000  3.245000 1.920000 3.415000 ;
      RECT 0.105000  2.660000 0.435000 3.245000 ;
      RECT 0.115000  0.085000 0.365000 0.790000 ;
      RECT 0.215000  0.960000 0.545000 1.630000 ;
      RECT 0.215000  1.630000 0.385000 2.320000 ;
      RECT 0.215000  2.320000 1.835000 2.490000 ;
      RECT 1.005000  2.660000 1.335000 3.245000 ;
      RECT 1.055000  0.085000 1.305000 0.810000 ;
      RECT 1.475000  0.350000 1.835000 0.810000 ;
      RECT 1.535000  2.490000 1.835000 2.980000 ;
      RECT 1.665000  0.810000 1.835000 2.320000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
  END
END sky130_fd_sc_hs__clkbuf_2
MACRO sky130_fd_sc_hs__clkbuf_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.880000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.231000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.055000 1.080000 2.455000 1.410000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.924000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.980000 1.750000 1.150000 ;
        RECT 0.535000 1.150000 0.705000 1.920000 ;
        RECT 0.535000 1.920000 1.795000 2.090000 ;
        RECT 0.535000 2.090000 0.815000 2.980000 ;
        RECT 0.560000 0.350000 0.890000 0.980000 ;
        RECT 1.420000 0.350000 1.750000 0.980000 ;
        RECT 1.465000 2.090000 1.795000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.880000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.880000 0.085000 ;
      RECT 0.000000  3.245000 2.880000 3.415000 ;
      RECT 0.115000  1.820000 0.365000 3.245000 ;
      RECT 0.130000  0.085000 0.380000 0.810000 ;
      RECT 0.875000  1.350000 1.885000 1.580000 ;
      RECT 0.875000  1.580000 2.795000 1.750000 ;
      RECT 1.015000  2.260000 1.265000 3.245000 ;
      RECT 1.070000  0.085000 1.240000 0.810000 ;
      RECT 1.920000  0.085000 2.250000 0.810000 ;
      RECT 1.995000  1.920000 2.245000 3.245000 ;
      RECT 2.415000  1.750000 2.795000 2.980000 ;
      RECT 2.420000  0.480000 2.795000 0.810000 ;
      RECT 2.625000  0.810000 2.795000 1.580000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
  END
END sky130_fd_sc_hs__clkbuf_4
MACRO sky130_fd_sc_hs__clkbuf_8
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.462000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.095000 1.780000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.841700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.615000 0.350000 1.945000 0.850000 ;
        RECT 1.615000 0.850000 4.880000 1.020000 ;
        RECT 1.615000 1.690000 5.155000 1.860000 ;
        RECT 1.615000 1.860000 1.880000 2.980000 ;
        RECT 2.585000 1.860000 2.845000 2.980000 ;
        RECT 2.615000 0.350000 2.865000 0.850000 ;
        RECT 3.415000 1.860000 3.680000 2.980000 ;
        RECT 3.555000 0.350000 3.725000 0.850000 ;
        RECT 4.385000 1.860000 4.645000 2.980000 ;
        RECT 4.485000 0.350000 4.655000 0.850000 ;
        RECT 4.710000 1.020000 4.880000 1.180000 ;
        RECT 4.710000 1.180000 5.155000 1.690000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.280000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.245000 5.280000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 0.810000 ;
      RECT 0.115000  1.950000 0.445000 3.245000 ;
      RECT 0.615000  0.350000 0.945000 0.980000 ;
      RECT 0.615000  0.980000 1.445000 1.150000 ;
      RECT 0.615000  1.950000 1.445000 2.120000 ;
      RECT 0.615000  2.120000 0.945000 2.980000 ;
      RECT 1.115000  0.085000 1.445000 0.810000 ;
      RECT 1.115000  2.290000 1.445000 3.245000 ;
      RECT 1.275000  1.150000 1.445000 1.190000 ;
      RECT 1.275000  1.190000 4.515000 1.520000 ;
      RECT 1.275000  1.520000 1.445000 1.950000 ;
      RECT 2.065000  2.030000 2.395000 3.245000 ;
      RECT 2.115000  0.085000 2.445000 0.680000 ;
      RECT 3.045000  0.085000 3.375000 0.680000 ;
      RECT 3.045000  2.030000 3.215000 3.245000 ;
      RECT 3.865000  2.030000 4.195000 3.245000 ;
      RECT 3.905000  0.085000 4.305000 0.680000 ;
      RECT 4.830000  2.030000 5.160000 3.245000 ;
      RECT 4.835000  0.085000 5.165000 0.680000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
  END
END sky130_fd_sc_hs__clkbuf_8
MACRO sky130_fd_sc_hs__clkdlyinv3sd1_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.880000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.231000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.190000 0.730000 1.860000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.424900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.435000 0.355000 2.795000 0.755000 ;
        RECT 2.435000 1.815000 2.795000 3.060000 ;
        RECT 2.530000 0.755000 2.795000 1.815000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.880000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.880000 0.085000 ;
      RECT 0.000000  3.245000 2.880000 3.415000 ;
      RECT 0.095000  0.305000 0.410000 0.820000 ;
      RECT 0.095000  0.820000 1.305000 1.020000 ;
      RECT 0.095000  2.030000 1.305000 2.205000 ;
      RECT 0.095000  2.205000 0.400000 2.725000 ;
      RECT 0.575000  2.380000 0.905000 3.245000 ;
      RECT 0.585000  0.085000 0.915000 0.650000 ;
      RECT 0.975000  1.020000 1.305000 2.030000 ;
      RECT 1.415000  2.650000 1.745000 2.900000 ;
      RECT 1.475000  0.305000 1.720000 1.295000 ;
      RECT 1.475000  1.295000 2.360000 1.625000 ;
      RECT 1.475000  1.625000 1.745000 2.650000 ;
      RECT 1.935000  0.085000 2.265000 0.750000 ;
      RECT 1.935000  1.900000 2.265000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
  END
END sky130_fd_sc_hs__clkdlyinv3sd1_1
MACRO sky130_fd_sc_hs__clkdlyinv3sd2_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.880000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.231000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.190000 0.730000 1.860000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.424900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.435000 0.355000 2.795000 0.755000 ;
        RECT 2.435000 1.815000 2.795000 3.060000 ;
        RECT 2.530000 0.755000 2.795000 1.815000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.880000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.880000 0.085000 ;
      RECT 0.000000  3.245000 2.880000 3.415000 ;
      RECT 0.095000  0.305000 0.410000 0.820000 ;
      RECT 0.095000  0.820000 1.305000 1.020000 ;
      RECT 0.095000  2.030000 1.305000 2.205000 ;
      RECT 0.095000  2.205000 0.400000 2.725000 ;
      RECT 0.575000  2.380000 0.905000 3.245000 ;
      RECT 0.585000  0.085000 0.915000 0.650000 ;
      RECT 0.975000  1.020000 1.305000 2.030000 ;
      RECT 1.415000  2.650000 1.745000 2.900000 ;
      RECT 1.475000  0.305000 1.720000 1.295000 ;
      RECT 1.475000  1.295000 2.360000 1.625000 ;
      RECT 1.475000  1.625000 1.745000 2.650000 ;
      RECT 1.935000  0.085000 2.265000 0.750000 ;
      RECT 1.935000  1.900000 2.265000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
  END
END sky130_fd_sc_hs__clkdlyinv3sd2_1
MACRO sky130_fd_sc_hs__clkdlyinv3sd3_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.880000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.231000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.190000 0.730000 1.860000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.424900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.435000 0.355000 2.795000 0.755000 ;
        RECT 2.435000 1.815000 2.795000 3.060000 ;
        RECT 2.530000 0.755000 2.795000 1.815000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.880000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.880000 0.085000 ;
      RECT 0.000000  3.245000 2.880000 3.415000 ;
      RECT 0.095000  0.305000 0.410000 0.820000 ;
      RECT 0.095000  0.820000 1.305000 1.020000 ;
      RECT 0.095000  2.030000 1.305000 2.205000 ;
      RECT 0.095000  2.205000 0.400000 2.725000 ;
      RECT 0.575000  2.380000 0.905000 3.245000 ;
      RECT 0.585000  0.085000 0.915000 0.650000 ;
      RECT 0.975000  1.020000 1.305000 2.030000 ;
      RECT 1.415000  2.650000 1.745000 2.900000 ;
      RECT 1.475000  0.305000 1.720000 1.295000 ;
      RECT 1.475000  1.295000 2.360000 1.625000 ;
      RECT 1.475000  1.625000 1.745000 2.650000 ;
      RECT 1.935000  0.085000 2.265000 0.750000 ;
      RECT 1.935000  1.900000 2.265000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
  END
END sky130_fd_sc_hs__clkdlyinv3sd3_1
MACRO sky130_fd_sc_hs__clkdlyinv5sd1_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.231000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.190000 0.730000 1.860000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.424900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.830000 0.355000 5.190000 0.755000 ;
        RECT 4.830000 1.900000 5.190000 3.060000 ;
        RECT 4.925000 0.755000 5.190000 1.900000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.280000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.245000 5.280000 3.415000 ;
      RECT 0.095000  0.305000 0.410000 0.820000 ;
      RECT 0.095000  0.820000 1.305000 1.020000 ;
      RECT 0.095000  2.030000 1.305000 2.205000 ;
      RECT 0.095000  2.205000 0.400000 2.725000 ;
      RECT 0.575000  2.380000 0.905000 3.245000 ;
      RECT 0.585000  0.085000 0.915000 0.650000 ;
      RECT 0.975000  1.020000 1.305000 2.030000 ;
      RECT 1.415000  2.650000 1.745000 2.900000 ;
      RECT 1.475000  0.305000 1.720000 1.140000 ;
      RECT 1.475000  1.140000 2.510000 1.470000 ;
      RECT 1.475000  1.470000 1.745000 2.650000 ;
      RECT 1.915000  0.085000 2.265000 0.745000 ;
      RECT 1.915000  1.940000 2.265000 3.245000 ;
      RECT 2.800000  0.415000 2.970000 1.220000 ;
      RECT 2.800000  1.220000 4.005000 1.390000 ;
      RECT 2.800000  1.390000 2.970000 2.980000 ;
      RECT 3.370000  0.400000 3.700000 0.880000 ;
      RECT 3.370000  0.880000 4.700000 0.925000 ;
      RECT 3.370000  0.925000 4.755000 1.050000 ;
      RECT 3.415000  1.560000 4.755000 1.730000 ;
      RECT 3.415000  1.730000 3.655000 2.980000 ;
      RECT 4.330000  0.085000 4.660000 0.670000 ;
      RECT 4.330000  1.900000 4.660000 3.245000 ;
      RECT 4.530000  1.050000 4.755000 1.560000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
  END
END sky130_fd_sc_hs__clkdlyinv5sd1_1
MACRO sky130_fd_sc_hs__clkdlyinv5sd2_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.231000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.190000 0.730000 1.860000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.424900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.830000 0.355000 5.190000 0.755000 ;
        RECT 4.830000 1.900000 5.190000 3.060000 ;
        RECT 4.925000 0.755000 5.190000 1.900000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.280000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.245000 5.280000 3.415000 ;
      RECT 0.095000  0.305000 0.410000 0.820000 ;
      RECT 0.095000  0.820000 1.305000 1.020000 ;
      RECT 0.095000  2.030000 1.305000 2.205000 ;
      RECT 0.095000  2.205000 0.400000 2.725000 ;
      RECT 0.575000  2.380000 0.905000 3.245000 ;
      RECT 0.585000  0.085000 0.915000 0.650000 ;
      RECT 0.975000  1.020000 1.305000 2.030000 ;
      RECT 1.415000  2.650000 1.745000 2.900000 ;
      RECT 1.475000  0.305000 1.720000 1.140000 ;
      RECT 1.475000  1.140000 2.510000 1.470000 ;
      RECT 1.475000  1.470000 1.745000 2.650000 ;
      RECT 1.915000  0.085000 2.265000 0.745000 ;
      RECT 1.915000  1.940000 2.265000 3.245000 ;
      RECT 2.800000  0.415000 2.970000 1.220000 ;
      RECT 2.800000  1.220000 4.005000 1.390000 ;
      RECT 2.800000  1.390000 2.970000 2.980000 ;
      RECT 3.370000  0.400000 3.700000 0.880000 ;
      RECT 3.370000  0.880000 4.700000 0.925000 ;
      RECT 3.370000  0.925000 4.755000 1.050000 ;
      RECT 3.415000  1.560000 4.755000 1.730000 ;
      RECT 3.415000  1.730000 3.655000 2.980000 ;
      RECT 4.330000  0.085000 4.660000 0.670000 ;
      RECT 4.330000  1.900000 4.660000 3.245000 ;
      RECT 4.530000  1.050000 4.755000 1.560000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
  END
END sky130_fd_sc_hs__clkdlyinv5sd2_1
MACRO sky130_fd_sc_hs__clkdlyinv5sd3_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.231000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.190000 0.730000 1.860000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.424900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.830000 0.355000 5.190000 0.755000 ;
        RECT 4.830000 1.900000 5.190000 3.060000 ;
        RECT 4.925000 0.755000 5.190000 1.900000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.280000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.245000 5.280000 3.415000 ;
      RECT 0.095000  0.305000 0.410000 0.820000 ;
      RECT 0.095000  0.820000 1.305000 1.020000 ;
      RECT 0.095000  2.030000 1.305000 2.205000 ;
      RECT 0.095000  2.205000 0.400000 2.725000 ;
      RECT 0.575000  2.380000 0.905000 3.245000 ;
      RECT 0.585000  0.085000 0.915000 0.650000 ;
      RECT 0.975000  1.020000 1.305000 2.030000 ;
      RECT 1.415000  2.650000 1.745000 2.900000 ;
      RECT 1.475000  0.305000 1.720000 1.140000 ;
      RECT 1.475000  1.140000 2.510000 1.470000 ;
      RECT 1.475000  1.470000 1.745000 2.650000 ;
      RECT 1.915000  0.085000 2.265000 0.745000 ;
      RECT 1.915000  1.940000 2.265000 3.245000 ;
      RECT 2.800000  0.415000 2.970000 1.220000 ;
      RECT 2.800000  1.220000 4.005000 1.390000 ;
      RECT 2.800000  1.390000 2.970000 2.980000 ;
      RECT 3.370000  0.400000 3.700000 0.880000 ;
      RECT 3.370000  0.880000 4.700000 0.925000 ;
      RECT 3.370000  0.925000 4.755000 1.050000 ;
      RECT 3.415000  1.560000 4.755000 1.730000 ;
      RECT 3.415000  1.730000 3.655000 2.980000 ;
      RECT 4.330000  0.085000 4.660000 0.670000 ;
      RECT 4.330000  1.900000 4.660000 3.245000 ;
      RECT 4.530000  1.050000 4.755000 1.560000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
  END
END sky130_fd_sc_hs__clkdlyinv5sd3_1
MACRO sky130_fd_sc_hs__clkinv_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.440000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 0.755000 1.780000 ;
        RECT 0.425000 0.920000 0.755000 1.180000 ;
        RECT 0.425000 1.780000 0.755000 1.930000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.477350 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.555000 2.100000 1.325000 2.430000 ;
        RECT 0.555000 2.430000 0.835000 2.955000 ;
        RECT 0.615000 0.350000 1.325000 0.680000 ;
        RECT 1.085000 0.680000 1.325000 2.100000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 1.440000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 1.440000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.440000 0.085000 ;
      RECT 0.000000  3.245000 1.440000 3.415000 ;
      RECT 0.105000  2.100000 0.355000 3.245000 ;
      RECT 0.115000  0.085000 0.445000 0.750000 ;
      RECT 1.005000  2.600000 1.335000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
  END
END sky130_fd_sc_hs__clkinv_1
MACRO sky130_fd_sc_hs__clkinv_16
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.52000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  5.040000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.985000 1.180000 10.935000 1.410000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  5.040000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.575000 1.920000 10.935000 2.150000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.520000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 11.520000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.520000 0.085000 ;
      RECT  0.000000  3.245000 11.520000 3.415000 ;
      RECT  0.115000  0.085000  0.445000 0.840000 ;
      RECT  0.115000  1.900000  0.445000 3.245000 ;
      RECT  0.615000  0.380000  0.805000 0.775000 ;
      RECT  0.625000  0.775000  0.805000 1.820000 ;
      RECT  0.625000  1.820000  0.815000 2.980000 ;
      RECT  0.975000  0.085000  1.260000 0.840000 ;
      RECT  0.975000  1.150000  1.295000 1.650000 ;
      RECT  1.015000  1.820000  1.265000 3.245000 ;
      RECT  1.440000  0.380000  1.700000 0.775000 ;
      RECT  1.465000  0.775000  1.695000 1.885000 ;
      RECT  1.465000  1.885000  1.795000 2.980000 ;
      RECT  1.865000  1.150000  2.195000 1.650000 ;
      RECT  1.885000  0.085000  2.165000 0.840000 ;
      RECT  1.995000  1.820000  2.165000 3.245000 ;
      RECT  2.350000  0.380000  2.665000 0.775000 ;
      RECT  2.365000  0.775000  2.665000 1.885000 ;
      RECT  2.365000  1.885000  2.695000 2.980000 ;
      RECT  2.835000  1.150000  3.165000 1.650000 ;
      RECT  2.845000  0.085000  3.095000 0.840000 ;
      RECT  2.895000  1.820000  3.065000 3.245000 ;
      RECT  3.300000  0.380000  3.595000 0.775000 ;
      RECT  3.335000  0.775000  3.595000 2.980000 ;
      RECT  3.765000  0.085000  4.095000 0.840000 ;
      RECT  3.765000  1.150000  4.095000 1.650000 ;
      RECT  3.795000  1.820000  3.965000 3.245000 ;
      RECT  4.165000  1.850000  4.525000 1.900000 ;
      RECT  4.165000  1.900000  4.495000 2.980000 ;
      RECT  4.265000  0.380000  4.525000 1.850000 ;
      RECT  4.695000  1.820000  4.865000 3.245000 ;
      RECT  4.755000  1.150000  5.085000 1.650000 ;
      RECT  4.765000  0.085000  5.085000 0.840000 ;
      RECT  5.065000  1.850000  5.425000 2.010000 ;
      RECT  5.065000  2.010000  5.395000 2.980000 ;
      RECT  5.255000  0.380000  5.525000 0.775000 ;
      RECT  5.255000  0.775000  5.425000 1.850000 ;
      RECT  5.595000  1.150000  5.925000 1.650000 ;
      RECT  5.595000  1.820000  5.845000 3.245000 ;
      RECT  5.695000  0.085000  5.980000 0.840000 ;
      RECT  6.015000  1.820000  6.330000 2.980000 ;
      RECT  6.095000  1.010000  6.340000 1.760000 ;
      RECT  6.095000  1.760000  6.330000 1.820000 ;
      RECT  6.160000  0.380000  6.385000 0.785000 ;
      RECT  6.160000  0.785000  6.340000 1.010000 ;
      RECT  6.510000  1.820000  6.795000 3.245000 ;
      RECT  6.545000  1.150000  6.875000 1.650000 ;
      RECT  6.555000  0.085000  6.875000 0.840000 ;
      RECT  7.045000  0.380000  7.290000 2.980000 ;
      RECT  7.475000  1.820000  7.805000 3.245000 ;
      RECT  7.485000  0.085000  9.825000 0.710000 ;
      RECT  7.525000  1.150000 10.915000 1.650000 ;
      RECT  8.005000  1.820000  8.175000 2.980000 ;
      RECT  8.375000  1.820000  8.625000 3.245000 ;
      RECT  8.905000  1.820000  9.075000 2.980000 ;
      RECT  9.275000  1.820000  9.605000 3.245000 ;
      RECT  9.805000  1.820000  9.975000 2.980000 ;
      RECT 10.175000  1.820000 10.505000 3.245000 ;
      RECT 10.705000  1.820000 10.875000 2.980000 ;
      RECT 11.075000  1.820000 11.405000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  1.950000  0.805000 2.120000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.045000  1.210000  1.215000 1.380000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.545000  1.950000  1.715000 2.120000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  1.945000  1.210000  2.115000 1.380000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.445000  1.950000  2.615000 2.120000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  2.915000  1.210000  3.085000 1.380000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.375000  1.950000  3.545000 2.120000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.845000  1.210000  4.015000 1.380000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.245000  1.950000  4.415000 2.120000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.835000  1.210000  5.005000 1.380000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.145000  1.950000  5.315000 2.120000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.675000  1.210000  5.845000 1.380000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.095000  1.950000  6.265000 2.120000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.625000  1.210000  6.795000 1.380000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.075000  1.950000  7.245000 2.120000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.745000  1.210000  7.915000 1.380000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.005000  1.950000  8.175000 2.120000 ;
      RECT  8.105000  1.210000  8.275000 1.380000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.465000  1.210000  8.635000 1.380000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  8.825000  1.210000  8.995000 1.380000 ;
      RECT  8.905000  1.950000  9.075000 2.120000 ;
      RECT  9.185000  1.210000  9.355000 1.380000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.545000  1.210000  9.715000 1.380000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT  9.805000  1.950000  9.975000 2.120000 ;
      RECT  9.905000  1.210000 10.075000 1.380000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.265000  1.210000 10.435000 1.380000 ;
      RECT 10.625000  1.210000 10.795000 1.380000 ;
      RECT 10.705000  1.950000 10.875000 2.120000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
  END
END sky130_fd_sc_hs__clkinv_16
MACRO sky130_fd_sc_hs__clkinv_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.920000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.315000 1.780000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.994000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.120000 1.950000 1.795000 2.120000 ;
        RECT 0.120000 2.120000 0.450000 2.980000 ;
        RECT 0.615000 0.510000 1.305000 1.010000 ;
        RECT 0.615000 1.010000 1.795000 1.180000 ;
        RECT 1.020000 2.120000 1.350000 2.980000 ;
        RECT 1.565000 1.180000 1.795000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 1.920000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 1.920000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.920000 0.085000 ;
      RECT 0.000000  3.245000 1.920000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 0.840000 ;
      RECT 0.650000  2.290000 0.820000 3.245000 ;
      RECT 1.475000  0.085000 1.805000 0.840000 ;
      RECT 1.550000  2.290000 1.800000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
  END
END sky130_fd_sc_hs__clkinv_2
MACRO sky130_fd_sc_hs__clkinv_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.350000 2.755000 1.780000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  1.432200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.265000 1.010000 3.235000 1.180000 ;
        RECT 0.265000 1.180000 0.435000 1.950000 ;
        RECT 0.265000 1.950000 3.235000 2.120000 ;
        RECT 0.565000 2.120000 0.895000 2.980000 ;
        RECT 0.990000 0.455000 1.745000 1.010000 ;
        RECT 1.465000 2.120000 1.795000 2.980000 ;
        RECT 2.415000 0.380000 2.745000 1.010000 ;
        RECT 2.415000 2.120000 2.745000 2.980000 ;
        RECT 3.005000 1.180000 3.235000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.115000  0.085000 0.820000 0.710000 ;
      RECT 0.115000  2.290000 0.365000 3.245000 ;
      RECT 1.095000  2.290000 1.265000 3.245000 ;
      RECT 1.915000  0.085000 2.245000 0.840000 ;
      RECT 1.995000  2.290000 2.245000 3.245000 ;
      RECT 2.915000  0.085000 3.245000 0.840000 ;
      RECT 2.915000  2.290000 3.245000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__clkinv_4
MACRO sky130_fd_sc_hs__clkinv_8
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  2.520000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.625000 1.350000 5.715000 1.780000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  3.242400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.285000 1.010000 6.115000 1.180000 ;
        RECT 0.285000 1.180000 0.455000 1.950000 ;
        RECT 0.285000 1.950000 6.115000 2.120000 ;
        RECT 0.590000 2.120000 0.920000 2.980000 ;
        RECT 0.615000 0.460000 2.625000 1.010000 ;
        RECT 1.540000 2.120000 1.870000 2.980000 ;
        RECT 2.490000 2.120000 2.820000 2.980000 ;
        RECT 3.295000 0.445000 3.625000 1.010000 ;
        RECT 3.440000 2.120000 3.770000 2.980000 ;
        RECT 4.295000 0.445000 4.625000 1.010000 ;
        RECT 4.390000 2.120000 4.720000 2.980000 ;
        RECT 5.295000 0.445000 5.625000 1.010000 ;
        RECT 5.340000 2.120000 5.670000 2.980000 ;
        RECT 5.885000 1.180000 6.115000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.240000 0.085000 ;
      RECT 0.000000  3.245000 6.240000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 0.775000 ;
      RECT 0.115000  2.290000 0.390000 3.245000 ;
      RECT 1.120000  2.290000 1.370000 3.245000 ;
      RECT 2.070000  2.290000 2.320000 3.245000 ;
      RECT 2.795000  0.085000 3.125000 0.775000 ;
      RECT 3.020000  2.290000 3.270000 3.245000 ;
      RECT 3.795000  0.085000 4.125000 0.775000 ;
      RECT 3.970000  2.290000 4.220000 3.245000 ;
      RECT 4.795000  0.085000 5.125000 0.775000 ;
      RECT 4.920000  2.290000 5.170000 3.245000 ;
      RECT 5.795000  0.085000 6.125000 0.775000 ;
      RECT 5.870000  2.290000 6.120000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
  END
END sky130_fd_sc_hs__clkinv_8
MACRO sky130_fd_sc_hs__conb_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.440000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN HI
    ANTENNAPARTIALMETALSIDEAREA  0.182000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.615000 0.845000 ;
        RECT 0.085000 0.845000 0.395000 2.335000 ;
    END
  END HI
  PIN LO
    ANTENNAPARTIALMETALSIDEAREA  0.182000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.825000 2.485000 1.355000 3.075000 ;
        RECT 1.055000 0.995000 1.355000 2.485000 ;
    END
  END LO
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 1.440000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 1.440000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.440000 0.085000 ;
      RECT 0.000000  3.245000 1.440000 3.415000 ;
      RECT 0.285000  2.505000 0.615000 3.245000 ;
      RECT 0.825000  0.085000 1.155000 0.825000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
  END
END sky130_fd_sc_hs__conb_1
MACRO sky130_fd_sc_hs__decap_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.920000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 1.920000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 1.920000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.920000 0.085000 ;
      RECT 0.000000  3.245000 1.920000 3.415000 ;
      RECT 0.240000  0.085000 0.855000 0.715000 ;
      RECT 0.240000  2.670000 0.490000 3.245000 ;
      RECT 0.605000  0.715000 0.855000 1.585000 ;
      RECT 1.065000  1.250000 1.315000 2.670000 ;
      RECT 1.065000  2.670000 1.680000 3.245000 ;
      RECT 1.425000  0.085000 1.680000 0.715000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
  END
END sky130_fd_sc_hs__decap_4
MACRO sky130_fd_sc_hs__decap_8
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.565000  0.085000 1.130000 0.810000 ;
      RECT 0.565000  2.285000 0.815000 3.245000 ;
      RECT 0.800000  0.810000 1.130000 1.585000 ;
      RECT 1.460000  1.250000 2.395000 3.245000 ;
      RECT 1.765000  0.085000 2.095000 0.805000 ;
      RECT 2.670000  0.085000 3.290000 0.810000 ;
      RECT 2.670000  0.810000 3.075000 1.585000 ;
      RECT 3.050000  2.295000 3.300000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__decap_8
MACRO sky130_fd_sc_hs__dfbbn_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.44000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.925000 1.180000 2.755000 1.510000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.519000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.005000 0.350000 13.340000 2.980000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.513400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.555000 0.405000 11.925000 1.150000 ;
        RECT 11.575000 1.820000 11.925000 2.980000 ;
        RECT 11.755000 1.150000 11.925000 1.820000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.685000 1.350000 11.015000 1.780000 ;
    END
  END RESET_B
  PIN SET_B
    ANTENNAPARTIALMETALSIDEAREA  2.541000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 5.375000 1.920000 5.665000 1.965000 ;
        RECT 5.375000 1.965000 9.025000 2.105000 ;
        RECT 5.375000 2.105000 5.665000 2.150000 ;
        RECT 8.735000 1.920000 9.025000 1.965000 ;
        RECT 8.735000 2.105000 9.025000 2.150000 ;
    END
  END SET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.495000 1.780000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 13.440000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 13.440000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.440000 0.085000 ;
      RECT  0.000000  3.245000 13.440000 3.415000 ;
      RECT  0.105000  1.950000  0.835000 2.120000 ;
      RECT  0.105000  2.120000  0.435000 2.980000 ;
      RECT  0.115000  0.350000  0.365000 0.960000 ;
      RECT  0.115000  0.960000  0.835000 1.130000 ;
      RECT  0.545000  0.085000  0.875000 0.790000 ;
      RECT  0.635000  2.290000  0.805000 3.245000 ;
      RECT  0.665000  1.130000  0.835000 1.300000 ;
      RECT  0.665000  1.300000  1.075000 1.630000 ;
      RECT  0.665000  1.630000  0.835000 1.950000 ;
      RECT  1.005000  1.820000  1.415000 2.905000 ;
      RECT  1.005000  2.905000  2.125000 3.075000 ;
      RECT  1.055000  0.350000  1.415000 1.130000 ;
      RECT  1.245000  1.130000  1.415000 1.820000 ;
      RECT  1.585000  0.575000  1.865000 0.840000 ;
      RECT  1.585000  0.840000  2.750000 1.010000 ;
      RECT  1.585000  1.010000  1.755000 2.405000 ;
      RECT  1.585000  2.405000  1.785000 2.735000 ;
      RECT  1.955000  1.685000  3.240000 1.855000 ;
      RECT  1.955000  1.855000  2.125000 2.905000 ;
      RECT  2.045000  0.085000  2.410000 0.670000 ;
      RECT  2.295000  2.525000  2.465000 3.245000 ;
      RECT  2.370000  2.025000  2.805000 2.355000 ;
      RECT  2.580000  0.255000  4.145000 0.425000 ;
      RECT  2.580000  0.425000  2.750000 0.840000 ;
      RECT  2.635000  2.355000  2.805000 2.905000 ;
      RECT  2.635000  2.905000  4.530000 3.075000 ;
      RECT  2.950000  0.595000  3.280000 0.785000 ;
      RECT  2.950000  0.785000  3.805000 0.955000 ;
      RECT  2.975000  1.125000  3.465000 1.455000 ;
      RECT  2.975000  1.455000  3.240000 1.685000 ;
      RECT  2.975000  1.855000  3.240000 2.355000 ;
      RECT  3.090000  2.565000  3.580000 2.735000 ;
      RECT  3.410000  1.625000  4.135000 1.795000 ;
      RECT  3.410000  1.795000  3.580000 2.565000 ;
      RECT  3.460000  0.425000  4.145000 0.615000 ;
      RECT  3.635000  0.955000  3.805000 1.395000 ;
      RECT  3.635000  1.395000  4.135000 1.625000 ;
      RECT  3.750000  1.965000  4.475000 2.135000 ;
      RECT  3.750000  2.135000  4.000000 2.735000 ;
      RECT  3.975000  0.615000  4.145000 0.995000 ;
      RECT  3.975000  0.995000  4.475000 1.165000 ;
      RECT  4.200000  2.305000  4.815000 2.320000 ;
      RECT  4.200000  2.320000  6.450000 2.490000 ;
      RECT  4.200000  2.490000  4.530000 2.905000 ;
      RECT  4.305000  1.165000  4.475000 1.965000 ;
      RECT  4.315000  0.255000  5.645000 0.425000 ;
      RECT  4.315000  0.425000  4.645000 0.825000 ;
      RECT  4.645000  0.995000  5.145000 1.165000 ;
      RECT  4.645000  1.165000  4.815000 2.305000 ;
      RECT  4.815000  0.715000  5.145000 0.995000 ;
      RECT  4.985000  1.335000  6.485000 1.505000 ;
      RECT  4.985000  1.505000  5.265000 1.665000 ;
      RECT  5.040000  2.660000  5.370000 3.245000 ;
      RECT  5.315000  0.425000  5.645000 1.035000 ;
      RECT  5.435000  1.675000  5.850000 1.960000 ;
      RECT  5.435000  1.960000  5.635000 2.150000 ;
      RECT  5.570000  2.490000  5.820000 2.980000 ;
      RECT  5.815000  0.085000  6.145000 1.035000 ;
      RECT  6.020000  2.660000  6.350000 3.245000 ;
      RECT  6.120000  1.675000  6.450000 2.320000 ;
      RECT  6.315000  0.340000  8.545000 0.510000 ;
      RECT  6.315000  0.510000  6.485000 1.335000 ;
      RECT  6.710000  1.180000  7.865000 1.560000 ;
      RECT  6.710000  1.560000  7.075000 1.930000 ;
      RECT  6.720000  0.680000  8.205000 1.010000 ;
      RECT  6.860000  2.100000  7.415000 2.980000 ;
      RECT  7.245000  1.730000  8.560000 1.900000 ;
      RECT  7.245000  1.900000  7.415000 2.100000 ;
      RECT  7.890000  2.070000  8.220000 2.630000 ;
      RECT  7.890000  2.630000 10.320000 2.800000 ;
      RECT  7.905000  2.970000  8.270000 3.245000 ;
      RECT  8.035000  1.010000  8.205000 1.730000 ;
      RECT  8.375000  0.510000  8.545000 0.935000 ;
      RECT  8.375000  0.935000 10.890000 1.105000 ;
      RECT  8.390000  1.900000  8.560000 2.290000 ;
      RECT  8.390000  2.290000  9.400000 2.460000 ;
      RECT  8.500000  2.800000  8.830000 2.980000 ;
      RECT  8.715000  0.085000  8.885000 0.765000 ;
      RECT  8.730000  1.275000  9.060000 2.120000 ;
      RECT  9.035000  2.970000  9.365000 3.245000 ;
      RECT  9.065000  0.255000 10.360000 0.425000 ;
      RECT  9.065000  0.425000  9.315000 0.765000 ;
      RECT  9.230000  1.950000 10.170000 2.120000 ;
      RECT  9.230000  2.120000  9.400000 2.290000 ;
      RECT  9.300000  1.105000  9.630000 1.560000 ;
      RECT  9.495000  0.595000 11.385000 0.765000 ;
      RECT  9.840000  1.420000 10.170000 1.950000 ;
      RECT  9.990000  2.290000 11.385000 2.460000 ;
      RECT  9.990000  2.460000 10.320000 2.630000 ;
      RECT  9.990000  2.800000 10.320000 2.980000 ;
      RECT 10.345000  1.105000 10.515000 1.950000 ;
      RECT 10.345000  1.950000 10.850000 2.120000 ;
      RECT 11.045000  2.630000 11.375000 3.245000 ;
      RECT 11.055000  0.085000 11.385000 0.425000 ;
      RECT 11.215000  0.765000 11.385000 1.320000 ;
      RECT 11.215000  1.320000 11.585000 1.650000 ;
      RECT 11.215000  1.650000 11.385000 2.290000 ;
      RECT 12.110000  0.350000 12.360000 1.255000 ;
      RECT 12.110000  1.255000 12.835000 1.585000 ;
      RECT 12.110000  1.585000 12.360000 2.910000 ;
      RECT 12.555000  1.820000 12.805000 3.245000 ;
      RECT 12.580000  0.085000 12.830000 0.810000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  1.210000  3.205000 1.380000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  1.950000  5.605000 2.120000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  1.210000  7.045000 1.380000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  1.950000  8.965000 2.120000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
    LAYER met1 ;
      RECT 2.975000 1.180000 3.265000 1.225000 ;
      RECT 2.975000 1.225000 7.105000 1.365000 ;
      RECT 2.975000 1.365000 3.265000 1.410000 ;
      RECT 6.815000 1.180000 7.105000 1.225000 ;
      RECT 6.815000 1.365000 7.105000 1.410000 ;
  END
END sky130_fd_sc_hs__dfbbn_1
MACRO sky130_fd_sc_hs__dfbbn_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.40000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.955000 1.180000 2.755000 1.510000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.515000 1.770000 14.035000 1.940000 ;
        RECT 13.515000 1.940000 13.845000 2.980000 ;
        RECT 13.540000 0.350000 13.800000 0.850000 ;
        RECT 13.540000 0.850000 14.035000 1.100000 ;
        RECT 13.865000 1.100000 14.035000 1.770000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.630000 0.440000 11.985000 1.180000 ;
        RECT 11.645000 1.850000 11.985000 2.020000 ;
        RECT 11.645000 2.020000 11.815000 2.980000 ;
        RECT 11.815000 1.180000 11.985000 1.850000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.715000 1.350000 11.115000 1.780000 ;
    END
  END RESET_B
  PIN SET_B
    ANTENNAPARTIALMETALSIDEAREA  2.541000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 5.375000 1.920000 5.665000 1.965000 ;
        RECT 5.375000 1.965000 9.025000 2.105000 ;
        RECT 5.375000 2.105000 5.665000 2.150000 ;
        RECT 8.735000 1.920000 9.025000 1.965000 ;
        RECT 8.735000 2.105000 9.025000 2.150000 ;
    END
  END SET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.495000 1.780000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 14.400000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 14.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.400000 0.085000 ;
      RECT  0.000000  3.245000 14.400000 3.415000 ;
      RECT  0.105000  1.950000  0.835000 2.120000 ;
      RECT  0.105000  2.120000  0.435000 2.980000 ;
      RECT  0.115000  0.350000  0.365000 0.960000 ;
      RECT  0.115000  0.960000  0.835000 1.130000 ;
      RECT  0.545000  0.085000  0.875000 0.790000 ;
      RECT  0.635000  2.290000  0.805000 3.245000 ;
      RECT  0.665000  1.130000  0.835000 1.300000 ;
      RECT  0.665000  1.300000  1.105000 1.630000 ;
      RECT  0.665000  1.630000  0.835000 1.950000 ;
      RECT  1.005000  1.820000  1.445000 2.905000 ;
      RECT  1.005000  2.905000  2.125000 3.075000 ;
      RECT  1.055000  0.350000  1.445000 1.130000 ;
      RECT  1.275000  1.130000  1.445000 1.820000 ;
      RECT  1.615000  0.575000  1.865000 0.840000 ;
      RECT  1.615000  0.840000  2.780000 1.010000 ;
      RECT  1.615000  1.010000  1.785000 2.735000 ;
      RECT  1.955000  1.685000  3.230000 1.855000 ;
      RECT  1.955000  1.855000  2.125000 2.905000 ;
      RECT  2.045000  0.085000  2.440000 0.670000 ;
      RECT  2.295000  2.525000  2.465000 3.245000 ;
      RECT  2.365000  2.025000  2.805000 2.355000 ;
      RECT  2.610000  0.255000  4.225000 0.425000 ;
      RECT  2.610000  0.425000  2.780000 0.840000 ;
      RECT  2.635000  2.355000  2.805000 2.905000 ;
      RECT  2.635000  2.905000  4.605000 3.075000 ;
      RECT  2.975000  1.855000  3.230000 2.355000 ;
      RECT  2.980000  0.595000  3.310000 0.785000 ;
      RECT  2.980000  0.785000  3.885000 0.955000 ;
      RECT  3.005000  1.125000  3.545000 1.455000 ;
      RECT  3.005000  1.455000  3.230000 1.685000 ;
      RECT  3.085000  2.565000  3.570000 2.735000 ;
      RECT  3.400000  1.625000  4.095000 1.795000 ;
      RECT  3.400000  1.795000  3.570000 2.565000 ;
      RECT  3.490000  0.425000  4.225000 0.615000 ;
      RECT  3.715000  0.955000  3.885000 1.465000 ;
      RECT  3.715000  1.465000  4.095000 1.625000 ;
      RECT  3.740000  1.965000  4.435000 2.135000 ;
      RECT  3.740000  2.135000  3.990000 2.735000 ;
      RECT  4.055000  0.615000  4.225000 1.125000 ;
      RECT  4.055000  1.125000  4.435000 1.295000 ;
      RECT  4.185000  2.305000  4.775000 2.320000 ;
      RECT  4.185000  2.320000  6.380000 2.490000 ;
      RECT  4.185000  2.490000  4.605000 2.905000 ;
      RECT  4.265000  1.295000  4.435000 1.965000 ;
      RECT  4.395000  0.265000  5.575000 0.435000 ;
      RECT  4.395000  0.435000  4.565000 0.955000 ;
      RECT  4.605000  1.125000  4.905000 1.295000 ;
      RECT  4.605000  1.295000  4.775000 2.305000 ;
      RECT  4.735000  0.605000  5.075000 1.120000 ;
      RECT  4.735000  1.120000  4.905000 1.125000 ;
      RECT  4.945000  1.610000  5.245000 1.940000 ;
      RECT  5.055000  2.660000  5.385000 3.245000 ;
      RECT  5.075000  1.290000  6.415000 1.460000 ;
      RECT  5.075000  1.460000  5.245000 1.610000 ;
      RECT  5.245000  0.435000  5.575000 1.025000 ;
      RECT  5.415000  1.630000  5.745000 2.150000 ;
      RECT  5.565000  2.490000  5.895000 2.980000 ;
      RECT  5.745000  0.085000  6.075000 1.025000 ;
      RECT  6.050000  1.630000  6.380000 2.320000 ;
      RECT  6.095000  2.660000  6.425000 3.245000 ;
      RECT  6.245000  0.340000  8.615000 0.510000 ;
      RECT  6.245000  0.510000  6.415000 1.290000 ;
      RECT  6.650000  0.680000  8.275000 1.010000 ;
      RECT  6.785000  1.180000  7.935000 1.410000 ;
      RECT  6.785000  1.410000  7.115000 1.910000 ;
      RECT  6.965000  2.100000  7.455000 2.980000 ;
      RECT  7.285000  1.720000  8.595000 1.890000 ;
      RECT  7.285000  1.890000  7.455000 2.100000 ;
      RECT  7.685000  1.410000  7.935000 1.550000 ;
      RECT  7.925000  2.060000  8.255000 2.630000 ;
      RECT  7.925000  2.630000 10.390000 2.800000 ;
      RECT  8.010000  2.970000  8.340000 3.245000 ;
      RECT  8.105000  1.010000  8.275000 1.720000 ;
      RECT  8.425000  1.890000  8.595000 2.290000 ;
      RECT  8.425000  2.290000  9.890000 2.460000 ;
      RECT  8.445000  0.510000  8.615000 1.010000 ;
      RECT  8.445000  1.010000 10.990000 1.180000 ;
      RECT  8.570000  2.800000  8.900000 2.980000 ;
      RECT  8.765000  1.450000  9.160000 1.780000 ;
      RECT  8.765000  1.780000  8.995000 2.120000 ;
      RECT  8.785000  0.085000  8.955000 0.840000 ;
      RECT  9.105000  2.970000  9.435000 3.245000 ;
      RECT  9.135000  0.255000 10.440000 0.425000 ;
      RECT  9.135000  0.425000  9.385000 0.840000 ;
      RECT  9.370000  1.180000  9.700000 1.550000 ;
      RECT  9.605000  0.595000  9.935000 0.670000 ;
      RECT  9.605000  0.670000 11.460000 0.840000 ;
      RECT  9.720000  1.720000 10.205000 1.890000 ;
      RECT  9.720000  1.890000  9.890000 2.290000 ;
      RECT  9.910000  1.470000 10.205000 1.720000 ;
      RECT 10.060000  2.290000 11.460000 2.460000 ;
      RECT 10.060000  2.460000 10.390000 2.630000 ;
      RECT 10.060000  2.800000 10.390000 2.980000 ;
      RECT 10.110000  0.425000 10.440000 0.500000 ;
      RECT 10.375000  1.180000 10.545000 1.950000 ;
      RECT 10.375000  1.950000 10.920000 2.120000 ;
      RECT 10.665000  0.085000 11.450000 0.500000 ;
      RECT 11.115000  2.630000 11.445000 3.245000 ;
      RECT 11.290000  0.840000 11.460000 1.350000 ;
      RECT 11.290000  1.350000 11.645000 1.680000 ;
      RECT 11.290000  1.680000 11.460000 2.290000 ;
      RECT 12.015000  2.190000 12.345000 3.245000 ;
      RECT 12.155000  0.085000 12.405000 1.260000 ;
      RECT 12.545000  1.820000 12.875000 2.860000 ;
      RECT 12.635000  0.350000 12.885000 1.270000 ;
      RECT 12.635000  1.270000 13.695000 1.600000 ;
      RECT 12.635000  1.600000 12.875000 1.820000 ;
      RECT 13.065000  1.820000 13.315000 3.245000 ;
      RECT 13.095000  0.085000 13.370000 1.050000 ;
      RECT 13.970000  0.085000 14.300000 0.680000 ;
      RECT 14.045000  2.110000 14.295000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  1.210000  3.205000 1.380000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  1.950000  5.605000 2.120000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  1.210000  7.045000 1.380000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  1.950000  8.965000 2.120000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
    LAYER met1 ;
      RECT 2.975000 1.180000 3.265000 1.225000 ;
      RECT 2.975000 1.225000 7.105000 1.365000 ;
      RECT 2.975000 1.365000 3.265000 1.410000 ;
      RECT 6.815000 1.180000 7.105000 1.225000 ;
      RECT 6.815000 1.365000 7.105000 1.410000 ;
  END
END sky130_fd_sc_hs__dfbbn_2
MACRO sky130_fd_sc_hs__dfbbp_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.96000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.960000 1.825000 2.290000 2.155000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.519000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.525000 0.350000 12.860000 2.980000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.518900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.065000 0.350000 11.460000 1.130000 ;
        RECT 11.120000 1.820000 11.460000 2.980000 ;
        RECT 11.290000 1.130000 11.460000 1.820000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.235000 0.980000 10.580000 1.650000 ;
    END
  END RESET_B
  PIN SET_B
    ANTENNAGATEAREA  0.470000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.230000 1.410000 4.560000 1.655000 ;
        RECT 4.360000 1.655000 4.530000 2.905000 ;
        RECT 4.360000 2.905000 5.330000 3.075000 ;
        RECT 5.160000 2.165000 6.210000 2.335000 ;
        RECT 5.160000 2.335000 5.330000 2.905000 ;
        RECT 6.040000 2.335000 6.210000 2.905000 ;
        RECT 6.040000 2.905000 7.450000 3.075000 ;
        RECT 7.280000 1.740000 8.570000 1.800000 ;
        RECT 7.280000 1.800000 8.515000 1.910000 ;
        RECT 7.280000 1.910000 7.450000 2.905000 ;
        RECT 8.240000 1.470000 8.570000 1.740000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.180000 0.805000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.960000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 12.960000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.960000 0.085000 ;
      RECT  0.000000  3.245000 12.960000 3.415000 ;
      RECT  0.085000  0.350000  0.445000 1.010000 ;
      RECT  0.085000  1.010000  0.255000 1.720000 ;
      RECT  0.085000  1.720000  1.145000 1.890000 ;
      RECT  0.085000  1.890000  0.535000 2.980000 ;
      RECT  0.615000  0.085000  0.945000 1.010000 ;
      RECT  0.705000  2.060000  1.035000 3.245000 ;
      RECT  0.975000  1.300000  1.145000 1.720000 ;
      RECT  1.125000  0.350000  1.485000 1.130000 ;
      RECT  1.315000  1.130000  1.485000 1.255000 ;
      RECT  1.315000  1.255000  2.615000 1.585000 ;
      RECT  1.315000  1.585000  1.565000 2.980000 ;
      RECT  1.655000  0.085000  1.905000 1.065000 ;
      RECT  1.805000  2.425000  2.410000 3.245000 ;
      RECT  2.085000  0.605000  2.335000 0.915000 ;
      RECT  2.085000  0.915000  2.955000 1.085000 ;
      RECT  2.575000  0.415000  3.295000 0.745000 ;
      RECT  2.580000  2.295000  2.955000 2.755000 ;
      RECT  2.785000  1.085000  2.955000 2.295000 ;
      RECT  3.125000  0.745000  3.295000 1.625000 ;
      RECT  3.125000  1.625000  4.060000 1.795000 ;
      RECT  3.125000  1.795000  3.430000 2.335000 ;
      RECT  3.465000  0.730000  5.335000 0.840000 ;
      RECT  3.465000  0.840000  6.020000 0.900000 ;
      RECT  3.465000  0.900000  3.720000 1.455000 ;
      RECT  3.560000  0.085000  4.155000 0.560000 ;
      RECT  3.890000  1.070000  4.915000 1.240000 ;
      RECT  3.890000  1.240000  4.060000 1.625000 ;
      RECT  3.940000  1.965000  4.190000 3.245000 ;
      RECT  4.415000  0.255000  5.840000 0.425000 ;
      RECT  4.415000  0.425000  4.825000 0.560000 ;
      RECT  4.700000  1.825000  6.020000 1.995000 ;
      RECT  4.700000  1.995000  4.950000 2.735000 ;
      RECT  4.745000  1.240000  4.915000 1.255000 ;
      RECT  4.745000  1.255000  5.100000 1.585000 ;
      RECT  5.015000  0.595000  5.335000 0.730000 ;
      RECT  5.085000  0.900000  6.020000 1.010000 ;
      RECT  5.310000  1.180000  5.640000 1.585000 ;
      RECT  5.500000  2.505000  5.870000 3.245000 ;
      RECT  5.510000  0.425000  5.840000 0.670000 ;
      RECT  5.850000  1.010000  6.020000 1.255000 ;
      RECT  5.850000  1.255000  6.180000 1.585000 ;
      RECT  5.850000  1.585000  6.020000 1.825000 ;
      RECT  6.060000  0.085000  6.430000 0.670000 ;
      RECT  6.190000  0.670000  6.430000 1.085000 ;
      RECT  6.440000  1.610000  6.770000 1.940000 ;
      RECT  6.540000  2.110000  7.110000 2.280000 ;
      RECT  6.540000  2.280000  6.870000 2.735000 ;
      RECT  6.600000  0.255000  7.670000 0.425000 ;
      RECT  6.600000  0.425000  6.770000 1.610000 ;
      RECT  6.940000  0.595000  7.175000 1.400000 ;
      RECT  6.940000  1.400000  8.070000 1.570000 ;
      RECT  6.940000  1.570000  7.110000 2.110000 ;
      RECT  7.345000  0.425000  7.670000 1.230000 ;
      RECT  7.620000  2.080000  9.385000 2.240000 ;
      RECT  7.620000  2.240000 10.950000 2.380000 ;
      RECT  7.620000  2.650000  8.420000 3.245000 ;
      RECT  7.900000  1.130000  9.045000 1.300000 ;
      RECT  7.900000  1.300000  8.070000 1.400000 ;
      RECT  8.085000  0.085000  8.415000 0.960000 ;
      RECT  8.585000  0.255000  9.725000 0.425000 ;
      RECT  8.585000  0.425000  8.915000 0.960000 ;
      RECT  8.685000  1.970000  9.385000 2.080000 ;
      RECT  8.685000  2.380000 10.950000 2.410000 ;
      RECT  8.685000  2.410000  8.935000 2.980000 ;
      RECT  8.780000  1.300000  9.045000 1.550000 ;
      RECT  9.085000  0.595000  9.385000 0.960000 ;
      RECT  9.215000  0.960000  9.385000 1.970000 ;
      RECT  9.470000  2.580000  9.800000 3.245000 ;
      RECT  9.555000  0.425000  9.725000 1.020000 ;
      RECT  9.710000  1.190000 10.065000 1.820000 ;
      RECT  9.710000  1.820000 10.405000 2.070000 ;
      RECT  9.895000  0.350000 10.385000 0.810000 ;
      RECT  9.895000  0.810000 10.065000 1.190000 ;
      RECT 10.565000  0.085000 10.895000 0.810000 ;
      RECT 10.590000  2.580000 10.920000 3.245000 ;
      RECT 10.780000  1.320000 11.120000 1.650000 ;
      RECT 10.780000  1.650000 10.950000 2.240000 ;
      RECT 11.640000  0.350000 11.875000 1.255000 ;
      RECT 11.640000  1.255000 12.355000 1.585000 ;
      RECT 11.640000  1.585000 11.810000 2.030000 ;
      RECT 11.640000  2.030000 11.890000 2.910000 ;
      RECT 12.055000  0.085000 12.305000 0.810000 ;
      RECT 12.075000  1.820000 12.325000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  1.210000  5.605000 1.380000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  1.210000  9.925000 1.380000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
    LAYER met1 ;
      RECT 5.375000 1.180000 5.665000 1.225000 ;
      RECT 5.375000 1.225000 9.985000 1.365000 ;
      RECT 5.375000 1.365000 5.665000 1.410000 ;
      RECT 9.695000 1.180000 9.985000 1.225000 ;
      RECT 9.695000 1.365000 9.985000 1.410000 ;
  END
END sky130_fd_sc_hs__dfbbp_1
MACRO sky130_fd_sc_hs__dfrbp_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.52000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.000000 0.520000 2.195000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.065000 0.350000 11.435000 1.130000 ;
        RECT 11.075000 1.820000 11.435000 2.980000 ;
        RECT 11.265000 1.130000 11.435000 1.820000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.951500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.260000 1.810000 9.950000 2.985000 ;
        RECT 9.560000 0.350000 9.950000 1.810000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.055000 1.920000 1.345000 1.965000 ;
        RECT 1.055000 1.965000 8.065000 2.105000 ;
        RECT 1.055000 2.105000 1.345000 2.150000 ;
        RECT 5.375000 1.920000 5.665000 1.965000 ;
        RECT 5.375000 2.105000 5.665000 2.150000 ;
        RECT 7.775000 1.920000 8.065000 1.965000 ;
        RECT 7.775000 2.105000 8.065000 2.150000 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.810000 1.310000 2.275000 1.695000 ;
        RECT 2.045000 1.695000 2.275000 1.780000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.520000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 11.520000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.520000 0.085000 ;
      RECT  0.000000  3.245000 11.520000 3.415000 ;
      RECT  0.115000  2.520000  0.365000 3.245000 ;
      RECT  0.170000  0.370000  0.500000 0.660000 ;
      RECT  0.170000  0.660000  0.860000 0.830000 ;
      RECT  0.565000  2.520000  3.345000 2.580000 ;
      RECT  0.565000  2.580000  0.890000 2.630000 ;
      RECT  0.565000  2.630000  0.845000 2.980000 ;
      RECT  0.690000  0.830000  0.860000 2.310000 ;
      RECT  0.690000  2.310000  1.425000 2.410000 ;
      RECT  0.690000  2.410000  1.530000 2.420000 ;
      RECT  0.690000  2.420000  3.345000 2.520000 ;
      RECT  1.015000  2.750000  1.345000 3.245000 ;
      RECT  1.030000  0.085000  1.280000 0.830000 ;
      RECT  1.030000  1.130000  1.300000 2.140000 ;
      RECT  1.405000  2.580000  1.965000 2.590000 ;
      RECT  1.470000  0.595000  1.920000 0.970000 ;
      RECT  1.470000  0.970000  2.560000 0.975000 ;
      RECT  1.470000  0.975000  2.775000 1.140000 ;
      RECT  1.470000  1.140000  1.640000 1.865000 ;
      RECT  1.470000  1.865000  1.825000 2.140000 ;
      RECT  1.595000  2.140000  1.825000 2.250000 ;
      RECT  1.890000  2.410000  3.345000 2.420000 ;
      RECT  2.025000  2.750000  2.355000 3.245000 ;
      RECT  2.090000  0.085000  2.420000 0.800000 ;
      RECT  2.445000  1.140000  2.775000 1.490000 ;
      RECT  2.445000  1.490000  2.805000 1.550000 ;
      RECT  2.475000  1.550000  2.805000 1.695000 ;
      RECT  2.475000  1.865000  3.500000 2.015000 ;
      RECT  2.475000  2.015000  3.050000 2.040000 ;
      RECT  2.475000  2.040000  3.025000 2.060000 ;
      RECT  2.475000  2.060000  3.020000 2.065000 ;
      RECT  2.475000  2.065000  3.000000 2.080000 ;
      RECT  2.475000  2.080000  2.975000 2.240000 ;
      RECT  2.610000  0.255000  4.520000 0.425000 ;
      RECT  2.610000  0.425000  3.115000 0.805000 ;
      RECT  2.915000  1.825000  3.500000 1.865000 ;
      RECT  2.945000  0.805000  3.115000 1.205000 ;
      RECT  2.945000  1.205000  3.160000 1.390000 ;
      RECT  2.945000  1.795000  3.500000 1.825000 ;
      RECT  2.975000  1.390000  3.160000 1.575000 ;
      RECT  2.975000  1.575000  3.500000 1.795000 ;
      RECT  3.065000  2.580000  3.345000 2.690000 ;
      RECT  3.145000  2.185000  3.840000 2.355000 ;
      RECT  3.145000  2.355000  3.345000 2.410000 ;
      RECT  3.285000  0.595000  3.535000 1.035000 ;
      RECT  3.330000  1.035000  3.535000 1.200000 ;
      RECT  3.330000  1.200000  3.840000 1.370000 ;
      RECT  3.515000  2.525000  4.270000 2.695000 ;
      RECT  3.670000  1.370000  3.840000 2.185000 ;
      RECT  3.705000  0.595000  4.180000 1.030000 ;
      RECT  4.010000  1.030000  4.180000 2.325000 ;
      RECT  4.010000  2.325000  5.325000 2.495000 ;
      RECT  4.010000  2.495000  4.270000 2.525000 ;
      RECT  4.350000  0.425000  4.520000 0.580000 ;
      RECT  4.350000  0.580000  6.255000 0.750000 ;
      RECT  4.350000  0.920000  5.915000 1.090000 ;
      RECT  4.350000  1.090000  4.630000 2.155000 ;
      RECT  4.440000  2.665000  4.785000 3.245000 ;
      RECT  4.890000  1.445000  5.560000 1.615000 ;
      RECT  4.890000  1.615000  5.060000 2.280000 ;
      RECT  4.890000  2.280000  5.105000 2.325000 ;
      RECT  4.945000  2.495000  5.325000 2.540000 ;
      RECT  4.990000  2.540000  5.325000 2.680000 ;
      RECT  4.995000  0.085000  5.325000 0.410000 ;
      RECT  5.230000  1.285000  5.560000 1.445000 ;
      RECT  5.230000  1.825000  5.610000 2.155000 ;
      RECT  5.745000  1.090000  5.915000 1.400000 ;
      RECT  5.745000  1.400000  6.480000 1.570000 ;
      RECT  5.780000  1.740000  6.030000 3.245000 ;
      RECT  6.085000  0.750000  6.255000 0.900000 ;
      RECT  6.085000  0.900000  6.820000 1.230000 ;
      RECT  6.230000  1.570000  6.480000 2.755000 ;
      RECT  6.425000  0.400000  7.160000 0.730000 ;
      RECT  6.650000  1.230000  6.820000 1.865000 ;
      RECT  6.650000  1.865000  7.325000 2.195000 ;
      RECT  6.700000  2.365000  7.665000 2.695000 ;
      RECT  6.990000  0.730000  7.160000 1.425000 ;
      RECT  6.990000  1.425000  8.630000 1.595000 ;
      RECT  7.430000  0.900000  8.970000 1.070000 ;
      RECT  7.430000  1.070000  7.760000 1.230000 ;
      RECT  7.495000  1.595000  7.665000 2.365000 ;
      RECT  7.535000  0.085000  7.995000 0.680000 ;
      RECT  7.835000  1.835000  8.300000 2.165000 ;
      RECT  7.835000  2.335000  8.060000 3.245000 ;
      RECT  8.260000  2.335000  8.640000 2.730000 ;
      RECT  8.330000  1.265000  8.630000 1.425000 ;
      RECT  8.470000  1.765000  8.970000 1.935000 ;
      RECT  8.470000  1.935000  8.640000 2.335000 ;
      RECT  8.485000  0.350000  8.970000 0.900000 ;
      RECT  8.800000  1.070000  8.970000 1.765000 ;
      RECT  8.810000  2.105000  9.025000 3.245000 ;
      RECT  9.140000  0.085000  9.390000 1.130000 ;
      RECT 10.190000  0.350000 10.440000 1.300000 ;
      RECT 10.190000  1.300000 11.095000 1.630000 ;
      RECT 10.190000  1.630000 10.440000 2.975000 ;
      RECT 10.610000  1.820000 10.905000 3.245000 ;
      RECT 10.645000  0.085000 10.895000 1.130000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  1.950000  1.285000 2.120000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  1.950000  5.605000 2.120000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  1.950000  8.005000 2.120000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
  END
END sky130_fd_sc_hs__dfrbp_1
MACRO sky130_fd_sc_hs__dfrbp_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.92000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.810000 0.515000 1.570000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.975000 1.820000 13.305000 2.980000 ;
        RECT 13.060000 0.330000 13.390000 1.130000 ;
        RECT 13.135000 1.130000 13.305000 1.820000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.895000 1.320000 11.875000 1.410000 ;
        RECT 10.895000 1.410000 11.725000 1.540000 ;
        RECT 10.895000 1.540000 11.065000 2.900000 ;
        RECT 11.195000 0.350000 11.455000 0.770000 ;
        RECT 11.195000 0.770000 11.875000 1.320000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.055000 1.550000 1.345000 1.595000 ;
        RECT 1.055000 1.595000 9.985000 1.735000 ;
        RECT 1.055000 1.735000 1.345000 1.780000 ;
        RECT 2.495000 1.550000 2.785000 1.595000 ;
        RECT 2.495000 1.735000 2.785000 1.780000 ;
        RECT 9.695000 1.550000 9.985000 1.595000 ;
        RECT 9.695000 1.735000 9.985000 1.780000 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.705000 1.180000 7.045000 1.670000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 13.920000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 13.920000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.920000 0.085000 ;
      RECT  0.000000  3.245000 13.920000 3.415000 ;
      RECT  0.115000  1.940000  0.510000 2.965000 ;
      RECT  0.115000  2.965000  1.435000 3.245000 ;
      RECT  0.325000  0.390000  0.855000 0.640000 ;
      RECT  0.680000  1.950000  1.010000 2.625000 ;
      RECT  0.680000  2.625000  1.775000 2.795000 ;
      RECT  0.685000  0.640000  0.855000 1.950000 ;
      RECT  1.025000  1.450000  1.315000 1.780000 ;
      RECT  1.145000  0.085000  1.475000 0.810000 ;
      RECT  1.485000  1.015000  3.095000 1.185000 ;
      RECT  1.485000  1.185000  1.655000 2.285000 ;
      RECT  1.485000  2.285000  1.970000 2.455000 ;
      RECT  1.605000  2.795000  1.775000 2.905000 ;
      RECT  1.605000  2.905000  2.775000 3.075000 ;
      RECT  1.645000  0.465000  1.975000 1.015000 ;
      RECT  1.825000  1.470000  2.155000 1.945000 ;
      RECT  1.825000  1.945000  4.120000 2.115000 ;
      RECT  2.185000  2.115000  2.435000 2.735000 ;
      RECT  2.205000  0.085000  2.535000 0.780000 ;
      RECT  2.385000  1.445000  2.755000 1.775000 ;
      RECT  2.605000  2.285000  3.535000 2.455000 ;
      RECT  2.605000  2.455000  2.775000 2.905000 ;
      RECT  2.705000  0.255000  5.235000 0.425000 ;
      RECT  2.705000  0.425000  2.875000 1.015000 ;
      RECT  2.925000  1.185000  3.095000 1.555000 ;
      RECT  2.925000  1.555000  3.255000 1.775000 ;
      RECT  2.945000  2.625000  3.195000 3.245000 ;
      RECT  3.045000  0.595000  4.895000 0.765000 ;
      RECT  3.345000  0.935000  4.475000 1.105000 ;
      RECT  3.345000  1.105000  3.715000 1.385000 ;
      RECT  3.365000  2.455000  3.535000 2.905000 ;
      RECT  3.365000  2.905000  4.460000 3.075000 ;
      RECT  3.790000  2.115000  4.120000 2.735000 ;
      RECT  3.885000  1.275000  4.135000 1.610000 ;
      RECT  3.885000  1.610000  4.120000 1.945000 ;
      RECT  4.290000  2.410000  4.475000 2.485000 ;
      RECT  4.290000  2.485000  4.960000 2.815000 ;
      RECT  4.290000  2.815000  4.460000 2.905000 ;
      RECT  4.305000  1.105000  4.475000 2.410000 ;
      RECT  4.645000  0.765000  4.895000 1.600000 ;
      RECT  4.645000  1.910000  5.785000 2.240000 ;
      RECT  5.065000  0.425000  5.235000 0.660000 ;
      RECT  5.065000  0.660000  6.195000 0.830000 ;
      RECT  5.095000  1.000000  5.425000 1.840000 ;
      RECT  5.095000  1.840000  5.785000 1.910000 ;
      RECT  5.425000  2.240000  5.785000 2.425000 ;
      RECT  5.425000  2.425000  7.505000 2.595000 ;
      RECT  5.425000  2.595000  5.785000 2.980000 ;
      RECT  5.595000  1.340000  6.535000 1.670000 ;
      RECT  5.605000  0.085000  5.855000 0.490000 ;
      RECT  5.990000  2.765000  6.500000 3.245000 ;
      RECT  6.025000  0.255000  8.780000 0.425000 ;
      RECT  6.025000  0.425000  6.195000 0.660000 ;
      RECT  6.095000  1.670000  6.265000 1.840000 ;
      RECT  6.095000  1.840000  7.505000 2.170000 ;
      RECT  6.365000  0.635000  6.960000 0.965000 ;
      RECT  6.365000  0.965000  6.535000 1.340000 ;
      RECT  6.705000  2.170000  7.035000 2.255000 ;
      RECT  7.215000  0.425000  7.385000 1.355000 ;
      RECT  7.215000  1.355000  7.880000 1.525000 ;
      RECT  7.315000  2.595000  7.505000 2.905000 ;
      RECT  7.315000  2.905000  8.220000 3.075000 ;
      RECT  7.555000  0.595000  9.235000 0.765000 ;
      RECT  7.555000  0.765000  7.725000 1.185000 ;
      RECT  7.710000  1.525000  7.880000 2.735000 ;
      RECT  7.905000  0.935000 10.335000 1.105000 ;
      RECT  8.050000  1.275000  8.555000 1.605000 ;
      RECT  8.050000  1.605000  8.220000 2.905000 ;
      RECT  8.390000  1.925000  8.895000 2.095000 ;
      RECT  8.390000  2.095000  8.640000 2.385000 ;
      RECT  8.725000  1.105000 10.335000 1.265000 ;
      RECT  8.725000  1.265000  8.895000 1.925000 ;
      RECT  8.985000  0.350000  9.235000 0.595000 ;
      RECT  9.065000  1.455000  9.330000 1.950000 ;
      RECT  9.065000  1.950000 10.675000 2.120000 ;
      RECT  9.265000  2.290000  9.625000 3.245000 ;
      RECT  9.415000  0.085000  9.745000 0.720000 ;
      RECT  9.540000  1.450000  9.955000 1.780000 ;
      RECT  9.830000  2.120000 10.160000 2.385000 ;
      RECT 10.205000  0.350000 10.675000 0.765000 ;
      RECT 10.365000  2.290000 10.695000 3.245000 ;
      RECT 10.505000  0.765000 10.675000 1.950000 ;
      RECT 10.845000  0.085000 11.015000 1.100000 ;
      RECT 11.265000  1.740000 11.595000 3.245000 ;
      RECT 11.625000  0.085000 11.965000 0.600000 ;
      RECT 11.895000  1.740000 12.305000 2.780000 ;
      RECT 12.135000  0.350000 12.430000 1.300000 ;
      RECT 12.135000  1.300000 12.965000 1.630000 ;
      RECT 12.135000  1.630000 12.305000 1.740000 ;
      RECT 12.475000  1.820000 12.805000 3.245000 ;
      RECT 12.630000  0.085000 12.880000 1.130000 ;
      RECT 13.475000  1.820000 13.805000 3.245000 ;
      RECT 13.560000  0.085000 13.820000 1.130000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  1.580000  1.285000 1.750000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  1.580000  2.725000 1.750000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  1.580000  9.925000 1.750000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
  END
END sky130_fd_sc_hs__dfrbp_2
MACRO sky130_fd_sc_hs__dfrtn_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.960000 0.370000 2.150000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.533800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.590000 0.440000 10.955000 1.150000 ;
        RECT 10.605000 1.820000 10.955000 2.980000 ;
        RECT 10.785000 1.150000 10.955000 1.820000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.055000 1.550000 1.345000 1.595000 ;
        RECT 1.055000 1.595000 8.545000 1.735000 ;
        RECT 1.055000 1.735000 1.345000 1.780000 ;
        RECT 4.895000 1.550000 5.185000 1.595000 ;
        RECT 4.895000 1.735000 5.185000 1.780000 ;
        RECT 8.255000 1.550000 8.545000 1.595000 ;
        RECT 8.255000 1.735000 8.545000 1.780000 ;
    END
  END RESET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.455000 1.180000 1.765000 1.650000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.040000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 11.040000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  3.245000 11.040000 3.415000 ;
      RECT  0.110000  2.520000  0.440000 3.245000 ;
      RECT  0.145000  0.350000  0.710000 0.790000 ;
      RECT  0.540000  0.790000  0.710000 2.180000 ;
      RECT  0.540000  2.180000  3.420000 2.350000 ;
      RECT  0.640000  2.350000  0.870000 2.980000 ;
      RECT  0.880000  1.245000  1.285000 1.780000 ;
      RECT  1.040000  2.520000  1.370000 3.245000 ;
      RECT  1.045000  0.085000  1.295000 0.810000 ;
      RECT  1.475000  0.350000  1.805000 0.665000 ;
      RECT  1.475000  0.665000  2.165000 1.010000 ;
      RECT  1.515000  1.820000  2.165000 2.010000 ;
      RECT  1.935000  1.010000  2.165000 1.820000 ;
      RECT  2.020000  0.085000  2.255000 0.465000 ;
      RECT  2.070000  2.520000  2.400000 3.245000 ;
      RECT  2.335000  0.625000  3.365000 0.655000 ;
      RECT  2.335000  0.655000  2.575000 0.685000 ;
      RECT  2.335000  0.685000  2.550000 0.705000 ;
      RECT  2.335000  0.705000  2.535000 0.725000 ;
      RECT  2.335000  0.725000  2.505000 2.180000 ;
      RECT  2.355000  0.605000  3.365000 0.625000 ;
      RECT  2.370000  0.595000  3.365000 0.605000 ;
      RECT  2.395000  0.565000  3.365000 0.595000 ;
      RECT  2.410000  0.545000  3.365000 0.565000 ;
      RECT  2.415000  0.525000  3.365000 0.545000 ;
      RECT  2.440000  0.485000  3.365000 0.525000 ;
      RECT  2.675000  0.825000  2.940000 1.245000 ;
      RECT  2.675000  1.245000  3.705000 2.010000 ;
      RECT  3.115000  0.655000  3.365000 1.075000 ;
      RECT  3.170000  2.350000  3.420000 2.735000 ;
      RECT  3.535000  0.255000  4.855000 0.465000 ;
      RECT  3.535000  0.465000  3.705000 1.245000 ;
      RECT  3.620000  2.180000  4.075000 2.735000 ;
      RECT  3.875000  0.635000  4.075000 1.970000 ;
      RECT  3.875000  1.970000  5.695000 2.140000 ;
      RECT  3.875000  2.140000  4.075000 2.180000 ;
      RECT  4.275000  1.130000  6.195000 1.300000 ;
      RECT  4.275000  1.300000  4.655000 1.775000 ;
      RECT  4.460000  2.310000  4.790000 3.245000 ;
      RECT  4.685000  0.465000  4.855000 0.790000 ;
      RECT  4.685000  0.790000  5.695000 0.960000 ;
      RECT  4.855000  1.470000  5.155000 1.800000 ;
      RECT  4.970000  2.140000  5.300000 2.735000 ;
      RECT  5.025000  0.085000  5.355000 0.620000 ;
      RECT  5.335000  1.470000  5.695000 1.970000 ;
      RECT  5.490000  2.360000  5.820000 3.245000 ;
      RECT  5.525000  0.255000  6.535000 0.425000 ;
      RECT  5.525000  0.425000  5.695000 0.790000 ;
      RECT  5.865000  0.595000  6.195000 1.130000 ;
      RECT  5.865000  1.300000  6.035000 1.970000 ;
      RECT  5.865000  1.970000  6.700000 2.140000 ;
      RECT  5.990000  2.140000  6.700000 2.980000 ;
      RECT  6.205000  1.470000  6.510000 1.630000 ;
      RECT  6.205000  1.630000  7.560000 1.800000 ;
      RECT  6.365000  0.425000  6.535000 1.125000 ;
      RECT  6.365000  1.125000  7.420000 1.295000 ;
      RECT  6.705000  0.625000  7.900000 0.955000 ;
      RECT  6.750000  1.295000  7.420000 1.455000 ;
      RECT  6.870000  2.535000  7.900000 2.705000 ;
      RECT  6.870000  2.705000  7.600000 2.865000 ;
      RECT  7.310000  1.800000  7.560000 2.365000 ;
      RECT  7.730000  0.955000  7.900000 1.125000 ;
      RECT  7.730000  1.125000  9.220000 1.295000 ;
      RECT  7.730000  1.295000  7.900000 2.535000 ;
      RECT  8.070000  1.965000  9.560000 2.135000 ;
      RECT  8.070000  2.135000  9.050000 2.335000 ;
      RECT  8.115000  0.085000  8.555000 0.905000 ;
      RECT  8.140000  2.520000  8.470000 3.245000 ;
      RECT  8.285000  1.465000  8.710000 1.795000 ;
      RECT  8.680000  2.335000  9.010000 2.980000 ;
      RECT  8.920000  1.295000  9.220000 1.795000 ;
      RECT  9.045000  0.575000  9.560000 0.955000 ;
      RECT  9.210000  2.520000  9.460000 3.245000 ;
      RECT  9.390000  0.955000  9.560000 1.965000 ;
      RECT  9.650000  2.305000  9.980000 2.980000 ;
      RECT  9.730000  0.530000  9.980000 1.320000 ;
      RECT  9.730000  1.320000 10.615000 1.650000 ;
      RECT  9.730000  1.650000  9.980000 2.305000 ;
      RECT 10.150000  2.100000 10.400000 3.245000 ;
      RECT 10.160000  0.085000 10.410000 1.130000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  1.580000  1.285000 1.750000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  1.580000  5.125000 1.750000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  1.580000  8.485000 1.750000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
  END
END sky130_fd_sc_hs__dfrtn_1
MACRO sky130_fd_sc_hs__dfrtp_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.000000 0.515000 2.170000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.591700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  9.725000 1.885000 10.425000 2.980000 ;
        RECT 10.165000 0.350000 10.495000 1.130000 ;
        RECT 10.165000 1.130000 10.425000 1.885000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.055000 1.920000 1.345000 1.965000 ;
        RECT 1.055000 1.965000 8.065000 2.105000 ;
        RECT 1.055000 2.105000 1.345000 2.150000 ;
        RECT 4.895000 1.920000 5.185000 1.965000 ;
        RECT 4.895000 2.105000 5.185000 2.150000 ;
        RECT 7.775000 1.920000 8.065000 1.965000 ;
        RECT 7.775000 2.105000 8.065000 2.150000 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.795000 1.310000 2.275000 1.775000 ;
        RECT 2.045000 1.775000 2.275000 1.780000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.040000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 11.040000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  3.245000 11.040000 3.415000 ;
      RECT  0.105000  2.520000  0.355000 3.245000 ;
      RECT  0.130000  0.370000  0.460000 0.660000 ;
      RECT  0.130000  0.660000  0.855000 0.830000 ;
      RECT  0.555000  2.520000  3.290000 2.560000 ;
      RECT  0.555000  2.560000  0.860000 2.605000 ;
      RECT  0.555000  2.605000  0.835000 2.640000 ;
      RECT  0.555000  2.640000  0.810000 2.980000 ;
      RECT  0.685000  0.830000  0.855000 2.310000 ;
      RECT  0.685000  2.310000  1.435000 2.335000 ;
      RECT  0.685000  2.335000  1.465000 2.360000 ;
      RECT  0.685000  2.360000  1.490000 2.375000 ;
      RECT  0.685000  2.375000  1.510000 2.390000 ;
      RECT  0.685000  2.390000  1.530000 2.410000 ;
      RECT  0.685000  2.410000  3.290000 2.520000 ;
      RECT  0.980000  2.730000  1.310000 3.245000 ;
      RECT  1.025000  1.130000  1.285000 2.140000 ;
      RECT  1.030000  0.085000  1.280000 0.830000 ;
      RECT  1.405000  2.560000  3.290000 2.570000 ;
      RECT  1.405000  2.570000  1.925000 2.575000 ;
      RECT  1.405000  2.575000  1.910000 2.580000 ;
      RECT  1.405000  2.580000  1.890000 2.585000 ;
      RECT  1.435000  2.585000  1.890000 2.590000 ;
      RECT  1.435000  2.590000  1.860000 2.610000 ;
      RECT  1.455000  0.350000  1.840000 0.970000 ;
      RECT  1.455000  0.970000  2.505000 0.975000 ;
      RECT  1.455000  0.975000  2.695000 1.140000 ;
      RECT  1.455000  1.140000  1.625000 1.945000 ;
      RECT  1.455000  1.945000  1.865000 2.140000 ;
      RECT  1.615000  2.140000  1.865000 2.205000 ;
      RECT  1.615000  2.205000  1.785000 2.240000 ;
      RECT  1.835000  2.405000  3.290000 2.410000 ;
      RECT  1.850000  2.400000  3.290000 2.405000 ;
      RECT  1.870000  2.390000  3.290000 2.400000 ;
      RECT  1.895000  2.375000  3.290000 2.390000 ;
      RECT  1.985000  2.740000  2.315000 3.245000 ;
      RECT  2.060000  0.085000  2.390000 0.800000 ;
      RECT  2.445000  1.140000  2.695000 1.490000 ;
      RECT  2.445000  1.490000  2.775000 1.695000 ;
      RECT  2.445000  1.865000  3.420000 1.985000 ;
      RECT  2.445000  1.985000  3.060000 2.035000 ;
      RECT  2.445000  2.035000  2.775000 2.205000 ;
      RECT  2.560000  0.330000  4.440000 0.500000 ;
      RECT  2.560000  0.500000  3.035000 0.805000 ;
      RECT  2.865000  0.805000  3.035000 1.195000 ;
      RECT  2.865000  1.195000  3.115000 1.345000 ;
      RECT  2.900000  1.820000  3.420000 1.865000 ;
      RECT  2.945000  1.345000  3.115000 1.560000 ;
      RECT  2.945000  1.560000  3.420000 1.820000 ;
      RECT  3.010000  2.205000  3.760000 2.325000 ;
      RECT  3.010000  2.325000  3.335000 2.370000 ;
      RECT  3.010000  2.370000  3.290000 2.375000 ;
      RECT  3.010000  2.570000  3.290000 2.725000 ;
      RECT  3.185000  2.155000  3.760000 2.205000 ;
      RECT  3.205000  0.670000  3.455000 1.045000 ;
      RECT  3.285000  1.045000  3.455000 1.220000 ;
      RECT  3.285000  1.220000  3.760000 1.390000 ;
      RECT  3.460000  2.495000  5.250000 2.570000 ;
      RECT  3.460000  2.570000  4.215000 2.725000 ;
      RECT  3.590000  1.390000  3.760000 2.155000 ;
      RECT  3.625000  0.670000  4.100000 1.050000 ;
      RECT  3.930000  1.050000  4.100000 2.400000 ;
      RECT  3.930000  2.400000  5.250000 2.495000 ;
      RECT  4.270000  0.500000  4.440000 0.565000 ;
      RECT  4.270000  0.565000  5.650000 0.735000 ;
      RECT  4.270000  0.905000  6.150000 1.075000 ;
      RECT  4.270000  1.075000  4.445000 2.125000 ;
      RECT  4.385000  2.740000  4.715000 3.245000 ;
      RECT  4.615000  1.245000  5.650000 1.575000 ;
      RECT  4.615000  1.575000  4.785000 2.320000 ;
      RECT  4.615000  2.320000  5.250000 2.400000 ;
      RECT  4.915000  0.085000  5.310000 0.395000 ;
      RECT  4.955000  1.795000  5.285000 2.150000 ;
      RECT  5.480000  0.255000  7.420000 0.425000 ;
      RECT  5.480000  0.425000  5.650000 0.565000 ;
      RECT  5.480000  1.745000  5.810000 3.245000 ;
      RECT  5.820000  0.665000  6.150000 0.905000 ;
      RECT  5.820000  1.075000  6.150000 1.130000 ;
      RECT  5.980000  1.130000  6.150000 1.865000 ;
      RECT  5.980000  1.865000  6.310000 2.755000 ;
      RECT  6.320000  0.595000  7.080000 0.845000 ;
      RECT  6.320000  0.845000  6.490000 1.515000 ;
      RECT  6.320000  1.515000  6.650000 1.685000 ;
      RECT  6.480000  1.685000  6.650000 2.475000 ;
      RECT  6.480000  2.475000  7.635000 2.805000 ;
      RECT  6.690000  1.015000  7.420000 1.345000 ;
      RECT  6.965000  1.345000  7.295000 2.305000 ;
      RECT  7.250000  0.425000  7.420000 1.015000 ;
      RECT  7.465000  1.515000  8.850000 1.685000 ;
      RECT  7.465000  1.685000  7.635000 2.475000 ;
      RECT  7.590000  1.015000  9.190000 1.185000 ;
      RECT  7.590000  1.185000  7.920000 1.345000 ;
      RECT  7.745000  0.085000  8.075000 0.845000 ;
      RECT  7.805000  1.920000  8.345000 2.255000 ;
      RECT  7.805000  2.445000  8.135000 3.245000 ;
      RECT  8.320000  2.445000  8.685000 2.905000 ;
      RECT  8.515000  1.855000  9.190000 2.025000 ;
      RECT  8.515000  2.025000  8.685000 2.445000 ;
      RECT  8.520000  1.355000  8.850000 1.515000 ;
      RECT  8.615000  0.385000  8.945000 1.015000 ;
      RECT  8.855000  2.195000  9.185000 3.245000 ;
      RECT  9.020000  1.185000  9.190000 1.855000 ;
      RECT  9.175000  0.085000  9.425000 0.845000 ;
      RECT  9.385000  1.385000  9.935000 1.715000 ;
      RECT  9.385000  1.715000  9.555000 2.905000 ;
      RECT  9.605000  0.350000  9.935000 1.385000 ;
      RECT 10.595000  1.820000 10.925000 3.245000 ;
      RECT 10.675000  0.085000 10.925000 1.130000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  1.950000  1.285000 2.120000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  1.950000  5.125000 2.120000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  1.950000  8.005000 2.120000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
  END
END sky130_fd_sc_hs__dfrtp_1
MACRO sky130_fd_sc_hs__dfrtp_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.52000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.000000 0.495000 2.170000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.650000 0.350000 10.980000 2.980000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.055000 1.920000 1.345000 1.965000 ;
        RECT 1.055000 1.965000 8.065000 2.105000 ;
        RECT 1.055000 2.105000 1.345000 2.150000 ;
        RECT 4.895000 1.920000 5.185000 1.965000 ;
        RECT 4.895000 2.105000 5.185000 2.150000 ;
        RECT 7.775000 1.920000 8.065000 1.965000 ;
        RECT 7.775000 2.105000 8.065000 2.150000 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.795000 1.320000 2.275000 1.730000 ;
        RECT 2.045000 1.730000 2.275000 1.780000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.520000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 11.520000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.520000 0.085000 ;
      RECT  0.000000  3.245000 11.520000 3.415000 ;
      RECT  0.105000  2.520000  0.435000 3.245000 ;
      RECT  0.130000  0.370000  0.460000 0.660000 ;
      RECT  0.130000  0.660000  0.835000 0.830000 ;
      RECT  0.635000  2.520000  3.325000 2.560000 ;
      RECT  0.635000  2.560000  0.890000 2.605000 ;
      RECT  0.635000  2.605000  0.870000 2.630000 ;
      RECT  0.635000  2.630000  0.835000 2.980000 ;
      RECT  0.665000  0.830000  0.835000 2.330000 ;
      RECT  0.665000  2.330000  2.340000 2.355000 ;
      RECT  0.665000  2.355000  2.360000 2.380000 ;
      RECT  0.665000  2.380000  2.385000 2.395000 ;
      RECT  0.665000  2.395000  2.405000 2.405000 ;
      RECT  0.665000  2.405000  2.420000 2.420000 ;
      RECT  0.665000  2.420000  2.440000 2.430000 ;
      RECT  0.665000  2.430000  2.460000 2.435000 ;
      RECT  0.665000  2.435000  2.470000 2.440000 ;
      RECT  0.665000  2.440000  2.485000 2.445000 ;
      RECT  0.665000  2.445000  3.325000 2.520000 ;
      RECT  1.005000  0.085000  1.285000 0.830000 ;
      RECT  1.005000  1.140000  1.285000 2.150000 ;
      RECT  1.015000  2.730000  1.345000 3.245000 ;
      RECT  1.405000  2.560000  3.325000 2.570000 ;
      RECT  1.455000  0.350000  1.875000 0.970000 ;
      RECT  1.455000  0.970000  2.540000 0.975000 ;
      RECT  1.455000  0.975000  2.685000 1.150000 ;
      RECT  1.455000  1.150000  1.625000 1.900000 ;
      RECT  1.455000  1.900000  1.865000 2.160000 ;
      RECT  1.955000  2.740000  2.285000 3.245000 ;
      RECT  2.095000  0.085000  2.425000 0.800000 ;
      RECT  2.330000  2.570000  3.325000 2.575000 ;
      RECT  2.345000  2.575000  3.325000 2.580000 ;
      RECT  2.355000  2.580000  3.325000 2.585000 ;
      RECT  2.365000  2.585000  3.325000 2.590000 ;
      RECT  2.375000  2.590000  3.325000 2.595000 ;
      RECT  2.390000  2.595000  3.325000 2.605000 ;
      RECT  2.405000  2.605000  3.325000 2.615000 ;
      RECT  2.445000  1.150000  2.685000 1.550000 ;
      RECT  2.515000  1.550000  2.685000 1.775000 ;
      RECT  2.515000  1.945000  3.425000 1.985000 ;
      RECT  2.515000  1.985000  3.095000 2.035000 ;
      RECT  2.515000  2.035000  3.010000 2.080000 ;
      RECT  2.515000  2.080000  2.940000 2.205000 ;
      RECT  2.515000  2.205000  2.775000 2.230000 ;
      RECT  2.530000  2.230000  2.775000 2.275000 ;
      RECT  2.595000  0.330000  4.475000 0.500000 ;
      RECT  2.595000  0.500000  3.070000 0.805000 ;
      RECT  2.810000  1.900000  3.425000 1.945000 ;
      RECT  2.865000  0.805000  3.070000 1.625000 ;
      RECT  2.865000  1.625000  3.425000 1.900000 ;
      RECT  2.945000  2.375000  3.370000 2.400000 ;
      RECT  2.945000  2.400000  3.325000 2.445000 ;
      RECT  3.045000  2.615000  3.325000 2.725000 ;
      RECT  3.110000  2.230000  3.765000 2.355000 ;
      RECT  3.110000  2.355000  3.370000 2.375000 ;
      RECT  3.200000  2.185000  3.765000 2.230000 ;
      RECT  3.240000  0.670000  3.490000 1.045000 ;
      RECT  3.320000  1.045000  3.490000 1.220000 ;
      RECT  3.320000  1.220000  3.765000 1.390000 ;
      RECT  3.495000  2.525000  5.285000 2.570000 ;
      RECT  3.495000  2.570000  4.250000 2.750000 ;
      RECT  3.595000  1.390000  3.765000 2.185000 ;
      RECT  3.660000  0.670000  4.105000 1.050000 ;
      RECT  3.935000  1.050000  4.105000 2.400000 ;
      RECT  3.935000  2.400000  5.285000 2.525000 ;
      RECT  4.275000  0.955000  6.185000 1.125000 ;
      RECT  4.275000  1.125000  4.445000 2.125000 ;
      RECT  4.305000  0.500000  4.475000 0.615000 ;
      RECT  4.305000  0.615000  5.685000 0.785000 ;
      RECT  4.420000  2.740000  4.750000 3.245000 ;
      RECT  4.615000  1.295000  5.685000 1.575000 ;
      RECT  4.615000  1.575000  4.785000 2.320000 ;
      RECT  4.615000  2.320000  5.285000 2.400000 ;
      RECT  4.920000  0.085000  5.345000 0.445000 ;
      RECT  4.955000  1.795000  5.285000 2.150000 ;
      RECT  5.515000  0.255000  7.455000 0.425000 ;
      RECT  5.515000  0.425000  5.685000 0.615000 ;
      RECT  5.515000  1.745000  5.845000 3.245000 ;
      RECT  5.855000  0.595000  6.185000 0.955000 ;
      RECT  5.855000  1.125000  6.185000 1.130000 ;
      RECT  6.015000  1.130000  6.185000 1.855000 ;
      RECT  6.015000  1.855000  6.345000 2.755000 ;
      RECT  6.355000  0.595000  7.115000 0.845000 ;
      RECT  6.355000  0.845000  6.525000 1.515000 ;
      RECT  6.355000  1.515000  6.685000 1.685000 ;
      RECT  6.515000  1.685000  6.685000 2.475000 ;
      RECT  6.515000  2.475000  7.625000 2.805000 ;
      RECT  6.725000  1.015000  7.455000 1.345000 ;
      RECT  6.955000  1.345000  7.285000 2.305000 ;
      RECT  7.285000  0.425000  7.455000 1.015000 ;
      RECT  7.455000  1.560000  9.035000 1.730000 ;
      RECT  7.455000  1.730000  7.625000 2.475000 ;
      RECT  7.625000  1.060000  7.955000 1.220000 ;
      RECT  7.625000  1.220000  9.375000 1.390000 ;
      RECT  7.770000  0.085000  8.190000 0.715000 ;
      RECT  7.795000  2.445000  8.125000 3.245000 ;
      RECT  7.805000  1.920000  8.395000 2.275000 ;
      RECT  8.295000  2.445000  8.885000 2.775000 ;
      RECT  8.680000  0.385000  9.010000 1.220000 ;
      RECT  8.705000  1.730000  9.035000 1.890000 ;
      RECT  8.715000  2.105000  9.375000 2.275000 ;
      RECT  8.715000  2.275000  8.885000 2.445000 ;
      RECT  9.090000  2.445000  9.420000 3.245000 ;
      RECT  9.205000  1.390000  9.375000 2.105000 ;
      RECT  9.230000  0.085000  9.480000 1.050000 ;
      RECT  9.590000  2.030000  9.920000 2.905000 ;
      RECT  9.660000  0.350000  9.990000 1.300000 ;
      RECT  9.660000  1.300000 10.190000 1.630000 ;
      RECT  9.660000  1.630000  9.920000 2.030000 ;
      RECT 10.150000  1.820000 10.480000 3.245000 ;
      RECT 10.220000  0.085000 10.470000 1.130000 ;
      RECT 11.155000  1.820000 11.405000 3.245000 ;
      RECT 11.160000  0.085000 11.410000 1.130000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  1.950000  1.285000 2.120000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  1.950000  5.125000 2.120000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  1.950000  8.005000 2.120000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
  END
END sky130_fd_sc_hs__dfrtp_2
MACRO sky130_fd_sc_hs__dfrtp_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.44000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.000000 0.515000 2.180000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.207100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.035000 1.800000 12.740000 1.970000 ;
        RECT 11.035000 1.970000 11.365000 2.980000 ;
        RECT 11.595000 0.365000 11.910000 0.880000 ;
        RECT 11.595000 0.880000 12.825000 1.130000 ;
        RECT 12.410000 1.610000 13.315000 1.780000 ;
        RECT 12.410000 1.780000 12.740000 1.800000 ;
        RECT 12.410000 1.970000 12.740000 2.980000 ;
        RECT 12.575000 0.350000 12.825000 0.880000 ;
        RECT 12.575000 1.130000 12.825000 1.270000 ;
        RECT 12.575000 1.270000 13.315000 1.610000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.055000 1.920000 1.345000 1.965000 ;
        RECT 1.055000 1.965000 9.025000 2.105000 ;
        RECT 1.055000 2.105000 1.345000 2.150000 ;
        RECT 5.375000 1.920000 5.665000 1.965000 ;
        RECT 5.375000 2.105000 5.665000 2.150000 ;
        RECT 8.735000 1.920000 9.025000 1.965000 ;
        RECT 8.735000 2.105000 9.025000 2.150000 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.795000 1.310000 2.275000 1.640000 ;
        RECT 1.845000 1.640000 2.275000 1.775000 ;
        RECT 2.045000 1.775000 2.275000 1.780000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 13.440000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 13.440000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.440000 0.085000 ;
      RECT  0.000000  3.245000 13.440000 3.415000 ;
      RECT  0.110000  2.520000  0.360000 3.245000 ;
      RECT  0.165000  0.370000  0.495000 0.660000 ;
      RECT  0.165000  0.660000  0.855000 0.830000 ;
      RECT  0.560000  2.520000  3.310000 2.580000 ;
      RECT  0.560000  2.580000  0.890000 2.605000 ;
      RECT  0.560000  2.605000  0.875000 2.615000 ;
      RECT  0.560000  2.615000  0.860000 2.640000 ;
      RECT  0.560000  2.640000  0.830000 2.980000 ;
      RECT  0.685000  0.830000  0.855000 2.410000 ;
      RECT  0.685000  2.410000  3.310000 2.520000 ;
      RECT  1.000000  2.750000  1.340000 3.245000 ;
      RECT  1.025000  1.130000  1.285000 2.140000 ;
      RECT  1.065000  0.085000  1.235000 0.830000 ;
      RECT  1.455000  0.350000  1.875000 0.970000 ;
      RECT  1.455000  0.970000  2.510000 0.975000 ;
      RECT  1.455000  0.975000  2.635000 1.140000 ;
      RECT  1.455000  1.140000  1.625000 1.945000 ;
      RECT  1.455000  1.945000  1.805000 2.240000 ;
      RECT  2.005000  2.750000  2.335000 3.245000 ;
      RECT  2.055000  0.085000  2.385000 0.800000 ;
      RECT  2.445000  1.140000  2.635000 1.550000 ;
      RECT  2.455000  1.550000  2.635000 1.775000 ;
      RECT  2.455000  1.945000  3.455000 2.015000 ;
      RECT  2.455000  2.015000  2.985000 2.055000 ;
      RECT  2.455000  2.055000  2.940000 2.240000 ;
      RECT  2.555000  0.330000  4.475000 0.500000 ;
      RECT  2.555000  0.500000  3.015000 0.805000 ;
      RECT  2.770000  1.905000  3.455000 1.945000 ;
      RECT  2.815000  0.805000  3.015000 1.560000 ;
      RECT  2.815000  1.560000  3.455000 1.905000 ;
      RECT  3.030000  2.580000  3.310000 2.755000 ;
      RECT  3.110000  2.185000  3.795000 2.355000 ;
      RECT  3.110000  2.355000  3.310000 2.410000 ;
      RECT  3.185000  0.670000  3.435000 1.220000 ;
      RECT  3.185000  1.220000  3.795000 1.390000 ;
      RECT  3.480000  2.525000  5.180000 2.570000 ;
      RECT  3.480000  2.570000  4.230000 2.755000 ;
      RECT  3.605000  0.670000  3.935000 0.880000 ;
      RECT  3.605000  0.880000  4.135000 1.050000 ;
      RECT  3.625000  1.390000  3.795000 2.185000 ;
      RECT  3.965000  1.050000  4.135000 2.400000 ;
      RECT  3.965000  2.400000  5.180000 2.525000 ;
      RECT  4.305000  0.500000  4.475000 0.540000 ;
      RECT  4.305000  0.540000  5.565000 0.710000 ;
      RECT  4.305000  0.880000  6.990000 1.050000 ;
      RECT  4.305000  1.050000  4.570000 2.105000 ;
      RECT  4.400000  2.740000  4.730000 3.245000 ;
      RECT  4.745000  1.220000  5.985000 1.500000 ;
      RECT  4.745000  1.500000  4.915000 2.295000 ;
      RECT  4.745000  2.295000  5.180000 2.400000 ;
      RECT  4.895000  0.085000  5.225000 0.370000 ;
      RECT  4.915000  2.570000  5.180000 2.755000 ;
      RECT  5.085000  1.670000  5.635000 2.120000 ;
      RECT  5.395000  0.255000  8.275000 0.425000 ;
      RECT  5.395000  0.425000  5.565000 0.540000 ;
      RECT  5.395000  2.290000  5.725000 2.405000 ;
      RECT  5.395000  2.405000  6.955000 2.575000 ;
      RECT  5.735000  0.720000  6.990000 0.880000 ;
      RECT  5.830000  2.745000  6.165000 3.245000 ;
      RECT  6.155000  1.050000  6.325000 1.940000 ;
      RECT  6.155000  1.940000  6.615000 2.235000 ;
      RECT  6.495000  1.260000  6.955000 1.590000 ;
      RECT  6.785000  1.590000  6.955000 2.405000 ;
      RECT  7.125000  2.475000  8.410000 2.805000 ;
      RECT  7.160000  0.595000  7.935000 0.845000 ;
      RECT  7.160000  0.845000  7.330000 2.475000 ;
      RECT  7.545000  1.015000  8.275000 1.345000 ;
      RECT  7.740000  1.345000  8.070000 2.305000 ;
      RECT  8.105000  0.425000  8.275000 1.015000 ;
      RECT  8.240000  1.535000  9.605000 1.705000 ;
      RECT  8.240000  1.705000  8.410000 2.475000 ;
      RECT  8.445000  1.035000  9.945000 1.205000 ;
      RECT  8.445000  1.205000  8.775000 1.365000 ;
      RECT  8.580000  2.445000  8.910000 3.245000 ;
      RECT  8.625000  0.085000  8.955000 0.845000 ;
      RECT  8.765000  1.920000  9.140000 2.275000 ;
      RECT  9.080000  2.445000  9.480000 2.905000 ;
      RECT  9.310000  1.875000  9.945000 2.045000 ;
      RECT  9.310000  2.045000  9.480000 2.445000 ;
      RECT  9.345000  1.375000  9.605000 1.535000 ;
      RECT  9.500000  0.385000  9.830000 1.035000 ;
      RECT  9.650000  2.445000  9.900000 3.245000 ;
      RECT  9.775000  1.205000  9.945000 1.875000 ;
      RECT 10.115000  0.085000 10.390000 1.130000 ;
      RECT 10.115000  1.460000 12.240000 1.630000 ;
      RECT 10.115000  1.630000 10.365000 2.905000 ;
      RECT 10.535000  2.025000 10.865000 3.245000 ;
      RECT 10.560000  0.350000 10.890000 1.300000 ;
      RECT 10.560000  1.300000 12.240000 1.460000 ;
      RECT 11.120000  0.085000 11.410000 1.130000 ;
      RECT 11.535000  2.140000 12.240000 3.245000 ;
      RECT 12.080000  0.085000 12.405000 0.710000 ;
      RECT 12.910000  1.950000 13.240000 3.245000 ;
      RECT 13.005000  0.085000 13.335000 1.100000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  1.950000  1.285000 2.120000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  1.950000  5.605000 2.120000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  1.950000  8.965000 2.120000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
  END
END sky130_fd_sc_hs__dfrtp_4
MACRO sky130_fd_sc_hs__dfsbp_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.475000 1.010000 0.805000 2.020000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.555000 0.350000 11.885000 1.050000 ;
        RECT 11.555000 1.820000 11.885000 2.980000 ;
        RECT 11.715000 1.050000 11.885000 1.820000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  9.985000 0.350000 10.315000 1.130000 ;
        RECT 10.120000 1.130000 10.315000 1.180000 ;
        RECT 10.120000 1.180000 10.435000 2.980000 ;
    END
  END Q_N
  PIN SET_B
    ANTENNAPARTIALMETALSIDEAREA  2.205000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 5.375000 1.550000 5.665000 1.595000 ;
        RECT 5.375000 1.595000 8.545000 1.735000 ;
        RECT 5.375000 1.735000 5.665000 1.780000 ;
        RECT 8.255000 1.550000 8.545000 1.595000 ;
        RECT 8.255000 1.735000 8.545000 1.780000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.315000 1.180000 1.795000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.000000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 12.000000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.000000 0.085000 ;
      RECT  0.000000  3.245000 12.000000 3.415000 ;
      RECT  0.115000  0.380000  0.365000 0.840000 ;
      RECT  0.115000  0.840000  0.285000 2.190000 ;
      RECT  0.115000  2.190000  2.695000 2.230000 ;
      RECT  0.115000  2.230000  1.795000 2.360000 ;
      RECT  0.115000  2.360000  0.365000 2.980000 ;
      RECT  0.545000  0.085000  0.795000 0.840000 ;
      RECT  0.565000  2.590000  0.895000 3.245000 ;
      RECT  0.975000  0.350000  1.435000 1.010000 ;
      RECT  0.975000  1.010000  1.145000 1.720000 ;
      RECT  0.975000  1.720000  2.355000 1.890000 ;
      RECT  0.975000  1.890000  1.455000 2.020000 ;
      RECT  1.575000  2.530000  1.905000 3.245000 ;
      RECT  1.605000  0.085000  1.865000 1.010000 ;
      RECT  1.625000  2.060000  2.695000 2.190000 ;
      RECT  2.025000  1.300000  2.355000 1.720000 ;
      RECT  2.045000  0.255000  3.195000 0.425000 ;
      RECT  2.045000  0.425000  2.295000 1.130000 ;
      RECT  2.105000  2.400000  2.355000 2.905000 ;
      RECT  2.105000  2.905000  3.875000 3.075000 ;
      RECT  2.525000  0.595000  2.855000 0.845000 ;
      RECT  2.525000  0.845000  2.695000 2.060000 ;
      RECT  2.525000  2.230000  2.695000 2.295000 ;
      RECT  2.525000  2.295000  3.005000 2.735000 ;
      RECT  2.865000  1.435000  3.195000 2.105000 ;
      RECT  3.025000  0.425000  3.195000 1.435000 ;
      RECT  3.175000  2.295000  3.535000 2.735000 ;
      RECT  3.365000  0.385000  3.615000 0.885000 ;
      RECT  3.365000  0.885000  4.285000 1.055000 ;
      RECT  3.365000  1.055000  3.535000 2.295000 ;
      RECT  3.705000  1.360000  3.945000 2.165000 ;
      RECT  3.705000  2.165000  4.780000 2.335000 ;
      RECT  3.705000  2.335000  3.875000 2.905000 ;
      RECT  4.045000  2.505000  4.440000 3.245000 ;
      RECT  4.105000  0.085000  4.435000 0.715000 ;
      RECT  4.115000  1.055000  4.285000 1.435000 ;
      RECT  4.115000  1.435000  5.235000 1.605000 ;
      RECT  4.230000  1.775000  5.200000 1.995000 ;
      RECT  4.455000  0.885000  4.775000 1.265000 ;
      RECT  4.605000  0.435000  5.180000 0.885000 ;
      RECT  4.610000  2.335000  4.780000 2.905000 ;
      RECT  4.610000  2.905000  5.540000 3.075000 ;
      RECT  4.950000  1.055000  5.235000 1.120000 ;
      RECT  4.950000  1.120000  6.265000 1.290000 ;
      RECT  4.950000  1.290000  5.235000 1.435000 ;
      RECT  4.950000  1.995000  5.200000 2.735000 ;
      RECT  5.370000  2.125000  6.035000 2.295000 ;
      RECT  5.370000  2.295000  5.540000 2.905000 ;
      RECT  5.405000  1.550000  5.695000 1.955000 ;
      RECT  5.710000  2.465000  6.050000 3.245000 ;
      RECT  5.855000  0.085000  6.185000 0.950000 ;
      RECT  5.865000  1.620000  6.605000 1.790000 ;
      RECT  5.865000  1.790000  6.035000 2.125000 ;
      RECT  5.935000  1.290000  6.265000 1.450000 ;
      RECT  6.435000  0.255000  7.560000 0.425000 ;
      RECT  6.435000  0.425000  6.605000 1.120000 ;
      RECT  6.435000  1.120000  6.880000 1.450000 ;
      RECT  6.435000  1.450000  6.605000 1.620000 ;
      RECT  6.760000  1.960000  7.010000 2.480000 ;
      RECT  6.760000  2.480000  7.900000 2.650000 ;
      RECT  6.760000  2.650000  7.450000 2.905000 ;
      RECT  6.775000  0.595000  7.220000 0.925000 ;
      RECT  6.840000  1.680000  7.220000 1.850000 ;
      RECT  6.840000  1.850000  7.010000 1.960000 ;
      RECT  7.050000  0.925000  7.220000 1.680000 ;
      RECT  7.230000  2.020000  7.560000 2.310000 ;
      RECT  7.390000  0.425000  7.560000 2.020000 ;
      RECT  7.730000  2.050000  9.395000 2.220000 ;
      RECT  7.730000  2.220000  8.770000 2.480000 ;
      RECT  7.770000  0.840000  9.735000 1.010000 ;
      RECT  7.770000  1.010000  8.100000 1.880000 ;
      RECT  8.065000  0.085000  8.755000 0.670000 ;
      RECT  8.070000  2.650000  8.240000 3.245000 ;
      RECT  8.285000  1.180000  8.670000 1.780000 ;
      RECT  8.440000  2.480000  8.770000 2.980000 ;
      RECT  8.925000  0.415000  9.255000 0.840000 ;
      RECT  9.000000  2.390000  9.735000 2.560000 ;
      RECT  9.000000  2.560000  9.330000 2.980000 ;
      RECT  9.065000  1.210000  9.395000 2.050000 ;
      RECT  9.485000  0.085000  9.815000 0.670000 ;
      RECT  9.560000  2.730000  9.910000 3.245000 ;
      RECT  9.565000  1.010000  9.735000 2.390000 ;
      RECT 10.545000  0.350000 10.875000 0.940000 ;
      RECT 10.680000  0.940000 10.875000 1.220000 ;
      RECT 10.680000  1.220000 11.540000 1.550000 ;
      RECT 10.680000  1.550000 10.850000 2.875000 ;
      RECT 11.050000  1.995000 11.380000 3.245000 ;
      RECT 11.055000  0.085000 11.385000 0.940000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  1.580000  5.605000 1.750000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  1.580000  8.485000 1.750000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
  END
END sky130_fd_sc_hs__dfsbp_1
MACRO sky130_fd_sc_hs__dfsbp_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.96000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.475000 0.980000 0.805000 1.990000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.065000 1.820000 12.425000 2.980000 ;
        RECT 12.085000 0.350000 12.425000 1.130000 ;
        RECT 12.255000 1.130000 12.425000 1.820000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.130000 1.820000 10.435000 2.970000 ;
        RECT 10.175000 0.350000 10.435000 1.820000 ;
    END
  END Q_N
  PIN SET_B
    ANTENNAPARTIALMETALSIDEAREA  2.205000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 5.375000 1.550000 5.665000 1.595000 ;
        RECT 5.375000 1.595000 8.545000 1.735000 ;
        RECT 5.375000 1.735000 5.665000 1.780000 ;
        RECT 8.255000 1.550000 8.545000 1.595000 ;
        RECT 8.255000 1.735000 8.545000 1.780000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.315000 1.180000 1.775000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.960000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 12.960000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.960000 0.085000 ;
      RECT  0.000000  3.245000 12.960000 3.415000 ;
      RECT  0.115000  0.350000  0.365000 0.810000 ;
      RECT  0.115000  0.810000  0.285000 2.190000 ;
      RECT  0.115000  2.190000  2.615000 2.230000 ;
      RECT  0.115000  2.230000  1.795000 2.360000 ;
      RECT  0.115000  2.360000  0.365000 2.980000 ;
      RECT  0.545000  0.085000  0.795000 0.810000 ;
      RECT  0.565000  2.530000  0.895000 3.245000 ;
      RECT  0.975000  0.350000  1.435000 1.010000 ;
      RECT  0.975000  1.010000  1.145000 1.720000 ;
      RECT  0.975000  1.720000  2.275000 1.890000 ;
      RECT  0.975000  1.890000  1.455000 2.020000 ;
      RECT  1.575000  2.530000  1.905000 3.245000 ;
      RECT  1.605000  0.085000  1.865000 1.010000 ;
      RECT  1.625000  2.060000  2.615000 2.190000 ;
      RECT  1.945000  1.300000  2.275000 1.720000 ;
      RECT  2.045000  0.255000  3.110000 0.425000 ;
      RECT  2.045000  0.425000  2.215000 1.130000 ;
      RECT  2.105000  2.400000  2.275000 2.905000 ;
      RECT  2.105000  2.905000  3.845000 3.075000 ;
      RECT  2.445000  0.595000  2.770000 0.925000 ;
      RECT  2.445000  0.925000  2.615000 2.060000 ;
      RECT  2.445000  2.230000  2.615000 2.295000 ;
      RECT  2.445000  2.295000  2.865000 2.735000 ;
      RECT  2.785000  1.435000  3.115000 2.105000 ;
      RECT  2.940000  0.425000  3.110000 1.435000 ;
      RECT  3.065000  2.295000  3.455000 2.735000 ;
      RECT  3.280000  0.465000  3.530000 0.925000 ;
      RECT  3.285000  0.925000  3.530000 1.095000 ;
      RECT  3.285000  1.095000  4.185000 1.265000 ;
      RECT  3.285000  1.265000  3.455000 2.295000 ;
      RECT  3.625000  1.435000  3.845000 2.395000 ;
      RECT  3.625000  2.395000  4.690000 2.565000 ;
      RECT  3.625000  2.565000  3.845000 2.905000 ;
      RECT  3.990000  0.085000  4.240000 0.845000 ;
      RECT  4.015000  1.265000  4.185000 1.515000 ;
      RECT  4.015000  1.515000  5.015000 1.685000 ;
      RECT  4.020000  2.735000  4.350000 3.245000 ;
      RECT  4.140000  1.855000  4.470000 2.055000 ;
      RECT  4.140000  2.055000  5.030000 2.225000 ;
      RECT  4.355000  1.015000  4.580000 1.345000 ;
      RECT  4.410000  0.350000  4.880000 1.015000 ;
      RECT  4.520000  2.565000  4.690000 2.905000 ;
      RECT  4.520000  2.905000  5.530000 3.075000 ;
      RECT  4.750000  1.240000  5.915000 1.410000 ;
      RECT  4.750000  1.410000  5.015000 1.515000 ;
      RECT  4.750000  1.685000  5.015000 1.885000 ;
      RECT  4.860000  2.225000  5.030000 2.295000 ;
      RECT  4.860000  2.295000  5.190000 2.735000 ;
      RECT  5.225000  1.580000  5.635000 2.020000 ;
      RECT  5.340000  0.085000  6.160000 0.680000 ;
      RECT  5.360000  2.190000  6.500000 2.360000 ;
      RECT  5.360000  2.360000  5.530000 2.905000 ;
      RECT  5.585000  1.120000  5.915000 1.240000 ;
      RECT  5.700000  2.530000  6.070000 3.245000 ;
      RECT  6.330000  0.280000  7.555000 0.450000 ;
      RECT  6.330000  0.450000  6.500000 1.120000 ;
      RECT  6.330000  1.120000  6.875000 1.450000 ;
      RECT  6.330000  1.450000  6.500000 2.190000 ;
      RECT  6.670000  0.620000  7.215000 0.950000 ;
      RECT  6.780000  1.680000  7.215000 1.850000 ;
      RECT  6.780000  1.850000  7.030000 2.480000 ;
      RECT  6.780000  2.480000  7.920000 2.650000 ;
      RECT  6.780000  2.650000  7.470000 2.980000 ;
      RECT  7.045000  0.950000  7.215000 1.680000 ;
      RECT  7.250000  2.020000  7.580000 2.310000 ;
      RECT  7.385000  0.450000  7.555000 2.020000 ;
      RECT  7.725000  0.840000  9.435000 1.010000 ;
      RECT  7.725000  1.010000  8.055000 1.780000 ;
      RECT  7.750000  1.950000  9.570000 2.120000 ;
      RECT  7.750000  2.120000  8.790000 2.480000 ;
      RECT  8.090000  2.650000  8.260000 3.245000 ;
      RECT  8.100000  0.085000  8.845000 0.670000 ;
      RECT  8.285000  1.180000  8.640000 1.780000 ;
      RECT  8.460000  2.480000  8.790000 2.915000 ;
      RECT  8.900000  1.350000  9.570000 1.950000 ;
      RECT  9.015000  2.290000  9.910000 2.460000 ;
      RECT  9.015000  2.460000  9.345000 2.620000 ;
      RECT  9.105000  0.635000  9.435000 0.840000 ;
      RECT  9.105000  1.010000  9.910000 1.180000 ;
      RECT  9.630000  2.630000  9.960000 3.245000 ;
      RECT  9.665000  0.085000  9.995000 0.840000 ;
      RECT  9.740000  1.180000  9.910000 2.290000 ;
      RECT 10.605000  0.085000 10.855000 1.130000 ;
      RECT 10.605000  1.820000 10.860000 3.245000 ;
      RECT 11.085000  0.350000 11.415000 1.300000 ;
      RECT 11.085000  1.300000 12.085000 1.630000 ;
      RECT 11.085000  1.630000 11.415000 2.860000 ;
      RECT 11.585000  0.085000 11.915000 1.030000 ;
      RECT 11.615000  1.820000 11.865000 3.245000 ;
      RECT 12.595000  0.085000 12.845000 1.130000 ;
      RECT 12.595000  1.820000 12.845000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  1.580000  5.605000 1.750000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  1.580000  8.485000 1.750000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
  END
END sky130_fd_sc_hs__dfsbp_2
MACRO sky130_fd_sc_hs__dfstp_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.475000 0.980000 0.805000 1.990000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.530100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.500000 0.350000 10.935000 1.050000 ;
        RECT 10.685000 1.050000 10.935000 2.980000 ;
    END
  END Q
  PIN SET_B
    ANTENNAPARTIALMETALSIDEAREA  2.205000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 5.375000 1.920000 5.665000 1.965000 ;
        RECT 5.375000 1.965000 8.545000 2.105000 ;
        RECT 5.375000 2.105000 5.665000 2.150000 ;
        RECT 8.255000 1.920000 8.545000 1.965000 ;
        RECT 8.255000 2.105000 8.545000 2.150000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.315000 1.180000 1.795000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.040000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 11.040000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  3.245000 11.040000 3.415000 ;
      RECT  0.105000  0.350000  0.365000 0.810000 ;
      RECT  0.105000  0.810000  0.275000 2.230000 ;
      RECT  0.105000  2.230000  1.760000 2.400000 ;
      RECT  0.105000  2.400000  0.355000 2.980000 ;
      RECT  0.545000  0.085000  0.795000 0.810000 ;
      RECT  0.555000  2.570000  0.885000 3.245000 ;
      RECT  0.975000  0.350000  1.435000 1.010000 ;
      RECT  0.975000  1.010000  1.145000 1.720000 ;
      RECT  0.975000  1.720000  2.315000 1.890000 ;
      RECT  0.975000  1.890000  1.420000 2.060000 ;
      RECT  1.540000  2.570000  1.870000 3.245000 ;
      RECT  1.590000  2.060000  2.660000 2.230000 ;
      RECT  1.615000  0.085000  1.785000 1.010000 ;
      RECT  1.965000  0.255000  3.075000 0.425000 ;
      RECT  1.965000  0.425000  2.295000 1.090000 ;
      RECT  1.985000  1.260000  2.315000 1.720000 ;
      RECT  2.070000  2.400000  2.320000 2.905000 ;
      RECT  2.070000  2.905000  3.755000 3.075000 ;
      RECT  2.485000  0.595000  2.735000 0.925000 ;
      RECT  2.485000  0.925000  2.660000 2.060000 ;
      RECT  2.490000  2.230000  2.660000 2.295000 ;
      RECT  2.490000  2.295000  2.910000 2.735000 ;
      RECT  2.830000  1.435000  3.075000 2.105000 ;
      RECT  2.905000  0.425000  3.075000 1.435000 ;
      RECT  3.080000  2.295000  3.415000 2.735000 ;
      RECT  3.245000  0.415000  3.575000 0.850000 ;
      RECT  3.245000  0.850000  4.095000 1.020000 ;
      RECT  3.245000  1.020000  3.415000 2.295000 ;
      RECT  3.585000  1.435000  3.755000 2.085000 ;
      RECT  3.585000  2.085000  4.570000 2.255000 ;
      RECT  3.585000  2.255000  3.755000 2.905000 ;
      RECT  3.925000  1.020000  4.095000 1.345000 ;
      RECT  3.925000  1.345000  6.065000 1.515000 ;
      RECT  3.950000  2.425000  4.230000 3.245000 ;
      RECT  4.055000  1.685000  4.385000 1.745000 ;
      RECT  4.055000  1.745000  4.910000 1.915000 ;
      RECT  4.065000  0.085000  4.455000 0.680000 ;
      RECT  4.265000  0.860000  5.010000 1.030000 ;
      RECT  4.265000  1.030000  4.625000 1.175000 ;
      RECT  4.400000  2.255000  4.570000 2.905000 ;
      RECT  4.400000  2.905000  5.365000 3.075000 ;
      RECT  4.625000  0.570000  5.010000 0.860000 ;
      RECT  4.740000  1.915000  4.910000 2.320000 ;
      RECT  4.740000  2.320000  5.025000 2.735000 ;
      RECT  4.805000  1.215000  6.065000 1.345000 ;
      RECT  4.805000  1.515000  6.065000 1.545000 ;
      RECT  5.080000  1.820000  5.635000 2.150000 ;
      RECT  5.195000  2.320000  5.975000 2.490000 ;
      RECT  5.195000  2.490000  5.365000 2.905000 ;
      RECT  5.535000  2.660000  5.785000 3.245000 ;
      RECT  5.620000  0.085000  5.950000 1.030000 ;
      RECT  5.805000  1.715000  6.405000 1.885000 ;
      RECT  5.805000  1.885000  5.975000 2.320000 ;
      RECT  6.235000  0.255000  7.325000 0.425000 ;
      RECT  6.235000  0.425000  6.405000 1.120000 ;
      RECT  6.235000  1.120000  6.645000 1.450000 ;
      RECT  6.235000  1.450000  6.405000 1.715000 ;
      RECT  6.475000  2.050000  6.810000 2.625000 ;
      RECT  6.475000  2.625000  7.600000 2.980000 ;
      RECT  6.575000  0.595000  6.985000 0.925000 ;
      RECT  6.575000  1.630000  6.985000 1.800000 ;
      RECT  6.575000  1.800000  6.810000 2.050000 ;
      RECT  6.815000  0.925000  6.985000 1.630000 ;
      RECT  6.980000  1.970000  7.325000 2.140000 ;
      RECT  6.980000  2.140000  7.260000 2.355000 ;
      RECT  7.155000  0.425000  7.325000 1.970000 ;
      RECT  7.430000  2.310000  9.105000 2.480000 ;
      RECT  7.430000  2.480000  7.600000 2.625000 ;
      RECT  7.495000  0.790000  9.260000 0.960000 ;
      RECT  7.495000  0.960000  7.730000 1.555000 ;
      RECT  7.770000  2.650000  7.940000 3.245000 ;
      RECT  7.870000  0.085000  8.760000 0.600000 ;
      RECT  8.140000  2.480000  8.470000 2.930000 ;
      RECT  8.185000  1.130000  8.515000 2.140000 ;
      RECT  8.665000  2.650000  8.915000 3.245000 ;
      RECT  8.775000  1.370000  9.105000 2.310000 ;
      RECT  8.930000  0.350000  9.260000 0.790000 ;
      RECT  9.090000  0.960000  9.260000 1.030000 ;
      RECT  9.090000  1.030000  9.445000 1.200000 ;
      RECT  9.115000  2.650000  9.445000 2.980000 ;
      RECT  9.275000  1.200000  9.445000 2.650000 ;
      RECT  9.490000  0.350000  9.820000 0.860000 ;
      RECT  9.635000  0.860000  9.820000 1.220000 ;
      RECT  9.635000  1.220000 10.515000 1.550000 ;
      RECT  9.635000  1.550000  9.965000 2.875000 ;
      RECT 10.000000  0.085000 10.330000 1.030000 ;
      RECT 10.155000  1.820000 10.485000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  1.950000  5.605000 2.120000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  1.950000  8.485000 2.120000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
  END
END sky130_fd_sc_hs__dfstp_1
MACRO sky130_fd_sc_hs__dfstp_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.475000 0.980000 0.805000 1.990000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.685000 1.820000 11.465000 2.150000 ;
        RECT 11.100000 0.350000 11.465000 1.130000 ;
        RECT 11.155000 2.150000 11.465000 2.980000 ;
        RECT 11.295000 1.130000 11.465000 1.820000 ;
    END
  END Q
  PIN SET_B
    ANTENNAPARTIALMETALSIDEAREA  1.869000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 5.855000 1.920000 6.145000 1.965000 ;
        RECT 5.855000 1.965000 8.545000 2.105000 ;
        RECT 5.855000 2.105000 6.145000 2.150000 ;
        RECT 8.255000 1.920000 8.545000 1.965000 ;
        RECT 8.255000 2.105000 8.545000 2.150000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.315000 1.180000 1.775000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.000000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 12.000000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.000000 0.085000 ;
      RECT  0.000000  3.245000 12.000000 3.415000 ;
      RECT  0.115000  0.395000  0.365000 0.765000 ;
      RECT  0.115000  0.765000  0.285000 2.190000 ;
      RECT  0.115000  2.190000  2.615000 2.230000 ;
      RECT  0.115000  2.230000  1.795000 2.360000 ;
      RECT  0.115000  2.360000  0.365000 2.980000 ;
      RECT  0.545000  0.085000  0.795000 0.765000 ;
      RECT  0.565000  2.530000  0.895000 3.245000 ;
      RECT  0.975000  0.350000  1.435000 1.010000 ;
      RECT  0.975000  1.010000  1.145000 1.720000 ;
      RECT  0.975000  1.720000  2.275000 1.890000 ;
      RECT  0.975000  1.890000  1.455000 2.020000 ;
      RECT  1.575000  2.530000  1.905000 3.245000 ;
      RECT  1.615000  0.085000  1.865000 1.010000 ;
      RECT  1.625000  2.060000  2.615000 2.190000 ;
      RECT  1.945000  1.300000  2.275000 1.720000 ;
      RECT  2.045000  0.255000  3.115000 0.425000 ;
      RECT  2.045000  0.425000  2.215000 1.130000 ;
      RECT  2.105000  2.400000  2.275000 2.890000 ;
      RECT  2.105000  2.890000  3.795000 3.060000 ;
      RECT  2.445000  0.595000  2.775000 0.925000 ;
      RECT  2.445000  0.925000  2.615000 2.060000 ;
      RECT  2.445000  2.230000  2.615000 2.260000 ;
      RECT  2.445000  2.260000  2.945000 2.720000 ;
      RECT  2.785000  1.380000  3.115000 2.050000 ;
      RECT  2.945000  0.425000  3.115000 1.380000 ;
      RECT  3.115000  2.260000  3.455000 2.720000 ;
      RECT  3.285000  0.400000  3.615000 1.040000 ;
      RECT  3.285000  1.040000  4.255000 1.210000 ;
      RECT  3.285000  1.210000  3.455000 2.260000 ;
      RECT  3.625000  1.380000  3.915000 2.240000 ;
      RECT  3.625000  2.240000  4.915000 2.410000 ;
      RECT  3.625000  2.410000  3.795000 2.890000 ;
      RECT  4.070000  2.580000  4.575000 2.910000 ;
      RECT  4.070000  2.910000  4.240000 3.245000 ;
      RECT  4.085000  1.210000  4.255000 1.400000 ;
      RECT  4.085000  1.400000  6.245000 1.570000 ;
      RECT  4.230000  1.740000  5.255000 2.070000 ;
      RECT  4.270000  0.085000  4.600000 0.710000 ;
      RECT  4.425000  0.880000  5.160000 1.050000 ;
      RECT  4.425000  1.050000  4.770000 1.230000 ;
      RECT  4.745000  2.410000  4.915000 2.890000 ;
      RECT  4.745000  2.890000  5.690000 3.060000 ;
      RECT  4.770000  0.570000  5.160000 0.880000 ;
      RECT  4.950000  1.220000  6.245000 1.400000 ;
      RECT  5.085000  2.070000  5.255000 2.320000 ;
      RECT  5.085000  2.320000  5.350000 2.720000 ;
      RECT  5.425000  1.790000  6.115000 2.150000 ;
      RECT  5.520000  2.320000  6.585000 2.490000 ;
      RECT  5.520000  2.490000  5.690000 2.890000 ;
      RECT  5.650000  0.085000  6.245000 1.030000 ;
      RECT  5.860000  2.660000  6.110000 3.245000 ;
      RECT  5.915000  1.215000  6.245000 1.220000 ;
      RECT  6.415000  0.280000  7.660000 0.450000 ;
      RECT  6.415000  0.450000  6.585000 1.120000 ;
      RECT  6.415000  1.120000  6.960000 1.450000 ;
      RECT  6.415000  1.450000  6.585000 2.320000 ;
      RECT  6.820000  1.620000  7.320000 1.790000 ;
      RECT  6.820000  1.790000  7.070000 2.550000 ;
      RECT  6.820000  2.550000  7.930000 2.730000 ;
      RECT  6.820000  2.730000  7.470000 2.980000 ;
      RECT  6.825000  0.620000  7.320000 0.950000 ;
      RECT  7.150000  0.950000  7.320000 1.620000 ;
      RECT  7.290000  1.980000  7.660000 2.150000 ;
      RECT  7.290000  2.150000  7.590000 2.380000 ;
      RECT  7.490000  0.450000  7.660000 1.980000 ;
      RECT  7.760000  2.320000  9.470000 2.490000 ;
      RECT  7.760000  2.490000  8.880000 2.550000 ;
      RECT  7.830000  1.070000  9.890000 1.240000 ;
      RECT  7.830000  1.240000  8.145000 2.130000 ;
      RECT  8.100000  2.720000  8.430000 3.245000 ;
      RECT  8.315000  1.480000  8.730000 2.150000 ;
      RECT  8.525000  0.085000  9.360000 0.900000 ;
      RECT  8.630000  2.550000  8.880000 2.980000 ;
      RECT  9.110000  2.660000  9.440000 3.245000 ;
      RECT  9.140000  1.615000  9.470000 2.320000 ;
      RECT  9.530000  0.635000  9.890000 1.070000 ;
      RECT  9.640000  1.240000  9.890000 2.980000 ;
      RECT 10.090000  0.450000 10.420000 1.300000 ;
      RECT 10.090000  1.300000 11.125000 1.630000 ;
      RECT 10.090000  1.630000 10.450000 2.860000 ;
      RECT 10.600000  0.085000 10.930000 1.130000 ;
      RECT 10.655000  2.320000 10.985000 3.245000 ;
      RECT 11.635000  0.085000 11.885000 1.130000 ;
      RECT 11.635000  1.820000 11.885000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  1.950000  6.085000 2.120000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  1.950000  8.485000 2.120000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
  END
END sky130_fd_sc_hs__dfstp_2
MACRO sky130_fd_sc_hs__dfstp_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.96000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.475000 0.980000 0.805000 1.990000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.119700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.680000 0.350000 11.010000 0.980000 ;
        RECT 10.680000 0.980000 12.835000 1.150000 ;
        RECT 11.175000 1.820000 12.835000 2.080000 ;
        RECT 11.175000 2.080000 11.455000 2.980000 ;
        RECT 12.015000 0.350000 12.345000 0.980000 ;
        RECT 12.125000 2.080000 12.835000 2.150000 ;
        RECT 12.125000 2.150000 12.355000 2.980000 ;
        RECT 12.605000 1.150000 12.835000 1.820000 ;
    END
  END Q
  PIN SET_B
    ANTENNAPARTIALMETALSIDEAREA  2.205000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 5.375000 1.550000 5.665000 1.595000 ;
        RECT 5.375000 1.595000 8.545000 1.735000 ;
        RECT 5.375000 1.735000 5.665000 1.780000 ;
        RECT 8.255000 1.550000 8.545000 1.595000 ;
        RECT 8.255000 1.735000 8.545000 1.780000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.315000 1.180000 1.775000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.960000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 12.960000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.960000 0.085000 ;
      RECT  0.000000  3.245000 12.960000 3.415000 ;
      RECT  0.115000  0.350000  0.365000 0.810000 ;
      RECT  0.115000  0.810000  0.285000 2.240000 ;
      RECT  0.115000  2.240000  1.795000 2.410000 ;
      RECT  0.115000  2.410000  0.365000 2.960000 ;
      RECT  0.545000  0.085000  0.795000 0.810000 ;
      RECT  0.565000  2.580000  0.895000 3.245000 ;
      RECT  0.975000  0.340000  1.435000 1.010000 ;
      RECT  0.975000  1.010000  1.145000 1.720000 ;
      RECT  0.975000  1.720000  2.275000 1.890000 ;
      RECT  0.975000  1.890000  1.455000 2.070000 ;
      RECT  1.575000  2.580000  1.905000 3.245000 ;
      RECT  1.615000  0.085000  1.865000 1.010000 ;
      RECT  1.625000  2.070000  2.615000 2.240000 ;
      RECT  1.945000  1.350000  2.275000 1.720000 ;
      RECT  2.045000  0.255000  3.115000 0.425000 ;
      RECT  2.045000  0.425000  2.215000 1.130000 ;
      RECT  2.105000  2.410000  2.275000 2.905000 ;
      RECT  2.105000  2.905000  3.795000 3.075000 ;
      RECT  2.445000  0.595000  2.775000 0.925000 ;
      RECT  2.445000  0.925000  2.615000 2.070000 ;
      RECT  2.445000  2.240000  2.615000 2.295000 ;
      RECT  2.445000  2.295000  2.945000 2.735000 ;
      RECT  2.785000  1.455000  3.115000 2.125000 ;
      RECT  2.945000  0.425000  3.115000 1.455000 ;
      RECT  3.115000  2.295000  3.455000 2.735000 ;
      RECT  3.285000  0.350000  3.535000 1.130000 ;
      RECT  3.285000  1.130000  4.135000 1.300000 ;
      RECT  3.285000  1.300000  3.455000 2.295000 ;
      RECT  3.625000  1.470000  3.795000 2.165000 ;
      RECT  3.625000  2.165000  4.685000 2.335000 ;
      RECT  3.625000  2.335000  3.795000 2.905000 ;
      RECT  3.965000  1.300000  4.135000 1.400000 ;
      RECT  3.965000  1.400000  5.025000 1.570000 ;
      RECT  3.985000  2.505000  4.345000 2.755000 ;
      RECT  3.985000  2.755000  4.155000 3.245000 ;
      RECT  4.025000  0.085000  4.420000 0.600000 ;
      RECT  4.115000  1.740000  5.025000 1.995000 ;
      RECT  4.305000  0.780000  5.050000 0.950000 ;
      RECT  4.305000  0.950000  4.590000 1.230000 ;
      RECT  4.515000  2.335000  4.685000 2.905000 ;
      RECT  4.515000  2.905000  5.510000 3.075000 ;
      RECT  4.590000  0.620000  5.050000 0.780000 ;
      RECT  4.770000  1.120000  5.025000 1.200000 ;
      RECT  4.770000  1.200000  6.135000 1.370000 ;
      RECT  4.770000  1.370000  5.025000 1.400000 ;
      RECT  4.855000  1.995000  5.025000 2.295000 ;
      RECT  4.855000  2.295000  5.170000 2.735000 ;
      RECT  5.195000  1.550000  5.635000 1.925000 ;
      RECT  5.340000  2.095000  6.475000 2.265000 ;
      RECT  5.340000  2.265000  5.510000 2.905000 ;
      RECT  5.670000  0.085000  6.000000 1.030000 ;
      RECT  5.680000  2.435000  5.940000 3.245000 ;
      RECT  5.805000  1.370000  6.135000 1.490000 ;
      RECT  6.305000  0.255000  7.375000 0.425000 ;
      RECT  6.305000  0.425000  6.475000 1.120000 ;
      RECT  6.305000  1.120000  6.695000 1.450000 ;
      RECT  6.305000  1.450000  6.475000 2.095000 ;
      RECT  6.590000  2.650000  7.265000 2.980000 ;
      RECT  6.645000  0.595000  7.035000 0.925000 ;
      RECT  6.670000  1.620000  7.035000 1.790000 ;
      RECT  6.670000  1.790000  6.840000 2.480000 ;
      RECT  6.670000  2.480000  7.715000 2.650000 ;
      RECT  6.865000  0.925000  7.035000 1.620000 ;
      RECT  7.045000  2.020000  7.375000 2.310000 ;
      RECT  7.205000  0.425000  7.375000 2.020000 ;
      RECT  7.545000  0.840000  9.450000 1.010000 ;
      RECT  7.545000  1.010000  7.875000 1.655000 ;
      RECT  7.545000  2.310000  9.110000 2.480000 ;
      RECT  7.885000  2.650000  8.055000 3.245000 ;
      RECT  7.935000  0.085000  8.950000 0.670000 ;
      RECT  8.185000  1.180000  8.515000 1.850000 ;
      RECT  8.255000  2.480000  8.585000 2.980000 ;
      RECT  8.780000  1.370000  9.110000 2.310000 ;
      RECT  8.780000  2.650000  9.030000 3.245000 ;
      RECT  9.120000  0.420000  9.450000 0.840000 ;
      RECT  9.230000  2.650000  9.560000 2.980000 ;
      RECT  9.280000  1.010000  9.450000 2.650000 ;
      RECT  9.680000  0.350000 10.010000 1.320000 ;
      RECT  9.680000  1.320000 11.995000 1.490000 ;
      RECT  9.755000  1.820000 10.005000 3.245000 ;
      RECT 10.180000  0.085000 10.510000 1.130000 ;
      RECT 10.205000  1.490000 11.995000 1.650000 ;
      RECT 10.205000  1.650000 10.535000 2.700000 ;
      RECT 10.725000  1.820000 11.005000 3.245000 ;
      RECT 11.180000  0.085000 11.845000 0.800000 ;
      RECT 11.625000  2.250000 11.955000 3.245000 ;
      RECT 12.515000  0.085000 12.845000 0.810000 ;
      RECT 12.525000  2.320000 12.855000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  1.580000  5.605000 1.750000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  1.580000  8.485000 1.750000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
  END
END sky130_fd_sc_hs__dfstp_4
MACRO sky130_fd_sc_hs__dfxbp_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.600000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.700000 2.025000 2.080000 2.355000 ;
        RECT 1.910000 1.125000 2.270000 1.780000 ;
        RECT 1.910000 1.780000 2.080000 2.025000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.530100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.640000 0.350000 8.070000 1.130000 ;
        RECT 7.665000 2.030000 8.070000 2.980000 ;
        RECT 7.900000 1.130000 8.070000 2.030000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.535700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.140000 0.350000 9.515000 1.130000 ;
        RECT 9.160000 1.820000 9.515000 2.980000 ;
        RECT 9.345000 1.130000 9.515000 1.820000 ;
    END
  END Q_N
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 0.500000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.600000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.600000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.600000 0.085000 ;
      RECT 0.000000  3.245000 9.600000 3.415000 ;
      RECT 0.110000  1.720000 0.840000 1.890000 ;
      RECT 0.110000  1.890000 0.360000 2.980000 ;
      RECT 0.115000  0.350000 0.445000 0.730000 ;
      RECT 0.115000  0.730000 2.545000 0.900000 ;
      RECT 0.115000  0.900000 0.445000 1.010000 ;
      RECT 0.560000  2.060000 0.810000 3.245000 ;
      RECT 0.625000  0.085000 1.005000 0.560000 ;
      RECT 0.670000  0.900000 1.090000 1.550000 ;
      RECT 0.670000  1.550000 0.840000 1.720000 ;
      RECT 1.010000  1.815000 1.435000 2.545000 ;
      RECT 1.010000  2.545000 2.225000 2.715000 ;
      RECT 1.010000  2.715000 1.340000 2.980000 ;
      RECT 1.265000  1.070000 1.595000 1.485000 ;
      RECT 1.265000  1.485000 1.740000 1.815000 ;
      RECT 1.555000  2.885000 1.885000 3.245000 ;
      RECT 1.855000  0.085000 2.205000 0.560000 ;
      RECT 2.055000  2.715000 4.470000 2.755000 ;
      RECT 2.055000  2.755000 3.290000 2.885000 ;
      RECT 2.250000  2.045000 2.610000 2.375000 ;
      RECT 2.375000  0.255000 3.655000 0.425000 ;
      RECT 2.375000  0.425000 2.545000 0.730000 ;
      RECT 2.440000  1.070000 2.885000 1.240000 ;
      RECT 2.440000  1.240000 2.610000 2.045000 ;
      RECT 2.715000  0.595000 2.885000 1.070000 ;
      RECT 2.780000  1.410000 3.315000 1.580000 ;
      RECT 2.780000  1.580000 2.950000 2.245000 ;
      RECT 2.780000  2.245000 4.280000 2.415000 ;
      RECT 2.780000  2.415000 2.950000 2.545000 ;
      RECT 3.065000  0.595000 3.315000 1.410000 ;
      RECT 3.120000  1.750000 3.655000 2.075000 ;
      RECT 3.120000  2.585000 4.470000 2.715000 ;
      RECT 3.485000  0.425000 3.655000 0.580000 ;
      RECT 3.485000  0.580000 5.715000 0.620000 ;
      RECT 3.485000  0.620000 4.650000 0.750000 ;
      RECT 3.485000  0.750000 3.655000 1.750000 ;
      RECT 3.740000  2.925000 4.130000 3.245000 ;
      RECT 3.825000  1.015000 4.900000 1.185000 ;
      RECT 3.825000  1.185000 4.620000 1.370000 ;
      RECT 3.980000  0.085000 4.310000 0.410000 ;
      RECT 4.020000  1.630000 4.280000 2.245000 ;
      RECT 4.300000  2.755000 4.470000 2.800000 ;
      RECT 4.300000  2.800000 5.150000 2.905000 ;
      RECT 4.300000  2.905000 5.990000 3.075000 ;
      RECT 4.450000  1.370000 4.620000 1.855000 ;
      RECT 4.450000  1.855000 4.810000 2.025000 ;
      RECT 4.480000  0.290000 5.715000 0.580000 ;
      RECT 4.570000  0.920000 4.900000 1.015000 ;
      RECT 4.640000  2.025000 4.810000 2.615000 ;
      RECT 4.790000  1.355000 5.150000 1.685000 ;
      RECT 4.980000  1.685000 5.150000 2.800000 ;
      RECT 5.125000  0.790000 5.590000 1.120000 ;
      RECT 5.320000  1.120000 5.590000 1.210000 ;
      RECT 5.320000  1.210000 7.130000 1.380000 ;
      RECT 5.320000  1.380000 5.490000 2.115000 ;
      RECT 5.320000  2.115000 5.570000 2.735000 ;
      RECT 5.660000  1.615000 5.990000 1.945000 ;
      RECT 5.820000  1.945000 5.990000 2.905000 ;
      RECT 6.080000  0.085000 6.410000 1.040000 ;
      RECT 6.165000  2.390000 6.495000 3.245000 ;
      RECT 6.230000  1.550000 6.560000 1.690000 ;
      RECT 6.230000  1.690000 7.730000 1.860000 ;
      RECT 6.230000  1.860000 7.040000 2.220000 ;
      RECT 6.640000  0.440000 6.970000 0.850000 ;
      RECT 6.640000  0.850000 7.470000 1.020000 ;
      RECT 6.710000  2.220000 7.040000 2.860000 ;
      RECT 6.800000  1.190000 7.130000 1.210000 ;
      RECT 6.800000  1.380000 7.130000 1.520000 ;
      RECT 7.140000  0.085000 7.470000 0.680000 ;
      RECT 7.240000  2.030000 7.490000 3.245000 ;
      RECT 7.300000  1.020000 7.470000 1.350000 ;
      RECT 7.300000  1.350000 7.730000 1.690000 ;
      RECT 8.280000  0.625000 8.530000 1.300000 ;
      RECT 8.280000  1.300000 9.175000 1.630000 ;
      RECT 8.280000  1.630000 8.455000 2.700000 ;
      RECT 8.655000  1.820000 8.985000 3.245000 ;
      RECT 8.710000  0.085000 8.960000 1.130000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
  END
END sky130_fd_sc_hs__dfxbp_1
MACRO sky130_fd_sc_hs__dfxbp_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.825000 2.025000 2.155000 2.355000 ;
        RECT 1.985000 1.125000 2.375000 1.780000 ;
        RECT 1.985000 1.780000 2.155000 2.025000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.145000 0.370000 8.450000 1.550000 ;
        RECT 8.145000 1.550000 8.515000 2.070000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.140000 1.820000 10.505000 2.980000 ;
        RECT 10.165000 0.350000 10.505000 1.130000 ;
        RECT 10.335000 1.130000 10.505000 1.820000 ;
    END
  END Q_N
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 0.585000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.040000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 11.040000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  3.245000 11.040000 3.415000 ;
      RECT  0.115000  0.350000  0.445000 0.730000 ;
      RECT  0.115000  0.730000  2.530000 0.900000 ;
      RECT  0.115000  0.900000  1.100000 1.010000 ;
      RECT  0.115000  1.720000  0.925000 1.890000 ;
      RECT  0.115000  1.890000  0.445000 2.980000 ;
      RECT  0.625000  0.085000  1.010000 0.560000 ;
      RECT  0.645000  2.060000  0.895000 3.245000 ;
      RECT  0.755000  1.010000  1.100000 1.550000 ;
      RECT  0.755000  1.550000  0.925000 1.720000 ;
      RECT  1.095000  1.815000  1.440000 2.625000 ;
      RECT  1.095000  2.625000  5.205000 2.795000 ;
      RECT  1.095000  2.795000  1.345000 2.980000 ;
      RECT  1.270000  1.070000  1.600000 1.485000 ;
      RECT  1.270000  1.485000  1.815000 1.815000 ;
      RECT  1.575000  2.965000  2.035000 3.245000 ;
      RECT  1.860000  0.085000  2.190000 0.560000 ;
      RECT  2.325000  2.205000  2.715000 2.455000 ;
      RECT  2.360000  0.255000  3.640000 0.425000 ;
      RECT  2.360000  0.425000  2.530000 0.730000 ;
      RECT  2.545000  1.070000  2.870000 1.240000 ;
      RECT  2.545000  1.240000  2.715000 2.205000 ;
      RECT  2.700000  0.595000  2.870000 1.070000 ;
      RECT  2.885000  1.410000  3.300000 1.580000 ;
      RECT  2.885000  1.580000  3.055000 2.285000 ;
      RECT  2.885000  2.285000  4.325000 2.455000 ;
      RECT  3.050000  0.595000  3.300000 1.410000 ;
      RECT  3.225000  1.750000  3.640000 2.065000 ;
      RECT  3.470000  0.425000  3.640000 0.780000 ;
      RECT  3.470000  0.780000  4.815000 0.950000 ;
      RECT  3.470000  0.950000  3.640000 1.750000 ;
      RECT  3.810000  1.120000  4.815000 1.450000 ;
      RECT  4.000000  2.965000  4.330000 3.245000 ;
      RECT  4.030000  0.085000  4.370000 0.610000 ;
      RECT  4.155000  1.630000  4.475000 1.960000 ;
      RECT  4.155000  1.960000  4.325000 2.285000 ;
      RECT  4.535000  2.180000  4.865000 2.455000 ;
      RECT  4.645000  0.255000  6.240000 0.530000 ;
      RECT  4.645000  0.530000  4.815000 0.780000 ;
      RECT  4.645000  1.450000  4.815000 2.180000 ;
      RECT  4.985000  1.120000  5.275000 1.450000 ;
      RECT  5.035000  1.450000  5.205000 2.625000 ;
      RECT  5.035000  2.795000  6.205000 2.965000 ;
      RECT  5.375000  1.620000  6.545000 1.670000 ;
      RECT  5.375000  1.670000  7.585000 1.790000 ;
      RECT  5.375000  1.790000  5.705000 2.625000 ;
      RECT  5.445000  0.530000  5.615000 1.170000 ;
      RECT  5.445000  1.170000  5.845000 1.450000 ;
      RECT  5.785000  0.700000  6.185000 0.950000 ;
      RECT  5.875000  1.960000  6.205000 2.795000 ;
      RECT  6.015000  0.950000  6.185000 1.620000 ;
      RECT  6.375000  1.790000  7.585000 1.960000 ;
      RECT  6.600000  2.375000  6.930000 3.245000 ;
      RECT  6.655000  0.085000  6.985000 1.000000 ;
      RECT  6.715000  1.170000  7.465000 1.330000 ;
      RECT  6.715000  1.330000  7.925000 1.500000 ;
      RECT  7.160000  2.130000  7.925000 2.240000 ;
      RECT  7.160000  2.240000  9.015000 2.410000 ;
      RECT  7.160000  2.410000  7.490000 2.980000 ;
      RECT  7.215000  0.370000  7.465000 1.170000 ;
      RECT  7.645000  0.085000  7.975000 1.150000 ;
      RECT  7.695000  2.580000  8.025000 3.245000 ;
      RECT  7.755000  1.500000  7.925000 2.130000 ;
      RECT  8.595000  2.580000  8.925000 3.245000 ;
      RECT  8.620000  0.085000  8.950000 1.150000 ;
      RECT  8.685000  1.320000  9.015000 2.240000 ;
      RECT  9.235000  0.540000  9.510000 1.300000 ;
      RECT  9.235000  1.300000 10.165000 1.630000 ;
      RECT  9.235000  1.630000  9.485000 2.860000 ;
      RECT  9.690000  1.820000  9.940000 3.245000 ;
      RECT  9.735000  0.085000  9.985000 1.130000 ;
      RECT 10.675000  0.085000 10.925000 1.130000 ;
      RECT 10.675000  1.820000 10.925000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
  END
END sky130_fd_sc_hs__dfxbp_2
MACRO sky130_fd_sc_hs__dfxtp_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.870000 2.025000 2.250000 2.355000 ;
        RECT 1.970000 1.125000 2.250000 2.025000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.715000 0.350000 8.075000 1.130000 ;
        RECT 7.715000 2.030000 8.075000 2.980000 ;
        RECT 7.905000 1.130000 8.075000 2.030000 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.505000 1.780000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.115000  0.350000 0.365000 0.960000 ;
      RECT 0.115000  0.960000 1.135000 1.130000 ;
      RECT 0.115000  1.950000 0.845000 2.120000 ;
      RECT 0.115000  2.120000 0.445000 2.980000 ;
      RECT 0.545000  0.085000 0.795000 0.790000 ;
      RECT 0.645000  2.290000 0.815000 3.245000 ;
      RECT 0.675000  1.130000 1.135000 1.550000 ;
      RECT 0.675000  1.550000 0.845000 1.950000 ;
      RECT 0.965000  0.255000 1.815000 0.425000 ;
      RECT 0.965000  0.425000 1.135000 0.960000 ;
      RECT 1.015000  1.820000 1.475000 2.625000 ;
      RECT 1.015000  2.625000 2.250000 2.795000 ;
      RECT 1.015000  2.795000 1.345000 2.980000 ;
      RECT 1.305000  0.595000 1.475000 1.350000 ;
      RECT 1.305000  1.350000 1.760000 1.680000 ;
      RECT 1.305000  1.680000 1.475000 1.820000 ;
      RECT 1.575000  2.965000 1.910000 3.245000 ;
      RECT 1.645000  0.425000 1.815000 0.730000 ;
      RECT 1.645000  0.730000 2.655000 0.900000 ;
      RECT 1.985000  0.085000 2.315000 0.560000 ;
      RECT 2.080000  2.795000 3.460000 2.965000 ;
      RECT 2.420000  1.070000 2.975000 1.240000 ;
      RECT 2.420000  1.240000 2.590000 2.625000 ;
      RECT 2.485000  0.275000 3.760000 0.445000 ;
      RECT 2.485000  0.445000 2.655000 0.730000 ;
      RECT 2.760000  1.410000 3.420000 1.580000 ;
      RECT 2.760000  1.580000 2.930000 2.285000 ;
      RECT 2.760000  2.285000 4.140000 2.455000 ;
      RECT 2.760000  2.455000 3.120000 2.625000 ;
      RECT 3.100000  1.750000 3.760000 2.080000 ;
      RECT 3.155000  0.615000 3.420000 1.410000 ;
      RECT 3.290000  2.625000 4.950000 2.795000 ;
      RECT 3.590000  0.445000 3.760000 0.690000 ;
      RECT 3.590000  0.690000 4.660000 0.860000 ;
      RECT 3.590000  0.860000 3.760000 1.750000 ;
      RECT 3.800000  2.965000 4.130000 3.245000 ;
      RECT 3.930000  1.030000 5.000000 1.200000 ;
      RECT 3.930000  1.200000 4.260000 1.415000 ;
      RECT 3.970000  1.625000 4.270000 1.955000 ;
      RECT 3.970000  1.955000 4.140000 2.285000 ;
      RECT 4.070000  0.085000 4.320000 0.520000 ;
      RECT 4.335000  2.125000 4.610000 2.455000 ;
      RECT 4.440000  1.200000 4.610000 2.125000 ;
      RECT 4.490000  0.255000 5.895000 0.425000 ;
      RECT 4.490000  0.425000 4.660000 0.690000 ;
      RECT 4.780000  1.370000 5.480000 1.540000 ;
      RECT 4.780000  1.540000 4.950000 2.625000 ;
      RECT 4.780000  2.795000 4.950000 2.905000 ;
      RECT 4.780000  2.905000 5.840000 3.075000 ;
      RECT 4.830000  0.595000 5.000000 1.030000 ;
      RECT 5.120000  1.710000 5.820000 1.880000 ;
      RECT 5.120000  1.880000 5.290000 2.735000 ;
      RECT 5.170000  1.150000 5.480000 1.370000 ;
      RECT 5.220000  0.730000 5.820000 0.980000 ;
      RECT 5.510000  2.050000 5.840000 2.905000 ;
      RECT 5.565000  0.425000 5.895000 0.510000 ;
      RECT 5.650000  0.980000 5.820000 1.230000 ;
      RECT 5.650000  1.230000 7.205000 1.400000 ;
      RECT 5.650000  1.400000 5.820000 1.710000 ;
      RECT 6.050000  1.570000 6.380000 1.690000 ;
      RECT 6.050000  1.690000 7.735000 1.860000 ;
      RECT 6.050000  1.860000 6.380000 2.240000 ;
      RECT 6.200000  2.520000 6.530000 3.245000 ;
      RECT 6.230000  0.085000 6.560000 1.060000 ;
      RECT 6.760000  1.860000 7.010000 2.700000 ;
      RECT 6.790000  0.350000 7.040000 0.850000 ;
      RECT 6.790000  0.850000 7.545000 1.020000 ;
      RECT 6.875000  1.190000 7.205000 1.230000 ;
      RECT 6.875000  1.400000 7.205000 1.520000 ;
      RECT 7.210000  2.030000 7.540000 3.245000 ;
      RECT 7.220000  0.085000 7.535000 0.680000 ;
      RECT 7.375000  1.020000 7.545000 1.350000 ;
      RECT 7.375000  1.350000 7.735000 1.690000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_hs__dfxtp_1
MACRO sky130_fd_sc_hs__dfxtp_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.725000 2.050000 2.055000 2.380000 ;
        RECT 1.885000 1.150000 2.275000 1.480000 ;
        RECT 1.885000 1.480000 2.055000 2.050000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.745000 2.030000 8.105000 2.980000 ;
        RECT 7.765000 0.350000 8.105000 1.130000 ;
        RECT 7.935000 1.130000 8.105000 2.030000 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.505000 1.780000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
      RECT 0.000000  3.245000 8.640000 3.415000 ;
      RECT 0.115000  0.350000 0.365000 0.960000 ;
      RECT 0.115000  0.960000 1.135000 1.130000 ;
      RECT 0.115000  1.950000 0.845000 2.120000 ;
      RECT 0.115000  2.120000 0.445000 2.980000 ;
      RECT 0.545000  0.085000 0.795000 0.790000 ;
      RECT 0.645000  2.290000 0.815000 3.245000 ;
      RECT 0.675000  1.130000 1.135000 1.550000 ;
      RECT 0.675000  1.550000 0.845000 1.950000 ;
      RECT 0.965000  0.255000 1.815000 0.425000 ;
      RECT 0.965000  0.425000 1.135000 0.960000 ;
      RECT 1.015000  1.720000 1.475000 2.625000 ;
      RECT 1.015000  2.625000 2.275000 2.755000 ;
      RECT 1.015000  2.755000 4.990000 2.795000 ;
      RECT 1.015000  2.795000 1.345000 2.980000 ;
      RECT 1.305000  0.595000 1.475000 1.350000 ;
      RECT 1.305000  1.350000 1.715000 1.720000 ;
      RECT 1.575000  2.965000 1.935000 3.245000 ;
      RECT 1.645000  0.425000 1.815000 0.810000 ;
      RECT 1.645000  0.810000 2.520000 0.980000 ;
      RECT 1.985000  0.085000 2.180000 0.640000 ;
      RECT 2.105000  2.795000 3.540000 2.925000 ;
      RECT 2.225000  1.650000 2.615000 1.820000 ;
      RECT 2.225000  1.820000 2.555000 2.455000 ;
      RECT 2.350000  0.255000 3.755000 0.425000 ;
      RECT 2.350000  0.425000 2.520000 0.810000 ;
      RECT 2.445000  1.150000 2.860000 1.320000 ;
      RECT 2.445000  1.320000 2.615000 1.650000 ;
      RECT 2.690000  0.595000 2.860000 1.150000 ;
      RECT 2.755000  2.125000 2.955000 2.255000 ;
      RECT 2.755000  2.255000 4.135000 2.425000 ;
      RECT 2.755000  2.425000 2.955000 2.585000 ;
      RECT 2.785000  1.490000 3.200000 1.660000 ;
      RECT 2.785000  1.660000 2.955000 2.125000 ;
      RECT 3.030000  0.615000 3.415000 0.945000 ;
      RECT 3.030000  0.945000 3.200000 1.490000 ;
      RECT 3.140000  1.830000 3.540000 2.085000 ;
      RECT 3.370000  1.285000 3.755000 1.455000 ;
      RECT 3.370000  1.455000 3.540000 1.830000 ;
      RECT 3.370000  2.625000 4.990000 2.755000 ;
      RECT 3.585000  0.425000 3.755000 0.690000 ;
      RECT 3.585000  0.690000 4.575000 0.860000 ;
      RECT 3.585000  0.860000 3.755000 1.285000 ;
      RECT 3.710000  2.965000 4.100000 3.245000 ;
      RECT 3.925000  1.030000 4.915000 1.200000 ;
      RECT 3.925000  1.200000 4.650000 1.415000 ;
      RECT 3.965000  1.625000 4.310000 1.955000 ;
      RECT 3.965000  1.955000 4.135000 2.255000 ;
      RECT 3.985000  0.085000 4.235000 0.520000 ;
      RECT 4.305000  2.125000 4.650000 2.455000 ;
      RECT 4.405000  0.255000 5.890000 0.425000 ;
      RECT 4.405000  0.425000 4.575000 0.690000 ;
      RECT 4.480000  1.415000 4.650000 2.125000 ;
      RECT 4.745000  0.595000 5.075000 0.945000 ;
      RECT 4.745000  0.945000 4.915000 1.030000 ;
      RECT 4.820000  1.370000 5.415000 1.540000 ;
      RECT 4.820000  1.540000 4.990000 2.625000 ;
      RECT 4.820000  2.795000 4.990000 2.905000 ;
      RECT 4.820000  2.905000 5.875000 3.075000 ;
      RECT 5.085000  1.150000 5.415000 1.370000 ;
      RECT 5.160000  1.710000 5.755000 1.880000 ;
      RECT 5.160000  1.880000 5.330000 2.735000 ;
      RECT 5.245000  0.695000 5.755000 0.945000 ;
      RECT 5.545000  2.050000 5.875000 2.905000 ;
      RECT 5.560000  0.425000 5.890000 0.510000 ;
      RECT 5.585000  0.945000 5.755000 1.230000 ;
      RECT 5.585000  1.230000 7.240000 1.400000 ;
      RECT 5.585000  1.400000 5.755000 1.710000 ;
      RECT 6.085000  1.570000 6.415000 1.690000 ;
      RECT 6.085000  1.690000 7.765000 1.860000 ;
      RECT 6.085000  1.860000 6.415000 2.240000 ;
      RECT 6.225000  0.085000 6.555000 1.060000 ;
      RECT 6.235000  2.520000 6.565000 3.245000 ;
      RECT 6.785000  0.350000 7.115000 0.850000 ;
      RECT 6.785000  0.850000 7.595000 1.020000 ;
      RECT 6.790000  1.860000 7.040000 2.860000 ;
      RECT 6.910000  1.190000 7.240000 1.230000 ;
      RECT 6.910000  1.400000 7.240000 1.520000 ;
      RECT 7.240000  2.030000 7.570000 3.245000 ;
      RECT 7.300000  0.085000 7.595000 0.680000 ;
      RECT 7.425000  1.020000 7.595000 1.350000 ;
      RECT 7.425000  1.350000 7.765000 1.690000 ;
      RECT 8.275000  0.085000 8.525000 1.130000 ;
      RECT 8.275000  1.820000 8.525000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
  END
END sky130_fd_sc_hs__dfxtp_2
MACRO sky130_fd_sc_hs__dfxtp_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.600000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.785000 2.025000 2.115000 2.355000 ;
        RECT 1.945000 1.125000 2.305000 1.780000 ;
        RECT 1.945000 1.780000 2.115000 2.025000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.116000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.805000 1.800000 9.035000 1.970000 ;
        RECT 7.805000 1.970000 8.135000 2.980000 ;
        RECT 7.820000 0.350000 8.150000 0.960000 ;
        RECT 7.820000 0.960000 9.035000 1.130000 ;
        RECT 8.700000 0.350000 9.035000 0.960000 ;
        RECT 8.705000 1.970000 9.035000 2.980000 ;
        RECT 8.865000 1.130000 9.035000 1.800000 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.505000 1.780000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.600000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.600000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.600000 0.085000 ;
      RECT 0.000000  3.245000 9.600000 3.415000 ;
      RECT 0.115000  0.350000 0.445000 0.960000 ;
      RECT 0.115000  0.960000 1.135000 1.130000 ;
      RECT 0.115000  1.950000 0.845000 2.120000 ;
      RECT 0.115000  2.120000 0.445000 2.980000 ;
      RECT 0.625000  0.085000 0.795000 0.790000 ;
      RECT 0.645000  2.290000 0.815000 3.245000 ;
      RECT 0.675000  1.130000 1.135000 1.550000 ;
      RECT 0.675000  1.550000 0.845000 1.950000 ;
      RECT 0.965000  0.255000 1.815000 0.425000 ;
      RECT 0.965000  0.425000 1.135000 0.960000 ;
      RECT 1.015000  1.820000 1.475000 2.525000 ;
      RECT 1.015000  2.525000 2.165000 2.695000 ;
      RECT 1.015000  2.695000 1.475000 2.980000 ;
      RECT 1.305000  0.595000 1.475000 1.220000 ;
      RECT 1.305000  1.220000 1.765000 1.550000 ;
      RECT 1.305000  1.550000 1.475000 1.820000 ;
      RECT 1.645000  0.425000 1.815000 0.730000 ;
      RECT 1.645000  0.730000 2.655000 0.900000 ;
      RECT 1.655000  2.865000 1.825000 3.245000 ;
      RECT 1.985000  0.085000 2.315000 0.560000 ;
      RECT 1.995000  2.695000 2.165000 2.905000 ;
      RECT 1.995000  2.905000 3.375000 3.075000 ;
      RECT 2.335000  1.950000 2.645000 2.120000 ;
      RECT 2.335000  2.120000 2.505000 2.735000 ;
      RECT 2.475000  1.070000 2.995000 1.240000 ;
      RECT 2.475000  1.240000 2.645000 1.950000 ;
      RECT 2.485000  0.255000 3.875000 0.425000 ;
      RECT 2.485000  0.425000 2.655000 0.730000 ;
      RECT 2.705000  2.485000 3.035000 2.735000 ;
      RECT 2.815000  1.410000 3.345000 1.580000 ;
      RECT 2.815000  1.580000 2.985000 2.250000 ;
      RECT 2.815000  2.250000 4.385000 2.420000 ;
      RECT 2.815000  2.420000 3.035000 2.485000 ;
      RECT 2.825000  0.595000 2.995000 1.070000 ;
      RECT 3.155000  1.750000 3.875000 2.080000 ;
      RECT 3.175000  0.620000 3.535000 0.950000 ;
      RECT 3.175000  0.950000 3.345000 1.410000 ;
      RECT 3.205000  2.590000 4.385000 2.760000 ;
      RECT 3.205000  2.760000 3.375000 2.905000 ;
      RECT 3.705000  0.425000 3.875000 0.690000 ;
      RECT 3.705000  0.690000 4.680000 0.860000 ;
      RECT 3.705000  0.860000 3.875000 1.750000 ;
      RECT 3.715000  2.930000 4.045000 3.245000 ;
      RECT 4.045000  1.030000 5.020000 1.200000 ;
      RECT 4.045000  1.200000 4.725000 1.370000 ;
      RECT 4.055000  1.630000 4.385000 2.250000 ;
      RECT 4.090000  0.085000 4.340000 0.520000 ;
      RECT 4.215000  2.760000 4.385000 2.905000 ;
      RECT 4.215000  2.905000 5.955000 3.075000 ;
      RECT 4.510000  0.255000 5.995000 0.425000 ;
      RECT 4.510000  0.425000 4.680000 0.690000 ;
      RECT 4.555000  1.370000 4.725000 2.735000 ;
      RECT 4.850000  0.595000 5.180000 0.950000 ;
      RECT 4.850000  0.950000 5.020000 1.030000 ;
      RECT 4.895000  1.370000 5.520000 1.540000 ;
      RECT 4.895000  1.540000 5.065000 2.905000 ;
      RECT 5.190000  1.150000 5.520000 1.370000 ;
      RECT 5.235000  1.710000 5.860000 1.880000 ;
      RECT 5.235000  1.880000 5.405000 2.735000 ;
      RECT 5.350000  0.720000 5.860000 0.970000 ;
      RECT 5.625000  2.050000 5.955000 2.905000 ;
      RECT 5.665000  0.425000 5.995000 0.510000 ;
      RECT 5.690000  0.970000 5.860000 1.140000 ;
      RECT 5.690000  1.140000 6.800000 1.220000 ;
      RECT 5.690000  1.220000 7.130000 1.310000 ;
      RECT 5.690000  1.310000 5.860000 1.710000 ;
      RECT 6.130000  1.480000 6.460000 1.720000 ;
      RECT 6.130000  1.720000 7.470000 1.810000 ;
      RECT 6.290000  1.810000 7.470000 1.890000 ;
      RECT 6.315000  2.450000 6.650000 3.245000 ;
      RECT 6.410000  0.085000 6.660000 0.970000 ;
      RECT 6.630000  1.310000 7.130000 1.390000 ;
      RECT 6.800000  1.390000 7.130000 1.550000 ;
      RECT 6.820000  1.890000 7.150000 2.980000 ;
      RECT 6.890000  0.350000 7.140000 0.880000 ;
      RECT 6.890000  0.880000 7.470000 0.970000 ;
      RECT 6.970000  0.970000 7.470000 1.050000 ;
      RECT 7.300000  1.050000 7.470000 1.300000 ;
      RECT 7.300000  1.300000 8.665000 1.630000 ;
      RECT 7.300000  1.630000 7.470000 1.720000 ;
      RECT 7.320000  0.085000 7.650000 0.710000 ;
      RECT 7.355000  2.060000 7.605000 3.245000 ;
      RECT 8.330000  0.085000 8.500000 0.790000 ;
      RECT 8.335000  2.140000 8.505000 3.245000 ;
      RECT 9.210000  0.085000 9.460000 1.130000 ;
      RECT 9.235000  1.820000 9.485000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
  END
END sky130_fd_sc_hs__dfxtp_4
MACRO sky130_fd_sc_hs__diode_2
  CLASS CORE ANTENNACELL ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.960000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN DIODE
    ANTENNADIFFAREA  0.641700 ;
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.265000 0.865000 3.065000 ;
    END
  END DIODE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 0.960000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 0.960000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.960000 0.085000 ;
      RECT 0.000000  3.245000 0.960000 3.415000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
  END
END sky130_fd_sc_hs__diode_2
MACRO sky130_fd_sc_hs__dlclkp_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN GATE
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.470000 1.335000 1.800000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.205000 1.550000 6.605000 2.980000 ;
        RECT 6.275000 0.350000 6.605000 1.550000 ;
    END
  END GCLK
  PIN CLK
    ANTENNAGATEAREA  0.459000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.475000 5.155000 1.805000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.720000 0.085000 ;
      RECT 0.000000  3.245000 6.720000 3.415000 ;
      RECT 0.095000  0.350000 0.445000 0.790000 ;
      RECT 0.095000  0.790000 1.215000 0.960000 ;
      RECT 0.095000  0.960000 0.445000 1.130000 ;
      RECT 0.095000  1.130000 0.265000 1.820000 ;
      RECT 0.095000  1.820000 0.445000 2.980000 ;
      RECT 0.435000  1.300000 0.785000 1.630000 ;
      RECT 0.615000  1.130000 1.555000 1.300000 ;
      RECT 0.615000  1.630000 0.785000 1.970000 ;
      RECT 0.615000  1.970000 1.555000 2.140000 ;
      RECT 0.615000  2.310000 0.945000 3.245000 ;
      RECT 0.625000  0.085000 0.875000 0.620000 ;
      RECT 1.045000  0.255000 2.955000 0.425000 ;
      RECT 1.045000  0.425000 1.215000 0.790000 ;
      RECT 1.385000  0.650000 2.260000 0.980000 ;
      RECT 1.385000  0.980000 1.555000 1.130000 ;
      RECT 1.385000  2.140000 1.555000 2.550000 ;
      RECT 1.385000  2.550000 2.285000 2.880000 ;
      RECT 1.725000  1.150000 1.995000 2.050000 ;
      RECT 1.725000  2.050000 3.200000 2.380000 ;
      RECT 2.205000  1.160000 3.775000 1.330000 ;
      RECT 2.205000  1.330000 2.535000 1.840000 ;
      RECT 2.625000  0.425000 2.955000 0.510000 ;
      RECT 2.750000  0.685000 3.295000 0.935000 ;
      RECT 2.835000  2.730000 3.165000 3.245000 ;
      RECT 3.030000  1.500000 3.435000 1.830000 ;
      RECT 3.030000  1.830000 3.200000 2.050000 ;
      RECT 3.030000  2.380000 3.200000 2.390000 ;
      RECT 3.030000  2.390000 4.260000 2.560000 ;
      RECT 3.125000  0.085000 3.295000 0.685000 ;
      RECT 3.370000  2.050000 3.775000 2.220000 ;
      RECT 3.465000  0.605000 3.775000 1.160000 ;
      RECT 3.605000  1.330000 3.775000 2.050000 ;
      RECT 3.945000  1.055000 4.205000 1.945000 ;
      RECT 3.945000  1.945000 4.260000 2.390000 ;
      RECT 3.945000  2.560000 4.260000 2.825000 ;
      RECT 4.385000  0.085000 4.715000 1.305000 ;
      RECT 4.430000  1.975000 4.760000 3.245000 ;
      RECT 4.930000  1.975000 5.535000 2.145000 ;
      RECT 4.930000  2.145000 5.260000 2.825000 ;
      RECT 5.285000  0.605000 5.615000 1.285000 ;
      RECT 5.365000  1.285000 5.615000 1.300000 ;
      RECT 5.365000  1.300000 6.035000 1.630000 ;
      RECT 5.365000  1.630000 5.535000 1.975000 ;
      RECT 5.705000  1.945000 6.035000 3.245000 ;
      RECT 5.845000  0.085000 6.095000 1.130000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
  END
END sky130_fd_sc_hs__dlclkp_1
MACRO sky130_fd_sc_hs__dlclkp_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN GATE
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.450000 1.335000 1.780000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.805000 0.440000 7.135000 2.980000 ;
    END
  END GCLK
  PIN CLK
    ANTENNAGATEAREA  0.498000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.550000 1.445000 5.220000 1.780000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.680000 0.085000 ;
      RECT 0.000000  3.245000 7.680000 3.415000 ;
      RECT 0.095000  0.350000 0.365000 0.770000 ;
      RECT 0.095000  0.770000 1.220000 0.940000 ;
      RECT 0.095000  0.940000 0.265000 1.820000 ;
      RECT 0.095000  1.820000 0.445000 2.980000 ;
      RECT 0.435000  1.110000 1.560000 1.280000 ;
      RECT 0.435000  1.280000 0.785000 1.550000 ;
      RECT 0.545000  0.085000 0.880000 0.600000 ;
      RECT 0.615000  1.550000 0.785000 1.950000 ;
      RECT 0.615000  1.950000 1.705000 2.120000 ;
      RECT 0.685000  2.290000 1.075000 3.245000 ;
      RECT 1.050000  0.255000 3.160000 0.425000 ;
      RECT 1.050000  0.425000 1.220000 0.770000 ;
      RECT 1.390000  0.620000 2.245000 0.950000 ;
      RECT 1.390000  0.950000 1.560000 1.110000 ;
      RECT 1.535000  2.120000 1.705000 2.550000 ;
      RECT 1.535000  2.550000 2.405000 2.880000 ;
      RECT 1.730000  1.120000 2.045000 1.450000 ;
      RECT 1.875000  1.450000 2.045000 2.050000 ;
      RECT 1.875000  2.050000 3.325000 2.220000 ;
      RECT 2.225000  2.220000 2.555000 2.380000 ;
      RECT 2.255000  1.215000 4.035000 1.385000 ;
      RECT 2.255000  1.385000 2.585000 1.840000 ;
      RECT 2.830000  0.425000 3.160000 0.585000 ;
      RECT 2.920000  0.755000 3.535000 1.005000 ;
      RECT 2.945000  2.650000 3.485000 3.245000 ;
      RECT 3.155000  1.555000 3.485000 1.885000 ;
      RECT 3.155000  1.885000 3.325000 2.050000 ;
      RECT 3.340000  0.085000 3.535000 0.755000 ;
      RECT 3.655000  1.385000 3.825000 2.100000 ;
      RECT 3.655000  2.100000 3.985000 2.980000 ;
      RECT 3.705000  0.605000 4.035000 1.215000 ;
      RECT 3.995000  1.555000 4.380000 1.885000 ;
      RECT 4.210000  0.575000 4.595000 1.275000 ;
      RECT 4.210000  1.275000 4.380000 1.555000 ;
      RECT 4.210000  1.885000 4.380000 2.075000 ;
      RECT 4.210000  2.075000 4.545000 2.955000 ;
      RECT 4.715000  2.075000 5.045000 3.245000 ;
      RECT 4.765000  0.085000 5.095000 1.275000 ;
      RECT 5.215000  1.950000 5.560000 2.955000 ;
      RECT 5.390000  0.940000 6.305000 1.610000 ;
      RECT 5.390000  1.610000 5.560000 1.950000 ;
      RECT 5.555000  0.575000 5.885000 0.940000 ;
      RECT 5.730000  1.950000 6.635000 3.245000 ;
      RECT 6.305000  0.085000 6.635000 0.770000 ;
      RECT 7.315000  0.085000 7.565000 1.220000 ;
      RECT 7.315000  1.820000 7.565000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
  END
END sky130_fd_sc_hs__dlclkp_2
MACRO sky130_fd_sc_hs__dlclkp_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN GATE
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.530000 1.430000 1.800000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  1.103200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.795000 1.550000 8.515000 1.720000 ;
        RECT 6.795000 1.720000 7.125000 2.980000 ;
        RECT 6.835000 0.350000 7.165000 1.210000 ;
        RECT 6.835000 1.210000 8.015000 1.380000 ;
        RECT 7.745000 1.720000 8.515000 1.780000 ;
        RECT 7.745000 1.780000 7.995000 2.980000 ;
        RECT 7.765000 0.350000 8.015000 1.210000 ;
        RECT 7.805000 1.380000 8.015000 1.550000 ;
    END
  END GCLK
  PIN CLK
    ANTENNAGATEAREA  0.516000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.400000 1.360000 5.070000 1.780000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
      RECT 0.000000  3.245000 8.640000 3.415000 ;
      RECT 0.115000  0.350000 0.365000 0.850000 ;
      RECT 0.115000  0.850000 1.265000 1.020000 ;
      RECT 0.115000  1.020000 0.365000 1.820000 ;
      RECT 0.115000  1.820000 0.540000 2.980000 ;
      RECT 0.535000  1.190000 1.605000 1.360000 ;
      RECT 0.535000  1.360000 0.880000 1.550000 ;
      RECT 0.550000  0.085000 0.925000 0.680000 ;
      RECT 0.710000  1.550000 0.880000 1.970000 ;
      RECT 0.710000  1.970000 1.605000 2.140000 ;
      RECT 0.785000  2.310000 1.160000 3.245000 ;
      RECT 1.095000  0.255000 3.145000 0.425000 ;
      RECT 1.095000  0.425000 1.265000 0.850000 ;
      RECT 1.435000  0.650000 2.330000 0.980000 ;
      RECT 1.435000  0.980000 1.605000 1.190000 ;
      RECT 1.435000  2.140000 1.605000 2.520000 ;
      RECT 1.435000  2.520000 2.485000 2.850000 ;
      RECT 1.775000  1.150000 2.065000 2.050000 ;
      RECT 1.775000  2.050000 3.475000 2.350000 ;
      RECT 2.305000  1.360000 4.155000 1.530000 ;
      RECT 2.305000  1.530000 2.635000 1.805000 ;
      RECT 2.815000  0.425000 3.145000 1.020000 ;
      RECT 2.815000  1.020000 5.430000 1.190000 ;
      RECT 3.110000  2.860000 3.440000 3.245000 ;
      RECT 3.305000  1.700000 3.655000 1.960000 ;
      RECT 3.305000  1.960000 3.475000 2.050000 ;
      RECT 3.305000  2.350000 3.475000 2.520000 ;
      RECT 3.305000  2.520000 4.535000 2.690000 ;
      RECT 3.315000  0.085000 3.645000 0.850000 ;
      RECT 3.645000  2.180000 3.995000 2.350000 ;
      RECT 3.815000  0.255000 4.610000 0.515000 ;
      RECT 3.825000  1.530000 4.155000 1.610000 ;
      RECT 3.825000  1.610000 3.995000 2.180000 ;
      RECT 4.205000  2.090000 4.535000 2.520000 ;
      RECT 4.205000  2.690000 4.535000 2.970000 ;
      RECT 4.280000  0.515000 4.610000 0.850000 ;
      RECT 4.740000  2.090000 5.070000 3.245000 ;
      RECT 4.780000  0.085000 5.110000 0.850000 ;
      RECT 5.240000  1.820000 6.350000 1.990000 ;
      RECT 5.240000  1.990000 5.570000 2.980000 ;
      RECT 5.260000  1.190000 5.430000 1.300000 ;
      RECT 5.260000  1.300000 5.805000 1.630000 ;
      RECT 5.600000  0.350000 5.975000 0.670000 ;
      RECT 5.600000  0.670000 6.350000 1.130000 ;
      RECT 5.740000  2.160000 6.625000 3.245000 ;
      RECT 5.975000  1.130000 6.350000 1.820000 ;
      RECT 6.160000  0.085000 6.655000 0.500000 ;
      RECT 7.295000  1.890000 7.545000 3.245000 ;
      RECT 7.335000  0.085000 7.585000 1.040000 ;
      RECT 8.195000  0.085000 8.525000 1.040000 ;
      RECT 8.195000  1.950000 8.525000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
  END
END sky130_fd_sc_hs__dlclkp_4
MACRO sky130_fd_sc_hs__dlrbn_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.435000 1.260000 0.835000 1.900000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.535700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.565000 0.350000 7.115000 1.050000 ;
        RECT 6.690000 1.720000 7.115000 2.850000 ;
        RECT 6.945000 1.050000 7.115000 1.720000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.195000 1.820000 8.530000 2.980000 ;
        RECT 8.245000 0.350000 8.530000 1.130000 ;
        RECT 8.360000 1.130000 8.530000 1.820000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.875000 1.180000 6.180000 1.550000 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.260000 1.335000 1.900000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
      RECT 0.000000  3.245000 8.640000 3.415000 ;
      RECT 0.095000  0.540000 0.450000 1.090000 ;
      RECT 0.095000  1.090000 0.265000 2.070000 ;
      RECT 0.095000  2.070000 1.235000 2.240000 ;
      RECT 0.095000  2.240000 0.365000 2.980000 ;
      RECT 0.565000  2.410000 0.895000 3.245000 ;
      RECT 0.630000  0.085000 0.960000 1.090000 ;
      RECT 1.065000  2.240000 1.235000 2.730000 ;
      RECT 1.065000  2.730000 2.015000 2.900000 ;
      RECT 1.130000  0.350000 1.675000 1.090000 ;
      RECT 1.405000  2.100000 1.675000 2.220000 ;
      RECT 1.405000  2.220000 2.555000 2.390000 ;
      RECT 1.405000  2.390000 1.675000 2.560000 ;
      RECT 1.505000  1.090000 1.675000 2.100000 ;
      RECT 1.845000  0.350000 2.175000 0.780000 ;
      RECT 1.845000  0.780000 4.205000 0.950000 ;
      RECT 1.845000  0.950000 2.175000 0.960000 ;
      RECT 1.845000  0.960000 2.015000 1.720000 ;
      RECT 1.845000  1.720000 2.215000 2.050000 ;
      RECT 1.845000  2.560000 2.910000 2.730000 ;
      RECT 2.185000  1.130000 3.610000 1.300000 ;
      RECT 2.185000  1.300000 2.555000 1.550000 ;
      RECT 2.345000  0.085000 2.915000 0.600000 ;
      RECT 2.385000  1.550000 2.555000 2.220000 ;
      RECT 2.505000  2.900000 2.835000 3.245000 ;
      RECT 2.740000  1.470000 3.070000 1.800000 ;
      RECT 2.740000  1.800000 2.910000 2.560000 ;
      RECT 3.120000  1.970000 3.450000 2.140000 ;
      RECT 3.120000  2.140000 3.290000 2.905000 ;
      RECT 3.120000  2.905000 4.290000 3.075000 ;
      RECT 3.280000  1.120000 3.610000 1.130000 ;
      RECT 3.280000  1.300000 3.610000 1.450000 ;
      RECT 3.280000  1.450000 3.450000 1.970000 ;
      RECT 3.405000  0.360000 4.545000 0.610000 ;
      RECT 3.460000  2.405000 3.790000 2.735000 ;
      RECT 3.620000  1.620000 4.725000 1.790000 ;
      RECT 3.620000  1.790000 3.790000 2.405000 ;
      RECT 3.875000  0.950000 4.205000 1.450000 ;
      RECT 3.960000  2.050000 4.290000 2.905000 ;
      RECT 4.375000  0.610000 4.545000 1.220000 ;
      RECT 4.375000  1.220000 5.120000 1.550000 ;
      RECT 4.375000  1.550000 4.725000 1.620000 ;
      RECT 4.530000  1.960000 5.945000 2.290000 ;
      RECT 4.680000  2.520000 5.445000 3.245000 ;
      RECT 4.730000  0.085000 4.980000 1.030000 ;
      RECT 5.210000  0.350000 5.460000 1.050000 ;
      RECT 5.290000  1.050000 5.460000 1.720000 ;
      RECT 5.290000  1.720000 6.520000 1.890000 ;
      RECT 5.290000  1.890000 5.945000 1.960000 ;
      RECT 5.615000  2.290000 5.945000 2.850000 ;
      RECT 6.030000  0.085000 6.360000 1.010000 ;
      RECT 6.115000  2.060000 6.445000 3.245000 ;
      RECT 6.350000  1.220000 6.775000 1.550000 ;
      RECT 6.350000  1.550000 6.520000 1.720000 ;
      RECT 7.285000  0.540000 7.560000 1.300000 ;
      RECT 7.285000  1.300000 8.190000 1.630000 ;
      RECT 7.285000  1.630000 7.535000 2.780000 ;
      RECT 7.745000  0.085000 8.075000 1.130000 ;
      RECT 7.745000  1.820000 8.010000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
  END
END sky130_fd_sc_hs__dlrbn_1
MACRO sky130_fd_sc_hs__dlrbn_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.260000 0.805000 1.930000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.260000 1.820000 6.590000 2.070000 ;
        RECT 6.285000 0.770000 6.615000 1.130000 ;
        RECT 6.285000 1.130000 6.455000 1.820000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.572800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.205000 0.880000 8.575000 1.050000 ;
        RECT 8.225000 1.820000 8.575000 2.980000 ;
        RECT 8.405000 1.050000 8.575000 1.820000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.570000 1.180000 6.115000 1.550000 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.975000 1.260000 1.285000 1.930000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.120000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.120000 0.085000 ;
      RECT 0.000000  3.245000 9.120000 3.415000 ;
      RECT 0.085000  0.540000 0.445000 1.090000 ;
      RECT 0.085000  1.090000 0.255000 2.100000 ;
      RECT 0.085000  2.100000 1.155000 2.270000 ;
      RECT 0.085000  2.270000 0.445000 2.980000 ;
      RECT 0.625000  0.085000 0.955000 1.090000 ;
      RECT 0.645000  2.440000 0.815000 3.245000 ;
      RECT 0.985000  2.270000 1.155000 2.650000 ;
      RECT 0.985000  2.650000 1.965000 2.820000 ;
      RECT 1.125000  0.350000 1.625000 1.090000 ;
      RECT 1.325000  2.100000 1.625000 2.140000 ;
      RECT 1.325000  2.140000 2.475000 2.310000 ;
      RECT 1.325000  2.310000 1.625000 2.480000 ;
      RECT 1.455000  1.090000 1.625000 2.100000 ;
      RECT 1.795000  0.350000 2.125000 0.780000 ;
      RECT 1.795000  0.780000 3.885000 0.950000 ;
      RECT 1.795000  0.950000 2.125000 0.960000 ;
      RECT 1.795000  0.960000 1.965000 1.720000 ;
      RECT 1.795000  1.720000 2.135000 1.970000 ;
      RECT 1.795000  2.480000 2.830000 2.650000 ;
      RECT 2.135000  1.130000 3.530000 1.300000 ;
      RECT 2.135000  1.300000 2.475000 1.550000 ;
      RECT 2.295000  0.085000 2.835000 0.600000 ;
      RECT 2.305000  1.550000 2.475000 2.140000 ;
      RECT 2.425000  2.820000 2.755000 3.245000 ;
      RECT 2.660000  1.470000 2.985000 1.800000 ;
      RECT 2.660000  1.800000 2.830000 2.480000 ;
      RECT 3.010000  1.970000 3.325000 2.140000 ;
      RECT 3.010000  2.140000 3.180000 2.905000 ;
      RECT 3.010000  2.905000 4.165000 3.075000 ;
      RECT 3.155000  1.120000 3.530000 1.130000 ;
      RECT 3.155000  1.300000 3.530000 1.450000 ;
      RECT 3.155000  1.450000 3.325000 1.970000 ;
      RECT 3.325000  0.360000 4.225000 0.610000 ;
      RECT 3.350000  2.405000 3.665000 2.735000 ;
      RECT 3.495000  1.710000 5.060000 1.880000 ;
      RECT 3.495000  1.880000 3.665000 2.405000 ;
      RECT 3.715000  0.950000 3.885000 1.225000 ;
      RECT 3.715000  1.225000 4.130000 1.540000 ;
      RECT 3.835000  2.050000 4.165000 2.905000 ;
      RECT 4.055000  0.610000 4.225000 0.885000 ;
      RECT 4.055000  0.885000 4.470000 1.055000 ;
      RECT 4.300000  1.055000 4.470000 1.710000 ;
      RECT 4.375000  2.050000 5.640000 2.240000 ;
      RECT 4.375000  2.240000 6.955000 2.350000 ;
      RECT 4.395000  0.085000 4.645000 0.715000 ;
      RECT 4.525000  2.650000 5.140000 3.245000 ;
      RECT 4.735000  1.350000 5.060000 1.710000 ;
      RECT 4.875000  0.350000 5.400000 1.130000 ;
      RECT 5.230000  1.130000 5.400000 1.820000 ;
      RECT 5.230000  1.820000 5.640000 2.050000 ;
      RECT 5.310000  2.350000 6.955000 2.410000 ;
      RECT 5.310000  2.410000 5.640000 2.980000 ;
      RECT 5.695000  0.085000 6.025000 1.010000 ;
      RECT 5.810000  2.580000 6.140000 3.245000 ;
      RECT 6.625000  1.320000 6.955000 1.650000 ;
      RECT 6.710000  2.580000 7.040000 3.245000 ;
      RECT 6.785000  0.085000 7.045000 1.050000 ;
      RECT 6.785000  1.650000 6.955000 2.240000 ;
      RECT 7.215000  0.350000 7.545000 1.220000 ;
      RECT 7.215000  1.220000 8.230000 1.550000 ;
      RECT 7.215000  1.550000 7.545000 2.860000 ;
      RECT 7.775000  0.085000 8.035000 1.050000 ;
      RECT 7.775000  1.820000 8.025000 3.245000 ;
      RECT 8.745000  0.085000 9.005000 1.130000 ;
      RECT 8.755000  1.820000 9.005000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
  END
END sky130_fd_sc_hs__dlrbn_2
MACRO sky130_fd_sc_hs__dlrbp_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.435000 1.450000 0.805000 1.780000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.130000 0.350000 6.460000 1.010000 ;
        RECT 6.130000 1.010000 6.670000 1.180000 ;
        RECT 6.200000 2.060000 6.670000 2.980000 ;
        RECT 6.500000 1.180000 6.670000 2.060000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.604200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.710000 0.350000 8.055000 1.040000 ;
        RECT 7.715000 1.820000 8.055000 2.980000 ;
        RECT 7.885000 1.040000 8.055000 1.820000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.425000 1.180000 5.795000 1.550000 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.975000 1.450000 1.305000 1.780000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.095000  0.690000 0.445000 1.280000 ;
      RECT 0.095000  1.280000 0.265000 1.970000 ;
      RECT 0.095000  1.970000 0.445000 2.390000 ;
      RECT 0.095000  2.390000 2.675000 2.560000 ;
      RECT 0.095000  2.560000 0.445000 2.850000 ;
      RECT 0.625000  0.085000 0.955000 1.280000 ;
      RECT 0.650000  2.730000 0.980000 3.245000 ;
      RECT 1.185000  0.500000 1.645000 0.580000 ;
      RECT 1.185000  0.580000 2.990000 0.750000 ;
      RECT 1.185000  0.750000 1.645000 1.280000 ;
      RECT 1.185000  1.970000 1.645000 2.220000 ;
      RECT 1.475000  1.280000 1.645000 1.420000 ;
      RECT 1.475000  1.420000 1.875000 1.750000 ;
      RECT 1.475000  1.750000 1.645000 1.970000 ;
      RECT 1.815000  1.940000 2.215000 2.220000 ;
      RECT 1.825000  0.920000 2.215000 1.130000 ;
      RECT 1.825000  1.130000 3.395000 1.250000 ;
      RECT 2.045000  1.250000 3.395000 1.300000 ;
      RECT 2.045000  1.300000 2.215000 1.940000 ;
      RECT 2.320000  0.085000 2.650000 0.410000 ;
      RECT 2.350000  2.730000 2.685000 3.245000 ;
      RECT 2.505000  1.470000 2.835000 1.800000 ;
      RECT 2.505000  1.800000 2.675000 2.390000 ;
      RECT 2.820000  0.255000 3.905000 0.510000 ;
      RECT 2.820000  0.510000 2.990000 0.580000 ;
      RECT 2.855000  1.970000 3.175000 2.140000 ;
      RECT 2.855000  2.140000 3.025000 2.905000 ;
      RECT 2.855000  2.905000 4.015000 3.075000 ;
      RECT 3.005000  1.300000 3.395000 1.480000 ;
      RECT 3.005000  1.480000 3.175000 1.970000 ;
      RECT 3.190000  0.710000 3.750000 0.960000 ;
      RECT 3.195000  2.405000 3.515000 2.735000 ;
      RECT 3.345000  1.650000 4.915000 1.820000 ;
      RECT 3.345000  1.820000 3.515000 2.405000 ;
      RECT 3.580000  0.960000 3.750000 1.650000 ;
      RECT 3.685000  2.050000 4.015000 2.905000 ;
      RECT 4.225000  1.990000 5.580000 2.320000 ;
      RECT 4.240000  0.085000 4.570000 1.060000 ;
      RECT 4.405000  2.650000 5.080000 3.245000 ;
      RECT 4.585000  1.350000 4.915000 1.650000 ;
      RECT 4.800000  0.350000 5.255000 1.130000 ;
      RECT 5.085000  1.130000 5.255000 1.720000 ;
      RECT 5.085000  1.720000 6.330000 1.890000 ;
      RECT 5.085000  1.890000 5.580000 1.990000 ;
      RECT 5.250000  2.320000 5.580000 2.980000 ;
      RECT 5.620000  0.085000 5.950000 1.010000 ;
      RECT 5.780000  2.060000 6.030000 3.245000 ;
      RECT 6.005000  1.350000 6.330000 1.720000 ;
      RECT 6.690000  0.350000 7.020000 0.840000 ;
      RECT 6.840000  0.840000 7.020000 1.320000 ;
      RECT 6.840000  1.320000 7.715000 1.650000 ;
      RECT 6.840000  1.650000 7.010000 2.980000 ;
      RECT 7.200000  0.085000 7.530000 0.940000 ;
      RECT 7.210000  2.100000 7.540000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_hs__dlrbp_1
MACRO sky130_fd_sc_hs__dlrbp_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.450000 0.805000 1.780000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.150000 0.350000 6.480000 0.960000 ;
        RECT 6.150000 0.960000 7.075000 1.130000 ;
        RECT 6.295000 1.800000 7.075000 1.970000 ;
        RECT 6.295000 1.970000 6.465000 2.980000 ;
        RECT 6.845000 1.130000 7.075000 1.800000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.225000 1.820000 8.585000 2.980000 ;
        RECT 8.245000 0.350000 8.585000 1.130000 ;
        RECT 8.415000 1.130000 8.585000 1.820000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.435000 1.180000 5.785000 1.550000 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.975000 1.180000 1.285000 1.550000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.120000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.120000 0.085000 ;
      RECT 0.000000  3.245000 9.120000 3.415000 ;
      RECT 0.085000  0.540000 0.445000 1.130000 ;
      RECT 0.085000  1.130000 0.255000 1.950000 ;
      RECT 0.085000  1.950000 0.445000 2.360000 ;
      RECT 0.085000  2.360000 2.805000 2.530000 ;
      RECT 0.085000  2.530000 0.445000 2.820000 ;
      RECT 0.625000  0.085000 0.955000 1.010000 ;
      RECT 0.650000  2.700000 0.980000 3.245000 ;
      RECT 1.125000  0.350000 1.625000 0.580000 ;
      RECT 1.125000  0.580000 2.980000 0.750000 ;
      RECT 1.125000  0.750000 1.625000 1.010000 ;
      RECT 1.185000  1.940000 1.625000 2.190000 ;
      RECT 1.455000  1.010000 1.625000 1.340000 ;
      RECT 1.455000  1.340000 1.865000 1.670000 ;
      RECT 1.455000  1.670000 1.625000 1.940000 ;
      RECT 1.795000  0.920000 2.205000 1.130000 ;
      RECT 1.795000  1.130000 3.385000 1.170000 ;
      RECT 1.795000  1.940000 2.205000 2.190000 ;
      RECT 2.035000  1.170000 3.385000 1.300000 ;
      RECT 2.035000  1.300000 2.205000 1.940000 ;
      RECT 2.305000  0.085000 2.640000 0.410000 ;
      RECT 2.330000  2.700000 2.695000 3.245000 ;
      RECT 2.485000  1.470000 2.805000 2.360000 ;
      RECT 2.810000  0.255000 3.895000 0.510000 ;
      RECT 2.810000  0.510000 2.980000 0.580000 ;
      RECT 2.975000  1.300000 3.385000 1.480000 ;
      RECT 2.975000  1.480000 3.145000 2.905000 ;
      RECT 2.975000  2.905000 4.035000 3.075000 ;
      RECT 3.180000  0.790000 3.740000 0.960000 ;
      RECT 3.315000  1.650000 4.925000 1.820000 ;
      RECT 3.315000  1.820000 3.485000 2.735000 ;
      RECT 3.570000  0.960000 3.740000 1.650000 ;
      RECT 3.705000  2.050000 4.035000 2.905000 ;
      RECT 4.230000  0.085000 4.560000 1.060000 ;
      RECT 4.245000  1.990000 5.565000 2.320000 ;
      RECT 4.425000  2.650000 5.065000 3.245000 ;
      RECT 4.605000  1.350000 4.925000 1.650000 ;
      RECT 4.790000  0.350000 5.265000 1.130000 ;
      RECT 5.095000  1.130000 5.265000 1.720000 ;
      RECT 5.095000  1.720000 6.125000 1.890000 ;
      RECT 5.095000  1.890000 5.565000 1.990000 ;
      RECT 5.235000  2.320000 5.565000 2.980000 ;
      RECT 5.610000  0.085000 5.940000 1.010000 ;
      RECT 5.735000  2.060000 6.065000 3.245000 ;
      RECT 5.955000  1.300000 6.650000 1.630000 ;
      RECT 5.955000  1.630000 6.125000 1.720000 ;
      RECT 6.650000  0.085000 6.980000 0.790000 ;
      RECT 6.665000  2.140000 6.995000 3.245000 ;
      RECT 7.245000  0.450000 7.575000 1.130000 ;
      RECT 7.245000  1.130000 7.555000 1.300000 ;
      RECT 7.245000  1.300000 8.245000 1.630000 ;
      RECT 7.245000  1.630000 7.555000 2.860000 ;
      RECT 7.725000  1.820000 8.055000 3.245000 ;
      RECT 7.745000  0.085000 8.075000 1.130000 ;
      RECT 8.755000  0.085000 9.005000 1.130000 ;
      RECT 8.755000  1.820000 9.005000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
  END
END sky130_fd_sc_hs__dlrbp_2
MACRO sky130_fd_sc_hs__dlrtn_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.435000 1.450000 0.835000 1.780000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.600500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.730000 0.350000 7.115000 1.130000 ;
        RECT 6.755000 1.820000 7.115000 2.980000 ;
        RECT 6.945000 1.130000 7.115000 1.820000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885000 1.180000 6.235000 1.550000 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.450000 1.335000 1.780000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.200000 0.085000 ;
      RECT 0.000000  3.245000 7.200000 3.415000 ;
      RECT 0.095000  0.580000 2.865000 0.750000 ;
      RECT 0.095000  0.750000 0.445000 1.250000 ;
      RECT 0.095000  1.250000 0.265000 1.950000 ;
      RECT 0.095000  1.950000 0.450000 2.830000 ;
      RECT 0.625000  0.085000 0.955000 0.410000 ;
      RECT 0.655000  1.950000 0.985000 3.245000 ;
      RECT 1.065000  0.920000 1.675000 1.250000 ;
      RECT 1.190000  1.950000 1.675000 2.520000 ;
      RECT 1.190000  2.520000 4.245000 2.690000 ;
      RECT 1.190000  2.690000 1.675000 2.830000 ;
      RECT 1.505000  1.250000 1.675000 1.340000 ;
      RECT 1.505000  1.340000 1.905000 1.670000 ;
      RECT 1.505000  1.670000 1.675000 1.950000 ;
      RECT 1.845000  0.920000 2.245000 1.170000 ;
      RECT 1.845000  1.840000 3.405000 2.010000 ;
      RECT 1.845000  2.010000 2.245000 2.350000 ;
      RECT 2.075000  1.170000 2.245000 1.840000 ;
      RECT 2.300000  2.860000 2.630000 3.245000 ;
      RECT 2.355000  0.085000 3.200000 0.410000 ;
      RECT 2.535000  0.750000 2.865000 1.590000 ;
      RECT 3.075000  1.190000 4.335000 1.520000 ;
      RECT 3.075000  1.520000 3.405000 1.840000 ;
      RECT 3.255000  2.180000 3.745000 2.350000 ;
      RECT 3.575000  1.690000 5.070000 1.860000 ;
      RECT 3.575000  1.860000 3.745000 2.180000 ;
      RECT 3.815000  0.350000 4.145000 0.850000 ;
      RECT 3.815000  0.850000 5.070000 1.020000 ;
      RECT 3.915000  2.030000 4.245000 2.520000 ;
      RECT 4.485000  2.030000 5.965000 2.360000 ;
      RECT 4.635000  2.530000 5.430000 3.245000 ;
      RECT 4.670000  0.085000 5.010000 0.680000 ;
      RECT 4.900000  1.020000 5.070000 1.300000 ;
      RECT 4.900000  1.300000 5.295000 1.630000 ;
      RECT 4.900000  1.630000 5.070000 1.690000 ;
      RECT 5.240000  0.350000 5.635000 1.130000 ;
      RECT 5.465000  1.130000 5.635000 1.720000 ;
      RECT 5.465000  1.720000 6.585000 1.890000 ;
      RECT 5.465000  1.890000 5.965000 2.030000 ;
      RECT 5.635000  2.360000 5.965000 2.860000 ;
      RECT 6.140000  0.085000 6.470000 1.010000 ;
      RECT 6.255000  2.060000 6.585000 3.245000 ;
      RECT 6.415000  1.320000 6.775000 1.650000 ;
      RECT 6.415000  1.650000 6.585000 1.720000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
  END
END sky130_fd_sc_hs__dlrtn_1
MACRO sky130_fd_sc_hs__dlrtn_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.435000 1.450000 0.835000 1.780000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.845000 1.820000 7.535000 2.980000 ;
        RECT 7.205000 0.350000 7.535000 1.470000 ;
        RECT 7.365000 1.470000 7.535000 1.820000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885000 1.180000 6.305000 1.550000 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.450000 1.335000 1.780000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.095000  0.580000 2.945000 0.750000 ;
      RECT 0.095000  0.750000 0.445000 1.250000 ;
      RECT 0.095000  1.250000 0.265000 1.950000 ;
      RECT 0.095000  1.950000 0.615000 2.830000 ;
      RECT 0.625000  0.085000 0.955000 0.410000 ;
      RECT 0.785000  1.950000 1.115000 3.245000 ;
      RECT 1.135000  0.920000 1.675000 1.250000 ;
      RECT 1.285000  1.950000 1.675000 2.520000 ;
      RECT 1.285000  2.520000 4.325000 2.690000 ;
      RECT 1.285000  2.690000 1.675000 2.830000 ;
      RECT 1.505000  1.250000 1.675000 1.340000 ;
      RECT 1.505000  1.340000 1.905000 1.670000 ;
      RECT 1.505000  1.670000 1.675000 1.950000 ;
      RECT 1.845000  0.920000 2.245000 1.170000 ;
      RECT 1.845000  1.840000 3.485000 2.010000 ;
      RECT 1.845000  2.010000 2.245000 2.350000 ;
      RECT 2.075000  1.170000 2.245000 1.840000 ;
      RECT 2.380000  0.085000 3.280000 0.410000 ;
      RECT 2.380000  2.860000 2.710000 3.245000 ;
      RECT 2.615000  0.750000 2.945000 1.590000 ;
      RECT 3.155000  1.190000 4.415000 1.520000 ;
      RECT 3.155000  1.520000 3.485000 1.840000 ;
      RECT 3.335000  2.180000 3.825000 2.350000 ;
      RECT 3.655000  1.690000 5.375000 1.860000 ;
      RECT 3.655000  1.860000 3.825000 2.180000 ;
      RECT 3.895000  0.350000 4.225000 0.850000 ;
      RECT 3.895000  0.850000 5.140000 1.020000 ;
      RECT 3.995000  2.030000 4.325000 2.520000 ;
      RECT 4.565000  2.030000 6.045000 2.360000 ;
      RECT 4.715000  2.630000 5.545000 3.245000 ;
      RECT 4.750000  0.085000 5.080000 0.680000 ;
      RECT 4.970000  1.020000 5.140000 1.350000 ;
      RECT 4.970000  1.350000 5.375000 1.690000 ;
      RECT 5.310000  0.350000 5.715000 1.130000 ;
      RECT 5.545000  1.130000 5.715000 1.720000 ;
      RECT 5.545000  1.720000 6.675000 1.890000 ;
      RECT 5.545000  1.890000 6.045000 2.030000 ;
      RECT 5.715000  2.360000 6.045000 2.980000 ;
      RECT 6.130000  0.085000 7.035000 1.010000 ;
      RECT 6.320000  2.060000 6.650000 3.245000 ;
      RECT 6.505000  1.320000 6.845000 1.650000 ;
      RECT 6.505000  1.650000 6.675000 1.720000 ;
      RECT 7.705000  0.085000 8.035000 1.130000 ;
      RECT 7.705000  1.820000 8.045000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_hs__dlrtn_2
MACRO sky130_fd_sc_hs__dlrtn_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.600000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.450000 0.805000 1.780000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.198400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.545000 1.960000 9.475000 1.970000 ;
        RECT 7.545000 1.970000 8.875000 2.130000 ;
        RECT 7.545000 2.130000 7.875000 2.980000 ;
        RECT 7.935000 0.360000 8.125000 0.960000 ;
        RECT 7.935000 0.960000 9.475000 1.130000 ;
        RECT 8.545000 1.800000 9.475000 1.960000 ;
        RECT 8.545000 2.130000 8.875000 2.980000 ;
        RECT 8.795000 0.360000 8.985000 0.800000 ;
        RECT 8.795000 0.800000 9.475000 0.960000 ;
        RECT 9.245000 1.130000 9.475000 1.800000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.444000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.320000 1.120000 7.555000 1.450000 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.975000 1.450000 1.290000 1.780000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.600000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.600000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.600000 0.085000 ;
      RECT 0.000000  3.245000 9.600000 3.415000 ;
      RECT 0.085000  0.660000 2.820000 0.830000 ;
      RECT 0.085000  0.830000 0.445000 1.250000 ;
      RECT 0.085000  1.250000 0.255000 1.950000 ;
      RECT 0.085000  1.950000 0.475000 2.830000 ;
      RECT 0.625000  0.085000 0.955000 0.490000 ;
      RECT 0.645000  1.950000 0.975000 3.245000 ;
      RECT 1.135000  1.000000 1.630000 1.250000 ;
      RECT 1.145000  1.950000 1.630000 2.600000 ;
      RECT 1.145000  2.600000 4.200000 2.770000 ;
      RECT 1.145000  2.770000 1.630000 2.830000 ;
      RECT 1.460000  1.250000 1.630000 1.420000 ;
      RECT 1.460000  1.420000 1.865000 1.750000 ;
      RECT 1.460000  1.750000 1.630000 1.950000 ;
      RECT 1.800000  1.000000 2.205000 1.250000 ;
      RECT 1.800000  1.920000 3.360000 2.090000 ;
      RECT 1.800000  2.090000 2.205000 2.430000 ;
      RECT 2.035000  1.250000 2.205000 1.920000 ;
      RECT 2.255000  2.940000 2.585000 3.245000 ;
      RECT 2.310000  0.085000 3.125000 0.490000 ;
      RECT 2.490000  0.830000 2.820000 1.670000 ;
      RECT 3.030000  1.190000 4.260000 1.520000 ;
      RECT 3.030000  1.520000 3.360000 1.920000 ;
      RECT 3.180000  2.260000 3.700000 2.430000 ;
      RECT 3.530000  1.690000 5.220000 1.860000 ;
      RECT 3.530000  1.860000 3.700000 2.260000 ;
      RECT 3.740000  0.400000 4.070000 0.850000 ;
      RECT 3.740000  0.850000 4.985000 1.020000 ;
      RECT 3.870000  2.030000 4.200000 2.600000 ;
      RECT 4.440000  2.030000 5.820000 2.360000 ;
      RECT 4.590000  2.630000 5.320000 3.245000 ;
      RECT 4.595000  0.085000 4.925000 0.680000 ;
      RECT 4.815000  1.020000 4.985000 1.120000 ;
      RECT 4.815000  1.120000 5.220000 1.690000 ;
      RECT 5.155000  0.255000 6.265000 0.425000 ;
      RECT 5.155000  0.425000 5.485000 0.950000 ;
      RECT 5.490000  1.620000 9.075000 1.630000 ;
      RECT 5.490000  1.630000 7.895000 1.790000 ;
      RECT 5.490000  1.790000 5.820000 2.030000 ;
      RECT 5.490000  2.360000 5.820000 2.960000 ;
      RECT 5.665000  0.595000 5.835000 1.620000 ;
      RECT 5.990000  2.080000 6.320000 3.245000 ;
      RECT 6.015000  0.425000 6.265000 0.770000 ;
      RECT 6.015000  0.770000 7.205000 0.950000 ;
      RECT 6.445000  0.085000 6.775000 0.600000 ;
      RECT 6.490000  1.790000 6.820000 2.960000 ;
      RECT 6.945000  0.355000 7.205000 0.770000 ;
      RECT 7.045000  2.080000 7.375000 3.245000 ;
      RECT 7.435000  0.085000 7.765000 0.950000 ;
      RECT 7.725000  1.300000 9.075000 1.620000 ;
      RECT 8.045000  2.300000 8.375000 3.245000 ;
      RECT 8.295000  0.085000 8.625000 0.790000 ;
      RECT 9.045000  2.140000 9.375000 3.245000 ;
      RECT 9.155000  0.085000 9.485000 0.630000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
  END
END sky130_fd_sc_hs__dlrtn_4
MACRO sky130_fd_sc_hs__dlrtp_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.300000 0.375000 1.780000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.100000 0.350000 6.635000 0.840000 ;
        RECT 6.275000 1.820000 6.635000 2.980000 ;
        RECT 6.465000 0.840000 6.635000 1.820000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.435000 1.350000 5.765000 1.780000 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.930000 1.450000 1.285000 1.780000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.720000 0.085000 ;
      RECT 0.000000  3.245000 6.720000 3.415000 ;
      RECT 0.115000  2.100000 0.715000 2.390000 ;
      RECT 0.115000  2.390000 2.695000 2.560000 ;
      RECT 0.115000  2.560000 0.445000 2.980000 ;
      RECT 0.220000  0.540000 0.715000 1.130000 ;
      RECT 0.545000  1.130000 0.715000 2.100000 ;
      RECT 0.615000  2.730000 0.945000 3.245000 ;
      RECT 0.885000  0.085000 1.055000 1.130000 ;
      RECT 1.150000  1.970000 1.625000 2.220000 ;
      RECT 1.235000  0.350000 1.625000 0.770000 ;
      RECT 1.235000  0.770000 3.020000 0.940000 ;
      RECT 1.235000  0.940000 1.625000 1.130000 ;
      RECT 1.455000  1.130000 1.625000 1.450000 ;
      RECT 1.455000  1.450000 1.830000 1.780000 ;
      RECT 1.455000  1.780000 1.625000 1.970000 ;
      RECT 1.795000  1.110000 3.325000 1.280000 ;
      RECT 1.795000  2.020000 2.170000 2.220000 ;
      RECT 2.000000  1.280000 2.170000 2.020000 ;
      RECT 2.295000  0.085000 2.680000 0.600000 ;
      RECT 2.330000  2.730000 2.705000 3.245000 ;
      RECT 2.525000  1.470000 2.855000 1.800000 ;
      RECT 2.525000  1.800000 2.695000 2.390000 ;
      RECT 2.850000  0.255000 4.005000 0.425000 ;
      RECT 2.850000  0.425000 3.020000 0.770000 ;
      RECT 2.905000  1.970000 3.195000 2.140000 ;
      RECT 2.905000  2.140000 3.075000 2.905000 ;
      RECT 2.905000  2.905000 4.045000 3.075000 ;
      RECT 3.025000  1.280000 3.325000 1.450000 ;
      RECT 3.025000  1.450000 3.195000 1.970000 ;
      RECT 3.190000  0.595000 3.665000 0.925000 ;
      RECT 3.245000  2.405000 3.535000 2.735000 ;
      RECT 3.365000  1.725000 4.925000 1.895000 ;
      RECT 3.365000  1.895000 3.535000 2.405000 ;
      RECT 3.495000  0.925000 3.665000 1.725000 ;
      RECT 3.715000  2.065000 4.045000 2.905000 ;
      RECT 3.835000  0.425000 4.005000 1.225000 ;
      RECT 3.835000  1.225000 4.095000 1.555000 ;
      RECT 4.210000  0.085000 4.540000 0.810000 ;
      RECT 4.305000  2.065000 5.575000 2.380000 ;
      RECT 4.435000  2.650000 5.075000 3.245000 ;
      RECT 4.665000  1.470000 4.925000 1.725000 ;
      RECT 4.770000  0.350000 5.100000 1.010000 ;
      RECT 4.770000  1.010000 6.295000 1.180000 ;
      RECT 5.095000  1.180000 5.265000 1.950000 ;
      RECT 5.095000  1.950000 5.575000 2.065000 ;
      RECT 5.245000  2.380000 5.575000 2.980000 ;
      RECT 5.590000  0.085000 5.920000 0.840000 ;
      RECT 5.745000  1.950000 6.075000 3.245000 ;
      RECT 5.975000  1.180000 6.295000 1.550000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
  END
END sky130_fd_sc_hs__dlrtp_1
MACRO sky130_fd_sc_hs__dlrtp_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.450000 0.515000 1.780000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.567400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.255000 0.350000 6.585000 0.960000 ;
        RECT 6.255000 0.960000 7.075000 1.130000 ;
        RECT 6.255000 2.060000 6.585000 2.980000 ;
        RECT 6.415000 1.800000 7.075000 1.970000 ;
        RECT 6.415000 1.970000 6.585000 2.060000 ;
        RECT 6.845000 1.130000 7.075000 1.800000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.435000 1.180000 5.840000 1.550000 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.025000 1.180000 1.285000 1.550000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.200000 0.085000 ;
      RECT 0.000000  3.245000 7.200000 3.415000 ;
      RECT 0.115000  1.950000 0.855000 2.440000 ;
      RECT 0.115000  2.440000 2.680000 2.610000 ;
      RECT 0.115000  2.610000 0.445000 2.820000 ;
      RECT 0.140000  0.540000 0.470000 1.110000 ;
      RECT 0.140000  1.110000 0.855000 1.280000 ;
      RECT 0.650000  0.085000 0.980000 0.940000 ;
      RECT 0.650000  2.780000 0.980000 3.245000 ;
      RECT 0.685000  1.280000 0.855000 1.950000 ;
      RECT 1.150000  0.350000 1.625000 0.580000 ;
      RECT 1.150000  0.580000 2.975000 0.750000 ;
      RECT 1.150000  0.750000 1.625000 1.010000 ;
      RECT 1.185000  1.940000 1.625000 2.270000 ;
      RECT 1.455000  1.010000 1.625000 1.420000 ;
      RECT 1.455000  1.420000 1.890000 1.750000 ;
      RECT 1.455000  1.750000 1.625000 1.940000 ;
      RECT 1.795000  0.920000 2.230000 1.080000 ;
      RECT 1.795000  1.080000 3.315000 1.250000 ;
      RECT 1.825000  1.940000 2.230000 2.270000 ;
      RECT 2.060000  1.250000 2.230000 1.940000 ;
      RECT 2.280000  2.780000 2.610000 3.245000 ;
      RECT 2.305000  0.085000 2.635000 0.410000 ;
      RECT 2.510000  1.440000 2.840000 1.770000 ;
      RECT 2.510000  1.770000 2.680000 2.440000 ;
      RECT 2.805000  0.255000 4.090000 0.425000 ;
      RECT 2.805000  0.425000 2.975000 0.580000 ;
      RECT 2.890000  1.940000 3.220000 2.110000 ;
      RECT 2.890000  2.110000 3.060000 2.905000 ;
      RECT 2.890000  2.905000 4.060000 3.075000 ;
      RECT 3.050000  1.250000 3.315000 1.450000 ;
      RECT 3.050000  1.450000 3.220000 1.940000 ;
      RECT 3.205000  0.595000 3.715000 0.845000 ;
      RECT 3.230000  2.405000 3.560000 2.735000 ;
      RECT 3.390000  1.760000 4.925000 1.930000 ;
      RECT 3.390000  1.930000 3.560000 2.405000 ;
      RECT 3.485000  0.845000 3.655000 1.760000 ;
      RECT 3.730000  2.100000 4.060000 2.905000 ;
      RECT 3.825000  1.260000 4.090000 1.590000 ;
      RECT 3.920000  0.425000 4.090000 1.260000 ;
      RECT 4.285000  0.085000 4.615000 0.845000 ;
      RECT 4.300000  2.100000 5.585000 2.380000 ;
      RECT 4.450000  2.650000 5.085000 3.245000 ;
      RECT 4.660000  1.350000 4.925000 1.760000 ;
      RECT 4.845000  0.350000 5.265000 1.130000 ;
      RECT 5.095000  1.130000 5.265000 1.720000 ;
      RECT 5.095000  1.720000 6.220000 1.890000 ;
      RECT 5.095000  1.890000 5.585000 2.100000 ;
      RECT 5.255000  2.380000 5.585000 2.980000 ;
      RECT 5.755000  0.085000 6.085000 1.010000 ;
      RECT 5.755000  2.060000 6.085000 3.245000 ;
      RECT 6.050000  1.300000 6.675000 1.630000 ;
      RECT 6.050000  1.630000 6.220000 1.720000 ;
      RECT 6.755000  0.085000 7.085000 0.790000 ;
      RECT 6.755000  2.140000 7.085000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
  END
END sky130_fd_sc_hs__dlrtp_2
MACRO sky130_fd_sc_hs__dlrtp_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.450000 0.515000 1.780000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.164800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.175000 1.800000 8.995000 1.970000 ;
        RECT 7.175000 1.970000 7.425000 2.980000 ;
        RECT 7.385000 0.365000 7.645000 0.880000 ;
        RECT 7.385000 0.880000 8.995000 1.130000 ;
        RECT 8.095000 1.970000 8.425000 2.980000 ;
        RECT 8.315000 0.365000 8.505000 0.880000 ;
        RECT 8.765000 1.130000 8.995000 1.800000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.444000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885000 1.120000 6.595000 1.450000 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.025000 1.450000 1.290000 1.780000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.120000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.120000 0.085000 ;
      RECT 0.000000  3.245000 9.120000 3.415000 ;
      RECT 0.115000  0.610000 0.445000 1.110000 ;
      RECT 0.115000  1.110000 0.855000 1.280000 ;
      RECT 0.115000  1.950000 0.855000 2.370000 ;
      RECT 0.115000  2.370000 2.665000 2.540000 ;
      RECT 0.115000  2.540000 0.445000 2.830000 ;
      RECT 0.650000  2.710000 0.980000 3.245000 ;
      RECT 0.680000  0.085000 1.010000 0.940000 ;
      RECT 0.685000  1.280000 0.855000 1.950000 ;
      RECT 1.185000  1.950000 1.630000 2.200000 ;
      RECT 1.240000  0.420000 1.630000 0.770000 ;
      RECT 1.240000  0.770000 3.005000 0.940000 ;
      RECT 1.240000  0.940000 1.630000 1.200000 ;
      RECT 1.460000  1.200000 1.630000 1.450000 ;
      RECT 1.460000  1.450000 1.900000 1.780000 ;
      RECT 1.460000  1.780000 1.630000 1.950000 ;
      RECT 1.800000  1.110000 3.340000 1.280000 ;
      RECT 1.800000  2.020000 2.240000 2.200000 ;
      RECT 2.070000  1.280000 2.240000 2.020000 ;
      RECT 2.335000  0.085000 2.665000 0.600000 ;
      RECT 2.335000  2.710000 2.665000 3.245000 ;
      RECT 2.495000  1.470000 2.785000 1.800000 ;
      RECT 2.495000  1.800000 2.665000 2.370000 ;
      RECT 2.835000  0.255000 4.020000 0.425000 ;
      RECT 2.835000  0.425000 3.005000 0.770000 ;
      RECT 2.845000  1.970000 3.125000 2.140000 ;
      RECT 2.845000  2.140000 3.015000 2.905000 ;
      RECT 2.845000  2.905000 3.985000 3.075000 ;
      RECT 2.955000  1.280000 3.340000 1.450000 ;
      RECT 2.955000  1.450000 3.125000 1.970000 ;
      RECT 3.175000  0.595000 3.680000 0.925000 ;
      RECT 3.185000  2.405000 3.465000 2.735000 ;
      RECT 3.295000  1.725000 5.020000 1.895000 ;
      RECT 3.295000  1.895000 3.465000 2.405000 ;
      RECT 3.510000  0.925000 3.680000 1.725000 ;
      RECT 3.655000  2.065000 3.985000 2.905000 ;
      RECT 3.850000  0.425000 4.020000 1.225000 ;
      RECT 3.850000  1.225000 4.150000 1.555000 ;
      RECT 4.190000  0.085000 4.440000 0.810000 ;
      RECT 4.195000  2.065000 5.440000 2.480000 ;
      RECT 4.345000  2.650000 4.905000 3.245000 ;
      RECT 4.670000  0.280000 5.785000 0.450000 ;
      RECT 4.670000  0.450000 5.000000 1.030000 ;
      RECT 4.720000  1.350000 5.020000 1.725000 ;
      RECT 5.110000  2.480000 5.440000 2.700000 ;
      RECT 5.180000  0.620000 5.360000 0.950000 ;
      RECT 5.190000  0.950000 5.360000 1.620000 ;
      RECT 5.190000  1.620000 8.595000 1.630000 ;
      RECT 5.190000  1.630000 6.935000 1.790000 ;
      RECT 5.190000  1.790000 5.440000 2.065000 ;
      RECT 5.535000  0.450000 5.785000 0.770000 ;
      RECT 5.535000  0.770000 6.725000 0.950000 ;
      RECT 5.610000  1.960000 5.940000 3.245000 ;
      RECT 5.965000  0.085000 6.295000 0.600000 ;
      RECT 6.110000  1.790000 6.440000 2.700000 ;
      RECT 6.465000  0.345000 6.725000 0.770000 ;
      RECT 6.645000  1.960000 6.975000 3.245000 ;
      RECT 6.765000  1.300000 8.595000 1.620000 ;
      RECT 6.955000  0.085000 7.215000 1.130000 ;
      RECT 7.595000  2.140000 7.925000 3.245000 ;
      RECT 7.815000  0.085000 8.145000 0.710000 ;
      RECT 8.595000  2.140000 8.925000 3.245000 ;
      RECT 8.675000  0.085000 9.005000 0.710000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
  END
END sky130_fd_sc_hs__dlrtp_4
MACRO sky130_fd_sc_hs__dlxbn_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.435000 1.260000 0.835000 1.930000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.524500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.765000 1.820000 6.130000 2.980000 ;
        RECT 5.790000 0.350000 6.130000 1.100000 ;
        RECT 5.960000 1.100000 6.130000 1.820000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.537600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.715000 0.350000 8.050000 2.980000 ;
    END
  END Q_N
  PIN GATE_N
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.690000 1.335000 2.150000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.095000  0.580000 2.865000 0.750000 ;
      RECT 0.095000  0.750000 0.445000 1.090000 ;
      RECT 0.095000  1.090000 0.265000 2.100000 ;
      RECT 0.095000  2.100000 0.545000 2.980000 ;
      RECT 0.625000  0.085000 0.955000 0.410000 ;
      RECT 0.735000  2.320000 1.065000 3.245000 ;
      RECT 1.135000  0.920000 1.465000 1.260000 ;
      RECT 1.135000  1.260000 1.905000 1.520000 ;
      RECT 1.235000  2.320000 1.675000 2.390000 ;
      RECT 1.235000  2.390000 4.145000 2.560000 ;
      RECT 1.235000  2.560000 1.565000 2.980000 ;
      RECT 1.505000  1.520000 1.675000 2.320000 ;
      RECT 1.695000  0.920000 2.245000 1.090000 ;
      RECT 1.845000  1.880000 2.910000 2.220000 ;
      RECT 2.075000  1.090000 2.245000 1.710000 ;
      RECT 2.075000  1.710000 3.340000 1.880000 ;
      RECT 2.340000  0.085000 2.675000 0.410000 ;
      RECT 2.380000  2.730000 2.710000 3.245000 ;
      RECT 2.535000  0.750000 2.865000 1.510000 ;
      RECT 3.035000  0.255000 4.260000 0.505000 ;
      RECT 3.035000  0.505000 3.205000 1.470000 ;
      RECT 3.035000  1.470000 3.340000 1.710000 ;
      RECT 3.260000  2.050000 3.805000 2.220000 ;
      RECT 3.375000  0.725000 4.135000 1.055000 ;
      RECT 3.510000  1.055000 4.135000 1.130000 ;
      RECT 3.510000  1.130000 5.220000 1.300000 ;
      RECT 3.510000  1.300000 3.680000 2.050000 ;
      RECT 3.850000  1.470000 4.145000 1.800000 ;
      RECT 3.975000  1.800000 4.145000 2.390000 ;
      RECT 4.315000  1.470000 4.645000 1.720000 ;
      RECT 4.315000  1.720000 5.560000 1.890000 ;
      RECT 4.480000  2.060000 5.020000 3.245000 ;
      RECT 4.705000  0.085000 5.035000 0.960000 ;
      RECT 4.890000  1.300000 5.220000 1.550000 ;
      RECT 5.205000  0.350000 5.560000 0.960000 ;
      RECT 5.220000  1.890000 5.560000 2.900000 ;
      RECT 5.390000  0.960000 5.560000 1.270000 ;
      RECT 5.390000  1.270000 5.790000 1.600000 ;
      RECT 5.390000  1.600000 5.560000 1.720000 ;
      RECT 6.300000  0.085000 6.550000 1.130000 ;
      RECT 6.300000  2.100000 6.550000 3.245000 ;
      RECT 6.720000  0.540000 7.060000 1.300000 ;
      RECT 6.720000  1.300000 7.500000 1.630000 ;
      RECT 6.720000  1.630000 7.065000 2.980000 ;
      RECT 7.265000  1.820000 7.515000 3.245000 ;
      RECT 7.290000  0.085000 7.540000 1.130000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_hs__dlxbn_1
MACRO sky130_fd_sc_hs__dlxbn_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.440000 1.450000 0.815000 1.780000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885000 0.850000 6.505000 1.130000 ;
        RECT 5.885000 1.130000 6.115000 1.800000 ;
        RECT 5.885000 1.800000 6.590000 2.070000 ;
        RECT 6.245000 0.355000 6.505000 0.850000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.225000 1.820000 8.555000 2.980000 ;
        RECT 8.245000 0.350000 8.495000 1.130000 ;
        RECT 8.325000 1.130000 8.495000 1.820000 ;
    END
  END Q_N
  PIN GATE_N
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.985000 1.695000 1.315000 2.150000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.120000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.120000 0.085000 ;
      RECT 0.000000  3.245000 9.120000 3.415000 ;
      RECT 0.100000  0.580000 2.845000 0.750000 ;
      RECT 0.100000  0.750000 0.445000 1.250000 ;
      RECT 0.100000  1.250000 0.270000 2.100000 ;
      RECT 0.100000  2.100000 0.445000 2.980000 ;
      RECT 0.625000  0.085000 0.955000 0.410000 ;
      RECT 0.650000  2.320000 0.980000 3.245000 ;
      RECT 1.135000  0.920000 1.465000 1.260000 ;
      RECT 1.135000  1.260000 1.885000 1.525000 ;
      RECT 1.150000  2.320000 1.655000 2.390000 ;
      RECT 1.150000  2.390000 4.275000 2.560000 ;
      RECT 1.150000  2.560000 1.485000 2.980000 ;
      RECT 1.485000  1.525000 1.655000 2.320000 ;
      RECT 1.695000  0.920000 2.225000 1.090000 ;
      RECT 1.825000  1.710000 3.385000 1.880000 ;
      RECT 1.825000  1.880000 2.155000 2.220000 ;
      RECT 2.055000  1.090000 2.225000 1.710000 ;
      RECT 2.285000  0.085000 2.640000 0.410000 ;
      RECT 2.360000  2.730000 2.690000 3.245000 ;
      RECT 2.515000  0.750000 2.845000 1.540000 ;
      RECT 3.015000  0.255000 4.265000 0.505000 ;
      RECT 3.015000  0.505000 3.185000 1.470000 ;
      RECT 3.015000  1.470000 3.385000 1.710000 ;
      RECT 3.230000  2.050000 3.935000 2.220000 ;
      RECT 3.355000  0.725000 4.070000 1.015000 ;
      RECT 3.355000  1.015000 5.315000 1.055000 ;
      RECT 3.555000  1.055000 5.315000 1.185000 ;
      RECT 3.555000  1.185000 3.725000 2.050000 ;
      RECT 3.895000  1.420000 4.275000 1.750000 ;
      RECT 4.105000  1.750000 4.275000 2.390000 ;
      RECT 4.445000  1.355000 4.775000 1.720000 ;
      RECT 4.445000  1.720000 5.655000 1.890000 ;
      RECT 4.630000  0.085000 5.015000 0.845000 ;
      RECT 4.670000  2.070000 5.080000 3.245000 ;
      RECT 4.985000  1.185000 5.315000 1.550000 ;
      RECT 5.185000  0.350000 5.655000 0.845000 ;
      RECT 5.250000  1.890000 5.655000 2.240000 ;
      RECT 5.250000  2.240000 6.955000 2.410000 ;
      RECT 5.250000  2.410000 5.655000 2.980000 ;
      RECT 5.485000  0.845000 5.655000 1.720000 ;
      RECT 5.825000  0.085000 6.075000 0.680000 ;
      RECT 5.890000  2.580000 6.140000 3.245000 ;
      RECT 6.285000  1.300000 6.955000 1.630000 ;
      RECT 6.675000  0.085000 7.005000 1.130000 ;
      RECT 6.710000  2.580000 7.040000 3.245000 ;
      RECT 6.785000  1.630000 6.955000 2.240000 ;
      RECT 7.185000  0.450000 7.515000 1.130000 ;
      RECT 7.215000  1.130000 7.515000 1.320000 ;
      RECT 7.215000  1.320000 8.155000 1.650000 ;
      RECT 7.215000  1.650000 7.545000 2.980000 ;
      RECT 7.745000  0.085000 8.075000 1.130000 ;
      RECT 7.775000  1.820000 8.025000 3.245000 ;
      RECT 8.675000  0.085000 9.005000 1.130000 ;
      RECT 8.755000  1.820000 9.005000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
  END
END sky130_fd_sc_hs__dlxbn_2
MACRO sky130_fd_sc_hs__dlxbp_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.435000 1.220000 0.835000 1.890000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.537600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.765000 1.820000 6.125000 2.980000 ;
        RECT 5.795000 0.370000 6.125000 1.150000 ;
        RECT 5.955000 1.150000 6.125000 1.820000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.535700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.715000 0.350000 8.050000 2.980000 ;
    END
  END Q_N
  PIN GATE
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.180000 1.335000 1.550000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.095000  0.540000 0.450000 1.050000 ;
      RECT 0.095000  1.050000 0.265000 2.060000 ;
      RECT 0.095000  2.060000 0.440000 2.545000 ;
      RECT 0.095000  2.545000 1.760000 2.715000 ;
      RECT 0.095000  2.715000 0.440000 2.925000 ;
      RECT 0.630000  0.085000 0.960000 1.010000 ;
      RECT 0.640000  2.885000 0.970000 3.245000 ;
      RECT 1.130000  0.350000 1.675000 0.580000 ;
      RECT 1.130000  0.580000 3.080000 0.750000 ;
      RECT 1.130000  0.750000 1.675000 1.010000 ;
      RECT 1.170000  1.720000 2.330000 1.890000 ;
      RECT 1.170000  1.890000 1.420000 2.375000 ;
      RECT 1.505000  1.010000 1.675000 1.470000 ;
      RECT 1.505000  1.470000 2.330000 1.720000 ;
      RECT 1.590000  2.060000 2.875000 2.230000 ;
      RECT 1.590000  2.230000 1.760000 2.545000 ;
      RECT 1.845000  0.920000 2.175000 1.020000 ;
      RECT 1.845000  1.020000 3.515000 1.190000 ;
      RECT 1.930000  2.400000 2.180000 2.440000 ;
      RECT 1.930000  2.440000 4.100000 2.610000 ;
      RECT 1.930000  2.610000 2.180000 2.820000 ;
      RECT 2.355000  0.085000 2.740000 0.410000 ;
      RECT 2.380000  2.780000 2.710000 3.245000 ;
      RECT 2.545000  1.470000 2.875000 2.060000 ;
      RECT 2.910000  0.255000 4.075000 0.510000 ;
      RECT 2.910000  0.510000 3.080000 0.580000 ;
      RECT 3.045000  1.190000 3.515000 1.480000 ;
      RECT 3.045000  1.480000 3.215000 2.440000 ;
      RECT 3.310000  0.680000 3.950000 0.850000 ;
      RECT 3.385000  1.650000 5.035000 1.820000 ;
      RECT 3.385000  1.820000 3.555000 2.270000 ;
      RECT 3.770000  2.050000 4.100000 2.440000 ;
      RECT 3.780000  0.850000 3.950000 1.650000 ;
      RECT 4.315000  1.990000 5.535000 2.320000 ;
      RECT 4.490000  2.545000 5.035000 3.245000 ;
      RECT 4.520000  0.085000 4.850000 1.060000 ;
      RECT 4.705000  1.240000 5.035000 1.650000 ;
      RECT 5.020000  0.350000 5.375000 1.070000 ;
      RECT 5.205000  1.070000 5.375000 1.320000 ;
      RECT 5.205000  1.320000 5.775000 1.650000 ;
      RECT 5.205000  1.650000 5.535000 1.990000 ;
      RECT 5.205000  2.320000 5.535000 2.980000 ;
      RECT 6.295000  0.085000 6.545000 1.150000 ;
      RECT 6.295000  2.100000 6.545000 3.245000 ;
      RECT 6.720000  0.560000 7.055000 1.320000 ;
      RECT 6.720000  1.320000 7.320000 1.650000 ;
      RECT 6.720000  1.650000 7.050000 2.980000 ;
      RECT 7.270000  1.820000 7.520000 3.245000 ;
      RECT 7.285000  0.085000 7.535000 1.130000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_hs__dlxbp_1
MACRO sky130_fd_sc_hs__dlxtn_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.435000 1.565000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.545000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.270000 0.350000 6.605000 2.980000 ;
    END
  END Q
  PIN GATE_N
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.945000 1.500000 1.315000 1.830000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.720000 0.085000 ;
      RECT 0.000000  3.245000 6.720000 3.415000 ;
      RECT 0.115000  0.555000 0.445000 0.660000 ;
      RECT 0.115000  0.660000 1.315000 0.830000 ;
      RECT 0.115000  0.830000 0.775000 1.010000 ;
      RECT 0.120000  1.735000 0.775000 1.905000 ;
      RECT 0.120000  1.905000 0.450000 2.955000 ;
      RECT 0.605000  1.010000 0.775000 1.735000 ;
      RECT 0.620000  2.075000 0.950000 3.245000 ;
      RECT 0.625000  0.085000 0.955000 0.490000 ;
      RECT 1.135000  1.000000 1.885000 1.330000 ;
      RECT 1.145000  0.255000 2.645000 0.425000 ;
      RECT 1.145000  0.425000 1.315000 0.660000 ;
      RECT 1.155000  2.075000 1.655000 2.440000 ;
      RECT 1.155000  2.440000 3.045000 2.610000 ;
      RECT 1.155000  2.610000 1.655000 2.955000 ;
      RECT 1.485000  0.760000 1.885000 1.000000 ;
      RECT 1.485000  1.330000 1.885000 1.770000 ;
      RECT 1.485000  1.770000 1.655000 2.075000 ;
      RECT 1.825000  1.940000 2.225000 2.270000 ;
      RECT 2.055000  0.595000 2.305000 1.725000 ;
      RECT 2.055000  1.725000 3.500000 1.895000 ;
      RECT 2.055000  1.895000 2.225000 1.940000 ;
      RECT 2.360000  2.780000 2.705000 3.245000 ;
      RECT 2.475000  0.425000 2.645000 1.225000 ;
      RECT 2.475000  1.225000 2.970000 1.555000 ;
      RECT 2.815000  0.085000 3.145000 1.055000 ;
      RECT 2.875000  2.610000 3.045000 2.905000 ;
      RECT 2.875000  2.905000 4.180000 3.075000 ;
      RECT 3.180000  1.470000 3.500000 1.725000 ;
      RECT 3.315000  0.255000 4.355000 0.585000 ;
      RECT 3.315000  0.585000 3.485000 1.470000 ;
      RECT 3.330000  2.065000 3.840000 2.735000 ;
      RECT 3.655000  0.805000 4.680000 1.055000 ;
      RECT 3.670000  1.055000 3.840000 2.065000 ;
      RECT 4.010000  1.455000 4.340000 1.785000 ;
      RECT 4.010000  1.785000 4.180000 2.905000 ;
      RECT 4.350000  2.025000 5.655000 2.355000 ;
      RECT 4.470000  2.525000 5.065000 3.245000 ;
      RECT 4.510000  1.055000 4.680000 1.305000 ;
      RECT 4.510000  1.305000 5.315000 1.635000 ;
      RECT 4.850000  0.085000 5.100000 1.135000 ;
      RECT 5.265000  1.940000 5.655000 2.025000 ;
      RECT 5.265000  2.355000 5.655000 2.980000 ;
      RECT 5.280000  0.455000 5.655000 1.135000 ;
      RECT 5.485000  1.135000 5.655000 1.300000 ;
      RECT 5.485000  1.300000 5.885000 1.630000 ;
      RECT 5.485000  1.630000 5.655000 1.940000 ;
      RECT 5.825000  1.820000 6.075000 3.245000 ;
      RECT 5.840000  0.085000 6.090000 1.130000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
  END
END sky130_fd_sc_hs__dlxtn_1
MACRO sky130_fd_sc_hs__dlxtn_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.455000 1.780000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.638000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.260000 1.920000 6.635000 2.890000 ;
        RECT 6.320000 0.350000 6.585000 1.125000 ;
        RECT 6.415000 1.125000 6.585000 1.920000 ;
    END
  END Q
  PIN GATE_N
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.985000 1.450000 1.315000 1.780000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.200000 0.085000 ;
      RECT 0.000000  3.245000 7.200000 3.415000 ;
      RECT 0.115000  0.580000 1.315000 0.750000 ;
      RECT 0.115000  0.750000 0.795000 1.130000 ;
      RECT 0.265000  1.950000 0.795000 2.120000 ;
      RECT 0.265000  2.120000 0.595000 2.980000 ;
      RECT 0.625000  0.085000 0.955000 0.410000 ;
      RECT 0.625000  1.130000 0.795000 1.950000 ;
      RECT 0.765000  2.290000 1.095000 3.245000 ;
      RECT 1.135000  0.920000 1.885000 1.170000 ;
      RECT 1.145000  0.255000 2.645000 0.425000 ;
      RECT 1.145000  0.425000 1.315000 0.580000 ;
      RECT 1.265000  2.100000 1.655000 2.440000 ;
      RECT 1.265000  2.440000 3.045000 2.610000 ;
      RECT 1.265000  2.610000 1.655000 2.980000 ;
      RECT 1.485000  0.760000 1.885000 0.920000 ;
      RECT 1.485000  1.170000 1.885000 1.770000 ;
      RECT 1.485000  1.770000 1.655000 2.100000 ;
      RECT 1.825000  1.940000 3.510000 1.970000 ;
      RECT 1.825000  1.970000 2.225000 2.270000 ;
      RECT 2.055000  0.595000 2.305000 1.800000 ;
      RECT 2.055000  1.800000 3.510000 1.940000 ;
      RECT 2.360000  2.780000 2.705000 3.245000 ;
      RECT 2.475000  0.425000 2.645000 1.300000 ;
      RECT 2.475000  1.300000 2.970000 1.630000 ;
      RECT 2.815000  0.085000 3.145000 1.055000 ;
      RECT 2.875000  2.610000 3.045000 2.905000 ;
      RECT 2.875000  2.905000 4.190000 3.075000 ;
      RECT 3.180000  1.470000 3.510000 1.800000 ;
      RECT 3.315000  0.255000 4.375000 0.585000 ;
      RECT 3.315000  0.585000 3.485000 1.470000 ;
      RECT 3.330000  2.140000 3.850000 2.735000 ;
      RECT 3.655000  0.805000 4.250000 1.055000 ;
      RECT 3.680000  1.055000 3.850000 2.140000 ;
      RECT 4.020000  1.485000 4.350000 1.815000 ;
      RECT 4.020000  1.815000 4.190000 2.905000 ;
      RECT 4.080000  1.055000 4.250000 1.145000 ;
      RECT 4.080000  1.145000 5.160000 1.295000 ;
      RECT 4.080000  1.295000 5.335000 1.315000 ;
      RECT 4.360000  2.025000 5.580000 2.355000 ;
      RECT 4.360000  2.625000 5.080000 3.245000 ;
      RECT 4.820000  0.085000 5.150000 0.975000 ;
      RECT 4.990000  1.315000 5.335000 1.625000 ;
      RECT 5.250000  1.795000 5.675000 1.965000 ;
      RECT 5.250000  1.965000 5.580000 2.025000 ;
      RECT 5.250000  2.355000 5.580000 2.955000 ;
      RECT 5.330000  0.355000 5.580000 0.955000 ;
      RECT 5.330000  0.955000 5.675000 1.125000 ;
      RECT 5.505000  1.125000 5.675000 1.295000 ;
      RECT 5.505000  1.295000 6.245000 1.625000 ;
      RECT 5.505000  1.625000 5.675000 1.795000 ;
      RECT 5.845000  0.085000 6.140000 1.125000 ;
      RECT 5.845000  1.820000 6.060000 3.245000 ;
      RECT 6.755000  0.085000 7.085000 1.130000 ;
      RECT 6.835000  1.820000 7.085000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
  END
END sky130_fd_sc_hs__dlxtn_2
MACRO sky130_fd_sc_hs__dlxtn_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.455000 1.780000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.270300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.265000 0.350000 6.615000 0.980000 ;
        RECT 6.265000 0.980000 8.035000 1.150000 ;
        RECT 6.315000 1.820000 8.035000 1.990000 ;
        RECT 6.315000 1.990000 6.645000 2.980000 ;
        RECT 7.295000 0.350000 7.545000 0.980000 ;
        RECT 7.315000 1.990000 8.035000 2.150000 ;
        RECT 7.315000 2.150000 7.545000 2.980000 ;
        RECT 7.805000 1.150000 8.035000 1.820000 ;
    END
  END Q
  PIN GATE_N
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.985000 1.500000 1.315000 1.830000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.115000  0.555000 0.445000 0.660000 ;
      RECT 0.115000  0.660000 1.315000 0.830000 ;
      RECT 0.115000  0.830000 0.795000 1.130000 ;
      RECT 0.135000  1.950000 0.795000 2.120000 ;
      RECT 0.135000  2.120000 0.465000 2.980000 ;
      RECT 0.625000  0.085000 0.955000 0.490000 ;
      RECT 0.625000  1.130000 0.795000 1.950000 ;
      RECT 0.635000  2.290000 0.965000 3.245000 ;
      RECT 1.135000  1.000000 1.885000 1.330000 ;
      RECT 1.135000  2.100000 1.655000 2.390000 ;
      RECT 1.135000  2.390000 3.160000 2.560000 ;
      RECT 1.135000  2.560000 1.655000 2.980000 ;
      RECT 1.145000  0.255000 2.645000 0.425000 ;
      RECT 1.145000  0.425000 1.315000 0.660000 ;
      RECT 1.485000  0.760000 1.885000 1.000000 ;
      RECT 1.485000  1.330000 1.885000 1.770000 ;
      RECT 1.485000  1.770000 1.655000 2.100000 ;
      RECT 1.825000  1.940000 2.225000 2.220000 ;
      RECT 2.055000  0.595000 2.305000 1.720000 ;
      RECT 2.055000  1.720000 3.540000 1.890000 ;
      RECT 2.055000  1.890000 2.225000 1.940000 ;
      RECT 2.360000  2.730000 2.820000 3.245000 ;
      RECT 2.475000  0.425000 2.645000 1.220000 ;
      RECT 2.475000  1.220000 3.000000 1.550000 ;
      RECT 2.815000  0.085000 3.145000 1.050000 ;
      RECT 2.990000  2.560000 3.160000 2.905000 ;
      RECT 2.990000  2.905000 4.220000 3.075000 ;
      RECT 3.210000  1.470000 3.540000 1.720000 ;
      RECT 3.315000  0.255000 4.445000 0.505000 ;
      RECT 3.315000  0.505000 3.485000 1.470000 ;
      RECT 3.360000  2.060000 3.880000 2.735000 ;
      RECT 3.655000  0.725000 4.720000 1.055000 ;
      RECT 3.710000  1.055000 3.880000 2.060000 ;
      RECT 4.050000  1.405000 4.380000 1.735000 ;
      RECT 4.050000  1.735000 4.220000 2.905000 ;
      RECT 4.390000  1.975000 5.830000 1.990000 ;
      RECT 4.390000  1.990000 5.645000 2.305000 ;
      RECT 4.390000  2.590000 5.145000 3.245000 ;
      RECT 4.550000  1.055000 4.720000 1.320000 ;
      RECT 4.550000  1.320000 5.490000 1.650000 ;
      RECT 4.890000  0.085000 5.140000 1.055000 ;
      RECT 5.315000  1.820000 5.830000 1.975000 ;
      RECT 5.315000  2.305000 5.645000 2.980000 ;
      RECT 5.320000  0.375000 5.570000 0.980000 ;
      RECT 5.320000  0.980000 5.830000 1.150000 ;
      RECT 5.660000  1.150000 5.830000 1.320000 ;
      RECT 5.660000  1.320000 7.490000 1.650000 ;
      RECT 5.660000  1.650000 5.830000 1.820000 ;
      RECT 5.750000  0.085000 6.080000 0.810000 ;
      RECT 5.815000  2.160000 6.145000 3.245000 ;
      RECT 6.785000  0.085000 7.115000 0.810000 ;
      RECT 6.815000  2.160000 7.145000 3.245000 ;
      RECT 7.715000  0.085000 8.045000 0.810000 ;
      RECT 7.715000  2.320000 8.045000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_hs__dlxtn_4
MACRO sky130_fd_sc_hs__dlxtp_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 0.595000 1.850000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.230000 1.820000 7.595000 2.980000 ;
        RECT 7.235000 0.390000 7.595000 1.150000 ;
        RECT 7.425000 1.150000 7.595000 1.820000 ;
    END
  END Q
  PIN GATE
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.365000 1.350000 6.715000 1.780000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.680000 0.085000 ;
      RECT 0.000000  3.245000 7.680000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 1.010000 ;
      RECT 0.115000  2.100000 0.445000 3.245000 ;
      RECT 0.615000  0.420000 0.945000 1.010000 ;
      RECT 0.645000  2.100000 0.945000 2.980000 ;
      RECT 0.775000  1.010000 0.945000 1.100000 ;
      RECT 0.775000  1.100000 1.165000 1.770000 ;
      RECT 0.775000  1.770000 0.945000 2.100000 ;
      RECT 1.125000  1.940000 1.455000 2.615000 ;
      RECT 1.125000  2.615000 2.335000 2.735000 ;
      RECT 1.125000  2.735000 2.970000 2.785000 ;
      RECT 1.125000  2.785000 1.455000 2.980000 ;
      RECT 1.175000  0.405000 1.505000 0.930000 ;
      RECT 1.335000  0.930000 1.505000 1.355000 ;
      RECT 1.335000  1.355000 2.345000 1.525000 ;
      RECT 1.660000  2.955000 1.995000 3.245000 ;
      RECT 1.675000  0.085000 2.005000 1.185000 ;
      RECT 2.080000  1.940000 2.330000 2.275000 ;
      RECT 2.080000  2.275000 2.675000 2.395000 ;
      RECT 2.080000  2.395000 3.310000 2.445000 ;
      RECT 2.165000  2.785000 2.970000 2.985000 ;
      RECT 2.175000  0.255000 4.815000 0.425000 ;
      RECT 2.175000  0.425000 2.505000 0.585000 ;
      RECT 2.175000  0.755000 3.895000 0.765000 ;
      RECT 2.175000  0.765000 2.845000 0.925000 ;
      RECT 2.175000  0.925000 2.345000 1.355000 ;
      RECT 2.505000  2.445000 3.310000 2.565000 ;
      RECT 2.515000  1.095000 4.395000 1.105000 ;
      RECT 2.515000  1.105000 3.355000 1.265000 ;
      RECT 2.515000  1.265000 2.685000 1.935000 ;
      RECT 2.515000  1.935000 3.015000 2.055000 ;
      RECT 2.515000  2.055000 3.420000 2.105000 ;
      RECT 2.675000  0.595000 3.895000 0.755000 ;
      RECT 2.845000  2.105000 3.420000 2.225000 ;
      RECT 2.855000  1.435000 3.355000 1.715000 ;
      RECT 2.855000  1.715000 3.760000 1.765000 ;
      RECT 3.015000  0.935000 4.395000 1.095000 ;
      RECT 3.140000  2.565000 3.310000 2.845000 ;
      RECT 3.140000  2.845000 4.040000 3.015000 ;
      RECT 3.185000  1.765000 3.760000 1.885000 ;
      RECT 3.525000  1.275000 4.100000 1.545000 ;
      RECT 3.590000  1.885000 3.760000 2.505000 ;
      RECT 3.590000  2.505000 6.525000 2.675000 ;
      RECT 3.930000  1.545000 4.100000 2.165000 ;
      RECT 3.930000  2.165000 5.625000 2.335000 ;
      RECT 4.065000  0.775000 4.395000 0.935000 ;
      RECT 4.270000  1.665000 4.815000 1.995000 ;
      RECT 4.565000  0.425000 4.815000 0.580000 ;
      RECT 4.565000  0.580000 7.065000 0.750000 ;
      RECT 4.565000  0.750000 4.815000 1.665000 ;
      RECT 4.840000  2.845000 5.170000 3.245000 ;
      RECT 4.995000  0.085000 5.325000 0.410000 ;
      RECT 5.340000  2.675000 6.525000 2.700000 ;
      RECT 5.375000  0.920000 5.835000 1.170000 ;
      RECT 5.375000  1.170000 5.625000 2.165000 ;
      RECT 5.845000  1.350000 6.175000 1.950000 ;
      RECT 5.845000  1.950000 6.525000 2.505000 ;
      RECT 6.005000  0.920000 6.410000 1.170000 ;
      RECT 6.005000  1.170000 6.175000 1.350000 ;
      RECT 6.590000  0.085000 7.055000 0.410000 ;
      RECT 6.730000  1.950000 7.060000 3.245000 ;
      RECT 6.895000  0.750000 7.065000 1.320000 ;
      RECT 6.895000  1.320000 7.255000 1.650000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
  END
END sky130_fd_sc_hs__dlxtp_1
MACRO sky130_fd_sc_hs__dlygate4sd1_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.190000 0.730000 1.860000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.509700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.325000 0.355000 3.740000 1.120000 ;
        RECT 3.325000 1.815000 3.740000 3.060000 ;
        RECT 3.450000 1.120000 3.740000 1.815000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.095000  0.305000 0.410000 0.820000 ;
      RECT 0.095000  0.820000 1.305000 1.020000 ;
      RECT 0.095000  2.030000 1.305000 2.205000 ;
      RECT 0.095000  2.205000 0.400000 2.725000 ;
      RECT 0.575000  2.380000 0.905000 3.245000 ;
      RECT 0.585000  0.085000 0.915000 0.650000 ;
      RECT 0.975000  1.020000 1.305000 2.030000 ;
      RECT 1.415000  0.305000 1.720000 0.635000 ;
      RECT 1.415000  2.395000 1.720000 2.725000 ;
      RECT 1.475000  0.635000 1.720000 1.380000 ;
      RECT 1.475000  1.380000 2.740000 1.610000 ;
      RECT 1.475000  1.610000 1.720000 2.395000 ;
      RECT 1.985000  0.710000 2.345000 1.040000 ;
      RECT 1.985000  1.040000 3.155000 1.210000 ;
      RECT 1.985000  1.825000 3.155000 1.995000 ;
      RECT 1.985000  1.995000 2.345000 2.190000 ;
      RECT 2.825000  0.085000 3.155000 0.870000 ;
      RECT 2.825000  2.165000 3.155000 3.245000 ;
      RECT 2.910000  1.210000 3.155000 1.295000 ;
      RECT 2.910000  1.295000 3.280000 1.625000 ;
      RECT 2.910000  1.625000 3.155000 1.825000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__dlygate4sd1_1
MACRO sky130_fd_sc_hs__dlygate4sd2_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.190000 0.730000 1.860000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.509700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.325000 0.355000 3.740000 1.120000 ;
        RECT 3.325000 1.815000 3.740000 3.060000 ;
        RECT 3.450000 1.120000 3.740000 1.815000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.095000  0.305000 0.410000 0.820000 ;
      RECT 0.095000  0.820000 1.305000 1.020000 ;
      RECT 0.095000  2.030000 1.305000 2.205000 ;
      RECT 0.095000  2.205000 0.400000 2.725000 ;
      RECT 0.575000  2.380000 0.905000 3.245000 ;
      RECT 0.585000  0.085000 0.915000 0.650000 ;
      RECT 0.975000  1.020000 1.305000 2.030000 ;
      RECT 1.415000  0.305000 1.720000 0.635000 ;
      RECT 1.415000  2.395000 1.720000 2.725000 ;
      RECT 1.475000  0.635000 1.720000 1.380000 ;
      RECT 1.475000  1.380000 2.740000 1.610000 ;
      RECT 1.475000  1.610000 1.720000 2.395000 ;
      RECT 1.985000  0.710000 2.345000 1.040000 ;
      RECT 1.985000  1.040000 3.155000 1.210000 ;
      RECT 1.985000  1.825000 3.155000 1.995000 ;
      RECT 1.985000  1.995000 2.345000 2.190000 ;
      RECT 2.825000  0.085000 3.155000 0.870000 ;
      RECT 2.825000  2.165000 3.155000 3.245000 ;
      RECT 2.910000  1.210000 3.155000 1.295000 ;
      RECT 2.910000  1.295000 3.280000 1.625000 ;
      RECT 2.910000  1.625000 3.155000 1.825000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__dlygate4sd2_1
MACRO sky130_fd_sc_hs__dlygate4sd3_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.190000 0.730000 1.860000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.509700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.325000 0.355000 3.740000 1.120000 ;
        RECT 3.325000 1.815000 3.740000 3.060000 ;
        RECT 3.450000 1.120000 3.740000 1.815000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.095000  0.305000 0.410000 0.820000 ;
      RECT 0.095000  0.820000 1.305000 1.020000 ;
      RECT 0.095000  2.030000 1.305000 2.205000 ;
      RECT 0.095000  2.205000 0.400000 2.725000 ;
      RECT 0.575000  2.380000 0.905000 3.245000 ;
      RECT 0.585000  0.085000 0.915000 0.650000 ;
      RECT 0.975000  1.020000 1.305000 2.030000 ;
      RECT 1.415000  0.305000 1.720000 0.635000 ;
      RECT 1.415000  2.395000 1.720000 2.725000 ;
      RECT 1.475000  0.635000 1.720000 1.380000 ;
      RECT 1.475000  1.380000 2.740000 1.610000 ;
      RECT 1.475000  1.610000 1.720000 2.395000 ;
      RECT 1.985000  0.710000 2.345000 1.040000 ;
      RECT 1.985000  1.040000 3.155000 1.210000 ;
      RECT 1.985000  1.825000 3.155000 1.995000 ;
      RECT 1.985000  1.995000 2.345000 2.190000 ;
      RECT 2.825000  0.085000 3.155000 0.870000 ;
      RECT 2.825000  2.165000 3.155000 3.245000 ;
      RECT 2.910000  1.210000 3.155000 1.295000 ;
      RECT 2.910000  1.295000 3.280000 1.625000 ;
      RECT 2.910000  1.625000 3.155000 1.825000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__dlygate4sd3_1
MACRO sky130_fd_sc_hs__dlymetal6s2s_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.355000 0.555000 1.765000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.504100 ;
    ANTENNAPARTIALMETALSIDEAREA  0.280000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.965000 1.920000 1.345000 2.320000 ;
        RECT 0.965000 2.320000 4.210000 2.490000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.100000  0.700000 0.395000 0.975000 ;
      RECT 0.100000  0.975000 0.895000 1.145000 ;
      RECT 0.100000  1.935000 0.895000 2.140000 ;
      RECT 0.100000  2.140000 0.430000 2.225000 ;
      RECT 0.590000  0.085000 0.920000 0.805000 ;
      RECT 0.590000  2.310000 0.885000 3.245000 ;
      RECT 0.725000  1.145000 0.895000 1.275000 ;
      RECT 0.725000  1.275000 1.040000 1.605000 ;
      RECT 0.725000  1.605000 0.895000 1.935000 ;
      RECT 1.065000  1.835000 1.380000 3.075000 ;
      RECT 1.090000  0.255000 1.380000 1.075000 ;
      RECT 1.210000  1.075000 1.380000 1.315000 ;
      RECT 1.210000  1.315000 1.995000 1.605000 ;
      RECT 1.210000  1.605000 1.380000 1.835000 ;
      RECT 1.550000  0.700000 1.835000 0.975000 ;
      RECT 1.550000  0.975000 2.335000 1.145000 ;
      RECT 1.550000  1.895000 2.335000 2.140000 ;
      RECT 1.550000  2.140000 1.870000 2.225000 ;
      RECT 2.030000  0.085000 2.360000 0.805000 ;
      RECT 2.100000  2.310000 2.395000 3.245000 ;
      RECT 2.165000  1.145000 2.335000 1.275000 ;
      RECT 2.165000  1.275000 2.525000 1.605000 ;
      RECT 2.165000  1.605000 2.335000 1.895000 ;
      RECT 2.505000  1.835000 2.865000 2.160000 ;
      RECT 2.530000  0.255000 2.865000 1.075000 ;
      RECT 2.565000  2.160000 2.865000 3.075000 ;
      RECT 2.695000  1.075000 2.865000 1.315000 ;
      RECT 2.695000  1.315000 3.435000 1.605000 ;
      RECT 2.695000  1.605000 2.865000 1.835000 ;
      RECT 3.060000  0.700000 3.275000 0.975000 ;
      RECT 3.060000  0.975000 3.775000 1.145000 ;
      RECT 3.070000  1.895000 3.805000 2.140000 ;
      RECT 3.070000  2.140000 3.400000 2.225000 ;
      RECT 3.470000  0.085000 3.800000 0.805000 ;
      RECT 3.585000  2.310000 3.880000 3.245000 ;
      RECT 3.605000  1.145000 3.775000 1.275000 ;
      RECT 3.605000  1.275000 4.010000 1.605000 ;
      RECT 3.605000  1.605000 3.805000 1.895000 ;
      RECT 3.970000  0.255000 4.350000 1.075000 ;
      RECT 3.975000  1.835000 4.350000 2.160000 ;
      RECT 4.050000  2.160000 4.350000 3.075000 ;
      RECT 4.180000  1.075000 4.350000 1.835000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  1.950000 1.285000 2.120000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  1.950000 2.725000 2.120000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  1.950000 4.165000 2.120000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
    LAYER met1 ;
      RECT 2.405000 1.920000 2.785000 2.150000 ;
      RECT 3.845000 1.920000 4.225000 2.150000 ;
  END
END sky130_fd_sc_hs__dlymetal6s2s_1
MACRO sky130_fd_sc_hs__dlymetal6s4s_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.355000 0.555000 1.765000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.504100 ;
    ANTENNAPARTIALMETALSIDEAREA  0.280000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.965000 2.320000 4.210000 2.490000 ;
        RECT 2.405000 1.920000 2.785000 2.320000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.100000  0.700000 0.395000 0.975000 ;
      RECT 0.100000  0.975000 0.895000 1.145000 ;
      RECT 0.100000  1.935000 0.895000 2.140000 ;
      RECT 0.100000  2.140000 0.430000 2.225000 ;
      RECT 0.590000  0.085000 0.920000 0.805000 ;
      RECT 0.590000  2.310000 0.885000 3.245000 ;
      RECT 0.725000  1.145000 0.895000 1.275000 ;
      RECT 0.725000  1.275000 1.040000 1.605000 ;
      RECT 0.725000  1.605000 0.895000 1.935000 ;
      RECT 1.065000  1.835000 1.380000 3.075000 ;
      RECT 1.090000  0.255000 1.380000 1.075000 ;
      RECT 1.210000  1.075000 1.380000 1.315000 ;
      RECT 1.210000  1.315000 1.995000 1.605000 ;
      RECT 1.210000  1.605000 1.380000 1.835000 ;
      RECT 1.550000  0.700000 1.835000 0.975000 ;
      RECT 1.550000  0.975000 2.335000 1.145000 ;
      RECT 1.550000  1.895000 2.335000 2.140000 ;
      RECT 1.550000  2.140000 1.870000 2.225000 ;
      RECT 2.030000  0.085000 2.360000 0.805000 ;
      RECT 2.100000  2.310000 2.395000 3.245000 ;
      RECT 2.165000  1.145000 2.335000 1.275000 ;
      RECT 2.165000  1.275000 2.525000 1.605000 ;
      RECT 2.165000  1.605000 2.335000 1.895000 ;
      RECT 2.505000  1.835000 2.865000 2.160000 ;
      RECT 2.530000  0.255000 2.865000 1.075000 ;
      RECT 2.565000  2.160000 2.865000 3.075000 ;
      RECT 2.695000  1.075000 2.865000 1.315000 ;
      RECT 2.695000  1.315000 3.435000 1.605000 ;
      RECT 2.695000  1.605000 2.865000 1.835000 ;
      RECT 3.060000  0.700000 3.275000 0.975000 ;
      RECT 3.060000  0.975000 3.775000 1.145000 ;
      RECT 3.070000  1.895000 3.805000 2.140000 ;
      RECT 3.070000  2.140000 3.400000 2.225000 ;
      RECT 3.470000  0.085000 3.800000 0.805000 ;
      RECT 3.585000  2.310000 3.880000 3.245000 ;
      RECT 3.605000  1.145000 3.775000 1.275000 ;
      RECT 3.605000  1.275000 4.010000 1.605000 ;
      RECT 3.605000  1.605000 3.805000 1.895000 ;
      RECT 3.970000  0.255000 4.350000 1.075000 ;
      RECT 3.975000  1.835000 4.350000 2.160000 ;
      RECT 4.050000  2.160000 4.350000 3.075000 ;
      RECT 4.180000  1.075000 4.350000 1.835000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  1.950000 1.285000 2.120000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  1.950000 2.725000 2.120000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  1.950000 4.165000 2.120000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
    LAYER met1 ;
      RECT 0.965000 1.920000 1.345000 2.150000 ;
      RECT 3.845000 1.920000 4.225000 2.150000 ;
  END
END sky130_fd_sc_hs__dlymetal6s4s_1
MACRO sky130_fd_sc_hs__dlymetal6s6s_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.355000 0.555000 1.765000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.504100 ;
    ANTENNAPARTIALMETALSIDEAREA  0.290500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.965000 2.320000 4.225000 2.490000 ;
        RECT 3.845000 1.920000 4.225000 2.320000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.100000  0.700000 0.395000 0.975000 ;
      RECT 0.100000  0.975000 0.895000 1.145000 ;
      RECT 0.100000  1.935000 0.895000 2.140000 ;
      RECT 0.100000  2.140000 0.430000 2.225000 ;
      RECT 0.590000  0.085000 0.920000 0.805000 ;
      RECT 0.590000  2.310000 0.885000 3.245000 ;
      RECT 0.725000  1.145000 0.895000 1.275000 ;
      RECT 0.725000  1.275000 1.040000 1.605000 ;
      RECT 0.725000  1.605000 0.895000 1.935000 ;
      RECT 1.065000  1.835000 1.380000 3.075000 ;
      RECT 1.090000  0.255000 1.380000 1.075000 ;
      RECT 1.210000  1.075000 1.380000 1.315000 ;
      RECT 1.210000  1.315000 1.995000 1.605000 ;
      RECT 1.210000  1.605000 1.380000 1.835000 ;
      RECT 1.550000  0.700000 1.835000 0.975000 ;
      RECT 1.550000  0.975000 2.335000 1.145000 ;
      RECT 1.550000  1.895000 2.335000 2.140000 ;
      RECT 1.550000  2.140000 1.870000 2.225000 ;
      RECT 2.030000  0.085000 2.360000 0.805000 ;
      RECT 2.100000  2.310000 2.395000 3.245000 ;
      RECT 2.165000  1.145000 2.335000 1.275000 ;
      RECT 2.165000  1.275000 2.525000 1.605000 ;
      RECT 2.165000  1.605000 2.335000 1.895000 ;
      RECT 2.505000  1.835000 2.865000 2.160000 ;
      RECT 2.530000  0.255000 2.865000 1.075000 ;
      RECT 2.565000  2.160000 2.865000 3.075000 ;
      RECT 2.695000  1.075000 2.865000 1.315000 ;
      RECT 2.695000  1.315000 3.435000 1.605000 ;
      RECT 2.695000  1.605000 2.865000 1.835000 ;
      RECT 3.060000  0.700000 3.275000 0.975000 ;
      RECT 3.060000  0.975000 3.775000 1.145000 ;
      RECT 3.070000  1.895000 3.805000 2.140000 ;
      RECT 3.070000  2.140000 3.400000 2.225000 ;
      RECT 3.470000  0.085000 3.800000 0.805000 ;
      RECT 3.585000  2.310000 3.880000 3.245000 ;
      RECT 3.605000  1.145000 3.775000 1.275000 ;
      RECT 3.605000  1.275000 4.010000 1.605000 ;
      RECT 3.605000  1.605000 3.805000 1.895000 ;
      RECT 3.970000  0.255000 4.350000 1.075000 ;
      RECT 3.975000  1.835000 4.350000 2.160000 ;
      RECT 4.050000  2.160000 4.350000 3.075000 ;
      RECT 4.180000  1.075000 4.350000 1.835000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  1.950000 1.285000 2.120000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  1.950000 2.725000 2.120000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  1.950000 4.165000 2.120000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
    LAYER met1 ;
      RECT 0.965000 1.920000 1.345000 2.150000 ;
      RECT 2.405000 1.920000 2.785000 2.150000 ;
  END
END sky130_fd_sc_hs__dlymetal6s6s_1
MACRO sky130_fd_sc_hs__ebufn_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.500000 1.795000 1.830000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.377000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.500000 0.835000 1.830000 ;
        RECT 0.665000 1.830000 0.835000 2.420000 ;
        RECT 0.665000 2.420000 2.195000 2.590000 ;
        RECT 1.865000 2.340000 2.195000 2.420000 ;
        RECT 1.865000 2.590000 2.195000 3.010000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.210000 0.350000 3.755000 1.130000 ;
        RECT 3.235000 1.820000 3.755000 2.980000 ;
        RECT 3.585000 1.130000 3.755000 1.820000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.085000  0.455000 0.530000 1.150000 ;
      RECT 0.085000  1.150000 2.200000 1.320000 ;
      RECT 0.085000  1.320000 0.255000 2.000000 ;
      RECT 0.085000  2.000000 0.445000 2.880000 ;
      RECT 0.650000  2.760000 0.980000 3.245000 ;
      RECT 0.700000  0.085000 0.985000 0.850000 ;
      RECT 1.155000  0.455000 1.450000 0.810000 ;
      RECT 1.155000  0.810000 2.660000 0.980000 ;
      RECT 1.185000  2.000000 2.135000 2.170000 ;
      RECT 1.185000  2.170000 1.695000 2.250000 ;
      RECT 1.870000  1.320000 2.200000 1.340000 ;
      RECT 1.965000  1.710000 3.065000 1.880000 ;
      RECT 1.965000  1.880000 2.135000 2.000000 ;
      RECT 2.365000  2.050000 2.695000 3.245000 ;
      RECT 2.390000  0.085000 2.720000 0.640000 ;
      RECT 2.460000  0.980000 2.660000 1.320000 ;
      RECT 2.460000  1.320000 3.415000 1.650000 ;
      RECT 2.460000  1.650000 3.065000 1.710000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__ebufn_1
MACRO sky130_fd_sc_hs__ebufn_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.350000 3.865000 1.780000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.582000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.965000 1.180000 3.295000 1.650000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.599200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.615000 0.875000 1.130000 ;
        RECT 0.535000 1.130000 0.705000 1.800000 ;
        RECT 0.535000 1.800000 1.795000 1.970000 ;
        RECT 0.645000 1.970000 1.795000 2.150000 ;
        RECT 0.645000 2.150000 0.975000 2.735000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  0.255000 1.375000 0.425000 ;
      RECT 0.115000  0.425000 0.365000 1.130000 ;
      RECT 0.145000  2.140000 0.475000 2.905000 ;
      RECT 0.145000  2.905000 1.475000 3.075000 ;
      RECT 0.875000  1.300000 2.135000 1.630000 ;
      RECT 1.045000  0.425000 1.375000 0.960000 ;
      RECT 1.045000  0.960000 2.225000 1.130000 ;
      RECT 1.145000  2.320000 1.475000 2.580000 ;
      RECT 1.145000  2.580000 2.545000 2.750000 ;
      RECT 1.145000  2.750000 1.475000 2.905000 ;
      RECT 1.545000  0.085000 1.795000 0.790000 ;
      RECT 1.680000  2.920000 2.010000 3.245000 ;
      RECT 1.965000  1.630000 2.135000 2.240000 ;
      RECT 1.965000  2.240000 4.205000 2.410000 ;
      RECT 1.975000  0.350000 2.225000 0.960000 ;
      RECT 2.215000  2.750000 2.545000 2.980000 ;
      RECT 2.395000  0.325000 3.170000 1.010000 ;
      RECT 2.395000  1.010000 2.725000 1.820000 ;
      RECT 2.395000  1.820000 3.105000 2.070000 ;
      RECT 3.225000  2.610000 3.705000 3.245000 ;
      RECT 3.340000  0.085000 3.670000 1.010000 ;
      RECT 3.840000  0.350000 4.205000 1.030000 ;
      RECT 3.875000  1.950000 4.205000 2.240000 ;
      RECT 3.875000  2.410000 4.205000 2.860000 ;
      RECT 4.035000  1.030000 4.205000 1.950000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__ebufn_2
MACRO sky130_fd_sc_hs__ebufn_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.300000 0.805000 1.780000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.951000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.975000 1.180000 1.285000 1.550000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  1.101200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.970000 1.820000 5.205000 1.990000 ;
        RECT 3.970000 1.990000 4.300000 2.735000 ;
        RECT 4.015000 0.595000 4.345000 0.980000 ;
        RECT 4.015000 0.980000 5.205000 1.150000 ;
        RECT 4.870000 1.990000 5.205000 2.735000 ;
        RECT 4.875000 0.595000 5.205000 0.980000 ;
        RECT 5.035000 1.150000 5.205000 1.820000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.085000  0.350000 0.405000 1.130000 ;
      RECT 0.085000  1.130000 0.255000 1.950000 ;
      RECT 0.085000  1.950000 0.365000 2.390000 ;
      RECT 0.085000  2.390000 1.630000 2.560000 ;
      RECT 0.085000  2.560000 0.365000 2.980000 ;
      RECT 0.565000  2.730000 0.920000 3.245000 ;
      RECT 0.585000  0.085000 0.915000 1.010000 ;
      RECT 1.040000  1.720000 1.775000 1.890000 ;
      RECT 1.040000  1.890000 1.290000 2.220000 ;
      RECT 1.095000  0.300000 1.775000 1.010000 ;
      RECT 1.455000  1.010000 1.775000 1.720000 ;
      RECT 1.460000  2.060000 2.530000 2.230000 ;
      RECT 1.460000  2.230000 1.630000 2.390000 ;
      RECT 1.800000  2.400000 2.870000 2.570000 ;
      RECT 1.800000  2.570000 1.970000 2.820000 ;
      RECT 1.945000  0.350000 2.115000 1.140000 ;
      RECT 1.945000  1.140000 3.835000 1.150000 ;
      RECT 1.945000  1.150000 2.975000 1.310000 ;
      RECT 2.170000  2.740000 2.500000 3.245000 ;
      RECT 2.295000  0.085000 2.625000 0.970000 ;
      RECT 2.360000  1.480000 4.830000 1.650000 ;
      RECT 2.360000  1.650000 2.530000 2.060000 ;
      RECT 2.700000  1.820000 3.770000 1.990000 ;
      RECT 2.700000  1.990000 2.870000 2.400000 ;
      RECT 2.700000  2.570000 2.870000 2.980000 ;
      RECT 2.805000  0.350000 2.975000 0.980000 ;
      RECT 2.805000  0.980000 3.835000 1.140000 ;
      RECT 3.070000  2.160000 3.320000 3.245000 ;
      RECT 3.155000  0.085000 3.405000 0.810000 ;
      RECT 3.520000  1.990000 3.770000 2.905000 ;
      RECT 3.520000  2.905000 5.650000 3.075000 ;
      RECT 3.585000  0.255000 5.655000 0.425000 ;
      RECT 3.585000  0.425000 3.835000 0.980000 ;
      RECT 3.820000  1.320000 4.830000 1.480000 ;
      RECT 4.470000  2.160000 4.700000 2.905000 ;
      RECT 4.525000  0.425000 4.695000 0.810000 ;
      RECT 5.400000  1.820000 5.650000 2.905000 ;
      RECT 5.405000  0.425000 5.655000 1.130000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_hs__ebufn_4
MACRO sky130_fd_sc_hs__ebufn_8
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.56000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.645000 1.180000 9.975000 1.550000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  1.623000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.265000 1.180000 9.475000 1.550000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  2.360500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.595000 0.875000 0.980000 ;
        RECT 0.545000 0.980000 3.760000 1.150000 ;
        RECT 0.545000 1.150000 0.835000 1.820000 ;
        RECT 0.545000 1.820000 3.700000 1.990000 ;
        RECT 0.545000 1.990000 0.900000 2.735000 ;
        RECT 1.430000 0.595000 1.760000 0.980000 ;
        RECT 1.520000 1.990000 1.850000 2.735000 ;
        RECT 2.420000 1.990000 2.750000 2.735000 ;
        RECT 2.430000 0.595000 2.760000 0.980000 ;
        RECT 3.370000 1.990000 3.700000 2.735000 ;
        RECT 3.430000 0.595000 3.760000 0.980000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.560000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.560000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 10.560000 0.085000 ;
      RECT  0.000000  3.245000 10.560000 3.415000 ;
      RECT  0.115000  0.255000  4.110000 0.425000 ;
      RECT  0.115000  0.425000  0.365000 1.130000 ;
      RECT  0.120000  1.820000  0.370000 2.905000 ;
      RECT  0.120000  2.905000  4.200000 3.075000 ;
      RECT  1.035000  1.320000  3.655000 1.480000 ;
      RECT  1.035000  1.480000  4.040000 1.650000 ;
      RECT  1.055000  0.425000  1.225000 0.810000 ;
      RECT  1.085000  2.160000  1.350000 2.905000 ;
      RECT  1.930000  0.425000  2.260000 0.810000 ;
      RECT  2.050000  2.160000  2.220000 2.905000 ;
      RECT  2.920000  2.160000  3.190000 2.905000 ;
      RECT  2.930000  0.425000  3.260000 0.810000 ;
      RECT  3.870000  1.650000  4.040000 2.050000 ;
      RECT  3.870000  2.050000  7.755000 2.220000 ;
      RECT  3.870000  2.390000  7.200000 2.560000 ;
      RECT  3.870000  2.560000  4.200000 2.905000 ;
      RECT  3.940000  0.425000  4.110000 1.140000 ;
      RECT  3.940000  1.140000  5.050000 1.300000 ;
      RECT  3.940000  1.300000  7.550000 1.310000 ;
      RECT  4.290000  0.085000  4.620000 0.970000 ;
      RECT  4.370000  2.730000  4.700000 3.245000 ;
      RECT  4.720000  1.310000  7.550000 1.470000 ;
      RECT  4.800000  0.350000  5.050000 1.140000 ;
      RECT  4.870000  2.560000  5.200000 2.980000 ;
      RECT  5.230000  0.085000  5.400000 1.130000 ;
      RECT  5.370000  2.730000  5.700000 3.245000 ;
      RECT  5.580000  0.350000  5.830000 1.300000 ;
      RECT  5.870000  2.560000  6.200000 2.980000 ;
      RECT  6.010000  0.085000  6.260000 1.130000 ;
      RECT  6.370000  2.730000  6.700000 3.245000 ;
      RECT  6.440000  0.350000  6.690000 1.300000 ;
      RECT  6.870000  0.085000  7.120000 1.130000 ;
      RECT  6.870000  2.560000  8.270000 2.730000 ;
      RECT  6.870000  2.730000  7.200000 2.980000 ;
      RECT  7.300000  0.350000  7.550000 1.300000 ;
      RECT  7.405000  2.900000  7.735000 3.245000 ;
      RECT  7.585000  2.220000  9.945000 2.390000 ;
      RECT  7.720000  0.340000  9.150000 0.670000 ;
      RECT  7.925000  0.670000  9.150000 1.010000 ;
      RECT  7.925000  1.010000  8.095000 1.800000 ;
      RECT  7.925000  1.800000  9.045000 2.050000 ;
      RECT  7.940000  2.730000  8.270000 2.980000 ;
      RECT  9.165000  2.560000  9.495000 3.245000 ;
      RECT  9.330000  0.085000  9.500000 1.010000 ;
      RECT  9.665000  1.720000 10.315000 1.890000 ;
      RECT  9.665000  1.890000  9.945000 2.220000 ;
      RECT  9.665000  2.390000  9.945000 2.980000 ;
      RECT  9.680000  0.340000  9.930000 0.840000 ;
      RECT  9.680000  0.840000 10.315000 1.010000 ;
      RECT 10.110000  0.085000 10.445000 0.600000 ;
      RECT 10.115000  2.060000 10.445000 3.245000 ;
      RECT 10.145000  1.010000 10.315000 1.720000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
  END
END sky130_fd_sc_hs__ebufn_8
MACRO sky130_fd_sc_hs__edfxbp_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.40000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.980000 0.835000 1.990000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.285000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.450000 1.905000 1.780000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.765000 0.620000 13.095000 1.000000 ;
        RECT 12.925000 1.000000 13.095000 1.820000 ;
        RECT 12.925000 1.820000 13.340000 2.980000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.955000 0.370000 14.315000 1.150000 ;
        RECT 13.990000 1.820000 14.315000 2.980000 ;
        RECT 14.145000 1.150000 14.315000 1.820000 ;
    END
  END Q_N
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.715000 1.180000 4.385000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 14.400000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 14.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.400000 0.085000 ;
      RECT  0.000000  3.245000 14.400000 3.415000 ;
      RECT  0.085000  0.420000  0.600000 0.750000 ;
      RECT  0.085000  0.750000  0.255000 2.290000 ;
      RECT  0.085000  2.290000  1.545000 2.460000 ;
      RECT  0.085000  2.460000  0.445000 2.980000 ;
      RECT  0.955000  2.630000  1.205000 3.245000 ;
      RECT  1.005000  1.110000  2.000000 1.280000 ;
      RECT  1.005000  1.280000  1.335000 1.950000 ;
      RECT  1.005000  1.950000  2.665000 2.120000 ;
      RECT  1.090000  0.085000  1.420000 0.810000 ;
      RECT  1.375000  2.460000  1.545000 2.905000 ;
      RECT  1.375000  2.905000  2.225000 3.075000 ;
      RECT  1.650000  0.480000  2.000000 1.110000 ;
      RECT  1.715000  2.120000  1.885000 2.735000 ;
      RECT  2.055000  2.290000  3.545000 2.310000 ;
      RECT  2.055000  2.310000  5.775000 2.460000 ;
      RECT  2.055000  2.460000  2.225000 2.905000 ;
      RECT  2.170000  0.085000  2.500000 0.810000 ;
      RECT  2.335000  0.980000  2.665000 1.950000 ;
      RECT  2.395000  2.630000  2.645000 3.245000 ;
      RECT  2.875000  0.980000  3.205000 1.990000 ;
      RECT  3.000000  0.350000  3.545000 0.810000 ;
      RECT  3.155000  2.460000  5.775000 2.480000 ;
      RECT  3.155000  2.480000  3.545000 2.960000 ;
      RECT  3.375000  0.810000  3.545000 2.290000 ;
      RECT  3.715000  0.085000  3.885000 1.010000 ;
      RECT  3.715000  2.650000  4.045000 3.245000 ;
      RECT  4.065000  0.350000  4.395000 0.840000 ;
      RECT  4.065000  0.840000  4.725000 1.010000 ;
      RECT  4.165000  1.810000  4.965000 2.140000 ;
      RECT  4.555000  1.010000  4.725000 1.810000 ;
      RECT  4.585000  0.085000  4.915000 0.670000 ;
      RECT  5.095000  0.255000  6.885000 0.425000 ;
      RECT  5.095000  0.425000  5.345000 1.130000 ;
      RECT  5.105000  2.650000  5.435000 3.245000 ;
      RECT  5.215000  1.300000  5.785000 1.470000 ;
      RECT  5.215000  1.470000  5.385000 2.310000 ;
      RECT  5.535000  0.595000  5.785000 1.300000 ;
      RECT  5.555000  1.810000  6.125000 1.970000 ;
      RECT  5.555000  1.970000  6.355000 2.140000 ;
      RECT  5.605000  2.480000  5.775000 2.890000 ;
      RECT  5.605000  2.890000  6.445000 3.060000 ;
      RECT  5.955000  0.425000  6.125000 1.810000 ;
      RECT  5.955000  2.140000  6.355000 2.380000 ;
      RECT  6.295000  0.595000  6.465000 1.515000 ;
      RECT  6.295000  1.515000  6.720000 1.685000 ;
      RECT  6.550000  1.685000  6.720000 1.740000 ;
      RECT  6.550000  1.740000  8.260000 1.910000 ;
      RECT  6.550000  1.910000  6.720000 2.550000 ;
      RECT  6.550000  2.550000  6.980000 2.720000 ;
      RECT  6.635000  0.425000  6.885000 0.965000 ;
      RECT  6.635000  0.965000  7.810000 1.135000 ;
      RECT  6.635000  1.135000  6.885000 1.345000 ;
      RECT  6.650000  2.720000  6.980000 2.980000 ;
      RECT  6.890000  2.080000  7.320000 2.380000 ;
      RECT  7.150000  2.380000  7.320000 2.545000 ;
      RECT  7.150000  2.545000  8.365000 2.715000 ;
      RECT  7.205000  1.305000  9.030000 1.475000 ;
      RECT  7.205000  1.475000  7.535000 1.570000 ;
      RECT  7.220000  0.085000  7.470000 0.795000 ;
      RECT  7.640000  0.255000  8.490000 0.425000 ;
      RECT  7.640000  0.425000  7.810000 0.965000 ;
      RECT  7.695000  2.885000  8.025000 3.245000 ;
      RECT  7.930000  1.645000  8.260000 1.740000 ;
      RECT  7.930000  1.910000  8.260000 1.955000 ;
      RECT  7.980000  0.595000  8.150000 1.305000 ;
      RECT  8.195000  2.715000  8.365000 2.755000 ;
      RECT  8.195000  2.755000  9.405000 2.925000 ;
      RECT  8.230000  2.125000  9.030000 2.375000 ;
      RECT  8.320000  0.425000  8.490000 0.965000 ;
      RECT  8.320000  0.965000  9.370000 1.120000 ;
      RECT  8.320000  1.120000 11.105000 1.135000 ;
      RECT  8.660000  0.085000  8.910000 0.770000 ;
      RECT  8.700000  1.475000  9.030000 2.125000 ;
      RECT  8.700000  2.375000  9.030000 2.585000 ;
      RECT  9.200000  1.135000 11.105000 1.290000 ;
      RECT  9.200000  1.290000 10.085000 1.450000 ;
      RECT  9.235000  1.620000 10.625000 1.790000 ;
      RECT  9.235000  1.790000  9.405000 2.755000 ;
      RECT  9.540000  0.620000 11.445000 0.950000 ;
      RECT  9.575000  1.960000  9.905000 3.245000 ;
      RECT 10.295000  1.460000 10.625000 1.620000 ;
      RECT 10.445000  1.985000 11.445000 2.155000 ;
      RECT 10.445000  2.155000 10.775000 2.980000 ;
      RECT 10.835000  1.290000 11.105000 1.800000 ;
      RECT 11.275000  0.950000 11.445000 1.155000 ;
      RECT 11.275000  1.155000 11.985000 1.485000 ;
      RECT 11.275000  1.485000 11.445000 1.985000 ;
      RECT 11.495000  2.325000 12.280000 3.245000 ;
      RECT 11.615000  1.725000 12.485000 1.805000 ;
      RECT 11.615000  1.805000 12.700000 2.120000 ;
      RECT 11.655000  0.085000 11.985000 0.985000 ;
      RECT 12.155000  0.255000 13.435000 0.425000 ;
      RECT 12.155000  0.425000 12.485000 1.725000 ;
      RECT 12.450000  2.120000 12.700000 2.845000 ;
      RECT 13.265000  0.425000 13.435000 1.320000 ;
      RECT 13.265000  1.320000 13.975000 1.650000 ;
      RECT 13.540000  1.820000 13.790000 3.245000 ;
      RECT 13.605000  0.085000 13.775000 1.150000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  1.580000  3.205000 1.750000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  1.580000 12.325000 1.750000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
    LAYER met1 ;
      RECT  2.975000 1.550000  3.265000 1.595000 ;
      RECT  2.975000 1.595000 12.385000 1.735000 ;
      RECT  2.975000 1.735000  3.265000 1.780000 ;
      RECT 12.095000 1.550000 12.385000 1.595000 ;
      RECT 12.095000 1.735000 12.385000 1.780000 ;
  END
END sky130_fd_sc_hs__edfxbp_1
MACRO sky130_fd_sc_hs__edfxtp_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.96000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.980000 0.805000 1.990000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.285000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.515000 1.110000 1.845000 1.440000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.518900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.015000 0.350000 12.345000 1.130000 ;
        RECT 12.075000 1.130000 12.345000 1.550000 ;
        RECT 12.075000 1.550000 12.405000 2.980000 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.450000 1.180000 3.780000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.960000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 12.960000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.960000 0.085000 ;
      RECT  0.000000  3.245000 12.960000 3.415000 ;
      RECT  0.085000  0.340000  0.530000 0.810000 ;
      RECT  0.085000  0.810000  0.255000 2.180000 ;
      RECT  0.085000  2.180000  1.535000 2.350000 ;
      RECT  0.085000  2.350000  0.435000 2.980000 ;
      RECT  0.945000  2.520000  1.195000 3.245000 ;
      RECT  0.975000  0.770000  1.820000 0.940000 ;
      RECT  0.975000  0.940000  1.305000 1.610000 ;
      RECT  0.975000  1.610000  2.385000 1.780000 ;
      RECT  0.975000  1.780000  1.305000 2.010000 ;
      RECT  1.020000  0.085000  1.350000 0.600000 ;
      RECT  1.365000  2.350000  1.535000 2.905000 ;
      RECT  1.365000  2.905000  2.215000 3.075000 ;
      RECT  1.570000  0.415000  1.820000 0.770000 ;
      RECT  1.705000  1.780000  1.875000 2.735000 ;
      RECT  2.000000  0.085000  2.330000 0.875000 ;
      RECT  2.045000  1.950000  3.270000 2.120000 ;
      RECT  2.045000  2.120000  2.215000 2.905000 ;
      RECT  2.055000  1.385000  2.385000 1.610000 ;
      RECT  2.385000  2.290000  2.635000 3.245000 ;
      RECT  2.555000  1.045000  2.930000 1.780000 ;
      RECT  2.790000  0.415000  3.270000 0.875000 ;
      RECT  3.100000  0.875000  3.270000 1.950000 ;
      RECT  3.100000  2.120000  3.475000 2.310000 ;
      RECT  3.100000  2.310000  5.610000 2.480000 ;
      RECT  3.100000  2.480000  3.475000 2.620000 ;
      RECT  3.440000  0.085000  3.610000 1.010000 ;
      RECT  3.670000  2.650000  4.000000 3.245000 ;
      RECT  3.790000  0.350000  4.120000 1.010000 ;
      RECT  3.950000  1.010000  4.120000 1.470000 ;
      RECT  3.950000  1.470000  4.900000 2.140000 ;
      RECT  4.335000  0.085000  4.585000 1.130000 ;
      RECT  4.765000  0.255000  6.960000 0.425000 ;
      RECT  4.765000  0.425000  5.095000 1.130000 ;
      RECT  5.020000  2.650000  5.270000 3.245000 ;
      RECT  5.130000  1.480000  5.655000 1.650000 ;
      RECT  5.130000  1.650000  5.300000 2.310000 ;
      RECT  5.325000  0.595000  5.655000 1.480000 ;
      RECT  5.440000  2.480000  5.610000 2.520000 ;
      RECT  5.440000  2.520000  6.245000 2.690000 ;
      RECT  5.470000  1.820000  5.995000 1.970000 ;
      RECT  5.470000  1.970000  6.245000 2.140000 ;
      RECT  5.825000  0.425000  5.995000 1.820000 ;
      RECT  5.825000  2.140000  6.245000 2.300000 ;
      RECT  5.995000  2.690000  6.245000 2.980000 ;
      RECT  6.165000  0.595000  6.620000 0.765000 ;
      RECT  6.165000  0.765000  6.335000 1.630000 ;
      RECT  6.165000  1.630000  8.030000 1.800000 ;
      RECT  6.415000  1.800000  6.585000 2.520000 ;
      RECT  6.415000  2.520000  6.775000 2.980000 ;
      RECT  6.505000  0.935000  7.760000 1.105000 ;
      RECT  6.505000  1.105000  6.960000 1.310000 ;
      RECT  6.755000  2.000000  7.115000 2.330000 ;
      RECT  6.790000  0.425000  6.960000 0.935000 ;
      RECT  6.945000  2.330000  7.115000 2.410000 ;
      RECT  6.945000  2.410000  9.800000 2.580000 ;
      RECT  7.130000  1.275000  8.940000 1.445000 ;
      RECT  7.130000  1.445000  7.460000 1.460000 ;
      RECT  7.170000  0.085000  7.420000 0.765000 ;
      RECT  7.410000  2.750000  7.740000 3.245000 ;
      RECT  7.590000  0.255000  8.440000 0.425000 ;
      RECT  7.590000  0.425000  7.760000 0.935000 ;
      RECT  7.700000  1.615000  8.030000 1.630000 ;
      RECT  7.700000  1.800000  8.030000 1.830000 ;
      RECT  7.930000  0.595000  8.100000 1.275000 ;
      RECT  7.945000  2.070000  8.440000 2.240000 ;
      RECT  8.270000  0.425000  8.440000 0.935000 ;
      RECT  8.270000  0.935000  9.280000 1.105000 ;
      RECT  8.270000  1.445000  8.940000 1.605000 ;
      RECT  8.270000  1.605000  8.440000 2.070000 ;
      RECT  8.505000  2.750000  8.835000 3.245000 ;
      RECT  8.610000  0.085000  8.860000 0.765000 ;
      RECT  9.110000  1.105000  9.280000 1.205000 ;
      RECT  9.110000  1.205000 10.605000 1.375000 ;
      RECT  9.110000  1.375000  9.460000 1.550000 ;
      RECT  9.450000  0.350000  9.780000 0.835000 ;
      RECT  9.450000  0.835000 10.945000 1.005000 ;
      RECT  9.630000  1.545000 10.065000 1.725000 ;
      RECT  9.630000  1.725000  9.800000 2.410000 ;
      RECT  9.970000  1.925000 10.405000 2.095000 ;
      RECT  9.970000  2.095000 10.220000 3.000000 ;
      RECT 10.235000  1.755000 10.945000 1.925000 ;
      RECT 10.275000  1.375000 10.605000 1.585000 ;
      RECT 10.350000  0.085000 11.310000 0.665000 ;
      RECT 10.665000  2.095000 11.885000 2.320000 ;
      RECT 10.775000  1.005000 11.505000 1.335000 ;
      RECT 10.775000  1.335000 10.945000 1.755000 ;
      RECT 10.845000  2.525000 11.385000 3.245000 ;
      RECT 11.490000  0.335000 11.845000 0.810000 ;
      RECT 11.555000  2.320000 11.885000 2.950000 ;
      RECT 11.645000  1.550000 11.885000 2.095000 ;
      RECT 11.675000  0.810000 11.845000 1.550000 ;
      RECT 12.515000  0.085000 12.845000 1.130000 ;
      RECT 12.605000  1.820000 12.855000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  1.580000  2.725000 1.750000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  1.580000 11.845000 1.750000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
    LAYER met1 ;
      RECT  2.495000 1.550000  2.785000 1.595000 ;
      RECT  2.495000 1.595000 11.905000 1.735000 ;
      RECT  2.495000 1.735000  2.785000 1.780000 ;
      RECT 11.615000 1.550000 11.905000 1.595000 ;
      RECT 11.615000 1.735000 11.905000 1.780000 ;
  END
END sky130_fd_sc_hs__edfxtp_1
MACRO sky130_fd_sc_hs__einvn_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.400000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.350000 1.975000 1.780000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.327000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455000 1.430000 1.315000 1.760000 ;
        RECT 1.085000 1.760000 1.315000 1.780000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.765000 1.950000 2.315000 2.980000 ;
        RECT 1.770000 0.480000 2.315000 1.180000 ;
        RECT 2.145000 1.180000 2.315000 1.950000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.400000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.400000 0.085000 ;
      RECT 0.000000  3.245000 2.400000 3.415000 ;
      RECT 0.110000  0.255000 0.780000 0.560000 ;
      RECT 0.110000  0.560000 0.770000 1.250000 ;
      RECT 0.110000  1.250000 0.280000 1.930000 ;
      RECT 0.110000  1.930000 0.720000 2.100000 ;
      RECT 0.390000  2.100000 0.720000 2.580000 ;
      RECT 0.925000  1.950000 1.255000 3.245000 ;
      RECT 0.950000  0.085000 1.280000 1.260000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
  END
END sky130_fd_sc_hs__einvn_1
MACRO sky130_fd_sc_hs__einvn_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925000 0.810000 3.255000 1.550000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.120000 0.550000 2.130000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.546900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.425000 0.770000 2.755000 1.130000 ;
        RECT 2.465000 1.130000 2.755000 1.820000 ;
        RECT 2.465000 1.820000 2.795000 2.735000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.110000  2.300000 0.360000 3.245000 ;
      RECT 0.130000  0.085000 0.380000 0.810000 ;
      RECT 0.560000  0.350000 0.890000 0.810000 ;
      RECT 0.560000  2.300000 0.890000 2.980000 ;
      RECT 0.720000  0.810000 0.890000 1.320000 ;
      RECT 0.720000  1.320000 1.160000 1.650000 ;
      RECT 0.720000  1.650000 0.890000 2.300000 ;
      RECT 1.115000  1.820000 2.295000 1.990000 ;
      RECT 1.115000  1.990000 1.400000 2.980000 ;
      RECT 1.135000  0.350000 1.385000 0.980000 ;
      RECT 1.135000  0.980000 2.245000 1.150000 ;
      RECT 1.565000  0.085000 1.895000 0.790000 ;
      RECT 1.580000  2.160000 1.815000 3.245000 ;
      RECT 2.015000  1.990000 2.295000 2.905000 ;
      RECT 2.015000  2.905000 3.245000 3.075000 ;
      RECT 2.075000  0.350000 3.200000 0.600000 ;
      RECT 2.075000  0.600000 2.245000 0.980000 ;
      RECT 2.965000  1.820000 3.245000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__einvn_2
MACRO sky130_fd_sc_hs__einvn_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.035000 1.180000 5.155000 1.550000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.951000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.455000 1.780000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.550000 3.815000 1.720000 ;
        RECT 3.485000 1.720000 4.715000 1.890000 ;
        RECT 3.485000 1.890000 3.815000 2.735000 ;
        RECT 3.615000 0.770000 4.655000 1.010000 ;
        RECT 3.615000 1.010000 3.865000 1.130000 ;
        RECT 3.615000 1.130000 3.815000 1.550000 ;
        RECT 4.385000 1.890000 4.715000 2.735000 ;
        RECT 4.485000 0.595000 4.655000 0.770000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.280000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.245000 5.280000 3.415000 ;
      RECT 0.115000  0.085000 0.365000 1.130000 ;
      RECT 0.175000  1.950000 0.425000 3.245000 ;
      RECT 0.545000  0.300000 1.295000 1.130000 ;
      RECT 0.625000  1.130000 1.295000 1.310000 ;
      RECT 0.625000  1.310000 0.955000 2.980000 ;
      RECT 1.185000  1.480000 3.285000 1.650000 ;
      RECT 1.185000  1.650000 1.435000 2.980000 ;
      RECT 1.465000  0.350000 1.635000 1.140000 ;
      RECT 1.465000  1.140000 3.435000 1.310000 ;
      RECT 1.635000  1.820000 1.885000 3.245000 ;
      RECT 1.815000  0.085000 2.145000 0.970000 ;
      RECT 2.085000  1.650000 2.335000 2.980000 ;
      RECT 2.325000  0.350000 2.495000 1.140000 ;
      RECT 2.535000  1.820000 2.865000 3.245000 ;
      RECT 2.675000  0.085000 3.005000 0.970000 ;
      RECT 3.035000  1.650000 3.285000 2.905000 ;
      RECT 3.035000  2.905000 5.165000 3.075000 ;
      RECT 3.185000  0.255000 5.165000 0.425000 ;
      RECT 3.185000  0.425000 4.305000 0.600000 ;
      RECT 3.185000  0.600000 3.435000 1.140000 ;
      RECT 4.015000  2.060000 4.185000 2.905000 ;
      RECT 4.835000  0.425000 5.165000 1.010000 ;
      RECT 4.915000  1.820000 5.165000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
  END
END sky130_fd_sc_hs__einvn_4
MACRO sky130_fd_sc_hs__einvn_8
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  2.232000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.995000 1.350000 8.995000 1.780000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  1.623000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.435000 1.630000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  2.332400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925000 1.550000 5.725000 1.780000 ;
        RECT 5.455000 0.770000 6.645000 1.010000 ;
        RECT 5.455000 1.010000 8.505000 1.130000 ;
        RECT 5.455000 1.130000 5.725000 1.550000 ;
        RECT 5.555000 1.780000 5.725000 1.950000 ;
        RECT 5.555000 1.950000 8.555000 2.120000 ;
        RECT 5.555000 2.120000 5.725000 2.735000 ;
        RECT 6.315000 1.130000 8.505000 1.180000 ;
        RECT 6.425000 2.120000 6.755000 2.735000 ;
        RECT 7.325000 0.615000 7.495000 1.010000 ;
        RECT 7.325000 2.120000 7.655000 2.735000 ;
        RECT 8.175000 0.615000 8.505000 1.010000 ;
        RECT 8.225000 2.120000 8.555000 2.735000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.120000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.120000 0.085000 ;
      RECT 0.000000  3.245000 9.120000 3.415000 ;
      RECT 0.115000  1.820000 0.445000 3.245000 ;
      RECT 0.175000  0.085000 0.505000 0.990000 ;
      RECT 0.615000  1.130000 1.355000 1.335000 ;
      RECT 0.615000  1.335000 0.945000 2.980000 ;
      RECT 0.685000  0.325000 1.355000 1.130000 ;
      RECT 1.175000  1.665000 4.495000 1.835000 ;
      RECT 1.175000  1.835000 1.425000 2.980000 ;
      RECT 1.525000  0.350000 1.695000 1.300000 ;
      RECT 1.525000  1.300000 5.275000 1.380000 ;
      RECT 1.525000  1.380000 4.415000 1.470000 ;
      RECT 1.625000  2.005000 1.955000 3.245000 ;
      RECT 1.875000  0.085000 2.125000 1.130000 ;
      RECT 2.125000  1.835000 2.375000 2.980000 ;
      RECT 2.305000  0.350000 2.555000 1.300000 ;
      RECT 2.575000  2.005000 2.905000 3.245000 ;
      RECT 2.735000  0.085000 3.065000 1.130000 ;
      RECT 3.075000  1.835000 3.325000 2.980000 ;
      RECT 3.235000  0.350000 3.485000 1.300000 ;
      RECT 3.525000  2.005000 3.855000 3.245000 ;
      RECT 3.665000  0.085000 3.995000 1.130000 ;
      RECT 4.025000  1.835000 4.495000 1.950000 ;
      RECT 4.025000  1.950000 5.355000 2.120000 ;
      RECT 4.025000  2.120000 4.355000 2.980000 ;
      RECT 4.165000  0.350000 4.415000 1.210000 ;
      RECT 4.165000  1.210000 5.275000 1.300000 ;
      RECT 4.525000  2.290000 4.855000 3.245000 ;
      RECT 4.595000  0.085000 4.925000 1.040000 ;
      RECT 5.025000  2.120000 5.355000 2.905000 ;
      RECT 5.025000  2.905000 9.005000 3.075000 ;
      RECT 5.105000  0.255000 9.005000 0.425000 ;
      RECT 5.105000  0.425000 7.145000 0.600000 ;
      RECT 5.105000  0.600000 5.275000 1.210000 ;
      RECT 5.925000  2.290000 6.255000 2.905000 ;
      RECT 6.815000  0.600000 7.145000 0.825000 ;
      RECT 6.955000  2.290000 7.125000 2.905000 ;
      RECT 7.675000  0.425000 8.005000 0.825000 ;
      RECT 7.855000  2.290000 8.025000 2.905000 ;
      RECT 8.675000  0.425000 9.005000 1.130000 ;
      RECT 8.755000  1.950000 9.005000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
  END
END sky130_fd_sc_hs__einvn_8
MACRO sky130_fd_sc_hs__einvp_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.400000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945000 1.300000 2.275000 1.780000 ;
    END
  END A
  PIN TE
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.445000 1.440000 1.315000 1.780000 ;
    END
  END TE
  PIN Z
    ANTENNADIFFAREA  0.505900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.605000 0.960000 2.285000 1.130000 ;
        RECT 1.605000 1.130000 1.775000 1.950000 ;
        RECT 1.605000 1.950000 2.285000 2.275000 ;
        RECT 1.955000 0.350000 2.285000 0.960000 ;
        RECT 1.955000 2.275000 2.285000 2.980000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.400000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.400000 0.085000 ;
      RECT 0.000000  3.245000 2.400000 3.415000 ;
      RECT 0.105000  0.410000 0.940000 1.060000 ;
      RECT 0.105000  1.060000 0.275000 2.010000 ;
      RECT 0.105000  2.010000 0.880000 2.745000 ;
      RECT 0.105000  2.745000 0.890000 3.075000 ;
      RECT 1.085000  2.020000 1.415000 3.245000 ;
      RECT 1.135000  0.085000 1.420000 1.130000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
  END
END sky130_fd_sc_hs__einvp_1
MACRO sky130_fd_sc_hs__einvp_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.435000 1.550000 ;
    END
  END A
  PIN TE
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.480000 0.260000 2.810000 0.670000 ;
    END
  END TE
  PIN Z
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.180000 0.920000 2.735000 ;
        RECT 0.670000 0.625000 0.920000 1.180000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.115000  1.820000 0.365000 2.905000 ;
      RECT 0.115000  2.905000 1.265000 3.075000 ;
      RECT 0.160000  0.255000 1.270000 0.425000 ;
      RECT 0.160000  0.425000 0.490000 1.010000 ;
      RECT 1.095000  1.480000 2.165000 1.650000 ;
      RECT 1.095000  1.650000 1.265000 2.905000 ;
      RECT 1.100000  0.425000 1.270000 1.140000 ;
      RECT 1.100000  1.140000 2.210000 1.310000 ;
      RECT 1.450000  0.085000 1.780000 0.970000 ;
      RECT 1.465000  1.820000 1.715000 3.245000 ;
      RECT 1.915000  1.650000 2.165000 2.980000 ;
      RECT 1.950000  0.350000 2.210000 1.140000 ;
      RECT 2.415000  0.840000 2.800000 1.140000 ;
      RECT 2.415000  1.140000 2.745000 2.980000 ;
      RECT 2.915000  2.300000 3.245000 3.245000 ;
      RECT 2.980000  0.085000 3.245000 1.010000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__einvp_2
MACRO sky130_fd_sc_hs__einvp_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.430000 1.780000 ;
    END
  END A
  PIN TE
    ANTENNAGATEAREA  0.723000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.980000 1.300000 5.650000 1.630000 ;
        RECT 5.405000 1.180000 5.650000 1.300000 ;
    END
  END TE
  PIN Z
    ANTENNADIFFAREA  1.221900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.615000 0.660000 0.945000 1.010000 ;
        RECT 0.615000 1.010000 1.945000 1.180000 ;
        RECT 0.615000 1.950000 1.895000 2.120000 ;
        RECT 0.615000 2.120000 0.945000 2.735000 ;
        RECT 1.565000 2.120000 1.895000 2.735000 ;
        RECT 1.615000 0.660000 1.945000 1.010000 ;
        RECT 1.615000 1.180000 1.895000 1.950000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.115000  0.255000 2.445000 0.425000 ;
      RECT 0.115000  0.425000 0.445000 1.130000 ;
      RECT 0.115000  1.950000 0.445000 2.905000 ;
      RECT 0.115000  2.905000 2.395000 3.075000 ;
      RECT 1.115000  0.425000 1.445000 0.800000 ;
      RECT 1.115000  2.290000 1.365000 2.905000 ;
      RECT 2.065000  1.640000 4.175000 1.810000 ;
      RECT 2.065000  1.810000 2.395000 2.905000 ;
      RECT 2.115000  0.425000 2.445000 1.300000 ;
      RECT 2.115000  1.300000 4.445000 1.470000 ;
      RECT 2.565000  1.980000 2.815000 3.245000 ;
      RECT 2.615000  0.085000 2.945000 1.130000 ;
      RECT 3.015000  1.810000 3.265000 2.980000 ;
      RECT 3.115000  0.350000 3.445000 1.300000 ;
      RECT 3.465000  1.980000 3.725000 3.245000 ;
      RECT 3.615000  0.085000 3.945000 1.130000 ;
      RECT 3.925000  1.810000 4.175000 2.980000 ;
      RECT 4.115000  0.350000 4.445000 1.300000 ;
      RECT 4.395000  1.640000 4.785000 1.820000 ;
      RECT 4.395000  1.820000 5.195000 2.980000 ;
      RECT 4.395000  2.980000 4.785000 2.990000 ;
      RECT 4.615000  0.350000 5.005000 1.130000 ;
      RECT 4.615000  1.130000 4.785000 1.640000 ;
      RECT 5.175000  0.085000 5.505000 1.010000 ;
      RECT 5.395000  1.820000 5.645000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_hs__einvp_4
MACRO sky130_fd_sc_hs__einvp_8
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  2.232000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.410000 1.180000 3.460000 1.550000 ;
    END
  END A
  PIN TE
    ANTENNAGATEAREA  1.167000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.435000 1.180000 8.995000 1.410000 ;
        RECT 8.435000 1.410000 8.765000 1.550000 ;
    END
  END TE
  PIN Z
    ANTENNADIFFAREA  2.328200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.560000 1.720000 4.195000 1.890000 ;
        RECT 0.560000 1.890000 0.890000 2.735000 ;
        RECT 0.625000 0.615000 0.875000 0.840000 ;
        RECT 0.625000 0.840000 3.875000 1.010000 ;
        RECT 1.460000 1.890000 1.790000 2.735000 ;
        RECT 1.545000 0.615000 1.875000 0.840000 ;
        RECT 2.360000 1.890000 2.690000 2.735000 ;
        RECT 2.545000 0.615000 2.875000 0.840000 ;
        RECT 3.260000 1.890000 3.590000 2.735000 ;
        RECT 3.545000 0.595000 3.875000 0.840000 ;
        RECT 3.705000 1.010000 3.875000 1.550000 ;
        RECT 3.705000 1.550000 4.195000 1.720000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.120000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.120000 0.085000 ;
      RECT 0.000000  3.245000 9.120000 3.415000 ;
      RECT 0.110000  1.820000 0.375000 2.905000 ;
      RECT 0.110000  2.905000 3.960000 3.075000 ;
      RECT 0.115000  0.255000 4.225000 0.425000 ;
      RECT 0.115000  0.425000 0.445000 1.010000 ;
      RECT 1.045000  0.425000 1.375000 0.670000 ;
      RECT 1.070000  2.060000 1.275000 2.905000 ;
      RECT 1.970000  2.060000 2.190000 2.905000 ;
      RECT 2.045000  0.425000 2.375000 0.670000 ;
      RECT 2.875000  2.060000 3.075000 2.905000 ;
      RECT 3.045000  0.425000 3.375000 0.670000 ;
      RECT 3.790000  2.060000 4.940000 2.230000 ;
      RECT 3.790000  2.230000 3.960000 2.905000 ;
      RECT 4.055000  0.425000 4.225000 1.210000 ;
      RECT 4.055000  1.210000 7.885000 1.380000 ;
      RECT 4.160000  2.400000 4.490000 3.245000 ;
      RECT 4.405000  0.085000 4.735000 1.040000 ;
      RECT 4.690000  1.550000 7.560000 1.720000 ;
      RECT 4.690000  1.720000 4.940000 2.060000 ;
      RECT 4.690000  2.230000 4.940000 2.980000 ;
      RECT 4.905000  0.350000 5.155000 1.210000 ;
      RECT 5.140000  1.890000 5.310000 3.245000 ;
      RECT 5.335000  0.085000 5.665000 1.040000 ;
      RECT 5.510000  1.720000 5.760000 2.980000 ;
      RECT 5.845000  0.350000 6.015000 1.210000 ;
      RECT 5.960000  1.890000 6.210000 3.245000 ;
      RECT 6.195000  0.085000 6.525000 1.040000 ;
      RECT 6.410000  1.720000 6.660000 2.980000 ;
      RECT 6.705000  0.350000 6.955000 1.210000 ;
      RECT 6.860000  1.890000 7.110000 3.245000 ;
      RECT 7.125000  0.085000 7.455000 1.040000 ;
      RECT 7.310000  1.720000 7.560000 2.980000 ;
      RECT 7.635000  0.350000 7.885000 1.210000 ;
      RECT 7.775000  1.615000 8.225000 1.820000 ;
      RECT 7.775000  1.820000 8.565000 2.965000 ;
      RECT 8.055000  0.350000 8.505000 1.010000 ;
      RECT 8.055000  1.010000 8.225000 1.615000 ;
      RECT 8.235000  2.965000 8.565000 2.980000 ;
      RECT 8.675000  0.085000 8.935000 1.010000 ;
      RECT 8.765000  1.820000 9.015000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
  END
END sky130_fd_sc_hs__einvp_8
MACRO sky130_fd_sc_hs__fa_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.984000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.885000 1.220000 1.215000 1.540000 ;
        RECT 1.045000 0.920000 4.710000 0.935000 ;
        RECT 1.045000 0.935000 5.980000 1.090000 ;
        RECT 1.045000 1.090000 1.215000 1.220000 ;
        RECT 3.300000 1.090000 3.630000 1.455000 ;
        RECT 4.380000 1.090000 5.980000 1.105000 ;
        RECT 4.380000 1.105000 4.710000 1.455000 ;
        RECT 5.810000 1.105000 5.980000 1.320000 ;
        RECT 5.810000 1.320000 6.210000 1.575000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.984000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.800000 1.320000 7.470000 1.780000 ;
    END
  END B
  PIN CIN
    ANTENNAPARTIALMETALSIDEAREA  2.604000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.535000 1.550000 1.825000 1.595000 ;
        RECT 1.535000 1.595000 5.185000 1.735000 ;
        RECT 1.535000 1.735000 1.825000 1.780000 ;
        RECT 3.935000 1.550000 4.225000 1.595000 ;
        RECT 3.935000 1.735000 4.225000 1.780000 ;
        RECT 4.895000 1.550000 5.185000 1.595000 ;
        RECT 4.895000 1.735000 5.185000 1.780000 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  0.519000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.210000 0.350000 8.540000 1.130000 ;
        RECT 8.285000 1.130000 8.540000 2.980000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.530100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.350000 0.365000 1.130000 ;
        RECT 0.085000 1.130000 0.255000 1.820000 ;
        RECT 0.085000 1.820000 0.355000 2.980000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
      RECT 0.000000  3.245000 8.640000 3.415000 ;
      RECT 0.425000  1.300000 0.705000 1.630000 ;
      RECT 0.535000  0.580000 2.270000 0.750000 ;
      RECT 0.535000  0.750000 0.705000 1.300000 ;
      RECT 0.535000  1.630000 0.705000 1.710000 ;
      RECT 0.535000  1.710000 1.225000 1.880000 ;
      RECT 0.555000  2.050000 0.885000 3.245000 ;
      RECT 0.625000  0.085000 0.980000 0.410000 ;
      RECT 1.055000  1.880000 1.225000 1.950000 ;
      RECT 1.055000  1.950000 2.410000 2.120000 ;
      RECT 1.565000  1.260000 2.115000 1.575000 ;
      RECT 1.565000  1.575000 1.795000 1.780000 ;
      RECT 1.940000  0.355000 2.270000 0.580000 ;
      RECT 2.080000  1.745000 2.410000 1.950000 ;
      RECT 2.080000  2.120000 2.410000 2.755000 ;
      RECT 2.325000  1.260000 2.750000 1.575000 ;
      RECT 2.480000  0.420000 2.890000 0.580000 ;
      RECT 2.480000  0.580000 3.910000 0.750000 ;
      RECT 2.580000  1.575000 2.750000 1.625000 ;
      RECT 2.580000  1.625000 3.200000 1.795000 ;
      RECT 2.610000  1.965000 2.860000 2.290000 ;
      RECT 2.610000  2.290000 3.930000 2.460000 ;
      RECT 2.610000  2.460000 2.860000 2.755000 ;
      RECT 3.030000  1.795000 3.200000 1.950000 ;
      RECT 3.030000  1.950000 5.495000 2.120000 ;
      RECT 3.070000  0.085000 3.400000 0.410000 ;
      RECT 3.080000  2.630000 3.410000 3.245000 ;
      RECT 3.580000  0.420000 3.910000 0.580000 ;
      RECT 3.600000  2.460000 3.930000 2.755000 ;
      RECT 3.840000  1.260000 4.195000 1.780000 ;
      RECT 4.080000  0.085000 4.555000 0.710000 ;
      RECT 4.105000  2.305000 4.435000 3.245000 ;
      RECT 4.925000  1.275000 5.640000 1.575000 ;
      RECT 4.925000  1.575000 5.155000 1.780000 ;
      RECT 5.045000  0.435000 5.375000 0.595000 ;
      RECT 5.045000  0.595000 6.320000 0.765000 ;
      RECT 5.070000  2.120000 5.495000 2.755000 ;
      RECT 5.325000  1.745000 6.550000 1.915000 ;
      RECT 5.325000  1.915000 5.495000 1.950000 ;
      RECT 5.555000  0.255000 6.660000 0.425000 ;
      RECT 5.665000  2.085000 7.320000 2.255000 ;
      RECT 5.665000  2.255000 5.950000 2.755000 ;
      RECT 6.120000  2.500000 6.825000 3.245000 ;
      RECT 6.150000  0.765000 6.320000 0.980000 ;
      RECT 6.150000  0.980000 8.040000 1.150000 ;
      RECT 6.380000  1.150000 6.550000 1.745000 ;
      RECT 6.490000  0.425000 6.660000 0.640000 ;
      RECT 6.490000  0.640000 7.590000 0.810000 ;
      RECT 6.830000  0.085000 7.080000 0.470000 ;
      RECT 6.990000  1.950000 7.320000 2.085000 ;
      RECT 7.000000  2.255000 7.320000 2.830000 ;
      RECT 7.260000  0.480000 7.590000 0.640000 ;
      RECT 7.710000  1.150000 8.040000 1.550000 ;
      RECT 7.755000  1.820000 8.085000 3.245000 ;
      RECT 7.780000  0.085000 8.030000 0.770000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  1.580000 1.765000 1.750000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  1.580000 4.165000 1.750000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  1.580000 5.125000 1.750000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
  END
END sky130_fd_sc_hs__fa_1
MACRO sky130_fd_sc_hs__fa_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAPARTIALMETALSIDEAREA  4.683000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.095000 1.550000 0.385000 1.595000 ;
        RECT 0.095000 1.595000 6.625000 1.735000 ;
        RECT 0.095000 1.735000 0.385000 1.780000 ;
        RECT 2.495000 1.550000 2.785000 1.595000 ;
        RECT 2.495000 1.735000 2.785000 1.780000 ;
        RECT 3.935000 1.550000 4.225000 1.595000 ;
        RECT 3.935000 1.735000 4.225000 1.780000 ;
        RECT 6.335000 1.550000 6.625000 1.595000 ;
        RECT 6.335000 1.735000 6.625000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.044000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.920000 0.835000 2.150000 ;
        RECT 0.665000 1.245000 1.165000 1.575000 ;
        RECT 0.665000 1.575000 0.835000 1.920000 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.783000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.715000 1.260000 2.225000 1.575000 ;
        RECT 2.055000 1.575000 2.225000 1.950000 ;
        RECT 2.055000 1.950000 4.535000 2.105000 ;
        RECT 2.055000 2.105000 4.195000 2.120000 ;
        RECT 3.215000 1.260000 3.545000 1.575000 ;
        RECT 3.375000 1.575000 3.545000 1.935000 ;
        RECT 3.375000 1.935000 4.535000 1.950000 ;
        RECT 3.375000 2.120000 4.195000 2.150000 ;
        RECT 4.365000 1.745000 5.635000 1.915000 ;
        RECT 4.365000 1.915000 4.535000 1.935000 ;
        RECT 5.305000 1.260000 5.635000 1.745000 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  0.649600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.985000 1.820000 7.555000 2.150000 ;
        RECT 7.105000 0.915000 7.555000 1.085000 ;
        RECT 7.385000 1.085000 7.555000 1.820000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.220000 1.820000 8.575000 2.980000 ;
        RECT 8.245000 0.375000 8.575000 1.150000 ;
        RECT 8.405000 1.150000 8.575000 1.820000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.120000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.120000 0.085000 ;
      RECT 0.000000  3.245000 9.120000 3.415000 ;
      RECT 0.095000  1.950000 0.425000 2.320000 ;
      RECT 0.095000  2.320000 1.545000 2.490000 ;
      RECT 0.095000  2.490000 0.445000 2.910000 ;
      RECT 0.105000  1.300000 0.435000 1.780000 ;
      RECT 0.115000  0.375000 0.445000 0.905000 ;
      RECT 0.115000  0.905000 1.205000 1.075000 ;
      RECT 0.115000  1.075000 0.445000 1.130000 ;
      RECT 0.615000  0.085000 0.865000 0.735000 ;
      RECT 0.615000  2.660000 1.010000 3.245000 ;
      RECT 1.035000  0.420000 1.810000 0.750000 ;
      RECT 1.035000  0.750000 1.205000 0.905000 ;
      RECT 1.215000  2.085000 1.545000 2.320000 ;
      RECT 1.215000  2.490000 1.545000 2.755000 ;
      RECT 1.375000  0.920000 6.935000 1.090000 ;
      RECT 1.375000  1.090000 1.545000 1.745000 ;
      RECT 1.375000  1.745000 1.885000 1.915000 ;
      RECT 1.715000  1.915000 1.885000 2.290000 ;
      RECT 1.715000  2.290000 2.185000 2.620000 ;
      RECT 1.980000  0.375000 2.310000 0.920000 ;
      RECT 2.525000  1.260000 3.005000 1.575000 ;
      RECT 2.525000  1.575000 2.755000 1.780000 ;
      RECT 2.800000  0.085000 3.310000 0.705000 ;
      RECT 2.825000  2.290000 3.155000 3.245000 ;
      RECT 3.405000  2.320000 4.825000 2.490000 ;
      RECT 3.405000  2.490000 3.735000 2.755000 ;
      RECT 3.480000  0.375000 3.810000 0.580000 ;
      RECT 3.480000  0.580000 4.970000 0.750000 ;
      RECT 3.905000  2.660000 4.290000 3.245000 ;
      RECT 3.965000  1.260000 4.525000 1.575000 ;
      RECT 3.965000  1.575000 4.195000 1.765000 ;
      RECT 3.990000  0.085000 4.320000 0.410000 ;
      RECT 4.495000  2.275000 4.825000 2.320000 ;
      RECT 4.495000  2.490000 4.825000 2.755000 ;
      RECT 4.500000  0.420000 4.970000 0.580000 ;
      RECT 4.765000  1.090000 5.095000 1.575000 ;
      RECT 5.005000  2.085000 5.335000 2.320000 ;
      RECT 5.005000  2.320000 8.050000 2.490000 ;
      RECT 5.005000  2.490000 5.335000 2.755000 ;
      RECT 5.140000  0.375000 5.470000 0.575000 ;
      RECT 5.140000  0.575000 8.050000 0.745000 ;
      RECT 5.140000  0.745000 5.470000 0.750000 ;
      RECT 6.265000  1.350000 6.595000 1.780000 ;
      RECT 6.470000  0.085000 6.925000 0.405000 ;
      RECT 6.535000  2.660000 6.865000 3.245000 ;
      RECT 6.765000  1.090000 6.935000 1.255000 ;
      RECT 6.765000  1.255000 7.165000 1.585000 ;
      RECT 7.530000  2.730000 8.050000 3.245000 ;
      RECT 7.615000  0.085000 8.065000 0.405000 ;
      RECT 7.880000  0.745000 8.050000 1.320000 ;
      RECT 7.880000  1.320000 8.235000 1.650000 ;
      RECT 7.880000  1.650000 8.050000 2.320000 ;
      RECT 8.750000  1.820000 9.000000 3.245000 ;
      RECT 8.755000  0.085000 9.005000 1.155000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  1.580000 0.325000 1.750000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  1.580000 2.725000 1.750000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  1.580000 4.165000 1.750000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  1.580000 6.565000 1.750000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
  END
END sky130_fd_sc_hs__fa_2
MACRO sky130_fd_sc_hs__fa_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.044000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.245000 0.835000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.044000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.345000 1.260000 1.835000 1.575000 ;
        RECT 1.665000 1.575000 1.835000 1.950000 ;
        RECT 1.665000 1.950000 2.650000 2.120000 ;
        RECT 2.480000 1.245000 2.810000 1.745000 ;
        RECT 2.480000 1.745000 6.595000 1.780000 ;
        RECT 2.480000 1.780000 6.085000 1.890000 ;
        RECT 2.480000 1.890000 4.620000 1.915000 ;
        RECT 2.480000 1.915000 2.650000 1.950000 ;
        RECT 3.950000 1.260000 4.280000 1.745000 ;
        RECT 4.450000 1.720000 6.595000 1.745000 ;
        RECT 5.915000 1.260000 6.340000 1.550000 ;
        RECT 5.915000 1.550000 6.595000 1.720000 ;
    END
  END B
  PIN CIN
    ANTENNAPARTIALMETALSIDEAREA  2.604000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2.015000 1.180000 2.305000 1.225000 ;
        RECT 2.015000 1.225000 5.665000 1.365000 ;
        RECT 2.015000 1.365000 2.305000 1.410000 ;
        RECT 2.975000 1.180000 3.265000 1.225000 ;
        RECT 2.975000 1.365000 3.265000 1.410000 ;
        RECT 5.375000 1.180000 5.665000 1.225000 ;
        RECT 5.375000 1.365000 5.665000 1.410000 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  9.145000 1.820000 10.435000 1.990000 ;
        RECT  9.145000 1.990000  9.475000 2.980000 ;
        RECT  9.305000 0.390000  9.555000 0.980000 ;
        RECT  9.305000 0.980000 10.425000 1.150000 ;
        RECT 10.095000 1.990000 10.435000 2.980000 ;
        RECT 10.165000 0.390000 10.425000 0.980000 ;
        RECT 10.165000 1.150000 10.425000 1.550000 ;
        RECT 10.165000 1.550000 10.435000 1.820000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.245000 1.840000 8.525000 2.010000 ;
        RECT 7.245000 2.010000 7.575000 2.980000 ;
        RECT 7.265000 0.920000 8.615000 1.170000 ;
        RECT 8.195000 2.010000 8.525000 2.980000 ;
        RECT 8.285000 1.170000 8.525000 1.840000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.040000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 11.040000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  3.245000 11.040000 3.415000 ;
      RECT  0.115000  0.350000  0.445000 0.580000 ;
      RECT  0.115000  0.580000  1.965000 0.670000 ;
      RECT  0.115000  0.670000  1.495000 0.750000 ;
      RECT  0.115000  0.750000  0.445000 1.075000 ;
      RECT  0.115000  1.950000  0.445000 2.085000 ;
      RECT  0.115000  2.085000  1.155000 2.255000 ;
      RECT  0.115000  2.255000  0.445000 2.980000 ;
      RECT  0.625000  0.085000  1.155000 0.410000 ;
      RECT  0.645000  2.425000  0.815000 3.245000 ;
      RECT  0.985000  2.255000  1.155000 2.630000 ;
      RECT  0.985000  2.630000  2.005000 2.960000 ;
      RECT  1.005000  0.920000  5.255000 1.010000 ;
      RECT  1.005000  1.010000  1.835000 1.090000 ;
      RECT  1.005000  1.090000  1.175000 1.745000 ;
      RECT  1.005000  1.745000  1.495000 1.915000 ;
      RECT  1.325000  0.350000  1.965000 0.580000 ;
      RECT  1.325000  1.915000  1.495000 2.290000 ;
      RECT  1.325000  2.290000  2.540000 2.460000 ;
      RECT  1.665000  0.840000  3.555000 0.920000 ;
      RECT  2.005000  1.180000  2.275000 1.780000 ;
      RECT  2.135000  0.350000  2.465000 0.840000 ;
      RECT  2.210000  2.460000  2.540000 2.755000 ;
      RECT  3.005000  1.180000  3.215000 1.260000 ;
      RECT  3.005000  1.260000  3.740000 1.575000 ;
      RECT  3.170000  2.085000  3.500000 3.245000 ;
      RECT  3.175000  0.085000  3.505000 0.670000 ;
      RECT  3.385000  1.010000  5.255000 1.090000 ;
      RECT  3.670000  2.085000  5.070000 2.255000 ;
      RECT  3.670000  2.255000  4.000000 2.755000 ;
      RECT  3.725000  0.350000  3.975000 0.580000 ;
      RECT  3.725000  0.580000  4.915000 0.750000 ;
      RECT  4.155000  0.085000  4.485000 0.410000 ;
      RECT  4.170000  2.425000  4.570000 3.245000 ;
      RECT  4.665000  0.350000  4.915000 0.580000 ;
      RECT  4.740000  2.255000  5.070000 2.755000 ;
      RECT  4.930000  1.090000  5.255000 1.220000 ;
      RECT  4.930000  1.220000  5.260000 1.550000 ;
      RECT  5.085000  0.255000  6.425000 0.425000 ;
      RECT  5.085000  0.425000  5.255000 0.920000 ;
      RECT  5.240000  2.060000  7.075000 2.120000 ;
      RECT  5.240000  2.120000  6.425000 2.230000 ;
      RECT  5.240000  2.230000  5.570000 2.755000 ;
      RECT  5.425000  0.595000  5.675000 0.840000 ;
      RECT  5.425000  0.840000  6.085000 0.920000 ;
      RECT  5.425000  0.920000  7.075000 1.010000 ;
      RECT  5.430000  1.180000  5.745000 1.550000 ;
      RECT  5.915000  1.010000  7.075000 1.090000 ;
      RECT  6.255000  0.425000  6.425000 0.580000 ;
      RECT  6.255000  0.580000  9.135000 0.750000 ;
      RECT  6.255000  1.950000  7.075000 2.060000 ;
      RECT  6.755000  0.085000  7.085000 0.410000 ;
      RECT  6.795000  2.290000  7.045000 3.245000 ;
      RECT  6.905000  1.090000  7.075000 1.340000 ;
      RECT  6.905000  1.340000  8.105000 1.670000 ;
      RECT  6.905000  1.670000  7.075000 1.950000 ;
      RECT  7.775000  0.085000  8.105000 0.410000 ;
      RECT  7.775000  2.180000  8.025000 3.245000 ;
      RECT  8.725000  1.820000  8.975000 3.245000 ;
      RECT  8.795000  0.085000  9.125000 0.410000 ;
      RECT  8.965000  0.750000  9.135000 1.320000 ;
      RECT  8.965000  1.320000  9.955000 1.650000 ;
      RECT  9.675000  2.160000  9.925000 3.245000 ;
      RECT  9.735000  0.085000  9.985000 0.810000 ;
      RECT 10.595000  0.085000 10.925000 1.170000 ;
      RECT 10.625000  1.820000 10.875000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  1.210000  2.245000 1.380000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  1.210000  3.205000 1.380000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  1.210000  5.605000 1.380000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
  END
END sky130_fd_sc_hs__fa_4
MACRO sky130_fd_sc_hs__fah_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.92000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAPARTIALMETALSIDEAREA  0.132000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.820000 1.470000 13.490000 1.800000 ;
    END
  END A
  PIN B
    ANTENNAPARTIALMETALSIDEAREA  0.072000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.145000 1.180000 9.475000 1.550000 ;
    END
  END B
  PIN CI
    ANTENNAPARTIALMETALSIDEAREA  0.072000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.410000 1.335000 1.780000 ;
    END
  END CI
  PIN COUT
    ANTENNADIFFAREA  0.674850 ;
    ANTENNAPARTIALMETALSIDEAREA  1.117000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.665000 0.730000 1.675000 0.900000 ;
        RECT 0.665000 0.900000 0.835000 1.950000 ;
        RECT 0.665000 1.950000 1.155000 2.120000 ;
        RECT 0.985000 2.120000 1.155000 2.905000 ;
        RECT 0.985000 2.905000 2.645000 3.075000 ;
        RECT 1.505000 0.400000 2.075000 0.730000 ;
        RECT 2.315000 2.875000 2.645000 2.905000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.537600 ;
    ANTENNAPARTIALMETALSIDEAREA  0.215000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 0.540000 0.445000 2.980000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 13.920000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 13.920000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.920000 0.085000 ;
      RECT  0.000000  3.245000 13.920000 3.415000 ;
      RECT  0.620000  0.085000  0.950000 0.560000 ;
      RECT  0.645000  2.290000  0.815000 3.245000 ;
      RECT  1.130000  1.070000  1.675000 1.240000 ;
      RECT  1.325000  1.950000  1.675000 2.535000 ;
      RECT  1.325000  2.535000  2.985000 2.625000 ;
      RECT  1.325000  2.625000  3.630000 2.705000 ;
      RECT  1.325000  2.705000  1.675000 2.735000 ;
      RECT  1.505000  1.240000  1.675000 1.950000 ;
      RECT  1.845000  0.900000  2.765000 1.070000 ;
      RECT  1.845000  1.070000  2.175000 2.195000 ;
      RECT  1.845000  2.195000  3.325000 2.285000 ;
      RECT  1.845000  2.285000  4.535000 2.365000 ;
      RECT  2.255000  0.085000  2.425000 0.730000 ;
      RECT  2.500000  1.240000  3.105000 1.410000 ;
      RECT  2.500000  1.410000  2.830000 1.635000 ;
      RECT  2.595000  0.255000  4.285000 0.425000 ;
      RECT  2.595000  0.425000  2.765000 0.900000 ;
      RECT  2.815000  2.705000  3.630000 2.795000 ;
      RECT  2.935000  0.595000  3.945000 0.765000 ;
      RECT  2.935000  0.765000  3.105000 1.240000 ;
      RECT  2.935000  2.965000  3.290000 3.245000 ;
      RECT  3.005000  1.580000  3.445000 1.855000 ;
      RECT  3.005000  1.855000  4.000000 2.025000 ;
      RECT  3.155000  2.365000  4.535000 2.455000 ;
      RECT  3.275000  0.935000  3.605000 1.185000 ;
      RECT  3.275000  1.185000  3.445000 1.580000 ;
      RECT  3.460000  2.795000  3.630000 2.905000 ;
      RECT  3.460000  2.905000  7.000000 3.075000 ;
      RECT  3.495000  2.025000  4.000000 2.115000 ;
      RECT  3.670000  1.435000  4.340000 1.595000 ;
      RECT  3.670000  1.595000  4.875000 1.685000 ;
      RECT  3.775000  0.765000  3.945000 1.095000 ;
      RECT  3.775000  1.095000  5.215000 1.265000 ;
      RECT  4.115000  0.425000  4.285000 0.755000 ;
      RECT  4.115000  0.755000  6.215000 0.765000 ;
      RECT  4.115000  0.765000  5.045000 0.925000 ;
      RECT  4.170000  1.685000  4.875000 1.765000 ;
      RECT  4.205000  2.100000  4.535000 2.285000 ;
      RECT  4.205000  2.455000  4.535000 2.735000 ;
      RECT  4.455000  0.255000  7.565000 0.425000 ;
      RECT  4.455000  0.425000  4.705000 0.585000 ;
      RECT  4.705000  1.765000  4.875000 2.730000 ;
      RECT  4.705000  2.730000  6.125000 2.905000 ;
      RECT  4.875000  0.595000  6.215000 0.755000 ;
      RECT  4.880000  1.265000  5.215000 1.425000 ;
      RECT  5.045000  1.425000  5.215000 2.320000 ;
      RECT  5.045000  2.320000  6.660000 2.490000 ;
      RECT  5.385000  0.935000  5.715000 1.035000 ;
      RECT  5.385000  1.035000  6.225000 1.205000 ;
      RECT  5.405000  1.375000  5.885000 1.705000 ;
      RECT  5.405000  1.705000  5.635000 2.150000 ;
      RECT  5.885000  0.765000  6.215000 0.865000 ;
      RECT  6.055000  1.205000  6.225000 1.950000 ;
      RECT  6.055000  1.950000  7.000000 2.120000 ;
      RECT  6.330000  2.290000  6.660000 2.320000 ;
      RECT  6.330000  2.490000  6.660000 2.640000 ;
      RECT  6.395000  0.670000  6.565000 1.550000 ;
      RECT  6.395000  1.550000  6.595000 1.780000 ;
      RECT  6.735000  0.710000  7.065000 1.380000 ;
      RECT  6.830000  2.120000  7.000000 2.905000 ;
      RECT  6.845000  1.380000  7.065000 1.550000 ;
      RECT  6.845000  1.550000  7.075000 1.780000 ;
      RECT  7.170000  1.950000  7.500000 2.925000 ;
      RECT  7.235000  0.425000  7.565000 0.620000 ;
      RECT  7.235000  0.620000 10.315000 0.790000 ;
      RECT  7.235000  0.790000  7.565000 1.130000 ;
      RECT  7.330000  1.130000  7.500000 1.950000 ;
      RECT  7.670000  1.765000  8.000000 3.245000 ;
      RECT  7.745000  0.085000  8.075000 0.450000 ;
      RECT  8.170000  0.960000  8.635000 1.210000 ;
      RECT  8.170000  1.210000  8.340000 1.880000 ;
      RECT  8.170000  1.880000  8.610000 2.905000 ;
      RECT  8.170000  2.905000 11.740000 3.075000 ;
      RECT  8.510000  1.380000  8.975000 1.710000 ;
      RECT  8.780000  1.880000  9.110000 2.565000 ;
      RECT  8.780000  2.565000 10.815000 2.735000 ;
      RECT  8.805000  0.790000  8.975000 1.380000 ;
      RECT  8.895000  0.255000 11.155000 0.425000 ;
      RECT  8.895000  0.425000  9.385000 0.450000 ;
      RECT  9.280000  1.805000 10.475000 2.395000 ;
      RECT  9.645000  0.960000  9.975000 1.805000 ;
      RECT 10.145000  0.790000 10.315000 1.220000 ;
      RECT 10.145000  1.220000 10.475000 1.550000 ;
      RECT 10.485000  0.595000 10.815000 1.050000 ;
      RECT 10.645000  1.050000 10.815000 2.565000 ;
      RECT 10.985000  0.425000 11.155000 1.550000 ;
      RECT 10.985000  1.550000 11.215000 1.780000 ;
      RECT 10.985000  1.780000 11.155000 2.735000 ;
      RECT 11.385000  1.130000 11.740000 2.905000 ;
      RECT 11.405000  0.350000 11.740000 1.130000 ;
      RECT 11.910000  0.790000 12.805000 0.960000 ;
      RECT 11.910000  0.960000 12.080000 1.720000 ;
      RECT 11.910000  1.720000 12.650000 1.940000 ;
      RECT 11.915000  0.085000 12.245000 0.620000 ;
      RECT 11.950000  2.110000 12.220000 2.330000 ;
      RECT 11.950000  2.330000 12.290000 3.245000 ;
      RECT 12.250000  1.130000 13.830000 1.300000 ;
      RECT 12.250000  1.300000 12.580000 1.550000 ;
      RECT 12.390000  1.940000 12.650000 1.970000 ;
      RECT 12.390000  1.970000 12.850000 2.160000 ;
      RECT 12.475000  0.350000 12.805000 0.790000 ;
      RECT 12.520000  2.160000 12.850000 2.980000 ;
      RECT 12.975000  0.085000 13.305000 0.960000 ;
      RECT 13.050000  1.970000 13.300000 3.245000 ;
      RECT 13.470000  1.970000 13.830000 2.980000 ;
      RECT 13.475000  0.350000 13.830000 1.130000 ;
      RECT 13.660000  1.300000 13.830000 1.970000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  1.580000  3.205000 1.750000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  1.950000  5.605000 2.120000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  1.580000  6.565000 1.750000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  1.580000  7.045000 1.750000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  8.840000  1.950000  9.010000 2.120000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT  9.885000  1.950000 10.055000 2.120000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.245000  1.950000 10.415000 2.120000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.015000  1.580000 11.185000 1.750000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.435000  1.950000 12.605000 2.120000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
    LAYER met1 ;
      RECT  2.975000 1.550000  3.265000 1.595000 ;
      RECT  2.975000 1.595000  6.625000 1.735000 ;
      RECT  2.975000 1.735000  3.265000 1.780000 ;
      RECT  5.375000 1.920000  5.665000 1.965000 ;
      RECT  5.375000 1.965000  9.070000 2.105000 ;
      RECT  5.375000 2.105000  5.665000 2.150000 ;
      RECT  6.335000 1.550000  6.625000 1.595000 ;
      RECT  6.335000 1.735000  6.625000 1.780000 ;
      RECT  6.815000 1.550000  7.105000 1.595000 ;
      RECT  6.815000 1.595000 11.245000 1.735000 ;
      RECT  6.815000 1.735000  7.105000 1.780000 ;
      RECT  8.780000 1.920000  9.070000 1.965000 ;
      RECT  8.780000 2.105000  9.070000 2.150000 ;
      RECT  9.825000 1.920000 10.475000 1.965000 ;
      RECT  9.825000 1.965000 12.665000 2.105000 ;
      RECT  9.825000 2.105000 10.475000 2.150000 ;
      RECT 10.955000 1.550000 11.245000 1.595000 ;
      RECT 10.955000 1.735000 11.245000 1.780000 ;
      RECT 12.375000 1.920000 12.665000 1.965000 ;
      RECT 12.375000 2.105000 12.665000 2.150000 ;
  END
END sky130_fd_sc_hs__fah_1
MACRO sky130_fd_sc_hs__fah_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.40000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.290000 2.045000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.723000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555000 1.355000 2.895000 2.150000 ;
        RECT 2.725000 0.595000 5.435000 0.765000 ;
        RECT 2.725000 0.765000 2.895000 1.355000 ;
        RECT 3.440000 1.630000 3.770000 1.960000 ;
        RECT 3.565000 0.765000 3.735000 1.630000 ;
        RECT 4.405000 0.765000 4.595000 1.605000 ;
        RECT 5.265000 0.765000 5.435000 0.920000 ;
        RECT 5.265000 0.920000 6.205000 1.090000 ;
        RECT 5.875000 1.090000 6.205000 1.185000 ;
    END
  END B
  PIN CI
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.450000 1.450000 11.875000 1.780000 ;
    END
  END CI
  PIN COUT
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.585000 0.350000 12.835000 1.550000 ;
        RECT 12.585000 1.550000 12.920000 2.200000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.561800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.515000 0.355000 13.785000 0.800000 ;
        RECT 13.515000 0.800000 14.275000 1.130000 ;
        RECT 13.570000 1.820000 13.875000 2.980000 ;
        RECT 13.705000 1.130000 14.275000 1.505000 ;
        RECT 13.705000 1.505000 13.875000 1.820000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 14.400000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 14.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.400000 0.085000 ;
      RECT  0.000000  3.245000 14.400000 3.415000 ;
      RECT  0.105000  2.160000  0.360000 3.245000 ;
      RECT  0.125000  1.180000  0.650000 1.470000 ;
      RECT  0.170000  0.085000  0.535000 0.790000 ;
      RECT  0.335000  1.470000  0.650000 1.820000 ;
      RECT  0.335000  1.820000  0.885000 1.990000 ;
      RECT  0.480000  0.960000  0.965000 1.130000 ;
      RECT  0.480000  1.130000  0.650000 1.180000 ;
      RECT  0.555000  1.990000  0.885000 2.980000 ;
      RECT  0.705000  0.350000  0.965000 0.960000 ;
      RECT  0.820000  1.300000  1.395000 1.630000 ;
      RECT  1.090000  1.630000  1.340000 2.980000 ;
      RECT  1.225000  0.505000  1.705000 1.120000 ;
      RECT  1.225000  1.120000  1.395000 1.300000 ;
      RECT  1.540000  1.950000  1.870000 3.245000 ;
      RECT  1.875000  0.085000  2.125000 0.845000 ;
      RECT  2.055000  2.015000  2.385000 2.890000 ;
      RECT  2.055000  2.890000  6.055000 3.060000 ;
      RECT  2.215000  1.015000  2.555000 1.185000 ;
      RECT  2.215000  1.185000  2.385000 2.015000 ;
      RECT  2.305000  0.255000  5.935000 0.425000 ;
      RECT  2.305000  0.425000  2.555000 1.015000 ;
      RECT  2.555000  2.390000  3.450000 2.550000 ;
      RECT  2.555000  2.550000  5.555000 2.720000 ;
      RECT  3.065000  0.935000  3.395000 1.185000 ;
      RECT  3.065000  1.185000  3.235000 2.390000 ;
      RECT  3.620000  2.130000  4.110000 2.380000 ;
      RECT  3.905000  0.935000  4.235000 1.185000 ;
      RECT  3.940000  1.185000  4.235000 1.410000 ;
      RECT  3.940000  1.410000  4.110000 2.130000 ;
      RECT  4.280000  2.100000  5.215000 2.350000 ;
      RECT  4.765000  0.935000  5.095000 1.260000 ;
      RECT  4.765000  1.260000  5.705000 1.355000 ;
      RECT  4.765000  1.355000  6.545000 1.430000 ;
      RECT  4.765000  1.430000  4.935000 2.100000 ;
      RECT  5.105000  1.600000  5.365000 1.760000 ;
      RECT  5.105000  1.760000  7.045000 1.930000 ;
      RECT  5.385000  2.100000  6.395000 2.240000 ;
      RECT  5.385000  2.240000  7.385000 2.270000 ;
      RECT  5.385000  2.270000  5.555000 2.550000 ;
      RECT  5.535000  1.430000  6.545000 1.525000 ;
      RECT  5.605000  0.425000  5.935000 0.750000 ;
      RECT  5.725000  2.440000  6.055000 2.890000 ;
      RECT  6.225000  2.270000  7.385000 2.410000 ;
      RECT  6.265000  2.580000  6.595000 3.245000 ;
      RECT  6.335000  0.085000  6.665000 0.680000 ;
      RECT  6.375000  0.850000  7.005000 1.020000 ;
      RECT  6.375000  1.020000  6.545000 1.355000 ;
      RECT  6.715000  1.190000  7.505000 1.360000 ;
      RECT  6.715000  1.360000  7.045000 1.760000 ;
      RECT  6.715000  1.930000  7.045000 2.070000 ;
      RECT  6.835000  0.255000  7.845000 0.425000 ;
      RECT  6.835000  0.425000  7.005000 0.850000 ;
      RECT  7.175000  0.630000  7.505000 1.190000 ;
      RECT  7.215000  1.630000  7.505000 1.960000 ;
      RECT  7.215000  1.960000  7.385000 2.240000 ;
      RECT  7.215000  2.410000  7.385000 2.905000 ;
      RECT  7.215000  2.905000  9.575000 3.075000 ;
      RECT  7.555000  2.130000  8.310000 2.735000 ;
      RECT  7.675000  0.425000  7.845000 1.275000 ;
      RECT  7.675000  1.275000  7.970000 1.945000 ;
      RECT  8.015000  0.390000  8.555000 0.640000 ;
      RECT  8.140000  0.640000  8.555000 1.040000 ;
      RECT  8.140000  1.040000  8.310000 2.130000 ;
      RECT  8.480000  1.225000  8.735000 2.905000 ;
      RECT  8.745000  0.255000 10.935000 0.425000 ;
      RECT  8.745000  0.425000  9.075000 1.055000 ;
      RECT  8.905000  1.055000  9.075000 2.130000 ;
      RECT  8.905000  2.130000  9.235000 2.735000 ;
      RECT  9.245000  0.595000 10.255000 0.765000 ;
      RECT  9.245000  0.765000  9.415000 1.630000 ;
      RECT  9.245000  1.630000  9.575000 1.960000 ;
      RECT  9.405000  1.960000  9.575000 2.905000 ;
      RECT  9.585000  0.935000  9.915000 1.185000 ;
      RECT  9.745000  1.185000  9.915000 2.100000 ;
      RECT  9.745000  2.100000 10.075000 2.600000 ;
      RECT  9.745000  2.600000 11.970000 2.770000 ;
      RECT  9.745000  2.770000 10.075000 2.980000 ;
      RECT 10.085000  0.765000 10.255000 1.355000 ;
      RECT 10.085000  1.355000 10.470000 1.685000 ;
      RECT 10.310000  2.130000 10.810000 2.430000 ;
      RECT 10.425000  0.595000 10.595000 1.015000 ;
      RECT 10.425000  1.015000 10.810000 1.185000 ;
      RECT 10.640000  1.185000 10.810000 2.130000 ;
      RECT 10.765000  0.425000 10.935000 0.675000 ;
      RECT 10.765000  0.675000 11.865000 0.845000 ;
      RECT 10.980000  0.845000 11.865000 1.055000 ;
      RECT 10.980000  1.055000 11.240000 1.950000 ;
      RECT 10.980000  1.950000 11.930000 2.200000 ;
      RECT 11.015000  2.940000 11.395000 3.245000 ;
      RECT 11.105000  0.085000 11.355000 0.505000 ;
      RECT 11.535000  0.375000 11.865000 0.675000 ;
      RECT 11.800000  2.370000 13.400000 2.540000 ;
      RECT 11.800000  2.540000 11.970000 2.600000 ;
      RECT 12.075000  0.085000 12.405000 0.640000 ;
      RECT 12.085000  0.810000 12.415000 1.550000 ;
      RECT 12.140000  2.710000 12.470000 3.245000 ;
      RECT 13.015000  0.085000 13.345000 1.130000 ;
      RECT 13.040000  2.710000 13.370000 3.245000 ;
      RECT 13.230000  1.300000 13.535000 1.630000 ;
      RECT 13.230000  1.630000 13.400000 2.370000 ;
      RECT 13.955000  0.085000 14.285000 0.630000 ;
      RECT 14.045000  1.820000 14.295000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  1.210000  0.325000 1.380000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  1.210000  4.165000 1.380000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  0.840000  8.485000 1.010000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  0.840000 12.325000 1.010000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
    LAYER met1 ;
      RECT  0.095000 1.180000  0.385000 1.225000 ;
      RECT  0.095000 1.225000  4.225000 1.365000 ;
      RECT  0.095000 1.365000  0.385000 1.410000 ;
      RECT  3.935000 1.180000  4.225000 1.225000 ;
      RECT  3.935000 1.365000  4.225000 1.410000 ;
      RECT  8.255000 0.810000  8.545000 0.855000 ;
      RECT  8.255000 0.855000 12.385000 0.995000 ;
      RECT  8.255000 0.995000  8.545000 1.040000 ;
      RECT 12.095000 0.810000 12.385000 0.855000 ;
      RECT 12.095000 0.995000 12.385000 1.040000 ;
  END
END sky130_fd_sc_hs__fah_2
MACRO sky130_fd_sc_hs__fah_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  15.36000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.510000 1.095000 1.800000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.723000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.675000 1.220000 4.925000 2.290000 ;
        RECT 4.675000 2.290000 5.155000 2.910000 ;
    END
  END B
  PIN CI
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.635000 1.350000 12.980000 1.780000 ;
    END
  END CI
  PIN COUT
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  9.890000 1.850000 11.395000 2.100000 ;
        RECT 10.475000 1.010000 11.785000 1.180000 ;
        RECT 10.960000 1.180000 11.785000 1.260000 ;
        RECT 10.960000 1.260000 11.395000 1.850000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  1.097600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.420000 1.850000 14.755000 2.020000 ;
        RECT 13.420000 2.020000 13.750000 2.980000 ;
        RECT 13.555000 0.480000 13.805000 1.010000 ;
        RECT 13.555000 1.010000 14.745000 1.180000 ;
        RECT 14.420000 2.020000 14.755000 2.980000 ;
        RECT 14.495000 0.480000 14.745000 1.010000 ;
        RECT 14.495000 1.180000 14.745000 1.850000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 15.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 15.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 15.360000 0.085000 ;
      RECT  0.000000  3.245000 15.360000 3.415000 ;
      RECT  0.085000  0.350000  0.365000 1.170000 ;
      RECT  0.085000  1.170000  1.665000 1.340000 ;
      RECT  0.085000  1.340000  0.255000 1.970000 ;
      RECT  0.085000  1.970000  0.365000 2.980000 ;
      RECT  0.545000  0.085000  0.795000 1.000000 ;
      RECT  0.565000  1.970000  0.815000 3.245000 ;
      RECT  0.975000  0.350000  1.305000 0.790000 ;
      RECT  0.975000  0.790000  2.135000 0.960000 ;
      RECT  0.975000  0.960000  2.005000 1.000000 ;
      RECT  1.015000  1.970000  1.345000 2.630000 ;
      RECT  1.015000  2.630000  3.495000 2.800000 ;
      RECT  1.015000  2.800000  1.345000 2.980000 ;
      RECT  1.335000  1.340000  1.665000 1.650000 ;
      RECT  1.535000  0.085000  1.795000 0.620000 ;
      RECT  1.575000  2.970000  1.915000 3.245000 ;
      RECT  1.835000  1.000000  2.005000 2.630000 ;
      RECT  1.965000  0.255000  3.415000 0.425000 ;
      RECT  1.965000  0.425000  2.135000 0.790000 ;
      RECT  2.175000  1.790000  2.505000 2.290000 ;
      RECT  2.175000  2.290000  4.505000 2.460000 ;
      RECT  2.305000  0.625000  2.475000 1.790000 ;
      RECT  2.655000  0.625000  2.985000 1.210000 ;
      RECT  2.655000  1.210000  3.545000 1.380000 ;
      RECT  2.705000  1.550000  3.205000 1.780000 ;
      RECT  2.705000  1.780000  2.960000 2.120000 ;
      RECT  3.155000  0.425000  3.415000 1.040000 ;
      RECT  3.165000  2.800000  3.495000 2.960000 ;
      RECT  3.375000  1.380000  3.545000 1.935000 ;
      RECT  3.375000  1.935000  4.030000 2.120000 ;
      RECT  3.715000  0.630000  3.885000 1.550000 ;
      RECT  3.715000  1.550000  4.165000 1.765000 ;
      RECT  4.055000  0.255000  4.385000 0.705000 ;
      RECT  4.055000  0.705000  5.405000 0.875000 ;
      RECT  4.065000  1.045000  4.505000 1.310000 ;
      RECT  4.230000  1.935000  4.505000 2.290000 ;
      RECT  4.230000  2.460000  4.505000 2.670000 ;
      RECT  4.335000  1.310000  4.505000 1.935000 ;
      RECT  4.585000  0.085000  4.915000 0.535000 ;
      RECT  5.095000  0.255000  8.195000 0.425000 ;
      RECT  5.095000  0.425000  5.405000 0.705000 ;
      RECT  5.095000  0.875000  5.405000 0.920000 ;
      RECT  5.095000  0.920000  5.265000 1.950000 ;
      RECT  5.095000  1.950000  6.025000 2.120000 ;
      RECT  5.325000  2.290000  5.655000 3.245000 ;
      RECT  5.435000  1.090000  5.805000 1.375000 ;
      RECT  5.435000  1.375000  5.635000 1.780000 ;
      RECT  5.855000  2.120000  6.025000 2.980000 ;
      RECT  5.875000  0.595000  6.205000 0.875000 ;
      RECT  5.885000  1.550000  6.145000 1.780000 ;
      RECT  5.975000  0.875000  6.145000 1.550000 ;
      RECT  6.195000  1.980000  6.485000 2.150000 ;
      RECT  6.195000  2.150000  6.365000 2.905000 ;
      RECT  6.195000  2.905000  8.715000 3.075000 ;
      RECT  6.315000  1.045000  7.195000 1.215000 ;
      RECT  6.315000  1.215000  6.485000 1.980000 ;
      RECT  6.375000  0.595000  8.535000 0.765000 ;
      RECT  6.375000  0.765000  6.705000 0.845000 ;
      RECT  6.535000  2.320000  7.535000 2.490000 ;
      RECT  6.535000  2.490000  6.785000 2.735000 ;
      RECT  6.655000  1.405000  7.075000 2.150000 ;
      RECT  6.865000  1.015000  7.195000 1.045000 ;
      RECT  6.990000  2.725000  7.875000 2.905000 ;
      RECT  7.365000  0.935000  8.875000 1.105000 ;
      RECT  7.365000  1.105000  7.685000 1.285000 ;
      RECT  7.365000  1.285000  7.535000 2.320000 ;
      RECT  7.705000  1.480000  8.875000 1.650000 ;
      RECT  7.705000  1.650000  7.875000 2.725000 ;
      RECT  8.045000  2.095000  8.375000 2.270000 ;
      RECT  8.045000  2.270000 12.125000 2.440000 ;
      RECT  8.045000  2.440000  8.375000 2.735000 ;
      RECT  8.205000  1.320000  8.875000 1.480000 ;
      RECT  8.365000  0.255000  9.895000 0.425000 ;
      RECT  8.365000  0.425000  8.535000 0.595000 ;
      RECT  8.545000  2.610000 12.715000 2.780000 ;
      RECT  8.545000  2.780000  8.715000 2.905000 ;
      RECT  8.580000  1.900000  9.215000 2.100000 ;
      RECT  8.705000  0.595000  9.555000 0.765000 ;
      RECT  8.705000  0.765000  8.875000 0.935000 ;
      RECT  9.045000  0.935000  9.215000 1.550000 ;
      RECT  9.045000  1.550000  9.475000 1.775000 ;
      RECT  9.045000  1.775000  9.215000 1.900000 ;
      RECT  9.115000  2.950000  9.685000 3.245000 ;
      RECT  9.385000  0.765000  9.555000 1.010000 ;
      RECT  9.385000  1.010000  9.950000 1.180000 ;
      RECT  9.725000  0.425000  9.895000 0.670000 ;
      RECT  9.725000  0.670000 13.385000 0.840000 ;
      RECT  9.780000  1.180000  9.950000 1.350000 ;
      RECT  9.780000  1.350000 10.710000 1.680000 ;
      RECT 10.065000  0.085000 10.315000 0.500000 ;
      RECT 10.425000  2.950000 10.755000 3.245000 ;
      RECT 10.965000  0.085000 11.295000 0.500000 ;
      RECT 11.495000  2.950000 12.125000 3.245000 ;
      RECT 11.955000  0.840000 12.125000 2.270000 ;
      RECT 11.965000  0.085000 12.295000 0.500000 ;
      RECT 12.295000  1.010000 12.855000 1.180000 ;
      RECT 12.295000  1.180000 12.465000 1.950000 ;
      RECT 12.295000  1.950000 12.715000 2.610000 ;
      RECT 12.295000  2.780000 12.715000 2.860000 ;
      RECT 12.920000  1.950000 13.250000 3.245000 ;
      RECT 13.035000  0.085000 13.375000 0.500000 ;
      RECT 13.215000  0.840000 13.385000 1.350000 ;
      RECT 13.215000  1.350000 14.325000 1.680000 ;
      RECT 13.920000  2.190000 14.250000 3.245000 ;
      RECT 13.985000  0.085000 14.315000 0.840000 ;
      RECT 14.915000  0.085000 15.245000 1.260000 ;
      RECT 14.950000  1.820000 15.200000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  1.580000  3.205000 1.750000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  1.950000  3.685000 2.120000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  1.580000  4.165000 1.750000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  1.580000  5.605000 1.750000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  1.580000  6.085000 1.750000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  1.950000  7.045000 2.120000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  1.580000  9.445000 1.750000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.245000 15.205000 3.415000 ;
    LAYER met1 ;
      RECT 2.975000 1.550000 3.265000 1.595000 ;
      RECT 2.975000 1.595000 5.665000 1.735000 ;
      RECT 2.975000 1.735000 3.265000 1.780000 ;
      RECT 3.455000 1.920000 3.745000 1.965000 ;
      RECT 3.455000 1.965000 7.105000 2.105000 ;
      RECT 3.455000 2.105000 3.745000 2.150000 ;
      RECT 3.935000 1.550000 4.225000 1.595000 ;
      RECT 3.935000 1.735000 4.225000 1.780000 ;
      RECT 5.375000 1.550000 5.665000 1.595000 ;
      RECT 5.375000 1.735000 5.665000 1.780000 ;
      RECT 5.855000 1.550000 6.145000 1.595000 ;
      RECT 5.855000 1.595000 9.505000 1.735000 ;
      RECT 5.855000 1.735000 6.145000 1.780000 ;
      RECT 6.815000 1.920000 7.105000 1.965000 ;
      RECT 6.815000 2.105000 7.105000 2.150000 ;
      RECT 9.215000 1.550000 9.505000 1.595000 ;
      RECT 9.215000 1.735000 9.505000 1.780000 ;
  END
END sky130_fd_sc_hs__fah_4
MACRO sky130_fd_sc_hs__fahcin_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.96000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 1.350000 0.835000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.723000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.875000 1.180000 5.205000 1.585000 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.525000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.705000 1.155000 9.035000 1.485000 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  1.959800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.640000 0.440000 8.035000 0.985000 ;
        RECT 6.640000 0.985000 7.070000 1.310000 ;
        RECT 6.820000 2.335000 7.615000 2.665000 ;
        RECT 6.900000 1.310000 7.070000 2.335000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.515000 0.440000 12.845000 0.840000 ;
        RECT 12.595000 0.840000 12.845000 2.980000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.960000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 12.960000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.960000 0.085000 ;
      RECT  0.000000  3.245000 12.960000 3.415000 ;
      RECT  0.120000  0.350000  0.450000 1.010000 ;
      RECT  0.120000  1.010000  1.290000 1.180000 ;
      RECT  0.120000  1.180000  0.375000 2.980000 ;
      RECT  0.575000  1.950000  0.825000 3.245000 ;
      RECT  0.620000  0.085000  0.950000 0.840000 ;
      RECT  1.005000  1.180000  1.290000 1.300000 ;
      RECT  1.005000  1.300000  1.445000 1.630000 ;
      RECT  1.005000  1.630000  1.175000 2.905000 ;
      RECT  1.005000  2.905000  3.935000 3.075000 ;
      RECT  1.120000  0.255000  2.835000 0.425000 ;
      RECT  1.120000  0.425000  1.290000 1.010000 ;
      RECT  1.345000  1.820000  1.835000 2.565000 ;
      RECT  1.345000  2.565000  2.980000 2.735000 ;
      RECT  1.475000  0.615000  1.835000 1.020000 ;
      RECT  1.615000  1.020000  1.835000 1.820000 ;
      RECT  2.045000  1.890000  2.415000 2.070000 ;
      RECT  2.045000  2.070000  2.485000 2.395000 ;
      RECT  2.165000  0.615000  2.415000 1.890000 ;
      RECT  2.585000  0.425000  2.835000 0.750000 ;
      RECT  2.655000  2.045000  2.980000 2.565000 ;
      RECT  2.810000  0.920000  3.175000 1.090000 ;
      RECT  2.810000  1.090000  2.980000 2.045000 ;
      RECT  3.005000  0.255000  3.945000 0.425000 ;
      RECT  3.005000  0.425000  3.175000 0.920000 ;
      RECT  3.185000  1.875000  3.515000 1.880000 ;
      RECT  3.185000  1.880000  4.275000 2.050000 ;
      RECT  3.185000  2.050000  3.515000 2.735000 ;
      RECT  3.345000  0.595000  3.515000 1.875000 ;
      RECT  3.685000  1.380000  4.285000 1.550000 ;
      RECT  3.685000  1.550000  3.990000 1.710000 ;
      RECT  3.685000  2.250000  3.935000 2.905000 ;
      RECT  3.695000  0.425000  3.945000 1.125000 ;
      RECT  4.105000  2.050000  4.275000 2.905000 ;
      RECT  4.105000  2.905000  5.045000 3.075000 ;
      RECT  4.115000  0.255000  5.295000 0.425000 ;
      RECT  4.115000  0.425000  4.285000 1.380000 ;
      RECT  4.445000  1.875000  4.705000 2.735000 ;
      RECT  4.455000  0.670000  4.705000 1.875000 ;
      RECT  4.875000  2.390000  6.650000 2.560000 ;
      RECT  4.875000  2.560000  5.045000 2.905000 ;
      RECT  4.955000  1.820000  5.800000 1.990000 ;
      RECT  4.955000  1.990000  5.285000 2.220000 ;
      RECT  4.965000  0.425000  5.295000 0.840000 ;
      RECT  4.965000  0.840000  5.800000 1.010000 ;
      RECT  5.405000  2.730000  5.765000 3.245000 ;
      RECT  5.465000  0.085000  5.970000 0.635000 ;
      RECT  5.630000  1.010000  5.800000 1.255000 ;
      RECT  5.630000  1.255000  5.970000 1.585000 ;
      RECT  5.630000  1.585000  5.800000 1.820000 ;
      RECT  5.970000  1.820000  6.310000 2.220000 ;
      RECT  6.140000  0.385000  6.470000 1.065000 ;
      RECT  6.140000  1.065000  6.310000 1.820000 ;
      RECT  6.150000  2.560000  6.650000 2.905000 ;
      RECT  6.150000  2.905000  8.715000 3.075000 ;
      RECT  6.480000  1.510000  6.730000 1.840000 ;
      RECT  6.480000  1.840000  6.650000 2.390000 ;
      RECT  7.240000  1.170000  7.555000 2.150000 ;
      RECT  7.745000  1.155000  8.035000 1.485000 ;
      RECT  7.785000  1.485000  7.955000 2.905000 ;
      RECT  8.125000  1.820000  8.375000 2.735000 ;
      RECT  8.205000  0.385000  8.535000 1.065000 ;
      RECT  8.205000  1.065000  8.375000 1.820000 ;
      RECT  8.545000  1.655000  9.385000 1.825000 ;
      RECT  8.545000  1.825000  8.715000 2.905000 ;
      RECT  8.705000  0.085000  9.045000 0.985000 ;
      RECT  8.885000  1.995000  9.055000 3.245000 ;
      RECT  9.215000  0.255000 10.575000 0.570000 ;
      RECT  9.215000  0.570000  9.385000 1.655000 ;
      RECT  9.255000  1.995000  9.725000 2.905000 ;
      RECT  9.255000  2.905000 11.975000 3.075000 ;
      RECT  9.555000  0.740000  9.885000 1.340000 ;
      RECT  9.555000  1.340000  9.725000 1.995000 ;
      RECT  9.895000  1.900000 10.065000 2.400000 ;
      RECT  9.895000  2.400000 11.635000 2.570000 ;
      RECT  9.895000  2.570000 10.065000 2.735000 ;
      RECT 10.070000  0.740000 10.915000 1.260000 ;
      RECT 10.265000  1.260000 10.515000 2.230000 ;
      RECT 10.685000  1.430000 11.015000 2.150000 ;
      RECT 10.745000  0.320000 11.755000 0.490000 ;
      RECT 10.745000  0.490000 10.915000 0.740000 ;
      RECT 10.800000  2.740000 11.155000 2.905000 ;
      RECT 11.085000  0.660000 11.415000 1.220000 ;
      RECT 11.085000  1.220000 11.365000 1.250000 ;
      RECT 11.195000  1.250000 11.365000 1.850000 ;
      RECT 11.195000  1.850000 11.635000 2.400000 ;
      RECT 11.385000  2.570000 11.635000 2.735000 ;
      RECT 11.535000  1.350000 11.975000 1.680000 ;
      RECT 11.585000  0.490000 11.755000 1.010000 ;
      RECT 11.585000  1.010000 12.425000 1.180000 ;
      RECT 11.805000  1.680000 11.975000 2.905000 ;
      RECT 11.925000  0.085000 12.345000 0.810000 ;
      RECT 12.145000  1.180000 12.425000 1.680000 ;
      RECT 12.145000  1.850000 12.395000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  1.950000  2.245000 2.120000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  1.950000  4.645000 2.120000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  1.950000  7.525000 2.120000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  1.950000 10.885000 2.120000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
    LAYER met1 ;
      RECT  2.015000 1.920000  2.305000 1.965000 ;
      RECT  2.015000 1.965000 10.945000 2.105000 ;
      RECT  2.015000 2.105000  2.305000 2.150000 ;
      RECT  4.415000 1.920000  4.705000 1.965000 ;
      RECT  4.415000 2.105000  4.705000 2.150000 ;
      RECT  7.295000 1.920000  7.585000 1.965000 ;
      RECT  7.295000 2.105000  7.585000 2.150000 ;
      RECT 10.655000 1.920000 10.945000 1.965000 ;
      RECT 10.655000 2.105000 10.945000 2.150000 ;
  END
END sky130_fd_sc_hs__fahcin_1
MACRO sky130_fd_sc_hs__fahcon_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.52000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.350000 0.805000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.969000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.180000 5.060000 1.550000 ;
    END
  END B
  PIN CI
    ANTENNAGATEAREA  0.525000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.675000 1.180000 8.005000 1.550000 ;
    END
  END CI
  PIN COUT_N
    ANTENNADIFFAREA  0.782600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.790000 2.085000 6.175000 2.255000 ;
        RECT 5.790000 2.255000 6.120000 2.965000 ;
        RECT 6.005000 1.210000 6.650000 1.380000 ;
        RECT 6.005000 1.380000 6.175000 2.085000 ;
        RECT 6.320000 0.350000 6.650000 1.210000 ;
    END
  END COUT_N
  PIN SUM
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.075000 1.820000 11.435000 2.980000 ;
        RECT 11.155000 0.350000 11.435000 1.130000 ;
        RECT 11.265000 1.130000 11.435000 1.820000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.520000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 11.520000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.520000 0.085000 ;
      RECT  0.000000  3.245000 11.520000 3.415000 ;
      RECT  0.085000  0.480000  0.365000 0.980000 ;
      RECT  0.085000  0.980000  1.245000 1.150000 ;
      RECT  0.085000  1.150000  1.180000 1.180000 ;
      RECT  0.085000  1.180000  0.255000 1.950000 ;
      RECT  0.085000  1.950000  0.485000 2.980000 ;
      RECT  0.545000  0.085000  0.715000 0.480000 ;
      RECT  0.545000  0.480000  0.905000 0.810000 ;
      RECT  0.655000  1.950000  0.985000 3.245000 ;
      RECT  0.975000  1.180000  1.180000 1.680000 ;
      RECT  1.075000  0.255000  2.615000 0.425000 ;
      RECT  1.075000  0.425000  1.245000 0.980000 ;
      RECT  1.190000  1.850000  1.520000 2.905000 ;
      RECT  1.190000  2.905000  3.810000 3.075000 ;
      RECT  1.350000  1.320000  1.745000 1.490000 ;
      RECT  1.350000  1.490000  1.520000 1.850000 ;
      RECT  1.415000  0.595000  1.745000 1.320000 ;
      RECT  1.690000  1.660000  2.095000 1.830000 ;
      RECT  1.690000  1.830000  1.860000 2.565000 ;
      RECT  1.690000  2.565000  3.260000 2.735000 ;
      RECT  1.925000  0.595000  2.275000 1.325000 ;
      RECT  1.925000  1.325000  2.095000 1.660000 ;
      RECT  2.030000  2.000000  2.200000 2.225000 ;
      RECT  2.030000  2.225000  3.275000 2.395000 ;
      RECT  2.400000  1.805000  2.775000 2.055000 ;
      RECT  2.445000  0.425000  2.615000 0.725000 ;
      RECT  2.445000  0.725000  2.775000 1.805000 ;
      RECT  2.785000  0.255000  4.735000 0.425000 ;
      RECT  2.785000  0.425000  3.115000 0.555000 ;
      RECT  2.945000  0.725000  3.275000 2.225000 ;
      RECT  3.460000  0.645000  3.810000 2.905000 ;
      RECT  4.040000  0.425000  4.735000 1.010000 ;
      RECT  4.040000  1.010000  4.210000 1.805000 ;
      RECT  4.040000  1.805000  4.375000 2.965000 ;
      RECT  4.545000  1.805000  4.875000 3.245000 ;
      RECT  4.905000  0.085000  5.155000 0.965000 ;
      RECT  5.100000  1.975000  5.430000 2.965000 ;
      RECT  5.230000  1.135000  5.495000 1.305000 ;
      RECT  5.230000  1.305000  5.400000 1.975000 ;
      RECT  5.325000  0.390000  6.150000 0.640000 ;
      RECT  5.325000  0.640000  5.495000 1.135000 ;
      RECT  5.570000  1.475000  5.835000 1.805000 ;
      RECT  5.665000  0.810000  6.115000 1.040000 ;
      RECT  5.665000  1.040000  5.835000 1.475000 ;
      RECT  6.345000  1.550000  6.610000 1.880000 ;
      RECT  6.345000  2.085000  7.475000 2.970000 ;
      RECT  6.820000  0.810000  7.075000 1.130000 ;
      RECT  6.820000  1.130000  7.135000 1.800000 ;
      RECT  7.245000  0.350000  7.575000 0.960000 ;
      RECT  7.305000  0.960000  7.475000 2.085000 ;
      RECT  7.645000  1.940000  7.815000 3.245000 ;
      RECT  7.745000  0.085000  7.995000 1.010000 ;
      RECT  8.015000  1.820000  8.345000 2.320000 ;
      RECT  8.015000  2.320000 10.030000 2.490000 ;
      RECT  8.015000  2.490000  8.345000 2.980000 ;
      RECT  8.175000  0.350000  8.515000 1.130000 ;
      RECT  8.175000  1.130000  8.345000 1.820000 ;
      RECT  8.515000  1.300000  8.765000 1.550000 ;
      RECT  8.515000  1.550000  8.965000 1.780000 ;
      RECT  8.575000  2.660000  8.905000 2.870000 ;
      RECT  8.575000  2.870000 10.455000 3.040000 ;
      RECT  8.775000  0.255000 10.325000 0.425000 ;
      RECT  8.775000  0.425000  9.105000 1.130000 ;
      RECT  8.935000  1.130000  9.105000 1.210000 ;
      RECT  8.935000  1.210000  9.305000 1.380000 ;
      RECT  9.135000  1.380000  9.305000 1.820000 ;
      RECT  9.135000  1.820000  9.360000 2.150000 ;
      RECT  9.275000  0.810000  9.645000 1.040000 ;
      RECT  9.475000  1.040000  9.645000 1.260000 ;
      RECT  9.475000  1.260000  9.690000 1.590000 ;
      RECT  9.560000  1.820000 10.030000 2.320000 ;
      RECT  9.560000  2.490000 10.030000 2.700000 ;
      RECT  9.815000  0.595000  9.985000 0.920000 ;
      RECT  9.815000  0.920000 10.625000 1.090000 ;
      RECT  9.860000  1.260000 10.285000 1.590000 ;
      RECT  9.860000  1.590000 10.030000 1.820000 ;
      RECT 10.155000  0.425000 10.325000 0.580000 ;
      RECT 10.155000  0.580000 10.980000 0.750000 ;
      RECT 10.200000  1.760000 10.625000 1.930000 ;
      RECT 10.200000  1.930000 10.455000 2.870000 ;
      RECT 10.455000  1.090000 10.625000 1.760000 ;
      RECT 10.495000  0.085000 10.895000 0.410000 ;
      RECT 10.650000  2.100000 10.900000 3.245000 ;
      RECT 10.810000  0.750000 10.980000 1.300000 ;
      RECT 10.810000  1.300000 11.095000 1.630000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  0.840000  2.245000 1.010000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  1.580000  3.205000 1.750000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  0.840000  6.085000 1.010000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  1.580000  6.565000 1.750000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  0.840000  7.045000 1.010000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  1.580000  8.965000 1.750000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  0.840000  9.445000 1.010000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
    LAYER met1 ;
      RECT 2.015000 0.810000 2.305000 0.855000 ;
      RECT 2.015000 0.855000 9.505000 0.995000 ;
      RECT 2.015000 0.995000 2.305000 1.040000 ;
      RECT 2.975000 1.550000 3.265000 1.595000 ;
      RECT 2.975000 1.595000 9.025000 1.735000 ;
      RECT 2.975000 1.735000 3.265000 1.780000 ;
      RECT 5.855000 0.810000 6.145000 0.855000 ;
      RECT 5.855000 0.995000 6.145000 1.040000 ;
      RECT 6.335000 1.550000 6.625000 1.595000 ;
      RECT 6.335000 1.735000 6.625000 1.780000 ;
      RECT 6.815000 0.810000 7.105000 0.855000 ;
      RECT 6.815000 0.995000 7.105000 1.040000 ;
      RECT 8.735000 1.550000 9.025000 1.595000 ;
      RECT 8.735000 1.735000 9.025000 1.780000 ;
      RECT 9.215000 0.810000 9.505000 0.855000 ;
      RECT 9.215000 0.995000 9.505000 1.040000 ;
  END
END sky130_fd_sc_hs__fahcon_1
MACRO sky130_fd_sc_hs__fill_1
  CLASS CORE SPACER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.480000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 0.480000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 0.480000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.480000 0.085000 ;
      RECT 0.000000  3.245000 0.480000 3.415000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
  END
END sky130_fd_sc_hs__fill_1
MACRO sky130_fd_sc_hs__fill_2
  CLASS CORE SPACER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.960000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 0.960000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 0.960000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.960000 0.085000 ;
      RECT 0.000000  3.245000 0.960000 3.415000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
  END
END sky130_fd_sc_hs__fill_2
MACRO sky130_fd_sc_hs__fill_4
  CLASS CORE SPACER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.920000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 1.920000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 1.920000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.920000 0.085000 ;
      RECT 0.000000  3.245000 1.920000 3.415000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
  END
END sky130_fd_sc_hs__fill_4
MACRO sky130_fd_sc_hs__fill_8
  CLASS CORE SPACER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__fill_8
MACRO sky130_fd_sc_hs__fill_diode_2
  CLASS CORE SPACER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.960000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 0.960000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 0.960000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.960000 0.085000 ;
      RECT 0.000000  3.245000 0.960000 3.415000 ;
      RECT 0.135000  0.085000 0.825000 0.580000 ;
      RECT 0.135000  2.750000 0.825000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
  END
END sky130_fd_sc_hs__fill_diode_2
MACRO sky130_fd_sc_hs__fill_diode_4
  CLASS CORE SPACER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.920000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 1.920000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 1.920000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.920000 0.085000 ;
      RECT 0.000000  3.245000 1.920000 3.415000 ;
      RECT 0.135000  0.085000 1.785000 0.580000 ;
      RECT 0.135000  2.750000 1.785000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
  END
END sky130_fd_sc_hs__fill_diode_4
MACRO sky130_fd_sc_hs__fill_diode_8
  CLASS CORE SPACER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.135000  0.085000 3.705000 0.580000 ;
      RECT 0.135000  2.750000 3.705000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__fill_diode_8
MACRO sky130_fd_sc_hs__ha_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.468000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.450000 0.255000 2.780000 0.670000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.468000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.765000 1.470000 2.095000 1.550000 ;
        RECT 1.765000 1.550000 3.300000 1.800000 ;
        RECT 2.970000 1.470000 3.300000 1.550000 ;
    END
  END B
  PIN COUT
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.310000 0.475000 4.715000 1.180000 ;
        RECT 4.310000 1.850000 4.715000 2.980000 ;
        RECT 4.545000 1.180000 4.715000 1.850000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.350000 0.445000 1.130000 ;
        RECT 0.115000 1.130000 0.355000 1.820000 ;
        RECT 0.115000 1.820000 0.445000 2.980000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.525000  1.300000 0.855000 1.630000 ;
      RECT 0.615000  2.650000 1.205000 3.245000 ;
      RECT 0.625000  0.085000 0.875000 0.795000 ;
      RECT 0.685000  1.130000 1.400000 1.300000 ;
      RECT 0.685000  1.630000 0.855000 2.310000 ;
      RECT 0.685000  2.310000 1.740000 2.480000 ;
      RECT 1.070000  0.910000 1.400000 1.130000 ;
      RECT 1.195000  1.470000 1.525000 1.970000 ;
      RECT 1.195000  1.970000 3.640000 2.140000 ;
      RECT 1.410000  2.480000 1.740000 2.800000 ;
      RECT 1.580000  0.630000 1.750000 1.130000 ;
      RECT 1.580000  1.130000 2.790000 1.300000 ;
      RECT 1.930000  0.085000 2.280000 0.960000 ;
      RECT 2.460000  0.840000 2.790000 1.130000 ;
      RECT 2.460000  1.300000 2.790000 1.355000 ;
      RECT 2.485000  2.310000 3.190000 3.245000 ;
      RECT 3.020000  0.575000 3.350000 1.085000 ;
      RECT 3.020000  1.085000 3.640000 1.255000 ;
      RECT 3.360000  2.140000 3.640000 2.980000 ;
      RECT 3.470000  1.255000 3.640000 1.350000 ;
      RECT 3.470000  1.350000 4.375000 1.680000 ;
      RECT 3.470000  1.680000 3.640000 1.970000 ;
      RECT 3.810000  0.085000 4.140000 1.180000 ;
      RECT 3.810000  2.100000 4.140000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_hs__ha_1
MACRO sky130_fd_sc_hs__ha_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.522000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.060000 1.450000 1.390000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.522000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.550000 1.630000 ;
        RECT 0.125000 1.630000 0.295000 2.320000 ;
        RECT 0.125000 2.320000 2.120000 2.520000 ;
        RECT 1.790000 1.450000 2.120000 2.320000 ;
    END
  END B
  PIN COUT
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.865000 1.820000 5.195000 2.170000 ;
        RECT 4.885000 0.350000 5.215000 1.130000 ;
        RECT 4.885000 1.130000 5.055000 1.820000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.580200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.820000 4.675000 2.170000 ;
        RECT 3.975000 0.880000 4.675000 1.050000 ;
        RECT 4.505000 1.050000 4.675000 1.820000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.115000  0.350000 0.445000 0.960000 ;
      RECT 0.115000  0.960000 0.890000 1.110000 ;
      RECT 0.115000  1.110000 2.460000 1.130000 ;
      RECT 0.115000  2.690000 0.445000 3.245000 ;
      RECT 0.565000  1.980000 0.895000 2.150000 ;
      RECT 0.720000  1.130000 2.460000 1.280000 ;
      RECT 0.720000  1.280000 0.890000 1.980000 ;
      RECT 0.935000  0.085000 1.265000 0.600000 ;
      RECT 1.015000  2.690000 1.400000 3.245000 ;
      RECT 1.365000  0.770000 2.465000 0.940000 ;
      RECT 1.795000  0.085000 2.125000 0.600000 ;
      RECT 2.290000  1.280000 3.035000 1.610000 ;
      RECT 2.290000  1.610000 2.460000 2.340000 ;
      RECT 2.290000  2.340000 5.555000 2.510000 ;
      RECT 2.295000  0.255000 3.315000 0.425000 ;
      RECT 2.295000  0.425000 2.465000 0.770000 ;
      RECT 2.630000  1.920000 3.490000 2.170000 ;
      RECT 2.635000  0.595000 2.805000 0.940000 ;
      RECT 2.635000  0.940000 3.490000 1.110000 ;
      RECT 2.985000  0.425000 3.315000 0.770000 ;
      RECT 3.080000  2.680000 3.845000 3.245000 ;
      RECT 3.320000  1.110000 3.490000 1.220000 ;
      RECT 3.320000  1.220000 4.330000 1.550000 ;
      RECT 3.320000  1.550000 3.490000 1.920000 ;
      RECT 3.545000  0.085000 3.875000 0.710000 ;
      RECT 4.415000  2.680000 4.745000 3.245000 ;
      RECT 4.455000  0.085000 4.705000 0.710000 ;
      RECT 5.225000  1.300000 5.555000 1.630000 ;
      RECT 5.315000  2.680000 5.645000 3.245000 ;
      RECT 5.385000  1.630000 5.555000 2.340000 ;
      RECT 5.395000  0.085000 5.645000 1.130000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_hs__ha_2
MACRO sky130_fd_sc_hs__ha_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.936000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.455000 1.315000 1.785000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.936000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.455000 2.275000 1.785000 ;
    END
  END B
  PIN COUT
    ANTENNADIFFAREA  1.265600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.220000 1.820000 7.555000 2.150000 ;
        RECT 6.350000 0.350000 6.600000 0.880000 ;
        RECT 6.350000 0.880000 7.555000 1.130000 ;
        RECT 7.210000 1.130000 7.555000 1.820000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  1.470100 ;
    ANTENNAPARTIALMETALSIDEAREA  0.861000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 8.735000 1.920000 9.025000 1.965000 ;
        RECT 8.735000 1.965000 9.985000 2.105000 ;
        RECT 8.735000 2.105000 9.025000 2.150000 ;
        RECT 9.695000 1.920000 9.985000 1.965000 ;
        RECT 9.695000 2.105000 9.985000 2.150000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.105000  1.955000  1.255000 2.125000 ;
      RECT 0.105000  2.125000  0.385000 2.965000 ;
      RECT 0.115000  0.605000  0.365000 1.115000 ;
      RECT 0.115000  1.115000  2.170000 1.285000 ;
      RECT 0.545000  0.085000  0.795000 0.945000 ;
      RECT 0.555000  2.295000  0.805000 3.245000 ;
      RECT 0.980000  0.605000  1.230000 1.115000 ;
      RECT 1.005000  2.125000  1.255000 2.905000 ;
      RECT 1.005000  2.905000  2.235000 3.075000 ;
      RECT 1.410000  0.085000  1.660000 0.945000 ;
      RECT 1.455000  1.955000  3.255000 2.125000 ;
      RECT 1.455000  2.125000  1.735000 2.735000 ;
      RECT 1.840000  0.265000  3.170000 0.435000 ;
      RECT 1.840000  0.435000  2.170000 1.115000 ;
      RECT 1.905000  2.295000  2.235000 2.905000 ;
      RECT 2.340000  0.605000  2.670000 1.285000 ;
      RECT 2.475000  2.405000  2.805000 3.245000 ;
      RECT 2.500000  1.285000  2.670000 1.905000 ;
      RECT 2.500000  1.905000  3.255000 1.955000 ;
      RECT 2.840000  0.435000  3.170000 1.235000 ;
      RECT 2.925000  2.125000  3.255000 2.165000 ;
      RECT 2.925000  2.165000  4.070000 2.235000 ;
      RECT 3.075000  1.405000  4.280000 1.575000 ;
      RECT 3.075000  1.575000  4.070000 1.735000 ;
      RECT 3.085000  2.235000  4.070000 2.320000 ;
      RECT 3.085000  2.320000  7.895000 2.335000 ;
      RECT 3.375000  2.505000  3.705000 3.245000 ;
      RECT 3.520000  0.315000  4.780000 0.485000 ;
      RECT 3.520000  0.485000  3.780000 1.235000 ;
      RECT 3.900000  1.735000  4.070000 1.745000 ;
      RECT 3.900000  1.745000  4.230000 1.820000 ;
      RECT 3.900000  1.820000  6.050000 1.995000 ;
      RECT 3.900000  2.335000  7.895000 2.490000 ;
      RECT 3.950000  0.655000  4.280000 1.405000 ;
      RECT 4.430000  2.660000  4.760000 3.245000 ;
      RECT 4.450000  0.485000  4.780000 1.425000 ;
      RECT 4.450000  1.425000  5.710000 1.595000 ;
      RECT 4.950000  0.085000  5.280000 1.255000 ;
      RECT 4.955000  1.995000  6.050000 2.150000 ;
      RECT 5.460000  0.575000  5.710000 1.425000 ;
      RECT 5.490000  2.660000  5.945000 3.245000 ;
      RECT 5.880000  1.320000  6.955000 1.650000 ;
      RECT 5.880000  1.650000  6.050000 1.820000 ;
      RECT 5.920000  0.085000  6.170000 1.130000 ;
      RECT 6.675000  2.660000  7.005000 3.245000 ;
      RECT 6.780000  0.085000  7.110000 0.710000 ;
      RECT 7.575000  2.660000  7.905000 3.245000 ;
      RECT 7.640000  0.085000  7.970000 0.710000 ;
      RECT 7.725000  1.320000  9.645000 1.650000 ;
      RECT 7.725000  1.650000  7.895000 2.320000 ;
      RECT 8.075000  1.820000  9.995000 2.150000 ;
      RECT 8.075000  2.150000  8.305000 2.980000 ;
      RECT 8.150000  0.350000  8.400000 0.980000 ;
      RECT 8.150000  0.980000  9.995000 1.150000 ;
      RECT 8.475000  2.320000  8.805000 3.245000 ;
      RECT 8.570000  0.085000  8.900000 0.810000 ;
      RECT 9.070000  0.350000  9.400000 0.980000 ;
      RECT 9.075000  2.150000  9.405000 2.980000 ;
      RECT 9.580000  0.085000  9.885000 0.810000 ;
      RECT 9.635000  2.320000  9.965000 3.245000 ;
      RECT 9.825000  1.150000  9.995000 1.820000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  1.950000 8.965000 2.120000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  1.950000 9.925000 2.120000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
  END
END sky130_fd_sc_hs__ha_4
MACRO sky130_fd_sc_hs__inv_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.440000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.815000 1.780000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985000 0.350000 1.315000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 1.440000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 1.440000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.440000 0.085000 ;
      RECT 0.000000  3.245000 1.440000 3.415000 ;
      RECT 0.485000  0.085000 0.815000 1.130000 ;
      RECT 0.485000  1.950000 0.815000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
  END
END sky130_fd_sc_hs__inv_1
MACRO sky130_fd_sc_hs__inv_16
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  4.464000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.085000 1.550000 7.070000 1.780000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  4.379200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.585000 1.920000 7.575000 2.150000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.115000  1.820000 0.365000 3.245000 ;
      RECT 0.185000  0.085000 0.445000 1.130000 ;
      RECT 0.565000  1.330000 0.885000 2.995000 ;
      RECT 0.615000  0.350000 0.945000 1.130000 ;
      RECT 0.615000  1.130000 0.885000 1.330000 ;
      RECT 1.055000  1.940000 1.345000 3.245000 ;
      RECT 1.070000  1.350000 1.380000 1.770000 ;
      RECT 1.115000  0.085000 1.375000 1.130000 ;
      RECT 1.515000  1.940000 1.845000 2.980000 ;
      RECT 1.555000  0.350000 1.845000 1.940000 ;
      RECT 2.020000  1.350000 2.310000 1.770000 ;
      RECT 2.025000  0.085000 2.305000 1.130000 ;
      RECT 2.045000  1.940000 2.295000 3.245000 ;
      RECT 2.465000  1.940000 2.795000 2.980000 ;
      RECT 2.485000  0.350000 2.795000 1.940000 ;
      RECT 2.970000  1.350000 3.245000 1.770000 ;
      RECT 2.975000  0.085000 3.245000 1.130000 ;
      RECT 2.995000  1.940000 3.245000 3.245000 ;
      RECT 3.415000  0.350000 3.710000 2.980000 ;
      RECT 3.885000  1.350000 4.165000 1.770000 ;
      RECT 3.890000  0.085000 4.150000 1.130000 ;
      RECT 3.915000  1.940000 4.150000 3.245000 ;
      RECT 4.340000  0.350000 4.595000 1.940000 ;
      RECT 4.340000  1.940000 4.630000 2.980000 ;
      RECT 4.765000  0.085000 5.025000 1.130000 ;
      RECT 4.770000  1.350000 5.085000 1.770000 ;
      RECT 4.810000  1.940000 5.095000 3.245000 ;
      RECT 5.215000  0.350000 5.525000 1.180000 ;
      RECT 5.265000  1.180000 5.525000 1.285000 ;
      RECT 5.265000  1.285000 5.580000 2.980000 ;
      RECT 5.705000  0.085000 6.025000 1.130000 ;
      RECT 5.755000  1.350000 6.090000 1.770000 ;
      RECT 5.765000  1.940000 6.095000 3.245000 ;
      RECT 6.195000  0.350000 6.525000 1.180000 ;
      RECT 6.265000  1.180000 6.525000 1.285000 ;
      RECT 6.265000  1.285000 6.595000 2.980000 ;
      RECT 6.705000  0.085000 7.045000 1.130000 ;
      RECT 6.765000  1.940000 7.095000 3.245000 ;
      RECT 6.770000  1.350000 7.090000 1.770000 ;
      RECT 7.215000  0.350000 7.545000 1.130000 ;
      RECT 7.265000  1.130000 7.545000 2.980000 ;
      RECT 7.715000  0.085000 8.045000 1.130000 ;
      RECT 7.735000  1.820000 8.045000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 0.645000  1.950000 0.815000 2.120000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.145000  1.580000 1.315000 1.750000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  1.950000 1.765000 2.120000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.085000  1.580000 2.255000 1.750000 ;
      RECT 2.545000  1.950000 2.715000 2.120000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.025000  1.580000 3.195000 1.750000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.495000  1.950000 3.665000 2.120000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.940000  1.580000 4.110000 1.750000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.395000  1.950000 4.565000 2.120000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.850000  1.580000 5.020000 1.750000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.345000  1.950000 5.515000 2.120000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.845000  1.580000 6.015000 1.750000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.345000  1.950000 6.515000 2.120000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.840000  1.580000 7.010000 1.750000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.345000  1.950000 7.515000 2.120000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_hs__inv_16
MACRO sky130_fd_sc_hs__inv_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.440000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.300000 0.435000 1.780000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.560000 0.350000 0.890000 1.130000 ;
        RECT 0.605000 1.130000 0.890000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 1.440000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 1.440000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.440000 0.085000 ;
      RECT 0.000000  3.245000 1.440000 3.415000 ;
      RECT 0.105000  1.950000 0.435000 3.245000 ;
      RECT 0.130000  0.085000 0.380000 1.130000 ;
      RECT 1.070000  0.085000 1.320000 1.130000 ;
      RECT 1.085000  1.820000 1.335000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
  END
END sky130_fd_sc_hs__inv_2
MACRO sky130_fd_sc_hs__inv_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.400000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.800000 1.780000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  1.116000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.600000 1.950000 2.275000 2.120000 ;
        RECT 0.600000 2.120000 0.930000 2.980000 ;
        RECT 0.615000 0.350000 0.865000 1.010000 ;
        RECT 0.615000 1.010000 2.275000 1.180000 ;
        RECT 1.500000 2.120000 1.830000 2.980000 ;
        RECT 1.605000 0.350000 1.775000 1.010000 ;
        RECT 2.045000 1.180000 2.275000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.400000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.400000 0.085000 ;
      RECT 0.000000  3.245000 2.400000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 1.130000 ;
      RECT 0.150000  1.950000 0.400000 3.245000 ;
      RECT 1.045000  0.085000 1.375000 0.840000 ;
      RECT 1.130000  2.290000 1.300000 3.245000 ;
      RECT 1.955000  0.085000 2.285000 0.840000 ;
      RECT 2.030000  2.290000 2.280000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
  END
END sky130_fd_sc_hs__inv_4
MACRO sky130_fd_sc_hs__inv_8
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  2.232000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.560000 1.350000 2.250000 1.780000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  2.172800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.560000 0.350000 0.810000 1.010000 ;
        RECT 0.560000 1.010000 2.680000 1.140000 ;
        RECT 0.560000 1.140000 4.195000 1.180000 ;
        RECT 0.565000 1.950000 2.665000 2.120000 ;
        RECT 0.565000 2.120000 0.815000 2.980000 ;
        RECT 1.500000 0.350000 1.670000 1.010000 ;
        RECT 1.515000 2.120000 1.845000 2.980000 ;
        RECT 2.350000 0.350000 2.680000 1.010000 ;
        RECT 2.420000 1.180000 4.195000 1.310000 ;
        RECT 2.495000 1.310000 4.195000 1.620000 ;
        RECT 2.495000 1.620000 2.665000 1.950000 ;
        RECT 2.495000 2.120000 2.665000 2.980000 ;
        RECT 3.350000 0.350000 3.610000 1.140000 ;
        RECT 3.365000 1.620000 3.695000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  1.820000 0.365000 3.245000 ;
      RECT 0.130000  0.085000 0.380000 1.130000 ;
      RECT 0.990000  0.085000 1.320000 0.840000 ;
      RECT 1.015000  2.290000 1.345000 3.245000 ;
      RECT 1.850000  0.085000 2.180000 0.840000 ;
      RECT 2.045000  2.290000 2.295000 3.245000 ;
      RECT 2.850000  0.085000 3.180000 0.970000 ;
      RECT 2.865000  1.820000 3.195000 3.245000 ;
      RECT 3.780000  0.085000 4.110000 0.970000 ;
      RECT 3.865000  1.820000 4.195000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__inv_8
MACRO sky130_fd_sc_hs__maj3_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.645000 0.255000 3.715000 0.570000 ;
        RECT 3.485000 0.570000 3.715000 0.670000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.430000 1.685000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.285000 1.430000 3.575000 1.760000 ;
        RECT 2.285000 1.760000 2.755000 1.780000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.538500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.480000 0.445000 1.180000 ;
        RECT 0.085000 1.180000 0.255000 1.850000 ;
        RECT 0.085000 1.850000 0.490000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.425000  1.350000 0.785000 1.680000 ;
      RECT 0.615000  0.085000 0.990000 0.910000 ;
      RECT 0.615000  1.090000 3.700000 1.260000 ;
      RECT 0.615000  1.260000 0.785000 1.350000 ;
      RECT 0.660000  1.950000 0.990000 3.245000 ;
      RECT 1.480000  0.580000 1.810000 1.090000 ;
      RECT 1.565000  1.950000 3.725000 2.120000 ;
      RECT 1.565000  2.120000 1.895000 2.940000 ;
      RECT 1.895000  1.260000 2.065000 1.950000 ;
      RECT 2.305000  0.085000 2.475000 0.740000 ;
      RECT 2.305000  0.740000 2.850000 0.910000 ;
      RECT 2.435000  2.290000 2.840000 3.245000 ;
      RECT 3.370000  0.840000 3.700000 1.090000 ;
      RECT 3.395000  1.930000 3.725000 1.950000 ;
      RECT 3.395000  2.120000 3.725000 2.940000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__maj3_1
MACRO sky130_fd_sc_hs__maj3_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.522000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 1.180000 1.795000 1.550000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.522000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.305000 1.245000 2.975000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.522000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.215000 1.245000 3.715000 1.300000 ;
        RECT 3.215000 1.300000 4.535000 1.630000 ;
        RECT 3.215000 1.630000 3.715000 1.780000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.555000 0.350000 0.895000 1.130000 ;
        RECT 0.555000 1.130000 0.725000 1.820000 ;
        RECT 0.555000 1.820000 0.915000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.135000  0.085000 0.385000 1.130000 ;
      RECT 0.135000  1.820000 0.385000 3.245000 ;
      RECT 0.895000  1.320000 1.255000 1.650000 ;
      RECT 1.075000  0.085000 1.795000 1.010000 ;
      RECT 1.085000  1.650000 1.255000 1.780000 ;
      RECT 1.085000  1.780000 2.135000 1.950000 ;
      RECT 1.085000  2.120000 1.780000 3.245000 ;
      RECT 1.965000  0.350000 2.760000 0.905000 ;
      RECT 1.965000  0.905000 4.660000 1.075000 ;
      RECT 1.965000  1.075000 2.135000 1.780000 ;
      RECT 1.965000  1.950000 4.685000 2.120000 ;
      RECT 1.965000  2.120000 2.785000 2.755000 ;
      RECT 3.340000  0.085000 3.840000 0.680000 ;
      RECT 3.485000  2.290000 3.815000 3.245000 ;
      RECT 4.330000  0.350000 4.660000 0.905000 ;
      RECT 4.330000  1.075000 4.660000 1.130000 ;
      RECT 4.355000  1.820000 4.685000 1.950000 ;
      RECT 4.355000  2.120000 4.685000 2.860000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_hs__maj3_2
MACRO sky130_fd_sc_hs__maj3_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.984000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.800000 1.470000 2.275000 1.800000 ;
        RECT 2.105000 1.800000 2.275000 1.875000 ;
        RECT 2.105000 1.875000 4.570000 2.045000 ;
        RECT 4.240000 1.470000 4.570000 1.875000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.984000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.135000 1.130000 3.235000 1.300000 ;
        RECT 1.135000 1.300000 1.465000 1.705000 ;
        RECT 2.525000 1.300000 3.235000 1.705000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.984000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.130000 4.925000 1.300000 ;
        RECT 3.485000 1.300000 4.010000 1.705000 ;
        RECT 4.755000 1.300000 4.925000 1.470000 ;
        RECT 4.755000 1.470000 5.220000 1.800000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  1.116000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365000 1.845000 7.515000 2.015000 ;
        RECT 6.365000 2.015000 6.695000 2.980000 ;
        RECT 6.425000 0.475000 6.675000 1.005000 ;
        RECT 6.425000 1.005000 8.035000 1.175000 ;
        RECT 7.345000 1.480000 8.035000 1.650000 ;
        RECT 7.345000 1.650000 7.515000 1.845000 ;
        RECT 7.345000 2.015000 7.515000 2.980000 ;
        RECT 7.805000 1.175000 8.035000 1.480000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 1.285000 ;
      RECT 0.130000  1.940000 0.380000 3.245000 ;
      RECT 0.580000  2.215000 0.910000 2.905000 ;
      RECT 0.580000  2.905000 1.860000 3.075000 ;
      RECT 0.625000  0.265000 1.965000 0.435000 ;
      RECT 0.625000  0.435000 0.955000 0.620000 ;
      RECT 0.795000  0.790000 1.465000 0.960000 ;
      RECT 0.795000  0.960000 0.965000 1.875000 ;
      RECT 0.795000  1.875000 1.410000 2.045000 ;
      RECT 1.095000  2.045000 1.410000 2.215000 ;
      RECT 1.095000  2.215000 5.290000 2.385000 ;
      RECT 1.095000  2.385000 1.350000 2.735000 ;
      RECT 1.135000  0.605000 1.465000 0.790000 ;
      RECT 1.530000  2.555000 1.860000 2.905000 ;
      RECT 1.635000  0.435000 1.965000 0.960000 ;
      RECT 2.060000  2.555000 2.320000 3.245000 ;
      RECT 2.145000  0.085000 2.315000 0.960000 ;
      RECT 2.490000  2.555000 2.820000 2.905000 ;
      RECT 2.490000  2.905000 3.820000 3.075000 ;
      RECT 2.495000  0.265000 3.825000 0.435000 ;
      RECT 2.495000  0.435000 2.885000 0.935000 ;
      RECT 2.990000  2.385000 3.320000 2.735000 ;
      RECT 3.065000  0.605000 3.315000 0.790000 ;
      RECT 3.065000  0.790000 5.265000 0.960000 ;
      RECT 3.490000  2.555000 3.820000 2.905000 ;
      RECT 3.495000  0.435000 3.825000 0.620000 ;
      RECT 3.990000  2.555000 4.320000 3.245000 ;
      RECT 4.005000  0.085000 4.335000 0.620000 ;
      RECT 4.505000  0.255000 5.775000 0.425000 ;
      RECT 4.505000  0.425000 4.835000 0.620000 ;
      RECT 4.510000  2.555000 5.740000 2.725000 ;
      RECT 4.510000  2.725000 4.840000 2.980000 ;
      RECT 4.960000  1.970000 5.560000 2.140000 ;
      RECT 4.960000  2.140000 5.290000 2.215000 ;
      RECT 5.095000  0.595000 5.265000 0.790000 ;
      RECT 5.095000  0.960000 5.265000 1.130000 ;
      RECT 5.095000  1.130000 5.560000 1.300000 ;
      RECT 5.390000  1.300000 5.560000 1.345000 ;
      RECT 5.390000  1.345000 7.150000 1.675000 ;
      RECT 5.390000  1.675000 5.560000 1.970000 ;
      RECT 5.410000  2.725000 5.740000 2.980000 ;
      RECT 5.445000  0.425000 5.775000 0.960000 ;
      RECT 5.940000  1.940000 6.190000 3.245000 ;
      RECT 5.955000  0.085000 6.205000 1.175000 ;
      RECT 6.855000  0.085000 7.185000 0.835000 ;
      RECT 6.895000  2.185000 7.145000 3.245000 ;
      RECT 7.715000  0.085000 8.045000 0.835000 ;
      RECT 7.715000  1.820000 8.045000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_hs__maj3_4
MACRO sky130_fd_sc_hs__mux2_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.885000 1.180000 2.275000 1.550000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.345000 1.220000 1.685000 1.550000 ;
        RECT 1.515000 0.810000 2.785000 0.980000 ;
        RECT 1.515000 0.980000 1.685000 1.220000 ;
        RECT 2.455000 0.980000 2.785000 1.550000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.470000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.505000 1.350000 0.835000 1.780000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.795000 1.820000 4.235000 2.980000 ;
        RECT 3.865000 0.350000 4.235000 1.130000 ;
        RECT 4.065000 1.130000 4.235000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  0.540000 0.445000 1.130000 ;
      RECT 0.115000  1.130000 0.285000 1.950000 ;
      RECT 0.115000  1.950000 0.445000 2.060000 ;
      RECT 0.115000  2.060000 1.320000 2.230000 ;
      RECT 0.115000  2.230000 0.445000 2.700000 ;
      RECT 0.625000  0.085000 1.005000 0.680000 ;
      RECT 0.625000  0.680000 0.835000 1.130000 ;
      RECT 0.650000  2.400000 0.980000 3.245000 ;
      RECT 1.005000  0.850000 1.345000 1.020000 ;
      RECT 1.005000  1.020000 1.175000 1.720000 ;
      RECT 1.005000  1.720000 2.395000 1.890000 ;
      RECT 1.150000  2.230000 1.320000 2.905000 ;
      RECT 1.150000  2.905000 3.125000 3.075000 ;
      RECT 1.175000  0.390000 3.125000 0.640000 ;
      RECT 1.175000  0.640000 1.345000 0.850000 ;
      RECT 2.065000  1.890000 2.395000 2.735000 ;
      RECT 2.955000  0.640000 3.125000 0.980000 ;
      RECT 2.955000  0.980000 3.695000 1.150000 ;
      RECT 2.955000  1.320000 3.355000 1.650000 ;
      RECT 2.955000  1.650000 3.125000 2.905000 ;
      RECT 3.295000  0.085000 3.625000 0.810000 ;
      RECT 3.295000  1.820000 3.625000 3.245000 ;
      RECT 3.525000  1.150000 3.695000 1.300000 ;
      RECT 3.525000  1.300000 3.895000 1.630000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__mux2_1
MACRO sky130_fd_sc_hs__mux2_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.435000 1.550000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.180000 1.195000 1.550000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.470000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.715000 1.450000 2.385000 1.780000 ;
        RECT 2.215000 1.130000 3.455000 1.300000 ;
        RECT 2.215000 1.300000 2.385000 1.450000 ;
        RECT 3.125000 1.300000 3.455000 1.460000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 0.770000 4.665000 2.140000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.280000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.245000 5.280000 3.415000 ;
      RECT 0.115000  1.825000 0.445000 2.905000 ;
      RECT 0.115000  2.905000 1.905000 3.075000 ;
      RECT 0.170000  0.290000 2.750000 0.460000 ;
      RECT 0.170000  0.460000 0.500000 1.010000 ;
      RECT 0.620000  1.820000 1.535000 1.970000 ;
      RECT 0.620000  1.970000 3.165000 2.140000 ;
      RECT 0.620000  2.140000 0.840000 2.725000 ;
      RECT 0.670000  0.680000 1.535000 1.010000 ;
      RECT 1.015000  2.310000 2.825000 2.480000 ;
      RECT 1.015000  2.480000 1.345000 2.735000 ;
      RECT 1.365000  1.010000 1.535000 1.820000 ;
      RECT 1.575000  2.650000 1.905000 2.905000 ;
      RECT 1.715000  0.790000 3.170000 0.960000 ;
      RECT 1.715000  0.960000 2.045000 1.130000 ;
      RECT 2.075000  2.650000 2.405000 3.245000 ;
      RECT 2.420000  0.460000 2.750000 0.620000 ;
      RECT 2.555000  1.470000 2.885000 1.630000 ;
      RECT 2.555000  1.630000 3.795000 1.800000 ;
      RECT 2.575000  2.480000 2.825000 2.980000 ;
      RECT 2.995000  2.140000 3.165000 2.310000 ;
      RECT 2.995000  2.310000 5.165000 2.480000 ;
      RECT 3.000000  0.085000 3.170000 0.790000 ;
      RECT 3.335000  1.800000 3.795000 2.140000 ;
      RECT 3.340000  0.350000 3.670000 0.770000 ;
      RECT 3.340000  0.770000 3.795000 0.940000 ;
      RECT 3.625000  0.940000 3.795000 1.630000 ;
      RECT 3.840000  0.085000 4.230000 0.600000 ;
      RECT 3.870000  2.650000 4.210000 3.245000 ;
      RECT 4.780000  2.650000 5.165000 3.245000 ;
      RECT 4.835000  0.085000 5.165000 1.130000 ;
      RECT 4.835000  1.300000 5.165000 2.310000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
  END
END sky130_fd_sc_hs__mux2_2
MACRO sky130_fd_sc_hs__mux2_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.640000 1.450000 7.075000 1.780000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.325000 1.450000 8.175000 1.780000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.738000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.350000 0.835000 1.780000 ;
        RECT 0.665000 1.780000 0.835000 2.050000 ;
        RECT 0.665000 2.050000 1.675000 2.155000 ;
        RECT 0.665000 2.155000 3.165000 2.220000 ;
        RECT 1.505000 2.220000 3.165000 2.325000 ;
        RECT 2.995000 1.435000 3.745000 1.765000 ;
        RECT 2.995000 1.765000 3.165000 2.155000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  1.576550 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.370000 2.755000 1.710000 ;
        RECT 1.085000 1.710000 2.770000 1.880000 ;
        RECT 1.310000 0.370000 1.640000 1.370000 ;
        RECT 2.330000 0.370000 2.755000 1.370000 ;
        RECT 2.440000 1.880000 2.770000 1.985000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
      RECT 0.000000  3.245000 8.640000 3.415000 ;
      RECT 0.085000  0.470000 0.600000 1.150000 ;
      RECT 0.085000  1.150000 0.255000 1.950000 ;
      RECT 0.085000  1.950000 0.445000 2.390000 ;
      RECT 0.085000  2.390000 1.335000 2.495000 ;
      RECT 0.085000  2.495000 3.505000 2.560000 ;
      RECT 0.085000  2.560000 0.445000 2.860000 ;
      RECT 0.650000  2.730000 0.995000 3.245000 ;
      RECT 0.770000  0.085000 1.100000 1.150000 ;
      RECT 1.165000  2.560000 3.505000 2.665000 ;
      RECT 1.810000  0.085000 2.140000 1.070000 ;
      RECT 1.820000  2.835000 2.150000 3.245000 ;
      RECT 2.925000  0.085000 3.255000 1.255000 ;
      RECT 3.060000  2.835000 3.390000 3.245000 ;
      RECT 3.335000  1.935000 4.085000 2.105000 ;
      RECT 3.335000  2.105000 3.505000 2.495000 ;
      RECT 3.520000  0.575000 3.850000 1.095000 ;
      RECT 3.520000  1.095000 5.325000 1.110000 ;
      RECT 3.520000  1.110000 8.020000 1.265000 ;
      RECT 3.675000  2.275000 3.925000 2.435000 ;
      RECT 3.675000  2.435000 5.790000 2.605000 ;
      RECT 3.675000  2.605000 3.925000 2.975000 ;
      RECT 3.915000  1.435000 4.985000 1.765000 ;
      RECT 3.915000  1.765000 4.085000 1.935000 ;
      RECT 4.020000  0.085000 4.490000 0.905000 ;
      RECT 4.130000  2.775000 4.460000 3.245000 ;
      RECT 4.660000  0.575000 4.990000 0.755000 ;
      RECT 4.660000  0.755000 5.665000 0.770000 ;
      RECT 4.660000  0.770000 7.090000 0.925000 ;
      RECT 4.665000  1.935000 5.140000 2.095000 ;
      RECT 4.665000  2.095000 6.130000 2.265000 ;
      RECT 5.155000  1.265000 8.020000 1.280000 ;
      RECT 5.170000  0.085000 5.575000 0.585000 ;
      RECT 5.200000  2.775000 5.450000 3.245000 ;
      RECT 5.385000  1.450000 6.470000 1.780000 ;
      RECT 5.495000  0.925000 7.090000 0.940000 ;
      RECT 5.620000  2.605000 5.790000 2.710000 ;
      RECT 5.620000  2.710000 7.115000 2.980000 ;
      RECT 5.835000  0.255000 8.525000 0.425000 ;
      RECT 5.835000  0.425000 6.590000 0.600000 ;
      RECT 5.960000  2.265000 6.130000 2.370000 ;
      RECT 5.960000  2.370000 8.025000 2.540000 ;
      RECT 6.300000  1.780000 6.470000 1.950000 ;
      RECT 6.300000  1.950000 8.525000 2.200000 ;
      RECT 6.760000  0.595000 7.090000 0.770000 ;
      RECT 7.260000  0.425000 7.590000 0.940000 ;
      RECT 7.695000  2.540000 8.025000 2.980000 ;
      RECT 7.770000  0.595000 8.020000 1.110000 ;
      RECT 8.190000  0.425000 8.525000 1.030000 ;
      RECT 8.195000  2.200000 8.525000 2.980000 ;
      RECT 8.355000  1.030000 8.525000 1.950000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
  END
END sky130_fd_sc_hs__mux2_4
MACRO sky130_fd_sc_hs__mux2i_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.350000 2.865000 1.780000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.395000 1.180000 3.725000 1.550000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.488000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 0.550000 1.855000 ;
    END
  END S
  PIN Y
    ANTENNADIFFAREA  0.857700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.495000 0.705000 3.225000 1.035000 ;
        RECT 3.035000 1.035000 3.225000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.105000  2.100000 0.355000 3.245000 ;
      RECT 0.115000  0.085000 0.365000 0.905000 ;
      RECT 0.545000  0.405000 0.890000 0.905000 ;
      RECT 0.555000  2.100000 0.890000 2.980000 ;
      RECT 0.720000  0.905000 0.890000 1.350000 ;
      RECT 0.720000  1.350000 2.130000 1.520000 ;
      RECT 0.720000  1.520000 0.890000 2.100000 ;
      RECT 1.080000  1.820000 1.330000 1.950000 ;
      RECT 1.080000  1.950000 2.835000 2.120000 ;
      RECT 1.080000  2.120000 1.330000 2.980000 ;
      RECT 1.105000  0.350000 1.435000 1.010000 ;
      RECT 1.105000  1.010000 2.275000 1.180000 ;
      RECT 1.530000  2.290000 1.860000 3.245000 ;
      RECT 1.605000  0.085000 1.935000 0.840000 ;
      RECT 1.800000  1.520000 2.130000 1.680000 ;
      RECT 2.060000  2.290000 2.310000 2.905000 ;
      RECT 2.060000  2.905000 3.735000 3.075000 ;
      RECT 2.105000  0.350000 3.680000 0.520000 ;
      RECT 2.105000  0.520000 2.275000 1.010000 ;
      RECT 2.505000  2.120000 2.835000 2.735000 ;
      RECT 3.395000  0.520000 3.680000 1.010000 ;
      RECT 3.405000  1.820000 3.735000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__mux2i_1
MACRO sky130_fd_sc_hs__mux2i_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.180000 1.315000 1.550000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.535000 1.430000 3.235000 1.775000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.804000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.430000 4.675000 1.840000 ;
        RECT 4.350000 1.840000 5.810000 2.010000 ;
        RECT 5.480000 1.350000 5.810000 1.840000 ;
    END
  END S
  PIN Y
    ANTENNADIFFAREA  2.040950 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 2.910000 0.425000 ;
        RECT 0.085000 0.425000 0.450000 1.010000 ;
        RECT 0.085000 1.010000 0.255000 1.820000 ;
        RECT 0.085000 1.820000 0.445000 1.945000 ;
        RECT 0.085000 1.945000 2.845000 2.115000 ;
        RECT 0.085000 2.115000 0.445000 2.980000 ;
        RECT 2.580000 0.425000 2.910000 0.580000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.240000 0.085000 ;
      RECT 0.000000  3.245000 6.240000 3.415000 ;
      RECT 0.615000  2.285000 4.005000 2.340000 ;
      RECT 0.615000  2.340000 3.185000 2.455000 ;
      RECT 0.615000  2.455000 0.945000 2.980000 ;
      RECT 0.640000  0.595000 2.410000 0.750000 ;
      RECT 0.640000  0.750000 5.115000 0.765000 ;
      RECT 0.640000  0.765000 0.970000 1.010000 ;
      RECT 1.685000  2.625000 5.090000 2.680000 ;
      RECT 1.685000  2.680000 3.525000 2.795000 ;
      RECT 1.685000  2.795000 2.395000 2.955000 ;
      RECT 1.740000  0.935000 2.070000 1.090000 ;
      RECT 1.740000  1.090000 4.030000 1.260000 ;
      RECT 2.240000  0.765000 5.115000 0.830000 ;
      RECT 2.240000  0.830000 3.250000 0.920000 ;
      RECT 3.015000  2.010000 4.005000 2.285000 ;
      RECT 3.075000  2.965000 3.470000 3.245000 ;
      RECT 3.080000  0.660000 5.115000 0.750000 ;
      RECT 3.140000  0.085000 3.470000 0.490000 ;
      RECT 3.355000  2.510000 5.090000 2.625000 ;
      RECT 3.650000  1.000000 4.030000 1.090000 ;
      RECT 4.210000  0.085000 4.555000 0.490000 ;
      RECT 4.210000  2.850000 4.555000 3.245000 ;
      RECT 4.735000  0.500000 5.115000 0.660000 ;
      RECT 4.760000  2.180000 5.090000 2.510000 ;
      RECT 4.760000  2.680000 5.090000 2.980000 ;
      RECT 4.910000  1.010000 6.150000 1.180000 ;
      RECT 4.910000  1.180000 5.240000 1.670000 ;
      RECT 5.260000  2.180000 5.590000 3.245000 ;
      RECT 5.285000  0.085000 5.615000 0.840000 ;
      RECT 5.795000  0.570000 6.150000 1.010000 ;
      RECT 5.795000  2.180000 6.150000 2.860000 ;
      RECT 5.980000  1.180000 6.150000 2.180000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
  END
END sky130_fd_sc_hs__mux2i_2
MACRO sky130_fd_sc_hs__mux2i_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.225000 1.350000 3.235000 1.680000 ;
        RECT 2.525000 1.680000 3.235000 1.780000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 1.350000 1.885000 1.780000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  1.479000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.080000 1.180000 9.475000 1.540000 ;
    END
  END S
  PIN Y
    ANTENNADIFFAREA  2.868700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.405000 0.365000 1.010000 ;
        RECT 0.115000 1.010000 4.085000 1.180000 ;
        RECT 0.115000 1.180000 0.365000 1.185000 ;
        RECT 0.115000 1.820000 0.365000 1.950000 ;
        RECT 0.115000 1.950000 4.245000 2.120000 ;
        RECT 0.115000 2.120000 0.365000 2.980000 ;
        RECT 1.055000 0.595000 1.225000 1.010000 ;
        RECT 1.095000 2.120000 1.265000 2.735000 ;
        RECT 1.915000 2.120000 2.245000 2.735000 ;
        RECT 1.920000 0.595000 2.250000 0.935000 ;
        RECT 1.920000 0.935000 4.085000 1.010000 ;
        RECT 2.915000 2.120000 3.245000 2.395000 ;
        RECT 3.485000 1.550000 4.245000 1.950000 ;
        RECT 3.915000 1.180000 4.085000 1.550000 ;
        RECT 3.915000 2.120000 4.245000 2.395000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.545000  0.255000  4.765000 0.425000 ;
      RECT 0.545000  0.425000  0.875000 0.840000 ;
      RECT 0.565000  2.290000  0.895000 2.905000 ;
      RECT 0.565000  2.905000  6.560000 3.075000 ;
      RECT 1.405000  0.425000  1.735000 0.840000 ;
      RECT 1.465000  2.290000  1.715000 2.905000 ;
      RECT 2.415000  2.290000  2.745000 2.565000 ;
      RECT 2.415000  2.565000  5.130000 2.735000 ;
      RECT 2.420000  0.595000  4.425000 0.765000 ;
      RECT 3.415000  2.290000  3.745000 2.565000 ;
      RECT 4.255000  0.765000  4.425000 1.000000 ;
      RECT 4.255000  1.000000  6.715000 1.170000 ;
      RECT 4.475000  1.840000  6.080000 2.050000 ;
      RECT 4.475000  2.050000  9.010000 2.220000 ;
      RECT 4.595000  0.425000  4.765000 0.660000 ;
      RECT 4.595000  0.660000  7.735000 0.750000 ;
      RECT 4.595000  0.750000  5.525000 0.830000 ;
      RECT 4.935000  0.085000  5.185000 0.490000 ;
      RECT 4.960000  2.390000  8.560000 2.560000 ;
      RECT 4.960000  2.560000  5.130000 2.565000 ;
      RECT 5.150000  1.340000  6.840000 1.670000 ;
      RECT 5.300000  2.730000  6.560000 2.905000 ;
      RECT 5.355000  0.580000  7.735000 0.660000 ;
      RECT 5.875000  0.085000  6.205000 0.410000 ;
      RECT 6.385000  0.920000  6.715000 1.000000 ;
      RECT 6.670000  1.670000  6.840000 1.710000 ;
      RECT 6.670000  1.710000  9.825000 1.880000 ;
      RECT 6.730000  2.730000  7.060000 3.245000 ;
      RECT 6.895000  0.085000  7.225000 0.410000 ;
      RECT 7.230000  2.560000  7.560000 2.980000 ;
      RECT 7.405000  0.390000  7.735000 0.580000 ;
      RECT 7.405000  0.750000  7.735000 0.840000 ;
      RECT 7.405000  0.840000  8.825000 1.010000 ;
      RECT 7.730000  2.730000  8.060000 3.245000 ;
      RECT 7.905000  0.085000  8.325000 0.640000 ;
      RECT 8.230000  2.560000  8.560000 2.980000 ;
      RECT 8.495000  0.390000  8.825000 0.840000 ;
      RECT 8.760000  2.220000  9.010000 3.245000 ;
      RECT 8.995000  0.085000  9.325000 1.010000 ;
      RECT 9.185000  1.880000  9.455000 2.700000 ;
      RECT 9.495000  0.390000  9.825000 1.010000 ;
      RECT 9.635000  2.050000  9.965000 3.245000 ;
      RECT 9.655000  1.010000  9.825000 1.710000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
  END
END sky130_fd_sc_hs__mux2i_4
MACRO sky130_fd_sc_hs__mux4_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.600000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.990000 1.215000 1.320000 1.780000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.000000 1.215000 3.330000 2.150000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.500000 1.215000 3.870000 2.150000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.850000 1.445000 6.180000 1.780000 ;
    END
  END A3
  PIN S0
    ANTENNAGATEAREA  0.738000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.450000 1.215000 0.820000 1.780000 ;
    END
  END S0
  PIN S1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.205000 1.350000 8.535000 1.780000 ;
    END
  END S1
  PIN X
    ANTENNADIFFAREA  0.558100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.080000 0.400000 9.485000 1.180000 ;
        RECT 9.220000 2.560000 9.485000 2.890000 ;
        RECT 9.245000 1.180000 9.485000 2.560000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.600000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.600000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.600000 0.085000 ;
      RECT 0.000000  3.245000 9.600000 3.415000 ;
      RECT 0.110000  0.350000 0.445000 0.860000 ;
      RECT 0.110000  0.860000 1.700000 1.030000 ;
      RECT 0.110000  1.030000 0.280000 1.950000 ;
      RECT 0.110000  1.950000 0.555000 2.880000 ;
      RECT 0.700000  0.085000 1.090000 0.680000 ;
      RECT 0.725000  1.950000 1.055000 3.245000 ;
      RECT 1.530000  0.255000 2.630000 0.425000 ;
      RECT 1.530000  0.425000 1.700000 0.860000 ;
      RECT 1.530000  1.030000 1.700000 1.200000 ;
      RECT 1.530000  1.200000 1.860000 1.530000 ;
      RECT 1.875000  0.595000 2.200000 1.030000 ;
      RECT 2.030000  1.030000 2.200000 1.685000 ;
      RECT 2.030000  1.685000 2.550000 2.335000 ;
      RECT 2.030000  2.335000 4.020000 2.505000 ;
      RECT 2.030000  2.505000 2.550000 2.725000 ;
      RECT 2.460000  0.425000 2.630000 0.875000 ;
      RECT 2.460000  0.875000 4.750000 1.045000 ;
      RECT 2.460000  1.045000 2.790000 1.450000 ;
      RECT 3.125000  0.085000 3.715000 0.680000 ;
      RECT 3.265000  2.675000 3.595000 3.245000 ;
      RECT 3.795000  2.505000 4.020000 2.905000 ;
      RECT 3.795000  2.905000 5.550000 3.075000 ;
      RECT 4.080000  1.045000 4.410000 1.450000 ;
      RECT 4.210000  0.375000 5.090000 0.705000 ;
      RECT 4.305000  1.995000 5.680000 2.165000 ;
      RECT 4.305000  2.165000 5.165000 2.735000 ;
      RECT 4.580000  1.045000 4.750000 1.445000 ;
      RECT 4.580000  1.445000 5.340000 1.775000 ;
      RECT 4.920000  0.705000 5.090000 1.105000 ;
      RECT 4.920000  1.105000 6.235000 1.275000 ;
      RECT 5.260000  0.085000 5.590000 0.935000 ;
      RECT 5.350000  2.335000 6.620000 2.505000 ;
      RECT 5.350000  2.505000 5.550000 2.905000 ;
      RECT 5.510000  1.275000 5.680000 1.995000 ;
      RECT 5.730000  2.675000 6.060000 3.245000 ;
      RECT 5.985000  0.265000 7.695000 0.435000 ;
      RECT 5.985000  0.435000 6.485000 0.445000 ;
      RECT 5.985000  0.445000 6.235000 1.105000 ;
      RECT 6.290000  1.950000 6.620000 2.335000 ;
      RECT 6.290000  2.505000 6.620000 2.980000 ;
      RECT 6.405000  0.615000 7.355000 0.785000 ;
      RECT 6.405000  0.785000 6.575000 1.950000 ;
      RECT 6.745000  0.955000 6.925000 1.115000 ;
      RECT 6.745000  1.115000 7.120000 1.285000 ;
      RECT 6.790000  1.285000 7.120000 2.905000 ;
      RECT 6.790000  2.905000 8.520000 3.075000 ;
      RECT 7.105000  0.605000 7.355000 0.615000 ;
      RECT 7.105000  0.785000 7.355000 0.935000 ;
      RECT 7.290000  1.105000 7.695000 1.275000 ;
      RECT 7.290000  1.275000 7.460000 1.945000 ;
      RECT 7.290000  1.945000 7.620000 2.735000 ;
      RECT 7.525000  0.435000 7.695000 1.105000 ;
      RECT 7.630000  1.445000 8.035000 1.775000 ;
      RECT 7.850000  1.775000 8.035000 1.950000 ;
      RECT 7.850000  1.950000 8.180000 2.735000 ;
      RECT 7.865000  0.500000 8.410000 1.180000 ;
      RECT 7.865000  1.180000 8.035000 1.445000 ;
      RECT 8.350000  1.950000 8.915000 2.120000 ;
      RECT 8.350000  2.120000 8.520000 2.905000 ;
      RECT 8.580000  0.085000 8.910000 1.180000 ;
      RECT 8.690000  2.290000 9.020000 3.245000 ;
      RECT 8.745000  1.350000 9.075000 1.680000 ;
      RECT 8.745000  1.680000 8.915000 1.950000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
  END
END sky130_fd_sc_hs__mux4_1
MACRO sky130_fd_sc_hs__mux4_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.56000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.315000 1.450000 3.685000 1.780000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.975000 1.450000 1.315000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.915000 1.180000 6.345000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.855000 1.450000 4.195000 1.780000 ;
    END
  END A3
  PIN S0
    ANTENNAGATEAREA  0.768000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.435000 1.180000 1.655000 1.260000 ;
        RECT 0.435000 1.260000 1.845000 1.280000 ;
        RECT 0.435000 1.280000 0.805000 1.550000 ;
        RECT 0.635000 1.110000 1.655000 1.180000 ;
        RECT 1.485000 0.420000 3.105000 0.590000 ;
        RECT 1.485000 0.590000 1.655000 1.110000 ;
        RECT 1.485000 1.280000 1.845000 1.590000 ;
        RECT 2.835000 0.590000 3.105000 1.110000 ;
        RECT 2.835000 1.110000 5.745000 1.280000 ;
        RECT 2.835000 1.280000 3.105000 1.780000 ;
        RECT 4.395000 1.280000 4.725000 1.550000 ;
        RECT 5.475000 1.280000 5.745000 1.750000 ;
    END
  END S0
  PIN S1
    ANTENNAGATEAREA  0.507000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.900000 1.450000 7.555000 1.780000 ;
    END
  END S1
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.650000 0.440000  9.980000 1.820000 ;
        RECT 9.650000 1.820000 10.000000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.560000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.560000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 10.560000 0.085000 ;
      RECT  0.000000  3.245000 10.560000 3.415000 ;
      RECT  0.095000  0.500000  0.465000 1.010000 ;
      RECT  0.095000  1.010000  0.265000 1.920000 ;
      RECT  0.095000  1.920000  0.585000 2.150000 ;
      RECT  0.255000  2.150000  0.585000 2.980000 ;
      RECT  0.755000  1.950000  1.085000 3.245000 ;
      RECT  0.820000  0.085000  1.150000 0.940000 ;
      RECT  1.850000  0.760000  2.665000 1.090000 ;
      RECT  2.045000  1.450000  2.325000 2.150000 ;
      RECT  2.495000  1.090000  2.665000 1.950000 ;
      RECT  2.495000  1.950000  4.285000 2.120000 ;
      RECT  2.495000  2.120000  3.445000 2.980000 ;
      RECT  3.445000  0.085000  3.925000 0.940000 ;
      RECT  3.615000  2.290000  3.945000 3.245000 ;
      RECT  4.115000  2.120000  4.285000 2.320000 ;
      RECT  4.115000  2.320000  5.605000 2.490000 ;
      RECT  4.530000  0.350000  5.105000 0.770000 ;
      RECT  4.530000  0.770000  8.015000 0.940000 ;
      RECT  4.925000  1.460000  5.265000 2.150000 ;
      RECT  5.055000  2.660000  5.945000 2.910000 ;
      RECT  5.435000  1.960000  7.080000 2.200000 ;
      RECT  5.435000  2.200000  5.605000 2.320000 ;
      RECT  5.775000  2.370000  7.980000 2.540000 ;
      RECT  5.775000  2.540000  5.945000 2.660000 ;
      RECT  6.140000  0.085000  6.470000 0.600000 ;
      RECT  6.165000  2.710000  6.495000 3.245000 ;
      RECT  6.560000  1.110000  7.955000 1.280000 ;
      RECT  6.560000  1.280000  6.730000 1.950000 ;
      RECT  6.560000  1.950000  7.080000 1.960000 ;
      RECT  6.690000  0.350000  6.940000 0.770000 ;
      RECT  7.120000  0.255000  9.130000 0.425000 ;
      RECT  7.120000  0.425000  7.450000 0.600000 ;
      RECT  7.200000  2.710000  7.530000 2.905000 ;
      RECT  7.200000  2.905000  9.130000 3.075000 ;
      RECT  7.650000  1.950000  7.980000 2.370000 ;
      RECT  7.725000  1.450000  8.450000 1.780000 ;
      RECT  7.810000  2.540000  7.980000 2.565000 ;
      RECT  7.810000  2.565000  8.790000 2.735000 ;
      RECT  7.845000  0.595000  8.790000 0.765000 ;
      RECT  7.845000  0.765000  8.015000 0.770000 ;
      RECT  8.185000  0.935000  8.450000 1.450000 ;
      RECT  8.200000  1.780000  8.450000 2.395000 ;
      RECT  8.620000  0.765000  8.790000 2.565000 ;
      RECT  8.960000  0.425000  9.130000 1.350000 ;
      RECT  8.960000  1.350000  9.385000 1.680000 ;
      RECT  8.960000  1.680000  9.130000 2.905000 ;
      RECT  9.300000  0.085000  9.470000 1.180000 ;
      RECT  9.300000  1.850000  9.470000 3.245000 ;
      RECT 10.160000  0.085000 10.410000 1.260000 ;
      RECT 10.200000  1.820000 10.450000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  1.950000  0.325000 2.120000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  1.950000  2.245000 2.120000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  1.950000  5.125000 2.120000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
    LAYER met1 ;
      RECT 0.095000 1.920000 0.385000 1.965000 ;
      RECT 0.095000 1.965000 5.185000 2.105000 ;
      RECT 0.095000 2.105000 0.385000 2.150000 ;
      RECT 2.015000 1.920000 2.305000 1.965000 ;
      RECT 2.015000 2.105000 2.305000 2.150000 ;
      RECT 4.895000 1.920000 5.185000 1.965000 ;
      RECT 4.895000 2.105000 5.185000 2.150000 ;
  END
END sky130_fd_sc_hs__mux4_2
MACRO sky130_fd_sc_hs__mux4_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  16.80000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.470000 2.355000 1.800000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.450000 0.890000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.765000 1.260000 9.475000 1.775000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.725000 1.445000 10.435000 1.775000 ;
    END
  END A3
  PIN S0
    ANTENNAGATEAREA  1.263000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.295000 1.435000 8.515000 1.775000 ;
    END
  END S0
  PIN S1
    ANTENNAGATEAREA  0.771000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.150000 1.275000 13.865000 1.300000 ;
        RECT 12.150000 1.300000 12.835000 1.780000 ;
        RECT 12.665000 1.130000 13.865000 1.275000 ;
        RECT 13.540000 1.300000 13.865000 1.550000 ;
    END
  END S1
  PIN X
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.875000 1.800000 16.675000 1.970000 ;
        RECT 14.875000 1.970000 15.205000 2.980000 ;
        RECT 15.065000 0.350000 15.315000 0.960000 ;
        RECT 15.065000 0.960000 16.675000 1.130000 ;
        RECT 15.825000 1.970000 16.155000 2.980000 ;
        RECT 15.925000 0.350000 16.175000 0.960000 ;
        RECT 16.445000 1.130000 16.675000 1.800000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 16.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 16.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 16.800000 0.085000 ;
      RECT  0.000000  3.245000 16.800000 3.415000 ;
      RECT  0.115000  0.085000  0.365000 1.030000 ;
      RECT  0.115000  1.030000  1.370000 1.280000 ;
      RECT  0.115000  1.950000  0.365000 3.245000 ;
      RECT  0.545000  0.275000  1.810000 0.470000 ;
      RECT  0.545000  0.470000  0.875000 0.860000 ;
      RECT  0.565000  1.950000  0.895000 1.970000 ;
      RECT  0.565000  1.970000  2.695000 2.140000 ;
      RECT  0.565000  2.140000  0.895000 2.980000 ;
      RECT  1.045000  0.640000  1.370000 1.030000 ;
      RECT  1.095000  2.310000  1.345000 3.245000 ;
      RECT  1.515000  2.310000  3.300000 2.480000 ;
      RECT  1.515000  2.480000  1.845000 2.980000 ;
      RECT  1.550000  0.960000  1.800000 1.130000 ;
      RECT  1.550000  1.130000  2.695000 1.260000 ;
      RECT  1.550000  1.260000  4.205000 1.300000 ;
      RECT  1.575000  0.470000  1.810000 0.620000 ;
      RECT  1.575000  0.620000  2.140000 0.790000 ;
      RECT  1.970000  0.790000  3.380000 0.960000 ;
      RECT  1.980000  0.085000  2.310000 0.450000 ;
      RECT  2.045000  2.650000  2.295000 3.245000 ;
      RECT  2.525000  1.300000  4.205000 1.430000 ;
      RECT  2.525000  1.600000  4.190000 1.770000 ;
      RECT  2.525000  1.770000  2.695000 1.970000 ;
      RECT  2.525000  2.650000  2.860000 2.905000 ;
      RECT  2.525000  2.905000  4.720000 3.075000 ;
      RECT  2.540000  0.255000  4.715000 0.425000 ;
      RECT  2.540000  0.425000  2.870000 0.620000 ;
      RECT  2.990000  1.940000  3.300000 2.310000 ;
      RECT  3.045000  2.480000  3.300000 2.735000 ;
      RECT  3.050000  0.595000  3.380000 0.790000 ;
      RECT  3.050000  0.960000  3.380000 1.090000 ;
      RECT  3.490000  1.940000  3.820000 2.905000 ;
      RECT  3.605000  0.425000  3.775000 1.090000 ;
      RECT  3.955000  0.595000  4.205000 1.260000 ;
      RECT  4.020000  1.770000  4.190000 2.735000 ;
      RECT  4.375000  0.425000  4.715000 1.180000 ;
      RECT  4.375000  1.180000  4.545000 1.920000 ;
      RECT  4.375000  1.920000  4.720000 2.905000 ;
      RECT  4.715000  1.350000  5.200000 1.365000 ;
      RECT  4.715000  1.365000  6.705000 1.535000 ;
      RECT  4.715000  1.535000  5.200000 1.680000 ;
      RECT  4.945000  0.350000  5.200000 1.350000 ;
      RECT  4.950000  1.680000  5.200000 2.980000 ;
      RECT  5.375000  0.085000  5.705000 1.130000 ;
      RECT  5.400000  1.820000  5.730000 3.245000 ;
      RECT  5.935000  0.585000  6.185000 1.025000 ;
      RECT  5.935000  1.025000  7.125000 1.195000 ;
      RECT  5.960000  1.865000  7.125000 1.945000 ;
      RECT  5.960000  1.945000 10.975000 2.035000 ;
      RECT  5.960000  2.035000  6.210000 2.905000 ;
      RECT  6.035000  1.535000  6.705000 1.695000 ;
      RECT  6.365000  0.255000  8.325000 0.425000 ;
      RECT  6.365000  0.425000  6.695000 0.855000 ;
      RECT  6.410000  2.205000  6.740000 2.905000 ;
      RECT  6.410000  2.905000  8.150000 3.075000 ;
      RECT  6.875000  0.595000  7.985000 0.765000 ;
      RECT  6.875000  0.765000  7.125000 1.025000 ;
      RECT  6.875000  1.195000  7.125000 1.265000 ;
      RECT  6.940000  1.265000  7.125000 1.865000 ;
      RECT  6.940000  2.035000 10.975000 2.115000 ;
      RECT  6.940000  2.115000  7.125000 2.735000 ;
      RECT  7.305000  0.935000  7.555000 1.095000 ;
      RECT  7.305000  1.095000  8.325000 1.265000 ;
      RECT  7.310000  2.285000  9.185000 2.455000 ;
      RECT  7.310000  2.455000  7.640000 2.735000 ;
      RECT  7.735000  0.765000  7.985000 0.925000 ;
      RECT  7.980000  2.625000 10.265000 2.795000 ;
      RECT  7.980000  2.795000  8.150000 2.905000 ;
      RECT  8.155000  0.425000  8.325000 0.580000 ;
      RECT  8.155000  0.580000  9.255000 0.750000 ;
      RECT  8.155000  0.920000 10.115000 1.090000 ;
      RECT  8.155000  1.090000  8.325000 1.095000 ;
      RECT  8.320000  2.965000  8.650000 3.245000 ;
      RECT  8.495000  0.085000  8.825000 0.410000 ;
      RECT  9.005000  0.350000  9.255000 0.580000 ;
      RECT  9.390000  2.965000  9.730000 3.245000 ;
      RECT  9.435000  0.085000  9.685000 0.750000 ;
      RECT  9.865000  0.350000 10.115000 0.920000 ;
      RECT  9.935000  2.285000 10.265000 2.625000 ;
      RECT  9.935000  2.795000 10.265000 2.980000 ;
      RECT 10.295000  0.085000 10.545000 1.030000 ;
      RECT 10.465000  2.285000 10.635000 3.245000 ;
      RECT 10.715000  0.255000 11.815000 0.425000 ;
      RECT 10.715000  0.425000 10.885000 1.945000 ;
      RECT 10.805000  2.115000 10.975000 2.905000 ;
      RECT 10.805000  2.905000 12.975000 3.075000 ;
      RECT 11.055000  0.595000 12.675000 0.620000 ;
      RECT 11.055000  0.620000 12.155000 0.765000 ;
      RECT 11.055000  0.765000 11.475000 1.030000 ;
      RECT 11.145000  1.030000 11.475000 2.565000 ;
      RECT 11.145000  2.565000 12.475000 2.735000 ;
      RECT 11.645000  0.935000 13.175000 0.960000 ;
      RECT 11.645000  0.960000 12.495000 1.105000 ;
      RECT 11.645000  1.105000 11.975000 2.395000 ;
      RECT 11.985000  0.255000 14.545000 0.425000 ;
      RECT 11.985000  0.425000 12.675000 0.595000 ;
      RECT 12.145000  1.950000 12.475000 2.060000 ;
      RECT 12.145000  2.060000 13.475000 2.230000 ;
      RECT 12.145000  2.230000 12.475000 2.565000 ;
      RECT 12.325000  0.790000 13.175000 0.935000 ;
      RECT 12.645000  2.400000 12.975000 2.905000 ;
      RECT 12.860000  0.595000 13.175000 0.790000 ;
      RECT 13.005000  1.470000 13.330000 1.720000 ;
      RECT 13.005000  1.720000 14.205000 1.890000 ;
      RECT 13.145000  2.230000 13.475000 2.980000 ;
      RECT 13.345000  0.425000 13.675000 0.960000 ;
      RECT 13.875000  1.890000 14.205000 2.980000 ;
      RECT 13.905000  0.595000 14.205000 0.960000 ;
      RECT 14.035000  0.960000 14.205000 1.720000 ;
      RECT 14.375000  0.425000 14.545000 1.300000 ;
      RECT 14.375000  1.300000 16.210000 1.630000 ;
      RECT 14.375000  1.820000 14.705000 3.245000 ;
      RECT 14.715000  0.085000 14.885000 1.130000 ;
      RECT 15.405000  2.140000 15.655000 3.245000 ;
      RECT 15.495000  0.085000 15.745000 0.790000 ;
      RECT 16.325000  2.140000 16.655000 3.245000 ;
      RECT 16.355000  0.085000 16.685000 0.790000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  1.950000  4.645000 2.120000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  1.950000 11.845000 2.120000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.245000 15.205000 3.415000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.245000 15.685000 3.415000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.245000 16.165000 3.415000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  3.245000 16.645000 3.415000 ;
    LAYER met1 ;
      RECT  4.415000 1.920000  4.705000 1.965000 ;
      RECT  4.415000 1.965000 11.905000 2.105000 ;
      RECT  4.415000 2.105000  4.705000 2.150000 ;
      RECT 11.615000 1.920000 11.905000 1.965000 ;
      RECT 11.615000 2.105000 11.905000 2.150000 ;
  END
END sky130_fd_sc_hs__mux4_4
MACRO sky130_fd_sc_hs__nand2_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.440000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.180000 1.335000 1.550000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.435000 1.550000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.546900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.180000 0.835000 2.980000 ;
        RECT 0.665000 0.840000 1.280000 1.010000 ;
        RECT 0.665000 1.010000 0.835000 1.180000 ;
        RECT 0.950000 0.350000 1.280000 0.840000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 1.440000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 1.440000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.440000 0.085000 ;
      RECT 0.000000  3.245000 1.440000 3.415000 ;
      RECT 0.105000  1.820000 0.435000 3.245000 ;
      RECT 0.130000  0.085000 0.460000 1.010000 ;
      RECT 1.005000  1.820000 1.335000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
  END
END sky130_fd_sc_hs__nand2_1
MACRO sky130_fd_sc_hs__nand2_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.400000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 1.350000 1.815000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.350000 1.315000 1.780000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.916200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.570000 1.950000 2.275000 2.120000 ;
        RECT 0.570000 2.120000 0.820000 2.980000 ;
        RECT 1.455000 0.595000 1.785000 1.010000 ;
        RECT 1.455000 1.010000 2.275000 1.180000 ;
        RECT 1.560000 2.120000 1.730000 2.980000 ;
        RECT 2.045000 1.180000 2.275000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.400000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.400000 0.085000 ;
      RECT 0.000000  3.245000 2.400000 3.415000 ;
      RECT 0.115000  0.350000 0.365000 1.010000 ;
      RECT 0.115000  1.010000 1.275000 1.180000 ;
      RECT 0.120000  1.820000 0.370000 3.245000 ;
      RECT 0.545000  0.085000 0.875000 0.840000 ;
      RECT 1.020000  2.290000 1.350000 3.245000 ;
      RECT 1.105000  0.255000 2.285000 0.425000 ;
      RECT 1.105000  0.425000 1.275000 1.010000 ;
      RECT 1.930000  2.290000 2.260000 3.245000 ;
      RECT 1.955000  0.425000 2.285000 0.840000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
  END
END sky130_fd_sc_hs__nand2_2
MACRO sky130_fd_sc_hs__nand2_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 1.350000 3.795000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.510000 1.350000 2.275000 1.680000 ;
        RECT 1.085000 1.680000 2.275000 1.780000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  3.286100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.615000 1.950000 4.195000 2.120000 ;
        RECT 0.615000 2.120000 1.660000 2.980000 ;
        RECT 2.330000 2.120000 3.705000 2.980000 ;
        RECT 2.335000 0.610000 2.665000 1.010000 ;
        RECT 2.335000 1.010000 4.195000 1.180000 ;
        RECT 3.335000 0.610000 3.705000 1.010000 ;
        RECT 3.965000 1.180000 4.195000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  0.350000 0.365000 1.010000 ;
      RECT 0.115000  1.010000 2.165000 1.180000 ;
      RECT 0.115000  1.850000 0.445000 3.245000 ;
      RECT 0.545000  0.085000 0.875000 0.805000 ;
      RECT 1.055000  0.350000 1.225000 1.010000 ;
      RECT 1.405000  0.085000 1.735000 0.805000 ;
      RECT 1.830000  2.290000 2.160000 3.245000 ;
      RECT 1.915000  0.255000 4.205000 0.425000 ;
      RECT 1.915000  0.425000 2.165000 1.010000 ;
      RECT 2.835000  0.425000 3.165000 0.805000 ;
      RECT 3.875000  0.425000 4.205000 0.805000 ;
      RECT 3.875000  2.290000 4.205000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__nand2_4
MACRO sky130_fd_sc_hs__nand2_8
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.560000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.185000 1.220000 7.555000 1.550000 ;
        RECT 5.965000 1.550000 7.555000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.560000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.350000 4.195000 1.780000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  2.284800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.140000 1.950000 4.710000 2.120000 ;
        RECT 2.140000 2.120000 2.470000 2.980000 ;
        RECT 4.335000 0.770000 7.895000 1.050000 ;
        RECT 4.335000 1.050000 4.710000 1.130000 ;
        RECT 4.380000 1.130000 4.710000 1.950000 ;
        RECT 4.380000 2.120000 4.710000 2.980000 ;
        RECT 5.940000 1.950000 7.895000 2.120000 ;
        RECT 5.940000 2.120000 6.270000 2.980000 ;
        RECT 7.320000 2.120000 7.550000 2.980000 ;
        RECT 7.725000 1.050000 7.895000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.105000  0.350000 0.355000 1.165000 ;
      RECT 0.105000  1.165000 4.155000 1.180000 ;
      RECT 0.105000  1.180000 1.860000 1.355000 ;
      RECT 0.535000  0.085000 0.865000 0.995000 ;
      RECT 0.660000  1.950000 1.970000 3.245000 ;
      RECT 1.035000  0.350000 1.225000 1.010000 ;
      RECT 1.035000  1.010000 4.155000 1.165000 ;
      RECT 1.395000  0.085000 1.725000 0.840000 ;
      RECT 1.895000  0.350000 2.155000 1.010000 ;
      RECT 2.325000  0.085000 2.905000 0.840000 ;
      RECT 2.640000  2.290000 4.210000 3.245000 ;
      RECT 3.075000  0.350000 3.305000 1.010000 ;
      RECT 3.475000  0.085000 3.805000 0.840000 ;
      RECT 3.985000  0.350000 8.045000 0.600000 ;
      RECT 3.985000  0.600000 4.155000 1.010000 ;
      RECT 4.880000  1.820000 5.210000 3.245000 ;
      RECT 5.440000  1.820000 5.770000 3.245000 ;
      RECT 6.440000  2.290000 7.150000 3.245000 ;
      RECT 7.720000  2.290000 8.050000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_hs__nand2_8
MACRO sky130_fd_sc_hs__nand2b_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.400000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.300000 0.835000 1.780000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015000 1.350000 1.345000 1.780000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.710200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 2.290000 2.255000 2.460000 ;
        RECT 1.085000 2.460000 1.565000 2.980000 ;
        RECT 1.855000 0.350000 2.255000 1.130000 ;
        RECT 2.085000 1.130000 2.255000 2.290000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.400000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.400000 0.085000 ;
      RECT 0.000000  3.245000 2.400000 3.415000 ;
      RECT 0.115000  0.540000 0.380000 0.960000 ;
      RECT 0.115000  0.960000 1.685000 1.130000 ;
      RECT 0.115000  1.950000 1.685000 2.120000 ;
      RECT 0.115000  2.120000 0.445000 2.700000 ;
      RECT 0.550000  0.085000 1.220000 0.790000 ;
      RECT 0.650000  2.290000 0.915000 3.245000 ;
      RECT 1.515000  1.130000 1.685000 1.300000 ;
      RECT 1.515000  1.300000 1.915000 1.630000 ;
      RECT 1.515000  1.630000 1.685000 1.950000 ;
      RECT 1.735000  2.650000 2.070000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
  END
END sky130_fd_sc_hs__nand2b_1
MACRO sky130_fd_sc_hs__nand2b_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 0.570000 1.780000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 1.350000 2.775000 1.780000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.879200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.645000 1.820000 2.275000 1.950000 ;
        RECT 1.645000 1.950000 2.795000 2.200000 ;
        RECT 1.700000 0.630000 1.870000 1.220000 ;
        RECT 1.700000 1.220000 2.275000 1.390000 ;
        RECT 2.045000 1.390000 2.275000 1.820000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.115000  0.350000 0.445000 1.010000 ;
      RECT 0.115000  1.010000 0.975000 1.140000 ;
      RECT 0.115000  1.140000 1.135000 1.180000 ;
      RECT 0.115000  1.950000 0.975000 2.120000 ;
      RECT 0.115000  2.120000 0.445000 2.860000 ;
      RECT 0.615000  0.085000 0.875000 0.840000 ;
      RECT 0.725000  2.290000 1.095000 3.245000 ;
      RECT 0.805000  1.180000 1.135000 1.470000 ;
      RECT 0.805000  1.470000 0.975000 1.950000 ;
      RECT 1.190000  0.255000 2.380000 0.425000 ;
      RECT 1.190000  0.425000 1.520000 0.970000 ;
      RECT 1.305000  0.970000 1.475000 2.370000 ;
      RECT 1.305000  2.370000 3.245000 2.540000 ;
      RECT 2.015000  2.710000 2.345000 3.245000 ;
      RECT 2.050000  0.425000 2.380000 1.050000 ;
      RECT 2.560000  0.085000 2.730000 1.130000 ;
      RECT 2.915000  0.350000 3.245000 1.130000 ;
      RECT 2.915000  2.710000 3.245000 3.245000 ;
      RECT 3.075000  1.130000 3.245000 2.370000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__nand2b_2
MACRO sky130_fd_sc_hs__nand2b_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.363000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.300000 1.115000 1.780000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.845000 1.300000 5.655000 1.630000 ;
        RECT 4.445000 1.630000 5.655000 1.780000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.634300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.625000 0.635000 1.885000 1.090000 ;
        RECT 1.625000 1.090000 3.655000 1.260000 ;
        RECT 2.265000 1.850000 4.195000 1.950000 ;
        RECT 2.265000 1.950000 5.145000 2.150000 ;
        RECT 2.265000 2.150000 2.875000 2.980000 ;
        RECT 2.555000 0.635000 2.880000 1.090000 ;
        RECT 3.285000 1.260000 3.655000 1.850000 ;
        RECT 4.815000 2.150000 5.145000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.135000  0.350000 0.385000 0.960000 ;
      RECT 0.135000  0.960000 1.455000 1.130000 ;
      RECT 0.435000  1.950000 1.060000 3.245000 ;
      RECT 0.565000  0.085000 0.895000 0.790000 ;
      RECT 1.195000  0.255000 3.380000 0.425000 ;
      RECT 1.195000  0.425000 1.455000 0.790000 ;
      RECT 1.230000  1.950000 1.560000 2.700000 ;
      RECT 1.285000  1.130000 1.455000 1.430000 ;
      RECT 1.285000  1.430000 3.075000 1.680000 ;
      RECT 1.285000  1.680000 1.455000 1.950000 ;
      RECT 1.765000  1.850000 2.095000 3.245000 ;
      RECT 2.055000  0.425000 2.385000 0.920000 ;
      RECT 3.045000  2.320000 4.645000 3.245000 ;
      RECT 3.050000  0.425000 3.380000 0.750000 ;
      RECT 3.050000  0.750000 4.310000 0.920000 ;
      RECT 3.550000  0.085000 3.880000 0.580000 ;
      RECT 3.980000  0.920000 4.310000 0.960000 ;
      RECT 3.980000  0.960000 5.645000 1.130000 ;
      RECT 4.050000  0.330000 4.310000 0.750000 ;
      RECT 4.480000  0.085000 5.145000 0.790000 ;
      RECT 5.315000  0.350000 5.645000 0.960000 ;
      RECT 5.315000  1.950000 5.600000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_hs__nand2b_4
MACRO sky130_fd_sc_hs__nand3_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.400000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.180000 1.915000 1.550000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015000 0.440000 1.345000 1.550000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.835000 1.550000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.877300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.720000 2.255000 1.890000 ;
        RECT 0.605000 1.890000 1.045000 2.980000 ;
        RECT 1.710000 0.350000 2.040000 0.840000 ;
        RECT 1.710000 0.840000 2.255000 1.010000 ;
        RECT 1.735000 1.890000 2.255000 2.980000 ;
        RECT 2.085000 1.010000 2.255000 1.720000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.400000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.400000 0.085000 ;
      RECT 0.000000  3.245000 2.400000 3.415000 ;
      RECT 0.185000  1.820000 0.435000 3.245000 ;
      RECT 0.320000  0.085000 0.650000 1.010000 ;
      RECT 1.215000  2.060000 1.545000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
  END
END sky130_fd_sc_hs__nand3_1
MACRO sky130_fd_sc_hs__nand3_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965000 1.430000 2.295000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.265000 1.430000 1.595000 1.550000 ;
        RECT 1.265000 1.550000 1.795000 1.680000 ;
        RECT 1.425000 1.680000 1.795000 1.950000 ;
        RECT 1.425000 1.950000 2.825000 2.120000 ;
        RECT 2.655000 1.320000 3.065000 1.650000 ;
        RECT 2.655000 1.650000 2.825000 1.950000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 0.735000 1.550000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  1.220800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565000 1.820000 1.095000 2.290000 ;
        RECT 0.565000 2.290000 2.795000 2.460000 ;
        RECT 0.565000 2.460000 0.895000 2.980000 ;
        RECT 0.925000 1.090000 2.275000 1.260000 ;
        RECT 0.925000 1.260000 1.095000 1.820000 ;
        RECT 1.515000 2.460000 1.845000 2.980000 ;
        RECT 1.945000 0.935000 2.275000 1.090000 ;
        RECT 2.525000 2.460000 2.795000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.100000  0.350000 0.350000 0.750000 ;
      RECT 0.100000  0.750000 3.260000 0.765000 ;
      RECT 0.100000  0.765000 1.370000 0.920000 ;
      RECT 0.100000  0.920000 0.430000 1.010000 ;
      RECT 0.115000  1.820000 0.365000 3.245000 ;
      RECT 0.530000  0.085000 0.860000 0.580000 ;
      RECT 1.040000  0.330000 1.210000 0.595000 ;
      RECT 1.040000  0.595000 3.260000 0.750000 ;
      RECT 1.065000  2.630000 1.315000 3.245000 ;
      RECT 1.455000  0.255000 2.765000 0.425000 ;
      RECT 2.015000  2.630000 2.345000 3.245000 ;
      RECT 2.930000  0.765000 3.260000 1.150000 ;
      RECT 2.945000  0.405000 3.260000 0.595000 ;
      RECT 2.995000  1.820000 3.245000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__nand3_2
MACRO sky130_fd_sc_hs__nand3_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525000 1.350000 1.535000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.130000 1.350000 3.715000 1.630000 ;
        RECT 2.560000 1.630000 3.715000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.140000 1.340000 6.115000 1.630000 ;
        RECT 4.495000 1.630000 6.115000 1.780000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  2.004800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.010000 1.725000 1.180000 ;
        RECT 0.125000 1.180000 0.355000 1.950000 ;
        RECT 0.125000 1.950000 4.290000 2.120000 ;
        RECT 0.535000 0.595000 0.865000 1.010000 ;
        RECT 0.615000 2.120000 1.365000 2.980000 ;
        RECT 1.395000 0.595000 1.725000 1.010000 ;
        RECT 2.035000 1.820000 2.365000 1.950000 ;
        RECT 2.035000 2.120000 2.365000 2.980000 ;
        RECT 3.960000 1.820000 4.290000 1.950000 ;
        RECT 3.960000 2.120000 4.290000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.240000 0.085000 ;
      RECT 0.000000  3.245000 6.240000 3.415000 ;
      RECT 0.105000  0.255000 3.875000 0.425000 ;
      RECT 0.105000  0.425000 0.355000 0.840000 ;
      RECT 0.115000  2.290000 0.445000 3.245000 ;
      RECT 1.045000  0.425000 1.215000 0.840000 ;
      RECT 1.535000  2.290000 1.865000 3.245000 ;
      RECT 1.905000  0.425000 2.075000 1.170000 ;
      RECT 2.255000  0.595000 2.585000 0.920000 ;
      RECT 2.255000  0.920000 5.625000 1.170000 ;
      RECT 2.535000  2.290000 3.790000 3.245000 ;
      RECT 2.755000  0.425000 2.945000 0.750000 ;
      RECT 3.115000  0.595000 3.445000 0.920000 ;
      RECT 3.615000  0.425000 3.875000 0.750000 ;
      RECT 4.085000  0.085000 4.415000 0.750000 ;
      RECT 4.460000  1.950000 5.765000 3.245000 ;
      RECT 4.585000  0.390000 4.775000 0.920000 ;
      RECT 4.945000  0.085000 5.275000 0.750000 ;
      RECT 5.455000  0.390000 5.625000 0.920000 ;
      RECT 5.805000  0.085000 6.135000 1.170000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
  END
END sky130_fd_sc_hs__nand3_4
MACRO sky130_fd_sc_hs__nand3b_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.880000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.445000 1.350000 0.835000 1.780000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.350000 1.915000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015000 1.350000 1.345000 1.780000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  1.006800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.305000 1.950000 2.795000 2.120000 ;
        RECT 1.305000 2.120000 1.635000 2.980000 ;
        RECT 2.250000 0.370000 2.795000 0.790000 ;
        RECT 2.305000 1.820000 2.795000 1.950000 ;
        RECT 2.305000 2.120000 2.795000 2.980000 ;
        RECT 2.425000 0.790000 2.795000 1.150000 ;
        RECT 2.625000 1.150000 2.795000 1.820000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.880000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.880000 0.085000 ;
      RECT 0.000000  3.245000 2.880000 3.415000 ;
      RECT 0.105000  0.560000 0.375000 0.980000 ;
      RECT 0.105000  0.980000 2.255000 1.150000 ;
      RECT 0.105000  1.150000 0.275000 1.950000 ;
      RECT 0.105000  1.950000 0.600000 2.700000 ;
      RECT 0.545000  0.085000 1.220000 0.810000 ;
      RECT 0.805000  1.950000 1.135000 3.245000 ;
      RECT 1.805000  2.290000 2.135000 3.245000 ;
      RECT 2.085000  1.150000 2.255000 1.320000 ;
      RECT 2.085000  1.320000 2.455000 1.650000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
  END
END sky130_fd_sc_hs__nand3b_1
MACRO sky130_fd_sc_hs__nand3b_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.450000 0.550000 1.780000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.350000 4.195000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.430000 1.795000 1.780000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  1.332800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.260000 1.950000 3.695000 2.120000 ;
        RECT 1.260000 2.120000 1.635000 2.980000 ;
        RECT 2.335000 2.120000 2.585000 2.980000 ;
        RECT 2.470000 1.010000 2.800000 1.180000 ;
        RECT 2.525000 1.180000 2.800000 1.950000 ;
        RECT 3.365000 2.120000 3.695000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.100000  0.450000 0.350000 1.090000 ;
      RECT 0.100000  1.090000 2.195000 1.260000 ;
      RECT 0.305000  1.950000 0.890000 2.120000 ;
      RECT 0.305000  2.120000 0.635000 2.980000 ;
      RECT 0.530000  0.085000 0.820000 0.910000 ;
      RECT 0.720000  1.260000 0.890000 1.950000 ;
      RECT 0.830000  2.290000 1.075000 3.245000 ;
      RECT 1.005000  0.330000 1.255000 0.750000 ;
      RECT 1.005000  0.750000 3.790000 0.840000 ;
      RECT 1.005000  0.840000 2.105000 0.920000 ;
      RECT 1.435000  0.085000 1.765000 0.580000 ;
      RECT 1.805000  2.290000 2.135000 3.245000 ;
      RECT 1.935000  0.670000 3.790000 0.750000 ;
      RECT 1.975000  0.330000 4.220000 0.500000 ;
      RECT 2.025000  1.260000 2.195000 1.350000 ;
      RECT 2.025000  1.350000 2.355000 1.680000 ;
      RECT 2.790000  2.290000 3.120000 3.245000 ;
      RECT 2.970000  0.840000 3.790000 1.180000 ;
      RECT 3.875000  1.950000 4.205000 3.245000 ;
      RECT 3.960000  0.500000 4.220000 1.180000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__nand3b_2
MACRO sky130_fd_sc_hs__nand3b_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.363000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.350000 1.095000 1.780000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.820000 1.180000 7.075000 1.650000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.765000 1.350000 3.235000 1.780000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  1.866500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.685000 1.950000 5.850000 2.140000 ;
        RECT 3.750000 1.820000 5.850000 1.950000 ;
        RECT 4.130000 0.800000 5.345000 1.130000 ;
        RECT 4.925000 0.770000 5.345000 0.800000 ;
        RECT 4.925000 1.130000 5.155000 1.820000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.680000 0.085000 ;
      RECT 0.000000  3.245000 7.680000 3.415000 ;
      RECT 0.085000  0.580000 1.790000 0.670000 ;
      RECT 0.085000  0.670000 2.970000 0.750000 ;
      RECT 0.085000  0.750000 0.255000 1.950000 ;
      RECT 0.085000  1.950000 0.785000 2.120000 ;
      RECT 0.115000  2.290000 0.445000 3.245000 ;
      RECT 0.425000  0.920000 0.755000 1.010000 ;
      RECT 0.425000  1.010000 3.770000 1.180000 ;
      RECT 0.615000  2.120000 0.785000 2.310000 ;
      RECT 0.615000  2.310000 6.230000 2.480000 ;
      RECT 0.935000  0.085000 1.280000 0.410000 ;
      RECT 0.955000  1.950000 1.435000 2.140000 ;
      RECT 1.265000  1.180000 1.435000 1.950000 ;
      RECT 1.460000  0.390000 1.790000 0.580000 ;
      RECT 1.460000  0.750000 2.970000 0.840000 ;
      RECT 1.490000  2.650000 2.565000 3.245000 ;
      RECT 1.970000  0.085000 2.460000 0.500000 ;
      RECT 2.640000  0.390000 2.970000 0.670000 ;
      RECT 3.135000  2.650000 3.630000 3.245000 ;
      RECT 3.140000  0.085000 3.470000 0.840000 ;
      RECT 3.600000  1.180000 3.770000 1.300000 ;
      RECT 3.600000  1.300000 4.610000 1.630000 ;
      RECT 3.700000  0.350000 7.565000 0.600000 ;
      RECT 3.700000  0.600000 4.030000 0.630000 ;
      RECT 4.580000  2.650000 5.400000 3.245000 ;
      RECT 5.515000  0.600000 7.565000 0.670000 ;
      RECT 5.945000  0.840000 7.415000 1.010000 ;
      RECT 5.970000  2.650000 7.565000 3.245000 ;
      RECT 6.060000  1.820000 7.415000 1.990000 ;
      RECT 6.060000  1.990000 6.230000 2.310000 ;
      RECT 6.400000  2.160000 7.565000 2.650000 ;
      RECT 7.245000  1.010000 7.415000 1.820000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
  END
END sky130_fd_sc_hs__nand3b_4
MACRO sky130_fd_sc_hs__nand4_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.880000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 1.180000 2.775000 1.550000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.715000 1.180000 2.275000 1.550000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.180000 1.475000 1.550000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.575000 1.180000 0.905000 1.550000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  0.936500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.235000 0.840000 2.740000 1.010000 ;
        RECT 0.235000 1.010000 0.405000 1.720000 ;
        RECT 0.235000 1.720000 1.205000 1.820000 ;
        RECT 0.235000 1.820000 2.265000 1.890000 ;
        RECT 0.875000 1.890000 2.265000 2.150000 ;
        RECT 0.875000 2.150000 1.205000 2.980000 ;
        RECT 1.935000 2.150000 2.265000 2.980000 ;
        RECT 2.410000 0.350000 2.740000 0.840000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.880000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.880000 0.085000 ;
      RECT 0.000000  3.245000 2.880000 3.415000 ;
      RECT 0.110000  0.085000 0.785000 0.600000 ;
      RECT 0.375000  2.060000 0.705000 3.245000 ;
      RECT 1.400000  2.320000 1.730000 3.245000 ;
      RECT 2.435000  1.820000 2.765000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
  END
END sky130_fd_sc_hs__nand4_1
MACRO sky130_fd_sc_hs__nand4_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.885000 1.350000 4.215000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.680000 1.350000 3.715000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.430000 1.350000 2.440000 1.780000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.090000 1.780000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.633200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.635000 1.950000 4.675000 2.120000 ;
        RECT 0.635000 2.120000 0.900000 2.980000 ;
        RECT 1.570000 2.120000 1.900000 2.980000 ;
        RECT 2.830000 2.120000 3.160000 2.980000 ;
        RECT 3.840000 2.120000 4.675000 2.150000 ;
        RECT 3.840000 2.150000 4.125000 2.980000 ;
        RECT 3.845000 0.645000 4.175000 1.010000 ;
        RECT 3.845000 1.010000 4.675000 1.180000 ;
        RECT 4.445000 1.180000 4.675000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.115000  0.350000 0.445000 1.010000 ;
      RECT 0.115000  1.010000 1.315000 1.180000 ;
      RECT 0.115000  1.950000 0.450000 3.245000 ;
      RECT 0.615000  0.085000 0.945000 0.840000 ;
      RECT 1.070000  2.290000 1.400000 3.245000 ;
      RECT 1.145000  0.255000 2.325000 0.425000 ;
      RECT 1.145000  0.425000 1.315000 1.010000 ;
      RECT 1.495000  0.595000 1.825000 1.010000 ;
      RECT 1.495000  1.010000 3.315000 1.180000 ;
      RECT 1.995000  0.425000 2.325000 0.840000 ;
      RECT 2.080000  2.290000 2.650000 3.245000 ;
      RECT 2.555000  0.255000 4.675000 0.425000 ;
      RECT 2.555000  0.425000 2.815000 0.840000 ;
      RECT 2.985000  0.645000 3.315000 1.010000 ;
      RECT 3.330000  2.290000 3.660000 3.245000 ;
      RECT 3.485000  0.425000 3.675000 1.130000 ;
      RECT 4.295000  2.320000 4.625000 3.245000 ;
      RECT 4.345000  0.425000 4.675000 0.840000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_hs__nand4_2
MACRO sky130_fd_sc_hs__nand4_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.735000 1.350000 8.085000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.350000 6.160000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.350000 4.195000 1.780000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 2.275000 1.780000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  3.321600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.820000 1.950000 8.515000 2.120000 ;
        RECT 1.820000 2.120000 2.150000 2.980000 ;
        RECT 2.820000 2.120000 3.430000 2.980000 ;
        RECT 4.670000 2.120000 5.280000 2.980000 ;
        RECT 6.745000 0.880000 8.515000 1.130000 ;
        RECT 6.815000 0.800000 7.005000 0.880000 ;
        RECT 7.320000 2.120000 8.010000 2.980000 ;
        RECT 7.755000 0.800000 7.945000 0.880000 ;
        RECT 8.285000 1.130000 8.515000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
      RECT 0.000000  3.245000 8.640000 3.415000 ;
      RECT 0.115000  0.350000 0.445000 1.010000 ;
      RECT 0.115000  1.010000 2.575000 1.180000 ;
      RECT 0.115000  1.950000 1.650000 3.245000 ;
      RECT 0.615000  0.085000 0.945000 0.840000 ;
      RECT 1.115000  0.350000 1.445000 1.010000 ;
      RECT 1.615000  0.085000 1.945000 0.840000 ;
      RECT 2.245000  0.350000 4.365000 0.680000 ;
      RECT 2.245000  0.680000 2.575000 1.010000 ;
      RECT 2.320000  2.290000 2.650000 3.245000 ;
      RECT 2.745000  0.850000 3.935000 0.880000 ;
      RECT 2.745000  0.880000 6.215000 1.130000 ;
      RECT 3.600000  2.290000 4.500000 3.245000 ;
      RECT 4.595000  0.350000 8.525000 0.520000 ;
      RECT 4.595000  0.520000 4.925000 0.710000 ;
      RECT 5.095000  0.800000 5.285000 0.880000 ;
      RECT 5.450000  2.290000 7.140000 3.245000 ;
      RECT 5.455000  0.520000 5.785000 0.710000 ;
      RECT 5.955000  0.800000 6.145000 0.880000 ;
      RECT 6.315000  0.520000 6.645000 0.710000 ;
      RECT 7.175000  0.520000 7.505000 0.710000 ;
      RECT 8.190000  2.290000 8.520000 3.245000 ;
      RECT 8.195000  0.520000 8.525000 0.710000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
  END
END sky130_fd_sc_hs__nand4_4
MACRO sky130_fd_sc_hs__nand4b_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.445000 1.180000 0.815000 1.550000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.180000 2.395000 1.550000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 1.180000 1.855000 1.550000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985000 1.180000 1.315000 1.550000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.012400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.285000 1.820000 3.275000 1.890000 ;
        RECT 1.285000 1.890000 2.635000 2.150000 ;
        RECT 1.285000 2.150000 1.615000 2.980000 ;
        RECT 1.615000 1.720000 3.275000 1.820000 ;
        RECT 2.285000 2.150000 2.635000 2.980000 ;
        RECT 2.905000 0.350000 3.275000 1.050000 ;
        RECT 3.105000 1.050000 3.275000 1.720000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.105000  0.680000 0.650000 0.840000 ;
      RECT 0.105000  0.840000 2.735000 1.010000 ;
      RECT 0.105000  1.010000 0.275000 1.820000 ;
      RECT 0.105000  1.820000 0.580000 2.700000 ;
      RECT 0.785000  1.820000 1.115000 3.245000 ;
      RECT 0.855000  0.085000 1.185000 0.670000 ;
      RECT 1.785000  2.320000 2.115000 3.245000 ;
      RECT 2.565000  1.010000 2.735000 1.220000 ;
      RECT 2.565000  1.220000 2.935000 1.550000 ;
      RECT 2.805000  2.060000 3.135000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__nand4b_1
MACRO sky130_fd_sc_hs__nand4b_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 0.985000 1.510000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.350000 2.590000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.350000 4.195000 1.780000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.350000 5.635000 1.780000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.573400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.535000 0.800000 1.895000 1.010000 ;
        RECT 1.535000 1.010000 3.235000 1.180000 ;
        RECT 1.550000 1.850000 1.825000 1.950000 ;
        RECT 1.550000 1.950000 5.190000 2.120000 ;
        RECT 1.550000 2.120000 1.825000 2.980000 ;
        RECT 2.760000 1.820000 3.235000 1.950000 ;
        RECT 2.760000 2.120000 3.090000 2.980000 ;
        RECT 3.005000 1.180000 3.235000 1.820000 ;
        RECT 3.760000 2.120000 4.090000 2.980000 ;
        RECT 4.860000 2.120000 5.190000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.115000  0.350000 0.365000 0.840000 ;
      RECT 0.115000  0.840000 1.325000 1.010000 ;
      RECT 0.505000  1.680000 1.325000 1.850000 ;
      RECT 0.505000  1.850000 0.835000 2.860000 ;
      RECT 0.545000  0.085000 0.875000 0.670000 ;
      RECT 1.040000  2.020000 1.370000 3.245000 ;
      RECT 1.105000  0.350000 2.325000 0.630000 ;
      RECT 1.155000  1.010000 1.325000 1.350000 ;
      RECT 1.155000  1.350000 1.720000 1.680000 ;
      RECT 1.995000  2.290000 2.590000 3.245000 ;
      RECT 2.075000  0.630000 2.325000 0.670000 ;
      RECT 2.075000  0.670000 3.345000 0.840000 ;
      RECT 2.505000  0.255000 4.335000 0.425000 ;
      RECT 2.505000  0.425000 2.835000 0.500000 ;
      RECT 3.015000  0.595000 3.345000 0.670000 ;
      RECT 3.260000  2.290000 3.590000 3.245000 ;
      RECT 3.575000  0.595000 3.825000 0.930000 ;
      RECT 3.575000  0.930000 5.645000 1.180000 ;
      RECT 4.005000  0.425000 4.335000 0.760000 ;
      RECT 4.320000  2.290000 4.650000 3.245000 ;
      RECT 4.505000  0.400000 4.695000 0.930000 ;
      RECT 4.865000  0.085000 5.195000 0.760000 ;
      RECT 5.360000  1.950000 5.645000 3.245000 ;
      RECT 5.395000  0.400000 5.645000 0.930000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_hs__nand4b_2
MACRO sky130_fd_sc_hs__nand4b_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.363000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.835000 1.780000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.130000 1.430000 4.140000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925000 1.350000 7.555000 1.780000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.805000 1.300000 9.015000 1.780000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  2.665600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.535000 0.880000 2.725000 1.090000 ;
        RECT 1.535000 1.090000 4.675000 1.130000 ;
        RECT 2.050000 1.850000 2.680000 1.950000 ;
        RECT 2.050000 1.950000 8.505000 2.120000 ;
        RECT 2.050000 2.120000 2.670000 2.980000 ;
        RECT 2.395000 0.595000 2.725000 0.880000 ;
        RECT 2.395000 1.130000 4.675000 1.260000 ;
        RECT 4.310000 1.820000 4.675000 1.950000 ;
        RECT 4.370000 2.120000 4.590000 2.980000 ;
        RECT 4.445000 1.260000 4.675000 1.820000 ;
        RECT 6.065000 2.120000 6.660000 2.980000 ;
        RECT 8.215000 2.120000 8.505000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.120000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.120000 0.085000 ;
      RECT 0.000000  3.245000 9.120000 3.415000 ;
      RECT 0.115000  0.770000 0.445000 0.960000 ;
      RECT 0.115000  0.960000 1.335000 1.130000 ;
      RECT 0.505000  1.950000 0.835000 3.245000 ;
      RECT 0.545000  0.085000 0.875000 0.600000 ;
      RECT 1.005000  1.130000 1.335000 1.430000 ;
      RECT 1.005000  1.430000 2.850000 1.680000 ;
      RECT 1.005000  1.680000 1.335000 2.700000 ;
      RECT 1.105000  0.255000 3.075000 0.425000 ;
      RECT 1.105000  0.425000 1.435000 0.710000 ;
      RECT 1.540000  1.850000 1.870000 3.245000 ;
      RECT 1.965000  0.425000 2.215000 0.710000 ;
      RECT 2.850000  2.290000 4.190000 3.245000 ;
      RECT 2.905000  0.425000 3.075000 0.750000 ;
      RECT 2.905000  0.750000 4.875000 0.920000 ;
      RECT 3.255000  0.330000 6.725000 0.580000 ;
      RECT 4.760000  2.290000 5.885000 3.245000 ;
      RECT 5.105000  0.770000 5.435000 0.960000 ;
      RECT 5.105000  0.960000 6.215000 1.010000 ;
      RECT 5.105000  1.010000 9.005000 1.130000 ;
      RECT 5.535000  0.580000 6.725000 0.600000 ;
      RECT 5.605000  0.600000 5.795000 0.710000 ;
      RECT 5.965000  0.770000 6.215000 0.960000 ;
      RECT 5.965000  1.130000 7.170000 1.180000 ;
      RECT 6.395000  0.600000 6.725000 0.840000 ;
      RECT 6.835000  2.290000 8.035000 3.245000 ;
      RECT 6.920000  0.350000 7.100000 0.960000 ;
      RECT 6.920000  0.960000 9.005000 1.010000 ;
      RECT 7.270000  0.085000 7.600000 0.780000 ;
      RECT 7.770000  0.350000 7.960000 0.960000 ;
      RECT 8.130000  0.085000 8.505000 0.780000 ;
      RECT 8.675000  0.350000 9.005000 0.960000 ;
      RECT 8.675000  1.950000 8.955000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
  END
END sky130_fd_sc_hs__nand4b_4
MACRO sky130_fd_sc_hs__nand4bb_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.255000 0.480000 0.670000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.470000 1.315000 1.800000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.985000 0.810000 3.315000 1.550000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.350000 3.885000 1.780000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.248650 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.675000 2.310000 3.095000 2.480000 ;
        RECT 1.675000 2.480000 2.005000 2.980000 ;
        RECT 1.720000 0.350000 3.655000 0.620000 ;
        RECT 2.525000 1.820000 3.095000 1.950000 ;
        RECT 2.525000 1.950000 4.225000 2.120000 ;
        RECT 2.525000 2.120000 3.095000 2.310000 ;
        RECT 2.765000 2.480000 3.095000 2.980000 ;
        RECT 3.485000 0.620000 3.655000 1.010000 ;
        RECT 3.485000 1.010000 4.225000 1.180000 ;
        RECT 3.765000 2.120000 4.225000 2.980000 ;
        RECT 4.055000 1.180000 4.225000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  0.840000 0.470000 1.130000 ;
      RECT 0.115000  1.130000 2.015000 1.300000 ;
      RECT 0.115000  1.300000 0.285000 1.970000 ;
      RECT 0.115000  1.970000 0.445000 2.850000 ;
      RECT 0.615000  1.970000 0.945000 3.245000 ;
      RECT 0.650000  0.085000 0.980000 0.960000 ;
      RECT 1.115000  1.970000 2.355000 2.140000 ;
      RECT 1.115000  2.140000 1.445000 2.850000 ;
      RECT 1.150000  0.630000 1.490000 0.790000 ;
      RECT 1.150000  0.790000 2.355000 0.960000 ;
      RECT 1.685000  1.300000 2.015000 1.550000 ;
      RECT 2.175000  2.650000 2.595000 3.245000 ;
      RECT 2.185000  0.960000 2.355000 1.220000 ;
      RECT 2.185000  1.220000 2.745000 1.550000 ;
      RECT 2.185000  1.550000 2.355000 1.970000 ;
      RECT 3.265000  2.290000 3.595000 3.245000 ;
      RECT 3.825000  0.085000 4.155000 0.840000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__nand4bb_1
MACRO sky130_fd_sc_hs__nand4bb_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.435000 1.300000 0.835000 1.780000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.180000 1.335000 1.510000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.350000 5.385000 1.780000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.625000 1.350000 6.595000 1.680000 ;
        RECT 6.365000 1.680000 6.595000 1.780000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.614500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.345000 0.670000 2.855000 0.840000 ;
        RECT 2.345000 1.820000 2.675000 1.850000 ;
        RECT 2.345000 1.850000 4.195000 1.950000 ;
        RECT 2.345000 1.950000 6.105000 2.020000 ;
        RECT 2.345000 2.020000 2.675000 2.980000 ;
        RECT 2.685000 0.840000 2.855000 1.090000 ;
        RECT 2.685000 1.090000 4.195000 1.260000 ;
        RECT 3.345000 2.020000 6.105000 2.120000 ;
        RECT 3.345000 2.120000 3.675000 2.980000 ;
        RECT 3.965000 1.260000 4.195000 1.850000 ;
        RECT 4.775000 2.120000 5.105000 2.980000 ;
        RECT 5.775000 1.850000 6.105000 1.950000 ;
        RECT 5.775000 2.120000 6.105000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.720000 0.085000 ;
      RECT 0.000000  3.245000 6.720000 3.415000 ;
      RECT 0.095000  0.350000 0.460000 1.030000 ;
      RECT 0.095000  1.030000 0.265000 1.950000 ;
      RECT 0.095000  1.950000 0.445000 2.240000 ;
      RECT 0.095000  2.240000 2.175000 2.410000 ;
      RECT 0.095000  2.410000 0.445000 2.860000 ;
      RECT 0.630000  0.085000 0.960000 1.010000 ;
      RECT 0.650000  2.580000 0.980000 3.245000 ;
      RECT 1.130000  0.350000 1.675000 1.010000 ;
      RECT 1.185000  1.820000 1.675000 2.070000 ;
      RECT 1.505000  1.010000 2.515000 1.180000 ;
      RECT 1.505000  1.180000 1.675000 1.820000 ;
      RECT 1.845000  0.330000 3.195000 0.500000 ;
      RECT 1.845000  0.500000 2.175000 0.840000 ;
      RECT 1.845000  1.350000 2.175000 2.240000 ;
      RECT 1.845000  2.580000 2.175000 3.245000 ;
      RECT 2.345000  1.180000 2.515000 1.430000 ;
      RECT 2.345000  1.430000 3.795000 1.600000 ;
      RECT 2.845000  2.190000 3.175000 3.245000 ;
      RECT 3.025000  0.500000 3.195000 0.750000 ;
      RECT 3.025000  0.750000 4.180000 0.920000 ;
      RECT 3.125000  1.600000 3.795000 1.680000 ;
      RECT 3.365000  0.255000 5.240000 0.425000 ;
      RECT 3.365000  0.425000 3.695000 0.580000 ;
      RECT 3.845000  2.290000 4.605000 3.245000 ;
      RECT 4.410000  0.620000 4.740000 1.010000 ;
      RECT 4.410000  1.010000 6.600000 1.180000 ;
      RECT 4.910000  0.425000 5.240000 0.815000 ;
      RECT 5.275000  2.290000 5.605000 3.245000 ;
      RECT 5.420000  0.350000 5.670000 1.010000 ;
      RECT 5.840000  0.085000 6.170000 0.815000 ;
      RECT 6.275000  1.950000 6.605000 3.245000 ;
      RECT 6.350000  0.350000 6.600000 1.010000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
  END
END sky130_fd_sc_hs__nand4bb_2
MACRO sky130_fd_sc_hs__nand4bb_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.363000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.440000 1.450000 0.835000 1.780000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.363000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 1.550000 1.795000 1.880000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.185000 1.320000 7.610000 1.650000 ;
        RECT 6.845000 1.650000 7.075000 1.780000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.265000 1.300000 9.955000 1.780000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  3.236100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.320000 0.595000 2.650000 0.870000 ;
        RECT 2.320000 0.870000 3.505000 1.040000 ;
        RECT 2.525000 2.060000 4.815000 2.230000 ;
        RECT 2.525000 2.230000 2.965000 2.990000 ;
        RECT 3.335000 0.595000 3.505000 0.870000 ;
        RECT 3.335000 1.040000 3.505000 1.090000 ;
        RECT 3.335000 1.090000 5.685000 1.260000 ;
        RECT 3.635000 2.230000 3.865000 2.990000 ;
        RECT 4.485000 1.850000 6.665000 1.950000 ;
        RECT 4.485000 1.950000 9.515000 1.990000 ;
        RECT 4.485000 1.990000 5.685000 2.020000 ;
        RECT 4.485000 2.020000 4.815000 2.060000 ;
        RECT 4.535000 2.230000 4.815000 2.980000 ;
        RECT 5.515000 1.260000 5.685000 1.820000 ;
        RECT 5.515000 1.820000 6.665000 1.850000 ;
        RECT 5.515000 2.020000 5.685000 2.980000 ;
        RECT 6.335000 1.990000 9.515000 2.120000 ;
        RECT 6.335000 2.120000 6.665000 2.980000 ;
        RECT 7.335000 1.820000 7.665000 1.950000 ;
        RECT 7.335000 2.120000 7.665000 2.980000 ;
        RECT 8.285000 2.120000 8.615000 2.980000 ;
        RECT 9.185000 2.120000 9.515000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.100000  0.550000  0.445000 0.660000 ;
      RECT 0.100000  0.660000  1.760000 0.830000 ;
      RECT 0.100000  0.830000  0.445000 1.280000 ;
      RECT 0.100000  1.280000  0.270000 1.950000 ;
      RECT 0.100000  1.950000  0.815000 2.120000 ;
      RECT 0.115000  2.290000  0.445000 3.245000 ;
      RECT 0.625000  0.085000  0.955000 0.490000 ;
      RECT 0.645000  2.120000  0.815000 2.980000 ;
      RECT 1.015000  2.390000  1.345000 3.245000 ;
      RECT 1.125000  1.000000  1.420000 1.330000 ;
      RECT 1.125000  1.330000  1.295000 2.050000 ;
      RECT 1.125000  2.050000  2.135000 2.220000 ;
      RECT 1.515000  2.220000  1.795000 2.980000 ;
      RECT 1.590000  0.830000  1.760000 1.210000 ;
      RECT 1.590000  1.210000  3.165000 1.380000 ;
      RECT 1.930000  0.255000  3.935000 0.425000 ;
      RECT 1.930000  0.425000  2.100000 1.040000 ;
      RECT 1.965000  1.720000  4.315000 1.890000 ;
      RECT 1.965000  1.890000  2.135000 2.050000 ;
      RECT 2.005000  2.390000  2.335000 3.245000 ;
      RECT 2.155000  1.380000  3.165000 1.550000 ;
      RECT 2.820000  0.425000  3.150000 0.700000 ;
      RECT 3.135000  2.400000  3.465000 3.245000 ;
      RECT 3.685000  0.425000  3.935000 0.750000 ;
      RECT 3.685000  0.750000  5.895000 0.920000 ;
      RECT 4.035000  2.400000  4.365000 3.245000 ;
      RECT 4.115000  0.255000  7.745000 0.425000 ;
      RECT 4.115000  0.425000  5.385000 0.580000 ;
      RECT 4.145000  1.430000  5.345000 1.680000 ;
      RECT 4.145000  1.680000  4.315000 1.720000 ;
      RECT 4.985000  2.190000  5.315000 3.245000 ;
      RECT 5.565000  0.595000  5.895000 0.750000 ;
      RECT 5.885000  2.160000  6.135000 3.245000 ;
      RECT 6.125000  0.595000  6.375000 0.980000 ;
      RECT 6.125000  0.980000  9.965000 1.130000 ;
      RECT 6.125000  1.130000  8.095000 1.150000 ;
      RECT 6.555000  0.425000  6.885000 0.810000 ;
      RECT 6.835000  2.290000  7.165000 3.245000 ;
      RECT 7.065000  0.595000  7.235000 0.980000 ;
      RECT 7.415000  0.425000  7.745000 0.810000 ;
      RECT 7.865000  2.290000  8.115000 3.245000 ;
      RECT 7.925000  0.350000  8.095000 0.960000 ;
      RECT 7.925000  0.960000  9.965000 0.980000 ;
      RECT 8.275000  0.085000  8.605000 0.790000 ;
      RECT 8.785000  0.350000  8.955000 0.960000 ;
      RECT 8.815000  2.290000  8.985000 3.245000 ;
      RECT 9.135000  0.085000  9.465000 0.790000 ;
      RECT 9.635000  0.350000  9.965000 0.960000 ;
      RECT 9.715000  1.950000  9.965000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
  END
END sky130_fd_sc_hs__nand4bb_4
MACRO sky130_fd_sc_hs__nor2_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.440000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.455000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985000 1.300000 1.315000 1.780000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.537600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565000 0.350000 0.815000 1.130000 ;
        RECT 0.645000 1.130000 0.815000 1.950000 ;
        RECT 0.645000 1.950000 1.315000 2.890000 ;
        RECT 0.985000 2.890000 1.315000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 1.440000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 1.440000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.440000 0.085000 ;
      RECT 0.000000  3.245000 1.440000 3.415000 ;
      RECT 0.115000  1.950000 0.445000 3.245000 ;
      RECT 0.135000  0.085000 0.385000 1.130000 ;
      RECT 0.995000  0.085000 1.325000 1.130000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
  END
END sky130_fd_sc_hs__nor2_1
MACRO sky130_fd_sc_hs__nor2_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.400000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.805000 0.255000 2.135000 0.440000 ;
        RECT 1.805000 0.440000 2.275000 1.410000 ;
        RECT 1.805000 1.410000 2.135000 1.605000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 1.180000 0.445000 1.550000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.820000 0.945000 2.735000 ;
        RECT 0.615000 0.350000 0.945000 1.820000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.400000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.400000 0.085000 ;
      RECT 0.000000  3.245000 2.400000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 1.010000 ;
      RECT 0.155000  1.820000 0.405000 2.905000 ;
      RECT 0.155000  2.905000 1.305000 3.075000 ;
      RECT 1.115000  0.085000 1.445000 1.130000 ;
      RECT 1.135000  1.775000 2.285000 1.945000 ;
      RECT 1.135000  1.945000 1.305000 2.905000 ;
      RECT 1.505000  2.115000 1.755000 3.245000 ;
      RECT 1.955000  1.945000 2.285000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
  END
END sky130_fd_sc_hs__nor2_2
MACRO sky130_fd_sc_hs__nor2_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 1.795000 1.550000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.180000 4.195000 1.550000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.793600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.640000 0.340000 1.690000 0.840000 ;
        RECT 0.640000 0.840000 2.690000 1.010000 ;
        RECT 2.360000 0.350000 2.690000 0.840000 ;
        RECT 2.360000 1.010000 2.690000 1.130000 ;
        RECT 2.365000 1.130000 2.690000 1.180000 ;
        RECT 2.365000 1.180000 2.755000 1.410000 ;
        RECT 2.365000 1.410000 2.695000 1.720000 ;
        RECT 2.365000 1.720000 3.695000 1.890000 ;
        RECT 2.365000 1.890000 2.695000 2.735000 ;
        RECT 3.365000 1.890000 3.695000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  0.085000 0.470000 1.010000 ;
      RECT 0.115000  1.720000 2.195000 1.890000 ;
      RECT 0.115000  1.890000 0.445000 2.980000 ;
      RECT 0.645000  2.060000 0.815000 3.245000 ;
      RECT 1.015000  1.890000 1.345000 2.980000 ;
      RECT 1.545000  2.060000 1.715000 3.245000 ;
      RECT 1.860000  0.085000 2.190000 0.670000 ;
      RECT 1.915000  1.890000 2.195000 2.905000 ;
      RECT 1.915000  2.905000 4.145000 3.075000 ;
      RECT 2.860000  0.085000 4.205000 1.010000 ;
      RECT 2.865000  2.060000 3.195000 2.905000 ;
      RECT 3.865000  1.820000 4.145000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__nor2_4
MACRO sky130_fd_sc_hs__nor2_8
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.788000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.350000 3.715000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.788000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.225000 0.300000 7.555000 1.310000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  2.839300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.860000 0.350000 2.190000 1.010000 ;
        RECT 1.860000 1.010000 5.275000 1.140000 ;
        RECT 1.860000 1.140000 6.275000 1.180000 ;
        RECT 3.260000 0.350000 3.590000 1.010000 ;
        RECT 4.260000 0.350000 5.275000 1.010000 ;
        RECT 4.260000 1.180000 6.275000 1.310000 ;
        RECT 4.415000 1.310000 6.275000 1.480000 ;
        RECT 4.415000 1.480000 7.545000 1.650000 ;
        RECT 4.415000 1.650000 5.695000 1.780000 ;
        RECT 4.415000 1.780000 4.745000 2.735000 ;
        RECT 5.365000 1.780000 5.695000 2.735000 ;
        RECT 5.945000 0.350000 6.275000 1.140000 ;
        RECT 6.265000 1.650000 6.595000 2.735000 ;
        RECT 7.215000 1.650000 7.545000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.115000  1.780000 1.315000 1.950000 ;
      RECT 0.115000  1.950000 0.445000 2.980000 ;
      RECT 0.615000  2.120000 0.945000 3.245000 ;
      RECT 0.650000  0.085000 1.690000 1.130000 ;
      RECT 1.145000  1.950000 4.245000 2.120000 ;
      RECT 1.145000  2.120000 1.315000 2.980000 ;
      RECT 1.515000  2.290000 1.845000 3.245000 ;
      RECT 2.045000  2.120000 2.295000 2.980000 ;
      RECT 2.360000  0.085000 3.090000 0.840000 ;
      RECT 2.465000  2.290000 2.795000 3.245000 ;
      RECT 2.995000  2.120000 3.245000 2.980000 ;
      RECT 3.415000  2.290000 3.745000 3.245000 ;
      RECT 3.760000  0.085000 4.090000 0.840000 ;
      RECT 3.915000  2.120000 4.245000 2.905000 ;
      RECT 3.915000  2.905000 8.045000 3.075000 ;
      RECT 4.925000  1.950000 5.185000 2.905000 ;
      RECT 5.445000  0.085000 5.775000 0.970000 ;
      RECT 5.875000  1.820000 6.080000 2.905000 ;
      RECT 6.445000  0.085000 6.775000 1.130000 ;
      RECT 6.775000  1.820000 7.035000 2.905000 ;
      RECT 7.715000  1.820000 8.045000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_hs__nor2_8
MACRO sky130_fd_sc_hs__nor2b_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.400000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.035000 1.180000 1.365000 1.550000 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.180000 0.440000 1.550000 ;
    END
  END B_N
  PIN Y
    ANTENNADIFFAREA  0.682700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.535000 0.350000 1.785000 0.980000 ;
        RECT 1.535000 0.980000 2.315000 1.150000 ;
        RECT 1.875000 1.820000 2.315000 2.980000 ;
        RECT 2.145000 1.150000 2.315000 1.820000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.400000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.400000 0.085000 ;
      RECT 0.000000  3.245000 2.400000 3.415000 ;
      RECT 0.255000  0.680000 0.780000 1.010000 ;
      RECT 0.315000  1.720000 1.705000 1.890000 ;
      RECT 0.315000  1.890000 0.645000 2.700000 ;
      RECT 0.610000  1.010000 0.780000 1.720000 ;
      RECT 0.925000  2.060000 1.255000 3.245000 ;
      RECT 0.950000  0.085000 1.280000 1.010000 ;
      RECT 1.535000  1.320000 1.975000 1.650000 ;
      RECT 1.535000  1.650000 1.705000 1.720000 ;
      RECT 1.955000  0.085000 2.230000 0.810000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
  END
END sky130_fd_sc_hs__nor2b_1
MACRO sky130_fd_sc_hs__nor2b_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.350000 2.755000 1.780000 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.530000 1.470000 0.860000 1.800000 ;
    END
  END B_N
  PIN Y
    ANTENNADIFFAREA  0.824400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 0.350000 1.815000 0.960000 ;
        RECT 1.645000 0.960000 2.745000 1.010000 ;
        RECT 1.645000 1.010000 3.235000 1.180000 ;
        RECT 1.645000 1.180000 1.820000 2.735000 ;
        RECT 2.495000 0.350000 2.745000 0.960000 ;
        RECT 3.005000 1.180000 3.235000 1.410000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.110000  0.450000 0.780000 1.130000 ;
      RECT 0.110000  1.130000 1.475000 1.300000 ;
      RECT 0.110000  1.300000 0.360000 2.980000 ;
      RECT 0.560000  1.970000 0.890000 3.245000 ;
      RECT 0.985000  0.085000 1.315000 0.960000 ;
      RECT 1.120000  1.820000 1.450000 2.905000 ;
      RECT 1.120000  2.905000 2.350000 3.075000 ;
      RECT 1.145000  1.300000 1.475000 1.550000 ;
      RECT 1.985000  0.085000 2.315000 0.790000 ;
      RECT 2.020000  1.950000 3.250000 2.120000 ;
      RECT 2.020000  2.120000 2.350000 2.905000 ;
      RECT 2.550000  2.290000 2.800000 3.245000 ;
      RECT 2.915000  0.085000 3.245000 0.840000 ;
      RECT 3.000000  1.820000 3.250000 1.950000 ;
      RECT 3.000000  2.120000 3.250000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__nor2b_2
MACRO sky130_fd_sc_hs__nor2b_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.790000 1.010000 3.975000 1.180000 ;
        RECT 0.790000 1.180000 1.795000 1.340000 ;
        RECT 1.085000 1.340000 1.795000 1.410000 ;
        RECT 3.645000 1.180000 3.975000 1.550000 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.363000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.750000 1.180000 5.155000 1.825000 ;
    END
  END B_N
  PIN Y
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.670000 3.810000 0.840000 ;
        RECT 0.125000 0.840000 0.355000 1.410000 ;
        RECT 0.185000 1.410000 0.355000 1.510000 ;
        RECT 0.185000 1.510000 0.705000 1.580000 ;
        RECT 0.185000 1.580000 2.055000 1.680000 ;
        RECT 0.535000 1.680000 2.055000 1.750000 ;
        RECT 1.885000 1.750000 2.055000 1.850000 ;
        RECT 1.885000 1.850000 2.165000 2.060000 ;
        RECT 1.885000 2.060000 3.145000 2.230000 ;
        RECT 1.885000 2.230000 2.165000 2.735000 ;
        RECT 2.060000 0.530000 2.390000 0.670000 ;
        RECT 2.895000 2.230000 3.145000 2.735000 ;
        RECT 3.560000 0.510000 3.810000 0.670000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.280000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.245000 5.280000 3.415000 ;
      RECT 0.115000  1.850000 0.365000 3.245000 ;
      RECT 0.565000  1.920000 1.715000 2.090000 ;
      RECT 0.565000  2.090000 0.895000 2.980000 ;
      RECT 1.095000  2.260000 1.265000 3.245000 ;
      RECT 1.465000  2.090000 1.715000 2.905000 ;
      RECT 1.465000  2.905000 3.645000 3.075000 ;
      RECT 1.550000  0.085000 1.880000 0.500000 ;
      RECT 2.225000  1.350000 3.225000 1.680000 ;
      RECT 2.365000  2.400000 2.695000 2.905000 ;
      RECT 2.570000  0.085000 3.380000 0.500000 ;
      RECT 3.055000  1.680000 3.225000 1.720000 ;
      RECT 3.055000  1.720000 4.580000 1.890000 ;
      RECT 3.315000  2.060000 3.645000 2.905000 ;
      RECT 3.815000  2.060000 4.145000 3.245000 ;
      RECT 3.990000  0.085000 4.240000 0.840000 ;
      RECT 4.350000  1.890000 4.580000 1.995000 ;
      RECT 4.350000  1.995000 4.680000 2.875000 ;
      RECT 4.410000  0.345000 5.165000 1.010000 ;
      RECT 4.410000  1.010000 4.580000 1.720000 ;
      RECT 4.880000  1.995000 5.130000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
  END
END sky130_fd_sc_hs__nor2b_4
MACRO sky130_fd_sc_hs__nor3_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.920000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.360000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.870000 1.300000 1.315000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 1.300000 1.815000 1.780000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.737300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.530000 0.880000 1.805000 1.130000 ;
        RECT 0.530000 1.130000 0.700000 1.950000 ;
        RECT 0.530000 1.950000 1.815000 2.120000 ;
        RECT 0.605000 2.120000 1.815000 2.980000 ;
        RECT 0.615000 0.365000 0.805000 0.880000 ;
        RECT 1.475000 0.350000 1.805000 0.880000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 1.920000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 1.920000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.920000 0.085000 ;
      RECT 0.000000  3.245000 1.920000 3.415000 ;
      RECT 0.105000  1.950000 0.355000 2.325000 ;
      RECT 0.105000  2.325000 0.435000 3.245000 ;
      RECT 0.115000  0.085000 0.445000 0.710000 ;
      RECT 0.115000  0.710000 0.360000 1.010000 ;
      RECT 0.975000  0.085000 1.305000 0.710000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
  END
END sky130_fd_sc_hs__nor3_1
MACRO sky130_fd_sc_hs__nor3_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.650000 0.310000 3.235000 0.980000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.305000 1.220000 1.635000 1.380000 ;
        RECT 1.305000 1.380000 3.255000 1.550000 ;
        RECT 2.925000 1.180000 3.255000 1.380000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.180000 0.975000 1.550000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.861900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.350000 0.445000 0.840000 ;
        RECT 0.115000 0.840000 1.980000 1.010000 ;
        RECT 0.115000 1.010000 0.355000 1.720000 ;
        RECT 0.115000 1.720000 0.945000 1.890000 ;
        RECT 0.615000 1.890000 0.945000 2.735000 ;
        RECT 1.650000 0.350000 1.980000 0.840000 ;
        RECT 1.650000 1.010000 1.980000 1.050000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.115000  2.060000 0.445000 2.905000 ;
      RECT 0.115000  2.905000 1.315000 3.075000 ;
      RECT 0.615000  0.085000 1.480000 0.650000 ;
      RECT 1.145000  1.720000 3.245000 1.890000 ;
      RECT 1.145000  1.890000 1.315000 2.905000 ;
      RECT 1.515000  2.060000 2.795000 2.230000 ;
      RECT 1.515000  2.230000 1.845000 2.990000 ;
      RECT 2.015000  2.400000 2.345000 3.245000 ;
      RECT 2.150000  0.085000 2.480000 1.130000 ;
      RECT 2.515000  2.230000 2.795000 2.990000 ;
      RECT 2.965000  1.890000 3.245000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__nor3_2
MACRO sky130_fd_sc_hs__nor3_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.350000 0.935000 1.920000 ;
        RECT 0.605000 1.920000 1.795000 2.170000 ;
        RECT 1.625000 2.170000 6.135000 2.190000 ;
        RECT 1.625000 2.190000 4.020000 2.340000 ;
        RECT 3.850000 2.020000 6.135000 2.170000 ;
        RECT 5.805000 0.330000 6.135000 2.020000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.310000 1.350000 4.965000 1.510000 ;
        RECT 1.310000 1.510000 2.755000 1.520000 ;
        RECT 1.310000 1.520000 1.640000 1.680000 ;
        RECT 2.045000 1.180000 4.965000 1.350000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.785000 0.340000 5.635000 0.670000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  1.674800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.350000 0.875000 1.010000 ;
        RECT 0.545000 1.010000 1.875000 1.180000 ;
        RECT 1.545000 0.350000 1.875000 0.840000 ;
        RECT 1.545000 0.840000 5.305000 1.010000 ;
        RECT 2.140000 1.750000 5.305000 1.850000 ;
        RECT 2.140000 1.850000 3.680000 2.000000 ;
        RECT 2.545000 0.350000 2.875000 0.840000 ;
        RECT 3.350000 1.680000 5.305000 1.750000 ;
        RECT 5.135000 1.010000 5.305000 1.680000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.720000 0.085000 ;
      RECT 0.000000  3.245000 6.720000 3.415000 ;
      RECT 0.110000  1.820000 0.360000 2.340000 ;
      RECT 0.110000  2.340000 1.340000 2.510000 ;
      RECT 0.110000  2.510000 0.360000 2.980000 ;
      RECT 0.115000  0.085000 0.365000 1.130000 ;
      RECT 0.560000  2.680000 0.890000 3.245000 ;
      RECT 1.045000  0.085000 1.375000 0.840000 ;
      RECT 1.090000  2.510000 6.615000 2.530000 ;
      RECT 1.090000  2.530000 4.735000 2.680000 ;
      RECT 1.090000  2.680000 1.340000 2.980000 ;
      RECT 1.540000  2.850000 4.285000 2.905000 ;
      RECT 1.540000  2.905000 5.265000 3.075000 ;
      RECT 2.045000  0.085000 2.375000 0.670000 ;
      RECT 3.055000  0.085000 3.365000 0.670000 ;
      RECT 4.485000  2.360000 6.615000 2.510000 ;
      RECT 4.485000  2.680000 4.735000 2.735000 ;
      RECT 4.935000  2.700000 5.265000 2.905000 ;
      RECT 5.465000  2.530000 5.635000 3.000000 ;
      RECT 5.835000  2.700000 6.165000 3.245000 ;
      RECT 6.365000  1.820000 6.615000 2.360000 ;
      RECT 6.365000  2.530000 6.615000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
  END
END sky130_fd_sc_hs__nor3_4
MACRO sky130_fd_sc_hs__nor3b_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.880000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985000 1.350000 1.315000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.555000 1.350000 1.885000 1.780000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.445000 1.180000 0.815000 1.550000 ;
    END
  END C_N
  PIN Y
    ANTENNADIFFAREA  0.778100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.330000 0.350000 1.660000 1.010000 ;
        RECT 1.330000 1.010000 2.795000 1.180000 ;
        RECT 2.275000 2.290000 2.795000 2.980000 ;
        RECT 2.330000 0.350000 2.795000 1.010000 ;
        RECT 2.625000 1.180000 2.795000 2.290000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.880000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.880000 0.085000 ;
      RECT 0.000000  3.245000 2.880000 3.415000 ;
      RECT 0.105000  0.680000 0.650000 1.010000 ;
      RECT 0.105000  1.010000 0.275000 1.820000 ;
      RECT 0.105000  1.820000 0.595000 1.950000 ;
      RECT 0.105000  1.950000 2.295000 2.120000 ;
      RECT 0.105000  2.120000 0.595000 2.700000 ;
      RECT 0.830000  0.085000 1.160000 1.010000 ;
      RECT 0.835000  2.290000 1.165000 3.245000 ;
      RECT 1.830000  0.085000 2.160000 0.840000 ;
      RECT 2.125000  1.350000 2.455000 1.680000 ;
      RECT 2.125000  1.680000 2.295000 1.950000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
  END
END sky130_fd_sc_hs__nor3b_1
MACRO sky130_fd_sc_hs__nor3b_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.350000 4.675000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.605000 1.350000 3.275000 1.780000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.450000 0.835000 1.780000 ;
    END
  END C_N
  PIN Y
    ANTENNADIFFAREA  1.005700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.120000 0.350000 1.395000 0.770000 ;
        RECT 1.120000 0.770000 2.695000 0.940000 ;
        RECT 1.565000 0.940000 2.695000 0.960000 ;
        RECT 1.565000 0.960000 4.185000 1.130000 ;
        RECT 1.640000 1.130000 1.810000 2.735000 ;
        RECT 2.505000 0.350000 2.695000 0.770000 ;
        RECT 3.925000 0.350000 4.185000 0.960000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.085000  0.350000 0.450000 1.110000 ;
      RECT 0.085000  1.110000 1.335000 1.280000 ;
      RECT 0.085000  1.280000 0.255000 1.950000 ;
      RECT 0.085000  1.950000 0.360000 2.980000 ;
      RECT 0.560000  1.950000 0.890000 3.245000 ;
      RECT 0.620000  0.085000 0.950000 0.940000 ;
      RECT 1.005000  1.280000 1.335000 1.550000 ;
      RECT 1.110000  1.820000 1.440000 2.905000 ;
      RECT 1.110000  2.905000 3.240000 3.075000 ;
      RECT 1.565000  0.085000 2.335000 0.600000 ;
      RECT 2.010000  1.820000 2.290000 2.905000 ;
      RECT 2.460000  1.950000 4.240000 2.120000 ;
      RECT 2.460000  2.120000 2.790000 2.735000 ;
      RECT 2.865000  0.085000 3.755000 0.770000 ;
      RECT 2.970000  2.290000 3.240000 2.905000 ;
      RECT 3.460000  2.290000 3.790000 3.245000 ;
      RECT 3.990000  2.120000 4.240000 2.980000 ;
      RECT 4.355000  0.085000 4.685000 1.130000 ;
      RECT 4.425000  1.950000 4.690000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_hs__nor3b_2
MACRO sky130_fd_sc_hs__nor3b_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.440000 1.220000 6.595000 1.550000 ;
        RECT 6.365000 1.180000 6.595000 1.220000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.815000 1.780000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.363000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.765000 1.180000 7.095000 1.550000 ;
    END
  END C_N
  PIN Y
    ANTENNADIFFAREA  1.985500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.615000 0.350000 0.945000 1.010000 ;
        RECT 0.615000 1.010000 5.935000 1.050000 ;
        RECT 0.615000 1.050000 3.805000 1.150000 ;
        RECT 0.615000 1.150000 2.275000 1.180000 ;
        RECT 1.615000 0.350000 1.945000 0.980000 ;
        RECT 1.615000 0.980000 5.935000 1.010000 ;
        RECT 2.045000 1.180000 2.275000 1.820000 ;
        RECT 2.045000 1.820000 3.720000 2.070000 ;
        RECT 2.625000 0.350000 2.795000 0.980000 ;
        RECT 3.475000 0.350000 3.805000 0.880000 ;
        RECT 3.475000 0.880000 5.935000 0.980000 ;
        RECT 4.475000 0.350000 4.805000 0.880000 ;
        RECT 5.605000 0.350000 5.935000 0.880000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.680000 0.085000 ;
      RECT 0.000000  3.245000 7.680000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 1.130000 ;
      RECT 0.115000  1.950000 0.445000 2.905000 ;
      RECT 0.115000  2.905000 2.370000 3.075000 ;
      RECT 0.615000  1.950000 1.870000 2.120000 ;
      RECT 0.615000  2.120000 0.945000 2.735000 ;
      RECT 1.115000  0.085000 1.445000 0.840000 ;
      RECT 1.145000  2.290000 1.315000 2.905000 ;
      RECT 1.525000  2.120000 1.870000 2.240000 ;
      RECT 1.525000  2.240000 5.100000 2.410000 ;
      RECT 1.525000  2.410000 1.855000 2.735000 ;
      RECT 2.040000  2.580000 4.170000 2.750000 ;
      RECT 2.040000  2.750000 2.370000 2.905000 ;
      RECT 2.115000  0.085000 2.445000 0.810000 ;
      RECT 2.580000  1.320000 4.195000 1.650000 ;
      RECT 2.940000  2.750000 3.270000 2.910000 ;
      RECT 2.975000  0.085000 3.305000 0.810000 ;
      RECT 3.840000  2.750000 4.170000 2.910000 ;
      RECT 3.890000  1.650000 4.195000 1.720000 ;
      RECT 3.890000  1.720000 7.565000 1.890000 ;
      RECT 3.975000  0.085000 4.305000 0.710000 ;
      RECT 4.400000  2.580000 4.730000 3.245000 ;
      RECT 4.795000  2.060000 6.080000 2.230000 ;
      RECT 4.795000  2.230000 5.100000 2.240000 ;
      RECT 4.930000  2.410000 5.100000 2.990000 ;
      RECT 4.975000  0.085000 5.435000 0.680000 ;
      RECT 5.300000  2.400000 5.630000 3.245000 ;
      RECT 5.810000  2.230000 6.080000 2.990000 ;
      RECT 6.105000  0.085000 6.435000 1.010000 ;
      RECT 6.250000  2.060000 6.580000 3.245000 ;
      RECT 6.605000  0.350000 7.565000 1.010000 ;
      RECT 6.785000  1.890000 7.055000 2.700000 ;
      RECT 7.235000  2.060000 7.565000 3.245000 ;
      RECT 7.395000  1.010000 7.565000 1.720000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
  END
END sky130_fd_sc_hs__nor3b_4
MACRO sky130_fd_sc_hs__nor4_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.880000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 0.540000 1.550000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.975000 1.350000 1.315000 2.890000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.545000 1.350000 1.875000 2.150000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.350000 2.445000 1.780000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  0.744800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.780000 0.350000 1.040000 1.010000 ;
        RECT 0.780000 1.010000 2.785000 1.180000 ;
        RECT 1.810000 0.350000 2.140000 1.010000 ;
        RECT 2.265000 1.950000 2.785000 2.980000 ;
        RECT 2.615000 1.180000 2.785000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.880000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.880000 0.085000 ;
      RECT 0.000000  3.245000 2.880000 3.415000 ;
      RECT 0.210000  0.085000 0.610000 1.010000 ;
      RECT 0.255000  1.820000 0.585000 3.245000 ;
      RECT 1.210000  0.085000 1.540000 0.840000 ;
      RECT 2.310000  0.085000 2.640000 0.840000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
  END
END sky130_fd_sc_hs__nor4_1
MACRO sky130_fd_sc_hs__nor4_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.095000 1.180000 3.715000 1.540000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.285000 1.320000 2.625000 1.650000 ;
        RECT 2.455000 1.650000 2.625000 1.710000 ;
        RECT 2.455000 1.710000 4.215000 1.880000 ;
        RECT 3.885000 0.280000 4.215000 1.710000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.170000 0.700000 1.320000 ;
        RECT 0.425000 1.320000 2.075000 1.500000 ;
        RECT 1.565000 1.500000 2.075000 1.650000 ;
        RECT 1.565000 1.650000 1.795000 2.150000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.330000 0.435000 0.660000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  0.808000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.830000 1.880000 0.980000 ;
        RECT 0.085000 0.980000 2.880000 1.000000 ;
        RECT 0.085000 1.000000 0.255000 1.670000 ;
        RECT 0.085000 1.670000 1.385000 1.840000 ;
        RECT 0.615000 1.840000 1.385000 2.150000 ;
        RECT 1.550000 0.350000 1.880000 0.830000 ;
        RECT 1.550000 1.000000 2.880000 1.150000 ;
        RECT 2.550000 0.350000 2.880000 0.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  2.010000 0.445000 2.320000 ;
      RECT 0.115000  2.320000 2.285000 2.490000 ;
      RECT 0.115000  2.490000 0.365000 3.000000 ;
      RECT 0.565000  2.660000 1.835000 2.980000 ;
      RECT 0.605000  0.085000 1.380000 0.600000 ;
      RECT 2.035000  1.820000 2.285000 2.050000 ;
      RECT 2.035000  2.050000 4.205000 2.220000 ;
      RECT 2.035000  2.220000 2.285000 2.320000 ;
      RECT 2.035000  2.490000 2.285000 2.980000 ;
      RECT 2.050000  0.085000 2.380000 0.810000 ;
      RECT 2.475000  2.390000 3.755000 2.560000 ;
      RECT 2.475000  2.560000 2.805000 3.000000 ;
      RECT 2.975000  2.730000 3.305000 3.245000 ;
      RECT 3.050000  0.085000 3.380000 1.010000 ;
      RECT 3.505000  2.560000 3.755000 3.000000 ;
      RECT 3.940000  2.220000 4.205000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__nor4_2
MACRO sky130_fd_sc_hs__nor4_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.045000 1.300000 8.515000 1.630000 ;
        RECT 7.805000 1.180000 8.515000 1.300000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.350000 6.595000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.435000 1.350000 3.785000 1.780000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525000 1.350000 1.875000 1.780000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  3.214400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.010000 7.570000 1.130000 ;
        RECT 0.125000 1.130000 4.590000 1.180000 ;
        RECT 0.125000 1.180000 0.355000 1.950000 ;
        RECT 0.125000 1.950000 1.895000 2.120000 ;
        RECT 0.615000 0.350000 1.740000 1.010000 ;
        RECT 0.615000 2.120000 0.945000 2.735000 ;
        RECT 1.565000 2.120000 1.895000 2.735000 ;
        RECT 2.410000 0.350000 3.590000 1.010000 ;
        RECT 4.260000 0.350000 4.590000 0.960000 ;
        RECT 4.260000 0.960000 7.860000 1.010000 ;
        RECT 7.240000 0.340000 7.860000 0.960000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
      RECT 0.000000  3.245000 8.640000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 0.840000 ;
      RECT 0.115000  2.290000 0.445000 2.905000 ;
      RECT 0.115000  2.905000 2.265000 3.075000 ;
      RECT 1.145000  2.290000 1.395000 2.905000 ;
      RECT 1.910000  0.085000 2.240000 0.840000 ;
      RECT 2.095000  1.820000 2.265000 1.950000 ;
      RECT 2.095000  1.950000 4.145000 2.120000 ;
      RECT 2.095000  2.120000 2.265000 2.905000 ;
      RECT 2.465000  2.290000 2.795000 2.905000 ;
      RECT 2.465000  2.905000 6.075000 3.075000 ;
      RECT 2.970000  2.120000 3.190000 2.735000 ;
      RECT 3.365000  2.290000 3.695000 2.905000 ;
      RECT 3.760000  0.085000 4.090000 0.840000 ;
      RECT 3.895000  2.120000 4.145000 2.735000 ;
      RECT 4.375000  1.950000 8.525000 2.120000 ;
      RECT 4.375000  2.120000 4.625000 2.735000 ;
      RECT 4.760000  0.085000 7.070000 0.790000 ;
      RECT 4.825000  2.300000 5.155000 2.905000 ;
      RECT 5.340000  2.120000 5.560000 2.735000 ;
      RECT 5.745000  2.300000 6.075000 2.905000 ;
      RECT 6.255000  2.120000 6.525000 2.980000 ;
      RECT 6.695000  2.290000 7.025000 3.245000 ;
      RECT 7.195000  2.120000 7.525000 2.980000 ;
      RECT 7.695000  2.290000 8.025000 3.245000 ;
      RECT 8.030000  0.085000 8.360000 1.010000 ;
      RECT 8.195000  1.820000 8.525000 1.950000 ;
      RECT 8.195000  2.120000 8.525000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
  END
END sky130_fd_sc_hs__nor4_4
MACRO sky130_fd_sc_hs__nor4b_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985000 1.350000 1.315000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 1.350000 1.855000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.350000 2.395000 1.780000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.445000 1.110000 0.815000 1.440000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  0.879200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.290000 0.350000 1.620000 1.010000 ;
        RECT 1.290000 1.010000 3.275000 1.180000 ;
        RECT 2.300000 0.350000 2.630000 1.010000 ;
        RECT 2.905000 1.850000 3.275000 2.980000 ;
        RECT 3.105000 1.180000 3.275000 1.850000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.105000  0.350000 0.620000 0.940000 ;
      RECT 0.105000  0.940000 0.275000 1.820000 ;
      RECT 0.105000  1.820000 0.595000 1.950000 ;
      RECT 0.105000  1.950000 2.735000 2.120000 ;
      RECT 0.105000  2.120000 0.595000 2.700000 ;
      RECT 0.790000  0.085000 1.120000 0.940000 ;
      RECT 0.835000  2.290000 1.165000 3.245000 ;
      RECT 1.790000  0.085000 2.120000 0.840000 ;
      RECT 2.565000  1.350000 2.935000 1.680000 ;
      RECT 2.565000  1.680000 2.735000 1.950000 ;
      RECT 2.800000  0.085000 3.130000 0.840000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__nor4b_1
MACRO sky130_fd_sc_hs__nor4b_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.350000 5.635000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.295000 1.350000 4.195000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.350000 2.755000 1.780000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 1.470000 0.865000 1.800000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  1.323900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.250000 0.330000 1.580000 0.790000 ;
        RECT 1.250000 0.790000 2.770000 0.960000 ;
        RECT 1.655000 1.820000 1.825000 1.950000 ;
        RECT 1.655000 1.950000 3.095000 2.120000 ;
        RECT 1.655000 2.120000 1.825000 2.735000 ;
        RECT 2.440000 0.350000 2.770000 0.790000 ;
        RECT 2.440000 0.960000 2.770000 1.010000 ;
        RECT 2.440000 1.010000 5.145000 1.180000 ;
        RECT 2.925000 1.180000 3.095000 1.950000 ;
        RECT 3.440000 0.350000 3.770000 1.010000 ;
        RECT 4.815000 0.350000 5.145000 1.010000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.115000  0.350000 0.580000 1.130000 ;
      RECT 0.115000  1.130000 1.775000 1.300000 ;
      RECT 0.115000  1.300000 0.365000 2.980000 ;
      RECT 0.565000  1.970000 0.895000 3.245000 ;
      RECT 0.750000  0.085000 1.080000 0.960000 ;
      RECT 1.105000  1.300000 1.775000 1.550000 ;
      RECT 1.125000  1.820000 1.455000 2.905000 ;
      RECT 1.125000  2.905000 2.275000 3.075000 ;
      RECT 1.750000  0.085000 2.270000 0.600000 ;
      RECT 2.025000  2.290000 3.255000 2.460000 ;
      RECT 2.025000  2.460000 2.275000 2.905000 ;
      RECT 2.475000  2.630000 2.805000 2.905000 ;
      RECT 2.475000  2.905000 4.265000 3.075000 ;
      RECT 2.940000  0.085000 3.270000 0.840000 ;
      RECT 3.005000  2.460000 3.255000 2.735000 ;
      RECT 3.485000  1.950000 5.625000 2.120000 ;
      RECT 3.485000  2.120000 3.735000 2.735000 ;
      RECT 3.935000  2.290000 4.265000 2.905000 ;
      RECT 3.940000  0.085000 4.645000 0.790000 ;
      RECT 4.465000  2.120000 4.635000 2.980000 ;
      RECT 4.835000  2.290000 5.165000 3.245000 ;
      RECT 5.315000  0.085000 5.645000 1.130000 ;
      RECT 5.375000  2.120000 5.625000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_hs__nor4b_2
MACRO sky130_fd_sc_hs__nor4b_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.805000 1.350000 9.475000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885000 1.350000 7.555000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.920000 1.350000 5.155000 1.780000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.363000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.920000 0.550000 1.930000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  2.440600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.570000 0.350000 1.820000 0.980000 ;
        RECT 1.570000 0.980000 2.830000 1.150000 ;
        RECT 2.025000 1.820000 3.305000 1.950000 ;
        RECT 2.025000 1.950000 5.635000 1.990000 ;
        RECT 2.025000 1.990000 2.355000 2.735000 ;
        RECT 2.500000 0.350000 2.830000 0.980000 ;
        RECT 2.500000 1.150000 2.830000 1.300000 ;
        RECT 2.500000 1.300000 3.750000 1.470000 ;
        RECT 2.975000 1.990000 5.635000 2.120000 ;
        RECT 2.975000 2.120000 3.305000 2.735000 ;
        RECT 3.500000 0.350000 3.750000 1.010000 ;
        RECT 3.500000 1.010000 9.465000 1.180000 ;
        RECT 3.500000 1.180000 3.750000 1.300000 ;
        RECT 4.905000 0.350000 5.235000 1.010000 ;
        RECT 5.405000 1.180000 5.635000 1.950000 ;
        RECT 6.250000 0.350000 6.580000 1.010000 ;
        RECT 7.250000 0.350000 7.580000 1.010000 ;
        RECT 8.275000 0.350000 8.525000 1.010000 ;
        RECT 9.215000 0.350000 9.465000 1.010000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.115000  2.100000  0.365000 3.245000 ;
      RECT 0.275000  0.420000  0.890000 0.750000 ;
      RECT 0.565000  2.100000  0.895000 2.980000 ;
      RECT 0.720000  0.750000  0.890000 1.320000 ;
      RECT 0.720000  1.320000  2.330000 1.650000 ;
      RECT 0.720000  1.650000  0.890000 2.100000 ;
      RECT 1.060000  0.085000  1.390000 1.130000 ;
      RECT 1.075000  2.100000  1.345000 3.245000 ;
      RECT 1.575000  1.820000  1.825000 2.905000 ;
      RECT 1.575000  2.905000  3.755000 3.075000 ;
      RECT 2.000000  0.085000  2.330000 0.790000 ;
      RECT 2.525000  2.160000  2.805000 2.905000 ;
      RECT 3.000000  0.085000  3.330000 1.130000 ;
      RECT 3.475000  2.320000  5.705000 2.460000 ;
      RECT 3.475000  2.460000  4.755000 2.490000 ;
      RECT 3.475000  2.490000  3.755000 2.905000 ;
      RECT 3.925000  2.660000  4.255000 2.905000 ;
      RECT 3.925000  2.905000  7.715000 3.075000 ;
      RECT 3.930000  0.085000  4.735000 0.840000 ;
      RECT 4.425000  2.290000  5.705000 2.320000 ;
      RECT 4.425000  2.490000  4.755000 2.720000 ;
      RECT 4.925000  2.630000  5.255000 2.905000 ;
      RECT 5.405000  0.085000  6.080000 0.840000 ;
      RECT 5.440000  2.460000  5.705000 2.540000 ;
      RECT 5.935000  1.950000  9.965000 2.120000 ;
      RECT 5.935000  2.120000  6.265000 2.735000 ;
      RECT 6.435000  2.290000  6.765000 2.905000 ;
      RECT 6.750000  0.085000  7.080000 0.805000 ;
      RECT 6.935000  2.120000  7.265000 2.735000 ;
      RECT 7.465000  2.290000  7.715000 2.905000 ;
      RECT 7.750000  0.085000  8.105000 0.805000 ;
      RECT 7.885000  2.120000  8.115000 2.980000 ;
      RECT 8.285000  2.290000  8.535000 3.245000 ;
      RECT 8.705000  0.085000  9.035000 0.805000 ;
      RECT 8.735000  2.120000  9.065000 2.980000 ;
      RECT 9.265000  2.290000  9.515000 3.245000 ;
      RECT 9.635000  0.085000  9.965000 1.130000 ;
      RECT 9.715000  1.820000  9.965000 1.950000 ;
      RECT 9.715000  2.120000  9.965000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
  END
END sky130_fd_sc_hs__nor4b_4
MACRO sky130_fd_sc_hs__nor4bb_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.075000 1.350000 1.405000 2.150000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.915000 1.350000 2.275000 1.780000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.435000 1.550000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.450000 4.345000 1.780000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  0.848400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.445000 0.350000 1.775000 0.880000 ;
        RECT 1.445000 0.880000 3.235000 1.050000 ;
        RECT 1.445000 1.050000 1.775000 1.130000 ;
        RECT 1.575000 1.130000 1.745000 2.060000 ;
        RECT 1.575000 2.060000 3.455000 2.390000 ;
        RECT 2.860000 0.350000 3.235000 0.880000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.115000  0.680000 0.775000 1.010000 ;
      RECT 0.115000  1.820000 0.775000 2.560000 ;
      RECT 0.115000  2.560000 3.795000 2.730000 ;
      RECT 0.605000  1.010000 0.775000 1.820000 ;
      RECT 0.650000  2.900000 1.345000 3.245000 ;
      RECT 0.945000  0.085000 1.275000 1.130000 ;
      RECT 1.945000  0.085000 2.690000 0.680000 ;
      RECT 2.485000  1.350000 2.815000 1.720000 ;
      RECT 2.485000  1.720000 3.795000 1.890000 ;
      RECT 3.070000  1.220000 4.685000 1.260000 ;
      RECT 3.070000  1.260000 3.740000 1.550000 ;
      RECT 3.405000  0.085000 4.175000 0.920000 ;
      RECT 3.570000  1.090000 4.685000 1.220000 ;
      RECT 3.625000  1.890000 3.795000 2.560000 ;
      RECT 3.965000  2.100000 4.185000 3.245000 ;
      RECT 4.355000  0.540000 4.685000 1.090000 ;
      RECT 4.355000  2.100000 4.685000 2.980000 ;
      RECT 4.515000  1.260000 4.685000 2.100000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_hs__nor4bb_1
MACRO sky130_fd_sc_hs__nor4bb_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.310000 1.350000 7.075000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.860000 1.350000 6.115000 1.635000 ;
        RECT 5.405000 1.635000 6.115000 1.780000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525000 1.470000 1.315000 1.800000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.495000 1.470000 1.825000 1.800000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  1.198100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.890000 0.350000 3.220000 0.670000 ;
        RECT 2.890000 0.670000 4.285000 0.840000 ;
        RECT 2.975000 1.850000 4.285000 2.020000 ;
        RECT 2.975000 2.020000 3.225000 2.735000 ;
        RECT 3.955000 0.350000 4.285000 0.670000 ;
        RECT 3.955000 0.840000 4.285000 1.010000 ;
        RECT 3.955000 1.010000 6.575000 1.180000 ;
        RECT 4.115000 1.180000 4.285000 1.550000 ;
        RECT 4.115000 1.550000 4.675000 1.780000 ;
        RECT 4.115000 1.780000 4.285000 1.850000 ;
        RECT 4.965000 0.350000 5.215000 1.010000 ;
        RECT 6.325000 0.350000 6.575000 1.010000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.200000 0.085000 ;
      RECT 0.000000  3.245000 7.200000 3.415000 ;
      RECT 0.115000  1.130000 0.815000 1.300000 ;
      RECT 0.115000  1.300000 0.285000 1.970000 ;
      RECT 0.115000  1.970000 0.445000 2.980000 ;
      RECT 0.485000  0.360000 0.815000 0.710000 ;
      RECT 0.485000  0.710000 2.665000 0.880000 ;
      RECT 0.485000  0.880000 0.815000 1.130000 ;
      RECT 0.615000  1.970000 1.715000 3.245000 ;
      RECT 0.990000  0.085000 1.515000 0.540000 ;
      RECT 1.620000  1.050000 2.325000 1.300000 ;
      RECT 1.885000  1.970000 2.325000 2.140000 ;
      RECT 1.885000  2.140000 2.215000 2.980000 ;
      RECT 2.155000  1.300000 2.325000 1.350000 ;
      RECT 2.155000  1.350000 3.165000 1.680000 ;
      RECT 2.155000  1.680000 2.325000 1.970000 ;
      RECT 2.195000  0.085000 2.710000 0.540000 ;
      RECT 2.495000  0.880000 2.665000 1.010000 ;
      RECT 2.495000  1.010000 3.785000 1.180000 ;
      RECT 2.495000  1.850000 2.775000 2.905000 ;
      RECT 2.495000  2.905000 3.725000 3.075000 ;
      RECT 3.395000  2.190000 4.675000 2.360000 ;
      RECT 3.395000  2.360000 3.725000 2.905000 ;
      RECT 3.400000  0.085000 3.775000 0.500000 ;
      RECT 3.615000  1.180000 3.785000 1.350000 ;
      RECT 3.615000  1.350000 3.945000 1.680000 ;
      RECT 3.895000  2.530000 4.175000 2.905000 ;
      RECT 3.895000  2.905000 5.685000 3.075000 ;
      RECT 4.345000  2.360000 4.675000 2.735000 ;
      RECT 4.455000  0.085000 4.785000 0.840000 ;
      RECT 4.905000  1.820000 5.155000 1.950000 ;
      RECT 4.905000  1.950000 7.085000 2.120000 ;
      RECT 4.905000  2.120000 5.155000 2.735000 ;
      RECT 5.355000  2.290000 5.685000 2.905000 ;
      RECT 5.385000  0.085000 6.155000 0.840000 ;
      RECT 5.855000  2.120000 6.185000 2.980000 ;
      RECT 6.385000  2.290000 6.555000 3.245000 ;
      RECT 6.755000  0.085000 7.085000 1.130000 ;
      RECT 6.755000  2.120000 7.085000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
  END
END sky130_fd_sc_hs__nor4bb_2
MACRO sky130_fd_sc_hs__nor4bb_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 1.180000 2.495000 1.540000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.265000 1.320000 1.315000 1.650000 ;
        RECT 1.085000 1.650000 1.315000 1.710000 ;
        RECT 1.085000 1.710000 2.890000 1.880000 ;
        RECT 2.720000 1.255000 3.920000 1.585000 ;
        RECT 2.720000 1.585000 2.890000 1.710000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.363000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.095000 1.530000 9.955000 1.860000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.363000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.125000 1.450000 10.455000 1.780000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  2.544200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.615000 0.350000 0.945000 0.840000 ;
        RECT 0.615000 0.840000 2.915000 0.915000 ;
        RECT 0.615000 0.915000 5.775000 1.010000 ;
        RECT 0.615000 1.010000 0.945000 1.130000 ;
        RECT 1.615000 0.350000 1.945000 0.840000 ;
        RECT 2.665000 0.350000 2.915000 0.840000 ;
        RECT 2.665000 1.010000 5.775000 1.085000 ;
        RECT 3.595000 0.350000 3.845000 0.915000 ;
        RECT 4.515000 0.350000 4.845000 0.915000 ;
        RECT 5.525000 0.350000 5.775000 0.915000 ;
        RECT 5.525000 1.085000 5.775000 1.300000 ;
        RECT 5.525000 1.300000 6.615000 1.470000 ;
        RECT 5.990000 1.470000 6.320000 1.725000 ;
        RECT 5.990000 1.725000 7.230000 2.055000 ;
        RECT 6.445000 0.350000 6.775000 0.885000 ;
        RECT 6.445000 0.885000 8.035000 1.055000 ;
        RECT 6.445000 1.055000 6.615000 1.300000 ;
        RECT 7.705000 0.350000 8.035000 0.885000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.040000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 11.040000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  3.245000 11.040000 3.415000 ;
      RECT  0.115000  0.085000  0.445000 1.130000 ;
      RECT  0.115000  1.820000  0.445000 2.050000 ;
      RECT  0.115000  2.050000  3.390000 2.220000 ;
      RECT  0.115000  2.220000  0.445000 2.980000 ;
      RECT  0.615000  2.390000  2.885000 2.560000 ;
      RECT  0.615000  2.560000  0.945000 2.980000 ;
      RECT  1.115000  0.085000  1.445000 0.670000 ;
      RECT  1.115000  2.730000  1.445000 3.245000 ;
      RECT  1.645000  2.560000  1.895000 2.980000 ;
      RECT  2.065000  2.730000  2.435000 3.245000 ;
      RECT  2.115000  0.085000  2.445000 0.670000 ;
      RECT  2.635000  2.560000  2.885000 2.905000 ;
      RECT  2.635000  2.905000  3.890000 3.075000 ;
      RECT  3.060000  1.755000  4.260000 1.925000 ;
      RECT  3.060000  1.925000  3.390000 2.050000 ;
      RECT  3.060000  2.220000  3.390000 2.735000 ;
      RECT  3.085000  0.085000  3.415000 0.745000 ;
      RECT  3.560000  2.095000  3.890000 2.905000 ;
      RECT  4.015000  0.085000  4.345000 0.745000 ;
      RECT  4.090000  1.925000  4.260000 2.905000 ;
      RECT  4.090000  2.905000  8.490000 3.075000 ;
      RECT  4.345000  1.255000  5.355000 1.585000 ;
      RECT  4.470000  1.755000  4.800000 2.565000 ;
      RECT  4.470000  2.565000  8.035000 2.735000 ;
      RECT  5.015000  0.085000  5.345000 0.745000 ;
      RECT  5.185000  1.585000  5.355000 2.225000 ;
      RECT  5.185000  2.225000  7.570000 2.395000 ;
      RECT  5.945000  0.085000  6.275000 1.130000 ;
      RECT  6.785000  1.225000  8.375000 1.555000 ;
      RECT  6.945000  0.085000  7.535000 0.680000 ;
      RECT  7.400000  1.725000  8.875000 1.895000 ;
      RECT  7.400000  1.895000  7.570000 2.225000 ;
      RECT  7.760000  2.065000  8.035000 2.565000 ;
      RECT  8.205000  0.085000  8.750000 0.680000 ;
      RECT  8.205000  0.850000  9.090000 1.020000 ;
      RECT  8.205000  1.020000  8.375000 1.225000 ;
      RECT  8.205000  2.065000  8.490000 2.905000 ;
      RECT  8.545000  1.190000  9.585000 1.360000 ;
      RECT  8.545000  1.360000  8.875000 1.725000 ;
      RECT  8.705000  1.895000  8.875000 2.030000 ;
      RECT  8.705000  2.030000  9.575000 2.200000 ;
      RECT  8.790000  2.370000  9.120000 3.245000 ;
      RECT  8.920000  0.255000  9.925000 0.425000 ;
      RECT  8.920000  0.425000  9.090000 0.850000 ;
      RECT  9.260000  0.670000  9.585000 1.190000 ;
      RECT  9.300000  2.200000  9.575000 2.980000 ;
      RECT  9.755000  0.425000  9.925000 1.110000 ;
      RECT  9.755000  1.110000 10.925000 1.280000 ;
      RECT  9.775000  2.100000  9.945000 3.245000 ;
      RECT 10.095000  0.085000 10.495000 0.940000 ;
      RECT 10.145000  1.950000 10.925000 2.120000 ;
      RECT 10.145000  2.120000 10.395000 2.980000 ;
      RECT 10.595000  2.290000 10.925000 3.245000 ;
      RECT 10.665000  0.350000 10.925000 1.110000 ;
      RECT 10.755000  1.280000 10.925000 1.950000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
  END
END sky130_fd_sc_hs__nor4bb_4
MACRO sky130_fd_sc_hs__o2111a_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405000 1.300000 3.735000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.715000 1.415000 3.235000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.415000 2.505000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.545000 0.440000 1.875000 1.900000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.550000 1.335000 1.880000 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.533900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.350000 0.355000 1.040000 ;
        RECT 0.095000 1.040000 0.265000 1.820000 ;
        RECT 0.095000 1.820000 0.445000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.435000  1.210000 1.330000 1.380000 ;
      RECT 0.435000  1.380000 0.785000 1.550000 ;
      RECT 0.535000  0.085000 0.865000 1.040000 ;
      RECT 0.615000  1.550000 0.785000 2.070000 ;
      RECT 0.615000  2.070000 2.865000 2.240000 ;
      RECT 0.615000  2.410000 0.945000 3.245000 ;
      RECT 1.080000  0.350000 1.330000 1.210000 ;
      RECT 1.195000  2.240000 2.865000 2.245000 ;
      RECT 1.195000  2.245000 1.525000 2.925000 ;
      RECT 1.740000  2.455000 2.290000 3.245000 ;
      RECT 2.380000  0.350000 2.710000 0.960000 ;
      RECT 2.380000  0.960000 3.710000 1.130000 ;
      RECT 2.535000  2.045000 2.865000 2.070000 ;
      RECT 2.535000  2.245000 2.865000 2.925000 ;
      RECT 2.880000  0.085000 3.210000 0.790000 ;
      RECT 3.380000  0.350000 3.710000 0.960000 ;
      RECT 3.405000  1.950000 3.735000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__o2111a_1
MACRO sky130_fd_sc_hs__o2111a_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.835000 1.550000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015000 1.180000 1.345000 1.550000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.180000 1.915000 1.550000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.155000 1.350000 2.755000 1.780000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925000 1.350000 3.255000 1.780000 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.855000 1.820000 4.185000 2.980000 ;
        RECT 3.910000 0.350000 4.240000 1.130000 ;
        RECT 4.015000 1.130000 4.185000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.250000  0.350000 0.580000 0.840000 ;
      RECT 0.250000  0.840000 1.720000 1.010000 ;
      RECT 0.295000  1.820000 0.625000 3.245000 ;
      RECT 0.750000  0.085000 1.220000 0.670000 ;
      RECT 1.285000  1.820000 1.615000 1.950000 ;
      RECT 1.285000  1.950000 3.685000 2.120000 ;
      RECT 1.285000  2.120000 1.615000 2.860000 ;
      RECT 1.390000  0.350000 1.720000 0.840000 ;
      RECT 1.785000  2.290000 2.115000 3.245000 ;
      RECT 2.375000  2.120000 2.705000 2.880000 ;
      RECT 2.850000  0.350000 3.180000 1.010000 ;
      RECT 2.850000  1.010000 3.685000 1.180000 ;
      RECT 2.875000  2.290000 3.685000 3.245000 ;
      RECT 3.410000  0.085000 3.740000 0.825000 ;
      RECT 3.515000  1.180000 3.685000 1.300000 ;
      RECT 3.515000  1.300000 3.845000 1.630000 ;
      RECT 3.515000  1.630000 3.685000 1.950000 ;
      RECT 4.355000  1.820000 4.685000 3.245000 ;
      RECT 4.420000  0.085000 4.685000 1.130000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_hs__o2111a_2
MACRO sky130_fd_sc_hs__o2111a_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.522000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.325000 1.450000 5.655000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.522000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.450000 5.155000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.474000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.985000 1.450000 3.315000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.474000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.450000 1.795000 1.780000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.474000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.450000 0.550000 1.780000 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  1.142400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.185000 0.350000 6.515000 1.010000 ;
        RECT 6.185000 1.010000 8.035000 1.180000 ;
        RECT 6.315000 1.850000 7.545000 2.180000 ;
        RECT 6.315000 2.180000 6.590000 2.980000 ;
        RECT 7.185000 0.350000 7.515000 1.010000 ;
        RECT 7.295000 1.480000 8.035000 1.650000 ;
        RECT 7.295000 1.650000 7.545000 1.850000 ;
        RECT 7.295000 2.180000 7.545000 2.980000 ;
        RECT 7.805000 1.180000 8.035000 1.480000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.115000  0.255000 2.250000 0.425000 ;
      RECT 0.115000  0.425000 1.230000 0.600000 ;
      RECT 0.115000  0.600000 0.380000 1.115000 ;
      RECT 0.115000  1.950000 6.145000 2.120000 ;
      RECT 0.115000  2.120000 0.445000 2.820000 ;
      RECT 0.550000  0.770000 0.890000 1.130000 ;
      RECT 0.615000  2.315000 0.945000 3.245000 ;
      RECT 0.720000  1.130000 0.890000 1.950000 ;
      RECT 1.060000  0.600000 1.230000 1.130000 ;
      RECT 1.115000  2.120000 1.445000 2.820000 ;
      RECT 1.410000  0.595000 1.740000 0.710000 ;
      RECT 1.410000  0.710000 3.125000 0.880000 ;
      RECT 1.410000  0.880000 1.740000 1.130000 ;
      RECT 1.615000  2.315000 1.945000 3.245000 ;
      RECT 1.920000  0.425000 2.250000 0.540000 ;
      RECT 2.150000  1.940000 2.480000 1.950000 ;
      RECT 2.150000  2.120000 2.480000 2.820000 ;
      RECT 2.365000  1.050000 3.555000 1.110000 ;
      RECT 2.365000  1.110000 5.505000 1.280000 ;
      RECT 2.365000  1.280000 2.775000 1.300000 ;
      RECT 2.685000  2.315000 3.015000 3.245000 ;
      RECT 2.875000  0.520000 3.125000 0.710000 ;
      RECT 3.220000  2.120000 3.550000 2.905000 ;
      RECT 3.220000  2.905000 4.550000 3.075000 ;
      RECT 3.305000  0.520000 3.555000 1.050000 ;
      RECT 3.720000  2.290000 5.610000 2.460000 ;
      RECT 3.720000  2.460000 4.050000 2.735000 ;
      RECT 3.735000  0.085000 4.065000 0.940000 ;
      RECT 4.220000  2.630000 4.550000 2.905000 ;
      RECT 4.235000  0.520000 4.565000 1.110000 ;
      RECT 4.780000  2.630000 5.110000 3.245000 ;
      RECT 4.825000  0.085000 5.155000 0.940000 ;
      RECT 5.280000  2.460000 5.610000 2.980000 ;
      RECT 5.335000  0.350000 5.505000 1.110000 ;
      RECT 5.685000  0.085000 6.015000 1.130000 ;
      RECT 5.815000  2.290000 6.145000 3.245000 ;
      RECT 5.975000  1.350000 7.125000 1.680000 ;
      RECT 5.975000  1.680000 6.145000 1.950000 ;
      RECT 6.685000  0.085000 7.015000 0.815000 ;
      RECT 6.765000  2.350000 7.095000 3.245000 ;
      RECT 7.685000  0.085000 8.015000 0.815000 ;
      RECT 7.715000  1.820000 8.045000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_hs__o2111a_4
MACRO sky130_fd_sc_hs__o2111ai_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925000 1.180000 3.255000 1.550000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.200000 1.180000 2.755000 1.550000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.595000 1.180000 1.990000 1.550000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 0.440000 1.425000 1.550000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.580000 1.180000 0.910000 1.550000 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  1.162500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.350000 0.785000 1.010000 ;
        RECT 0.115000 1.010000 0.285000 1.720000 ;
        RECT 0.115000 1.720000 2.315000 1.890000 ;
        RECT 0.880000 1.890000 1.315000 2.980000 ;
        RECT 1.985000 1.890000 2.315000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.380000  2.060000 0.710000 3.245000 ;
      RECT 1.485000  2.060000 1.815000 3.245000 ;
      RECT 1.825000  0.350000 2.155000 0.840000 ;
      RECT 1.825000  0.840000 3.245000 1.010000 ;
      RECT 2.325000  0.085000 2.745000 0.600000 ;
      RECT 2.890000  1.820000 3.220000 3.245000 ;
      RECT 2.915000  0.350000 3.245000 0.840000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__o2111ai_1
MACRO sky130_fd_sc_hs__o2111ai_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925000 1.350000 5.635000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.350000 4.675000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.350000 3.715000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.345000 1.300000 2.015000 1.630000 ;
        RECT 1.565000 1.180000 1.795000 1.300000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.435000 1.550000 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  1.551200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.180000 0.935000 1.800000 ;
        RECT 0.605000 1.800000 1.885000 1.950000 ;
        RECT 0.605000 1.950000 4.245000 1.970000 ;
        RECT 0.605000 1.970000 0.935000 2.980000 ;
        RECT 0.690000 0.595000 0.940000 1.130000 ;
        RECT 0.690000 1.130000 0.935000 1.180000 ;
        RECT 1.555000 1.970000 4.245000 2.120000 ;
        RECT 1.555000 2.120000 1.885000 2.980000 ;
        RECT 2.455000 2.120000 2.785000 2.980000 ;
        RECT 3.915000 2.120000 4.245000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.155000  1.820000 0.405000 3.245000 ;
      RECT 0.180000  0.255000 1.290000 0.425000 ;
      RECT 0.180000  0.425000 0.510000 1.010000 ;
      RECT 1.105000  2.140000 1.355000 3.245000 ;
      RECT 1.120000  0.425000 1.290000 0.840000 ;
      RECT 1.120000  0.840000 2.300000 1.010000 ;
      RECT 1.120000  1.010000 1.290000 1.130000 ;
      RECT 1.470000  0.255000 3.360000 0.425000 ;
      RECT 1.470000  0.425000 1.800000 0.670000 ;
      RECT 1.970000  0.595000 2.300000 0.840000 ;
      RECT 1.970000  1.010000 2.300000 1.130000 ;
      RECT 2.085000  2.290000 2.255000 3.245000 ;
      RECT 2.530000  0.595000 2.860000 1.010000 ;
      RECT 2.530000  1.010000 5.600000 1.180000 ;
      RECT 2.985000  2.290000 3.235000 3.245000 ;
      RECT 3.030000  0.425000 3.360000 0.840000 ;
      RECT 3.465000  2.290000 3.715000 2.905000 ;
      RECT 3.465000  2.905000 4.615000 3.075000 ;
      RECT 3.540000  0.350000 3.710000 1.010000 ;
      RECT 3.890000  0.085000 4.220000 0.840000 ;
      RECT 4.420000  0.350000 4.670000 1.010000 ;
      RECT 4.445000  1.950000 5.645000 2.120000 ;
      RECT 4.445000  2.120000 4.615000 2.905000 ;
      RECT 4.815000  2.290000 5.145000 3.245000 ;
      RECT 4.840000  0.085000 5.170000 0.840000 ;
      RECT 5.315000  2.120000 5.645000 2.980000 ;
      RECT 5.350000  0.350000 5.600000 1.010000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_hs__o2111ai_2
MACRO sky130_fd_sc_hs__o2111ai_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.285000 1.350000 7.635000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.805000 1.350000 9.490000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.350000 6.115000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.210000 1.300000 4.195000 1.630000 ;
        RECT 3.965000 1.630000 4.195000 1.780000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.350000 1.780000 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  3.411800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 1.950000 9.515000 1.970000 ;
        RECT 0.115000 1.970000 2.200000 2.120000 ;
        RECT 0.115000 2.120000 1.200000 2.980000 ;
        RECT 0.615000 0.770000 1.805000 1.130000 ;
        RECT 1.565000 1.130000 1.805000 1.550000 ;
        RECT 1.565000 1.550000 2.040000 1.780000 ;
        RECT 1.870000 1.780000 2.040000 1.800000 ;
        RECT 1.870000 1.800000 3.520000 1.950000 ;
        RECT 1.870000 2.120000 2.200000 2.980000 ;
        RECT 3.190000 1.970000 9.515000 2.120000 ;
        RECT 3.190000 2.120000 3.520000 2.980000 ;
        RECT 4.190000 2.120000 4.520000 2.980000 ;
        RECT 8.185000 2.120000 8.515000 2.735000 ;
        RECT 9.185000 2.120000 9.515000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.115000  0.350000  2.155000 0.600000 ;
      RECT 0.115000  0.600000  0.445000 1.130000 ;
      RECT 1.370000  2.290000  1.700000 3.245000 ;
      RECT 1.985000  0.600000  2.155000 0.815000 ;
      RECT 1.985000  0.815000  3.955000 1.130000 ;
      RECT 2.335000  0.350000  5.805000 0.645000 ;
      RECT 2.370000  2.140000  3.020000 3.245000 ;
      RECT 3.690000  2.290000  4.020000 3.245000 ;
      RECT 4.185000  0.815000  4.515000 0.850000 ;
      RECT 4.185000  0.850000  6.305000 1.010000 ;
      RECT 4.185000  1.010000  9.965000 1.130000 ;
      RECT 4.750000  2.290000  8.015000 2.460000 ;
      RECT 4.750000  2.460000  6.165000 2.980000 ;
      RECT 5.045000  1.130000  9.965000 1.180000 ;
      RECT 5.475000  0.645000  5.805000 0.680000 ;
      RECT 5.975000  0.350000  6.305000 0.850000 ;
      RECT 6.335000  2.630000  6.585000 3.245000 ;
      RECT 6.475000  0.085000  6.805000 0.820000 ;
      RECT 6.785000  2.460000  7.115000 2.980000 ;
      RECT 6.985000  0.350000  7.155000 1.010000 ;
      RECT 7.315000  2.630000  7.485000 3.245000 ;
      RECT 7.335000  0.085000  7.665000 0.820000 ;
      RECT 7.685000  2.460000  8.015000 2.905000 ;
      RECT 7.685000  2.905000  9.965000 3.075000 ;
      RECT 7.845000  0.350000  8.095000 1.010000 ;
      RECT 8.265000  0.085000  8.595000 0.820000 ;
      RECT 8.685000  2.290000  9.015000 2.905000 ;
      RECT 8.775000  0.350000  9.025000 1.010000 ;
      RECT 9.205000  0.085000  9.535000 0.820000 ;
      RECT 9.715000  0.350000  9.965000 1.010000 ;
      RECT 9.715000  1.820000  9.965000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
  END
END sky130_fd_sc_hs__o2111ai_4
MACRO sky130_fd_sc_hs__o211a_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.335000 1.470000 2.005000 1.800000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.325000 0.255000 3.715000 0.640000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.490000 3.335000 1.800000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.635000 1.490000 4.195000 1.800000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.350000 0.445000 1.130000 ;
        RECT 0.085000 1.130000 0.255000 1.820000 ;
        RECT 0.085000 1.820000 0.445000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.425000  1.320000 1.095000 1.650000 ;
      RECT 0.615000  0.085000 0.945000 1.130000 ;
      RECT 0.615000  2.310000 1.855000 3.245000 ;
      RECT 0.925000  1.650000 1.095000 1.970000 ;
      RECT 0.925000  1.970000 4.205000 2.140000 ;
      RECT 1.265000  0.660000 1.595000 1.130000 ;
      RECT 1.265000  1.130000 2.495000 1.300000 ;
      RECT 1.765000  0.085000 2.155000 0.925000 ;
      RECT 2.325000  0.810000 3.185000 0.980000 ;
      RECT 2.325000  0.980000 2.495000 1.130000 ;
      RECT 2.395000  1.940000 2.835000 1.970000 ;
      RECT 2.395000  2.140000 2.725000 2.980000 ;
      RECT 2.665000  1.150000 4.135000 1.320000 ;
      RECT 2.665000  1.320000 2.835000 1.940000 ;
      RECT 2.895000  2.310000 3.705000 3.245000 ;
      RECT 3.760000  0.835000 4.135000 1.150000 ;
      RECT 3.875000  2.140000 4.205000 2.980000 ;
      RECT 3.885000  0.660000 4.135000 0.835000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__o211a_1
MACRO sky130_fd_sc_hs__o211a_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965000 1.350000 2.295000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.335000 1.350000 1.795000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.350000 1.125000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.435000 1.550000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.895000 1.820000 3.225000 2.980000 ;
        RECT 2.980000 0.350000 3.235000 1.130000 ;
        RECT 3.005000 1.130000 3.235000 1.410000 ;
        RECT 3.005000 1.410000 3.225000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.105000  1.820000 0.435000 1.950000 ;
      RECT 0.105000  1.950000 2.675000 2.120000 ;
      RECT 0.105000  2.120000 0.435000 2.860000 ;
      RECT 0.130000  0.350000 0.775000 1.010000 ;
      RECT 0.605000  1.010000 2.675000 1.180000 ;
      RECT 0.605000  2.290000 0.935000 3.245000 ;
      RECT 1.025000  0.350000 1.355000 0.670000 ;
      RECT 1.025000  0.670000 2.350000 0.840000 ;
      RECT 1.105000  2.120000 1.435000 2.860000 ;
      RECT 1.525000  0.085000 1.775000 0.500000 ;
      RECT 2.020000  0.350000 2.350000 0.670000 ;
      RECT 2.025000  2.290000 2.725000 3.245000 ;
      RECT 2.505000  1.180000 2.675000 1.300000 ;
      RECT 2.505000  1.300000 2.835000 1.630000 ;
      RECT 2.505000  1.630000 2.675000 1.950000 ;
      RECT 2.550000  0.085000 2.800000 0.840000 ;
      RECT 3.395000  1.820000 3.725000 3.245000 ;
      RECT 3.410000  0.085000 3.740000 1.130000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__o211a_2
MACRO sky130_fd_sc_hs__o211a_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.075000 1.450000 6.595000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925000 1.450000 5.835000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.444000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505000 1.435000 2.835000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.444000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.450000 1.450000 3.780000 1.780000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.960000 1.760000 1.130000 ;
        RECT 0.125000 1.130000 0.355000 1.800000 ;
        RECT 0.125000 1.800000 1.945000 1.970000 ;
        RECT 0.580000 0.350000 0.830000 0.960000 ;
        RECT 0.615000 1.970000 0.945000 2.980000 ;
        RECT 1.510000 0.350000 1.760000 0.960000 ;
        RECT 1.615000 1.970000 1.945000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.720000 0.085000 ;
      RECT 0.000000  3.245000 6.720000 3.415000 ;
      RECT 0.115000  2.140000 0.445000 3.245000 ;
      RECT 0.150000  0.085000 0.400000 0.790000 ;
      RECT 0.615000  1.300000 2.285000 1.630000 ;
      RECT 1.010000  0.085000 1.340000 0.790000 ;
      RECT 1.115000  2.140000 1.445000 3.245000 ;
      RECT 1.940000  0.085000 2.270000 1.130000 ;
      RECT 2.115000  1.630000 2.285000 1.950000 ;
      RECT 2.115000  1.950000 5.655000 2.120000 ;
      RECT 2.115000  2.290000 2.445000 3.245000 ;
      RECT 2.530000  0.255000 4.650000 0.425000 ;
      RECT 2.530000  0.425000 2.780000 1.265000 ;
      RECT 2.775000  2.120000 3.105000 2.815000 ;
      RECT 3.040000  0.595000 4.220000 0.765000 ;
      RECT 3.040000  0.765000 3.210000 1.285000 ;
      RECT 3.275000  2.290000 3.605000 3.245000 ;
      RECT 3.390000  0.935000 3.720000 1.110000 ;
      RECT 3.390000  1.110000 4.120000 1.280000 ;
      RECT 3.790000  2.120000 4.120000 2.815000 ;
      RECT 3.890000  0.765000 4.220000 0.940000 ;
      RECT 3.950000  1.280000 4.120000 1.950000 ;
      RECT 4.325000  2.290000 4.655000 3.245000 ;
      RECT 4.400000  0.425000 4.650000 1.110000 ;
      RECT 4.400000  1.110000 6.605000 1.280000 ;
      RECT 4.400000  1.280000 4.650000 1.285000 ;
      RECT 4.825000  2.290000 5.155000 2.905000 ;
      RECT 4.825000  2.905000 6.105000 3.075000 ;
      RECT 4.830000  0.085000 5.175000 0.935000 ;
      RECT 5.325000  2.120000 5.655000 2.735000 ;
      RECT 5.345000  0.605000 5.595000 1.110000 ;
      RECT 5.775000  0.085000 6.105000 0.940000 ;
      RECT 5.855000  1.950000 6.105000 2.905000 ;
      RECT 6.275000  0.605000 6.605000 1.110000 ;
      RECT 6.275000  1.950000 6.605000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
  END
END sky130_fd_sc_hs__o211a_4
MACRO sky130_fd_sc_hs__o211ai_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.880000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.300000 0.435000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.550000 1.165000 1.630000 ;
        RECT 0.605000 1.630000 0.835000 2.890000 ;
        RECT 0.665000 1.300000 1.165000 1.550000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.405000 1.300000 1.795000 1.630000 ;
        RECT 1.565000 0.440000 1.795000 1.300000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975000 1.180000 2.305000 1.550000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.427600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.125000 1.800000 2.770000 1.970000 ;
        RECT 1.125000 1.970000 1.455000 2.980000 ;
        RECT 2.045000 0.440000 2.770000 1.010000 ;
        RECT 2.205000 1.970000 2.770000 2.980000 ;
        RECT 2.595000 1.010000 2.770000 1.800000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.880000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.880000 0.085000 ;
      RECT 0.000000  3.245000 2.880000 3.415000 ;
      RECT 0.115000  1.950000 0.365000 3.245000 ;
      RECT 0.135000  0.350000 0.465000 0.960000 ;
      RECT 0.135000  0.960000 1.395000 1.130000 ;
      RECT 0.635000  0.085000 0.965000 0.780000 ;
      RECT 1.145000  0.350000 1.395000 0.960000 ;
      RECT 1.705000  2.140000 2.035000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
  END
END sky130_fd_sc_hs__o211ai_1
MACRO sky130_fd_sc_hs__o211ai_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.685000 1.320000 4.695000 1.650000 ;
        RECT 4.365000 1.180000 4.695000 1.320000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.435000 1.320000 3.445000 1.650000 ;
        RECT 2.435000 1.650000 3.235000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.350000 2.015000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 0.550000 1.780000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.215200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.560000 0.595000 0.890000 1.180000 ;
        RECT 0.595000 1.950000 3.285000 2.120000 ;
        RECT 0.595000 2.120000 0.925000 2.980000 ;
        RECT 0.720000 1.180000 0.890000 1.950000 ;
        RECT 1.495000 2.120000 1.825000 2.980000 ;
        RECT 2.955000 2.120000 3.285000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.130000  0.255000 2.330000 0.425000 ;
      RECT 0.130000  0.425000 0.380000 1.180000 ;
      RECT 0.145000  1.950000 0.395000 3.245000 ;
      RECT 1.060000  0.425000 2.330000 0.730000 ;
      RECT 1.060000  0.730000 1.390000 1.180000 ;
      RECT 1.125000  2.290000 1.295000 3.245000 ;
      RECT 1.560000  0.900000 1.890000 0.980000 ;
      RECT 1.560000  0.980000 4.160000 1.150000 ;
      RECT 1.560000  1.150000 1.890000 1.180000 ;
      RECT 2.025000  2.290000 2.275000 3.245000 ;
      RECT 2.505000  2.290000 2.755000 2.905000 ;
      RECT 2.505000  2.905000 3.655000 3.075000 ;
      RECT 2.560000  0.085000 2.890000 0.795000 ;
      RECT 3.070000  0.350000 3.240000 0.980000 ;
      RECT 3.420000  0.085000 3.750000 0.795000 ;
      RECT 3.485000  1.820000 4.685000 1.990000 ;
      RECT 3.485000  1.990000 3.655000 2.905000 ;
      RECT 3.855000  2.160000 4.185000 3.245000 ;
      RECT 3.935000  0.350000 4.160000 0.980000 ;
      RECT 4.330000  0.085000 4.685000 1.010000 ;
      RECT 4.355000  1.990000 4.685000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_hs__o211ai_2
MACRO sky130_fd_sc_hs__o211ai_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.795000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.350000 4.195000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.350000 5.635000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.870000 1.350000 7.075000 1.780000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.915200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.430000 1.950000 8.035000 2.120000 ;
        RECT 2.430000 2.120000 2.760000 2.735000 ;
        RECT 3.380000 2.120000 3.710000 2.735000 ;
        RECT 4.940000 2.120000 5.270000 2.980000 ;
        RECT 5.940000 2.120000 6.270000 2.980000 ;
        RECT 6.505000 0.595000 6.675000 1.010000 ;
        RECT 6.505000 1.010000 7.545000 1.180000 ;
        RECT 7.365000 0.595000 7.545000 1.010000 ;
        RECT 7.365000 1.180000 7.545000 1.550000 ;
        RECT 7.365000 1.550000 8.035000 1.950000 ;
        RECT 7.545000 2.120000 8.035000 2.890000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.115000  0.350000 0.445000 1.010000 ;
      RECT 0.115000  1.010000 5.765000 1.180000 ;
      RECT 0.130000  1.950000 2.260000 2.120000 ;
      RECT 0.130000  2.120000 0.460000 2.980000 ;
      RECT 0.615000  0.085000 0.945000 0.840000 ;
      RECT 0.660000  2.290000 0.830000 3.245000 ;
      RECT 1.030000  2.120000 1.360000 2.980000 ;
      RECT 1.125000  0.350000 1.375000 1.010000 ;
      RECT 1.545000  0.085000 1.875000 0.840000 ;
      RECT 1.560000  2.290000 1.730000 3.245000 ;
      RECT 1.930000  2.120000 2.260000 2.905000 ;
      RECT 1.930000  2.905000 4.210000 3.075000 ;
      RECT 2.055000  0.350000 2.225000 1.010000 ;
      RECT 2.405000  0.085000 2.735000 0.840000 ;
      RECT 2.915000  0.350000 3.085000 1.010000 ;
      RECT 2.960000  2.290000 3.210000 2.905000 ;
      RECT 3.265000  0.085000 3.595000 0.840000 ;
      RECT 3.795000  0.350000 3.965000 0.820000 ;
      RECT 3.795000  0.820000 4.905000 1.010000 ;
      RECT 3.880000  2.290000 4.210000 2.905000 ;
      RECT 4.145000  0.255000 8.045000 0.425000 ;
      RECT 4.145000  0.425000 5.255000 0.650000 ;
      RECT 4.440000  2.290000 4.770000 3.245000 ;
      RECT 5.085000  0.650000 5.255000 0.840000 ;
      RECT 5.435000  0.595000 5.765000 1.010000 ;
      RECT 5.440000  2.290000 5.770000 3.245000 ;
      RECT 5.995000  0.425000 6.325000 1.180000 ;
      RECT 6.440000  2.290000 7.290000 3.245000 ;
      RECT 6.855000  0.425000 7.185000 0.840000 ;
      RECT 7.715000  0.425000 8.045000 1.180000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_hs__o211ai_4
MACRO sky130_fd_sc_hs__o21a_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.880000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 1.300000 2.775000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.715000 1.445000 2.275000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.445000 1.435000 1.780000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.350000 0.365000 1.820000 ;
        RECT 0.115000 1.820000 0.445000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.880000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.880000 0.085000 ;
      RECT 0.000000  3.245000 2.880000 3.415000 ;
      RECT 0.535000  1.105000 1.395000 1.275000 ;
      RECT 0.535000  1.275000 0.865000 1.550000 ;
      RECT 0.545000  0.085000 0.875000 0.935000 ;
      RECT 0.615000  2.290000 1.180000 3.245000 ;
      RECT 0.695000  1.550000 0.865000 1.950000 ;
      RECT 0.695000  1.950000 1.690000 2.120000 ;
      RECT 1.145000  0.350000 1.395000 1.105000 ;
      RECT 1.360000  2.120000 1.690000 2.795000 ;
      RECT 1.575000  0.350000 1.825000 0.960000 ;
      RECT 1.575000  0.960000 2.765000 1.130000 ;
      RECT 2.005000  0.085000 2.335000 0.790000 ;
      RECT 2.435000  1.950000 2.765000 3.245000 ;
      RECT 2.515000  0.350000 2.765000 0.960000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
  END
END sky130_fd_sc_hs__o21a_1
MACRO sky130_fd_sc_hs__o21a_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.835000 1.550000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055000 1.180000 1.385000 1.550000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.180000 1.955000 1.550000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.465000 1.720000 3.295000 1.890000 ;
        RECT 2.465000 1.890000 2.795000 2.980000 ;
        RECT 2.965000 0.350000 3.295000 1.720000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.250000  0.340000 0.580000 0.840000 ;
      RECT 0.250000  0.840000 1.735000 1.010000 ;
      RECT 0.335000  1.820000 0.665000 3.245000 ;
      RECT 0.750000  0.085000 1.235000 0.600000 ;
      RECT 1.325000  1.720000 2.295000 1.890000 ;
      RECT 1.325000  1.890000 1.655000 2.860000 ;
      RECT 1.405000  0.340000 1.735000 0.840000 ;
      RECT 1.905000  0.340000 2.295000 1.010000 ;
      RECT 1.965000  2.060000 2.295000 3.245000 ;
      RECT 2.125000  1.010000 2.295000 1.220000 ;
      RECT 2.125000  1.220000 2.645000 1.550000 ;
      RECT 2.125000  1.550000 2.295000 1.720000 ;
      RECT 2.465000  0.085000 2.795000 1.050000 ;
      RECT 2.965000  2.060000 3.295000 3.245000 ;
      RECT 3.475000  0.085000 3.725000 1.130000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__o21a_2
MACRO sky130_fd_sc_hs__o21a_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.795000 1.445000 2.275000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.835000 1.445000 1.505000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.444000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 1.515000 3.235000 1.780000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.815000 1.720000 5.635000 1.780000 ;
        RECT 3.815000 1.780000 5.145000 1.890000 ;
        RECT 3.815000 1.890000 4.145000 2.980000 ;
        RECT 3.990000 0.330000 4.240000 0.835000 ;
        RECT 3.990000 0.835000 5.135000 1.005000 ;
        RECT 4.815000 1.890000 5.145000 2.980000 ;
        RECT 4.965000 0.350000 5.135000 0.835000 ;
        RECT 4.965000 1.005000 5.135000 1.550000 ;
        RECT 4.965000 1.550000 5.635000 1.720000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.115000  0.605000 0.445000 1.105000 ;
      RECT 0.115000  1.105000 2.390000 1.275000 ;
      RECT 0.115000  1.275000 0.445000 1.285000 ;
      RECT 0.115000  1.915000 0.445000 3.245000 ;
      RECT 0.615000  0.085000 0.950000 0.935000 ;
      RECT 0.615000  1.950000 0.865000 2.905000 ;
      RECT 0.615000  2.905000 1.895000 3.075000 ;
      RECT 1.065000  1.950000 3.575000 2.120000 ;
      RECT 1.065000  2.120000 1.395000 2.735000 ;
      RECT 1.130000  0.605000 1.380000 1.105000 ;
      RECT 1.560000  0.085000 1.890000 0.935000 ;
      RECT 1.565000  2.290000 1.895000 2.905000 ;
      RECT 2.060000  0.265000 3.330000 0.435000 ;
      RECT 2.060000  0.435000 2.390000 1.105000 ;
      RECT 2.065000  2.290000 2.395000 3.245000 ;
      RECT 2.565000  2.120000 2.895000 2.795000 ;
      RECT 2.570000  0.605000 2.820000 1.175000 ;
      RECT 2.570000  1.175000 4.795000 1.345000 ;
      RECT 3.000000  0.435000 3.330000 1.005000 ;
      RECT 3.135000  2.300000 3.615000 3.245000 ;
      RECT 3.405000  1.345000 4.795000 1.550000 ;
      RECT 3.405000  1.550000 3.575000 1.950000 ;
      RECT 3.560000  0.085000 3.810000 1.005000 ;
      RECT 4.315000  2.060000 4.645000 3.245000 ;
      RECT 4.420000  0.085000 4.785000 0.665000 ;
      RECT 5.315000  0.085000 5.645000 1.130000 ;
      RECT 5.315000  1.950000 5.645000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_hs__o21a_4
MACRO sky130_fd_sc_hs__o21ai_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.400000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 0.555000 1.550000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 1.350000 1.395000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.350000 2.275000 1.780000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.828300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.725000 1.010000 2.285000 1.180000 ;
        RECT 0.725000 1.180000 0.895000 1.950000 ;
        RECT 0.725000 1.950000 1.545000 2.980000 ;
        RECT 1.955000 0.350000 2.285000 1.010000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.400000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.400000 0.085000 ;
      RECT 0.000000  3.245000 2.400000 3.415000 ;
      RECT 0.115000  0.350000 0.420000 0.670000 ;
      RECT 0.115000  0.670000 1.785000 0.840000 ;
      RECT 0.115000  0.840000 0.445000 1.010000 ;
      RECT 0.305000  1.820000 0.555000 3.245000 ;
      RECT 0.605000  0.085000 1.295000 0.500000 ;
      RECT 1.480000  0.350000 1.785000 0.670000 ;
      RECT 1.870000  1.950000 2.200000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
  END
END sky130_fd_sc_hs__o21ai_1
MACRO sky130_fd_sc_hs__o21ai_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.265000 1.350000 0.595000 1.950000 ;
        RECT 0.265000 1.950000 2.275000 2.120000 ;
        RECT 1.755000 1.350000 2.275000 1.950000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.845000 1.350000 1.515000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905000 1.180000 3.235000 1.550000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.961100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 2.290000 2.795000 2.460000 ;
        RECT 1.065000 2.460000 1.395000 2.735000 ;
        RECT 2.475000 0.715000 2.735000 1.130000 ;
        RECT 2.525000 1.130000 2.735000 1.820000 ;
        RECT 2.525000 1.820000 2.795000 2.290000 ;
        RECT 2.525000 2.460000 2.795000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.115000  0.350000 0.445000 1.010000 ;
      RECT 0.115000  1.010000 2.305000 1.180000 ;
      RECT 0.115000  2.290000 0.365000 3.245000 ;
      RECT 0.565000  2.290000 0.895000 2.905000 ;
      RECT 0.565000  2.905000 1.895000 3.075000 ;
      RECT 0.615000  0.085000 0.945000 0.830000 ;
      RECT 1.125000  0.350000 1.375000 1.010000 ;
      RECT 1.545000  0.085000 1.875000 0.830000 ;
      RECT 1.565000  2.630000 1.895000 2.905000 ;
      RECT 2.055000  0.350000 3.245000 0.520000 ;
      RECT 2.055000  0.520000 2.305000 1.010000 ;
      RECT 2.095000  2.630000 2.345000 3.245000 ;
      RECT 2.915000  0.520000 3.245000 1.010000 ;
      RECT 2.995000  1.820000 3.245000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__o21ai_2
MACRO sky130_fd_sc_hs__o21ai_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.445000 1.320000 1.795000 1.650000 ;
        RECT 1.085000 1.650000 1.795000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.350000 5.635000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.180000 3.165000 1.550000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.478400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.280000 0.595000 2.530000 0.840000 ;
        RECT 2.280000 0.840000 3.505000 1.010000 ;
        RECT 2.365000 1.820000 3.715000 1.950000 ;
        RECT 2.365000 1.950000 5.190000 2.120000 ;
        RECT 3.220000 0.595000 3.505000 0.840000 ;
        RECT 3.335000 1.010000 3.505000 1.550000 ;
        RECT 3.335000 1.550000 3.715000 1.820000 ;
        RECT 3.960000 2.120000 4.290000 2.735000 ;
        RECT 4.860000 2.120000 5.190000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.115000  0.350000 0.365000 0.980000 ;
      RECT 0.115000  0.980000 2.100000 1.010000 ;
      RECT 0.115000  1.010000 1.225000 1.150000 ;
      RECT 0.115000  1.820000 0.365000 3.245000 ;
      RECT 0.545000  0.085000 0.875000 0.810000 ;
      RECT 0.565000  1.820000 0.895000 1.950000 ;
      RECT 0.565000  1.950000 1.795000 2.120000 ;
      RECT 0.565000  2.120000 0.895000 2.980000 ;
      RECT 1.055000  0.350000 1.225000 0.840000 ;
      RECT 1.055000  0.840000 2.100000 0.980000 ;
      RECT 1.095000  2.290000 1.265000 3.245000 ;
      RECT 1.405000  0.085000 1.735000 0.670000 ;
      RECT 1.465000  2.120000 1.795000 2.290000 ;
      RECT 1.465000  2.290000 3.790000 2.460000 ;
      RECT 1.465000  2.460000 1.795000 2.980000 ;
      RECT 1.930000  0.255000 3.845000 0.425000 ;
      RECT 1.930000  0.425000 2.100000 0.840000 ;
      RECT 1.995000  2.630000 2.245000 3.245000 ;
      RECT 2.710000  0.425000 3.040000 0.670000 ;
      RECT 2.900000  2.630000 3.230000 3.245000 ;
      RECT 3.460000  2.460000 3.790000 2.905000 ;
      RECT 3.460000  2.905000 5.640000 3.075000 ;
      RECT 3.675000  0.425000 3.845000 1.010000 ;
      RECT 3.675000  1.010000 5.645000 1.180000 ;
      RECT 4.025000  0.085000 4.355000 0.840000 ;
      RECT 4.490000  2.290000 4.660000 2.905000 ;
      RECT 4.535000  0.350000 4.705000 1.010000 ;
      RECT 4.885000  0.085000 5.215000 0.840000 ;
      RECT 5.390000  1.950000 5.640000 2.905000 ;
      RECT 5.395000  0.350000 5.645000 1.010000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_hs__o21ai_4
MACRO sky130_fd_sc_hs__o21ba_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.130000 0.550000 1.800000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.835000 1.130000 1.315000 1.800000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.515000 1.180000 2.845000 1.550000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.390000 0.350000 3.755000 1.130000 ;
        RECT 3.395000 1.820000 3.755000 2.980000 ;
        RECT 3.585000 1.130000 3.755000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.115000  0.350000 0.445000 0.790000 ;
      RECT 0.115000  0.790000 1.445000 0.960000 ;
      RECT 0.115000  1.970000 0.445000 3.245000 ;
      RECT 0.615000  0.085000 0.945000 0.620000 ;
      RECT 1.055000  1.970000 1.785000 2.320000 ;
      RECT 1.055000  2.320000 3.225000 2.490000 ;
      RECT 1.055000  2.490000 1.385000 2.980000 ;
      RECT 1.115000  0.350000 1.445000 0.790000 ;
      RECT 1.555000  2.660000 1.885000 3.245000 ;
      RECT 1.615000  0.350000 1.945000 1.030000 ;
      RECT 1.615000  1.030000 1.785000 1.970000 ;
      RECT 1.975000  1.220000 2.305000 1.820000 ;
      RECT 1.975000  1.820000 2.690000 2.150000 ;
      RECT 2.135000  0.680000 2.720000 1.010000 ;
      RECT 2.135000  1.010000 2.305000 1.220000 ;
      RECT 2.890000  0.085000 3.220000 1.010000 ;
      RECT 2.895000  2.660000 3.225000 3.245000 ;
      RECT 3.055000  1.320000 3.415000 1.650000 ;
      RECT 3.055000  1.650000 3.225000 2.320000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__o21ba_1
MACRO sky130_fd_sc_hs__o21ba_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405000 1.180000 3.735000 1.550000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.720000 1.180000 3.235000 1.550000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.455000 1.780000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.010000 0.350000 1.340000 1.130000 ;
        RECT 1.010000 1.130000 1.180000 1.820000 ;
        RECT 1.010000 1.820000 1.440000 2.070000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.105000  0.455000 0.355000 0.960000 ;
      RECT 0.105000  0.960000 0.795000 1.130000 ;
      RECT 0.115000  1.950000 0.795000 2.240000 ;
      RECT 0.115000  2.240000 2.210000 2.410000 ;
      RECT 0.115000  2.410000 0.445000 2.700000 ;
      RECT 0.535000  0.085000 0.785000 0.790000 ;
      RECT 0.625000  1.130000 0.795000 1.950000 ;
      RECT 0.650000  2.580000 0.980000 3.245000 ;
      RECT 1.350000  1.300000 1.680000 1.630000 ;
      RECT 1.510000  1.010000 2.550000 1.180000 ;
      RECT 1.510000  1.180000 1.680000 1.300000 ;
      RECT 1.520000  0.085000 1.770000 0.820000 ;
      RECT 1.565000  2.580000 2.235000 3.245000 ;
      RECT 1.890000  1.350000 2.210000 2.240000 ;
      RECT 1.980000  0.350000 2.230000 1.010000 ;
      RECT 2.380000  1.180000 2.550000 1.820000 ;
      RECT 2.380000  1.820000 2.775000 2.410000 ;
      RECT 2.410000  0.350000 2.740000 0.670000 ;
      RECT 2.410000  0.670000 3.740000 0.840000 ;
      RECT 2.445000  2.410000 2.775000 2.860000 ;
      RECT 2.910000  0.085000 3.240000 0.500000 ;
      RECT 3.405000  1.820000 3.735000 3.245000 ;
      RECT 3.410000  0.350000 3.740000 0.670000 ;
      RECT 3.410000  0.840000 3.740000 1.010000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__o21ba_2
MACRO sky130_fd_sc_hs__o21ba_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.175000 1.450000 4.675000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.845000 1.450000 6.115000 1.780000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.180000 0.835000 1.550000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  1.093800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.550000 1.315000 1.820000 ;
        RECT 1.085000 1.820000 2.345000 2.220000 ;
        RECT 1.145000 0.350000 1.340000 0.950000 ;
        RECT 1.145000 0.950000 2.210000 1.120000 ;
        RECT 1.145000 1.120000 1.315000 1.550000 ;
        RECT 1.960000 0.350000 2.210000 0.950000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.240000 0.085000 ;
      RECT 0.000000  3.245000 6.240000 3.415000 ;
      RECT 0.085000  0.350000 0.475000 1.010000 ;
      RECT 0.085000  1.010000 0.255000 1.820000 ;
      RECT 0.085000  1.820000 0.445000 2.390000 ;
      RECT 0.085000  2.390000 3.320000 2.560000 ;
      RECT 0.085000  2.560000 0.445000 2.980000 ;
      RECT 0.615000  2.730000 0.995000 3.245000 ;
      RECT 0.645000  0.085000 0.975000 1.010000 ;
      RECT 1.485000  1.290000 3.830000 1.460000 ;
      RECT 1.485000  1.460000 2.980000 1.620000 ;
      RECT 1.530000  0.085000 1.780000 0.780000 ;
      RECT 1.565000  2.730000 1.895000 3.245000 ;
      RECT 2.390000  0.085000 2.640000 1.120000 ;
      RECT 2.465000  2.730000 3.205000 3.245000 ;
      RECT 2.810000  0.255000 3.830000 0.425000 ;
      RECT 2.810000  0.425000 2.980000 1.290000 ;
      RECT 3.150000  0.595000 3.320000 0.950000 ;
      RECT 3.150000  0.950000 4.330000 1.110000 ;
      RECT 3.150000  1.110000 6.125000 1.120000 ;
      RECT 3.150000  1.630000 3.490000 1.960000 ;
      RECT 3.150000  1.960000 3.320000 2.390000 ;
      RECT 3.490000  2.130000 5.145000 2.300000 ;
      RECT 3.490000  2.300000 3.740000 2.980000 ;
      RECT 3.500000  0.425000 3.830000 0.780000 ;
      RECT 3.660000  1.460000 3.830000 1.950000 ;
      RECT 3.660000  1.950000 5.145000 2.130000 ;
      RECT 3.945000  2.470000 4.275000 3.245000 ;
      RECT 4.000000  0.605000 4.330000 0.950000 ;
      RECT 4.000000  1.120000 6.125000 1.280000 ;
      RECT 4.445000  2.470000 4.775000 2.905000 ;
      RECT 4.445000  2.905000 5.675000 3.075000 ;
      RECT 4.500000  0.085000 4.750000 0.940000 ;
      RECT 4.930000  0.605000 5.180000 1.110000 ;
      RECT 4.975000  2.300000 5.145000 2.735000 ;
      RECT 5.345000  1.950000 5.675000 2.905000 ;
      RECT 5.360000  0.085000 5.610000 0.940000 ;
      RECT 5.790000  0.605000 6.125000 1.110000 ;
      RECT 5.875000  1.950000 6.125000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
  END
END sky130_fd_sc_hs__o21ba_4
MACRO sky130_fd_sc_hs__o21bai_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.880000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 1.300000 2.775000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.750000 1.300000 2.275000 1.630000 ;
        RECT 2.045000 1.630000 2.275000 2.890000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.450000 0.565000 1.780000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 0.350000 1.475000 1.130000 ;
        RECT 1.305000 1.130000 1.475000 1.820000 ;
        RECT 1.305000 1.820000 1.840000 1.990000 ;
        RECT 1.475000 1.990000 1.840000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.880000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.880000 0.085000 ;
      RECT 0.000000  3.245000 2.880000 3.415000 ;
      RECT 0.110000  0.350000 0.360000 1.110000 ;
      RECT 0.110000  1.110000 0.915000 1.280000 ;
      RECT 0.135000  1.950000 0.915000 2.120000 ;
      RECT 0.135000  2.120000 0.465000 2.980000 ;
      RECT 0.540000  0.085000 0.870000 0.940000 ;
      RECT 0.635000  2.290000 1.305000 3.245000 ;
      RECT 0.745000  1.280000 0.915000 1.300000 ;
      RECT 0.745000  1.300000 1.135000 1.630000 ;
      RECT 0.745000  1.630000 0.915000 1.950000 ;
      RECT 1.645000  0.350000 1.815000 0.960000 ;
      RECT 1.645000  0.960000 2.765000 1.130000 ;
      RECT 1.995000  0.085000 2.335000 0.680000 ;
      RECT 2.515000  0.350000 2.765000 0.960000 ;
      RECT 2.520000  1.950000 2.770000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
  END
END sky130_fd_sc_hs__o21bai_1
MACRO sky130_fd_sc_hs__o21bai_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.250000 1.350000 2.580000 1.950000 ;
        RECT 2.250000 1.950000 3.715000 2.120000 ;
        RECT 3.485000 1.320000 4.055000 1.650000 ;
        RECT 3.485000 1.650000 3.715000 1.950000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.820000 1.350000 3.235000 1.780000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.460000 1.350000 0.835000 1.780000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.879200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.530000 1.180000 1.865000 2.290000 ;
        RECT 1.530000 2.290000 3.220000 2.460000 ;
        RECT 1.530000 2.460000 1.780000 2.980000 ;
        RECT 1.615000 0.615000 1.865000 1.180000 ;
        RECT 3.050000 2.460000 3.220000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  0.350000 0.365000 1.010000 ;
      RECT 0.115000  1.010000 1.360000 1.180000 ;
      RECT 0.115000  1.180000 0.285000 1.950000 ;
      RECT 0.115000  1.950000 0.640000 2.860000 ;
      RECT 0.545000  0.085000 0.875000 0.840000 ;
      RECT 1.005000  1.820000 1.335000 3.245000 ;
      RECT 1.030000  1.180000 1.360000 1.550000 ;
      RECT 1.105000  0.255000 2.365000 0.425000 ;
      RECT 1.105000  0.425000 1.435000 0.840000 ;
      RECT 1.980000  2.650000 2.350000 3.245000 ;
      RECT 2.035000  0.425000 2.365000 1.010000 ;
      RECT 2.035000  1.010000 4.185000 1.150000 ;
      RECT 2.035000  1.150000 3.245000 1.180000 ;
      RECT 2.520000  2.630000 2.850000 2.905000 ;
      RECT 2.520000  2.905000 3.755000 3.075000 ;
      RECT 2.535000  0.085000 2.865000 0.840000 ;
      RECT 3.075000  0.350000 3.245000 0.980000 ;
      RECT 3.075000  0.980000 4.185000 1.010000 ;
      RECT 3.420000  2.290000 3.755000 2.905000 ;
      RECT 3.425000  0.085000 3.755000 0.810000 ;
      RECT 3.935000  0.350000 4.185000 0.980000 ;
      RECT 3.955000  1.820000 4.205000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__o21bai_2
MACRO sky130_fd_sc_hs__o21bai_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.795000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.350000 3.715000 1.780000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.363000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365000 1.450000 7.075000 1.780000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  1.855000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.370000 1.950000 5.625000 2.020000 ;
        RECT 2.370000 2.020000 4.710000 2.120000 ;
        RECT 2.370000 2.120000 2.620000 2.735000 ;
        RECT 3.320000 2.120000 3.650000 2.735000 ;
        RECT 3.965000 1.010000 5.595000 1.180000 ;
        RECT 3.965000 1.180000 4.195000 1.950000 ;
        RECT 4.265000 0.595000 4.595000 1.010000 ;
        RECT 4.380000 1.850000 5.625000 1.950000 ;
        RECT 4.380000 2.120000 4.710000 2.980000 ;
        RECT 5.265000 0.595000 5.595000 1.010000 ;
        RECT 5.295000 2.020000 5.625000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.200000 0.085000 ;
      RECT 0.000000  3.245000 7.200000 3.415000 ;
      RECT 0.115000  0.350000 0.365000 1.010000 ;
      RECT 0.115000  1.010000 3.075000 1.180000 ;
      RECT 0.120000  1.950000 2.170000 2.120000 ;
      RECT 0.120000  2.120000 0.370000 2.980000 ;
      RECT 0.545000  0.085000 0.875000 0.840000 ;
      RECT 0.570000  2.290000 0.820000 3.245000 ;
      RECT 1.020000  2.120000 1.270000 2.980000 ;
      RECT 1.105000  0.350000 1.275000 1.010000 ;
      RECT 1.455000  0.085000 1.785000 0.840000 ;
      RECT 1.470000  2.290000 1.800000 3.245000 ;
      RECT 1.965000  0.350000 2.135000 1.010000 ;
      RECT 2.000000  1.820000 2.170000 1.950000 ;
      RECT 2.000000  2.120000 2.170000 2.905000 ;
      RECT 2.000000  2.905000 4.150000 3.075000 ;
      RECT 2.315000  0.085000 2.645000 0.840000 ;
      RECT 2.820000  2.290000 3.150000 2.905000 ;
      RECT 2.825000  0.350000 3.075000 0.670000 ;
      RECT 2.825000  0.670000 4.095000 0.840000 ;
      RECT 2.825000  0.840000 3.075000 1.010000 ;
      RECT 3.255000  0.085000 3.585000 0.500000 ;
      RECT 3.765000  0.255000 6.095000 0.425000 ;
      RECT 3.765000  0.425000 4.095000 0.670000 ;
      RECT 3.820000  2.290000 4.150000 2.905000 ;
      RECT 4.370000  1.350000 5.965000 1.680000 ;
      RECT 4.765000  0.425000 5.095000 0.840000 ;
      RECT 4.910000  2.190000 5.080000 3.245000 ;
      RECT 5.765000  0.425000 6.095000 0.940000 ;
      RECT 5.795000  1.110000 6.575000 1.280000 ;
      RECT 5.795000  1.280000 5.965000 1.350000 ;
      RECT 5.795000  1.680000 5.965000 1.950000 ;
      RECT 5.795000  1.950000 6.555000 2.120000 ;
      RECT 5.855000  2.290000 6.105000 3.245000 ;
      RECT 6.305000  2.120000 6.555000 2.980000 ;
      RECT 6.325000  0.500000 6.575000 1.110000 ;
      RECT 6.755000  0.085000 7.085000 1.280000 ;
      RECT 6.755000  2.100000 7.085000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
  END
END sky130_fd_sc_hs__o21bai_4
MACRO sky130_fd_sc_hs__o221a_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.450000 1.335000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.450000 1.905000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925000 1.460000 3.255000 1.790000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.145000 1.450000 2.755000 1.780000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.120000 3.825000 1.790000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.350000 0.520000 1.130000 ;
        RECT 0.115000 1.130000 0.285000 1.820000 ;
        RECT 0.115000 1.820000 0.445000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.455000  1.320000 0.785000 1.650000 ;
      RECT 0.615000  1.650000 0.785000 1.950000 ;
      RECT 0.615000  1.950000 2.055000 1.960000 ;
      RECT 0.615000  1.960000 4.205000 2.120000 ;
      RECT 0.680000  2.290000 1.060000 3.245000 ;
      RECT 0.690000  0.085000 1.020000 1.130000 ;
      RECT 1.200000  0.450000 1.530000 1.110000 ;
      RECT 1.200000  1.110000 3.100000 1.280000 ;
      RECT 1.700000  0.085000 2.030000 0.940000 ;
      RECT 1.725000  2.120000 4.205000 2.130000 ;
      RECT 1.725000  2.130000 2.055000 2.980000 ;
      RECT 2.260000  0.255000 3.600000 0.425000 ;
      RECT 2.260000  0.425000 2.590000 0.940000 ;
      RECT 2.770000  0.595000 3.100000 1.110000 ;
      RECT 2.865000  2.300000 3.705000 3.245000 ;
      RECT 3.270000  0.425000 3.600000 0.950000 ;
      RECT 3.770000  0.360000 4.205000 0.950000 ;
      RECT 3.875000  2.130000 4.205000 2.980000 ;
      RECT 4.035000  0.950000 4.205000 1.960000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__o221a_1
MACRO sky130_fd_sc_hs__o221a_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.350000 3.385000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.485000 1.350000 2.815000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 1.350000 1.395000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.350000 2.275000 1.780000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.435000 1.550000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.790000 0.350000 4.265000 1.130000 ;
        RECT 3.905000 1.820000 4.265000 2.980000 ;
        RECT 4.095000 1.130000 4.265000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.115000  1.820000 0.775000 1.950000 ;
      RECT 0.115000  1.950000 3.735000 2.120000 ;
      RECT 0.115000  2.120000 0.445000 2.860000 ;
      RECT 0.370000  0.350000 0.775000 1.010000 ;
      RECT 0.605000  1.010000 0.775000 1.820000 ;
      RECT 0.615000  2.290000 1.525000 3.245000 ;
      RECT 0.945000  0.350000 2.130000 0.520000 ;
      RECT 0.945000  0.520000 1.115000 1.130000 ;
      RECT 1.295000  0.800000 1.620000 1.010000 ;
      RECT 1.295000  1.010000 3.120000 1.180000 ;
      RECT 1.800000  0.520000 2.130000 0.830000 ;
      RECT 2.065000  2.120000 2.395000 2.860000 ;
      RECT 2.360000  0.085000 2.690000 0.830000 ;
      RECT 2.870000  0.350000 3.120000 1.010000 ;
      RECT 3.290000  0.085000 3.620000 1.130000 ;
      RECT 3.405000  2.290000 3.735000 3.245000 ;
      RECT 3.565000  1.320000 3.925000 1.650000 ;
      RECT 3.565000  1.650000 3.735000 1.950000 ;
      RECT 4.435000  0.085000 4.685000 1.130000 ;
      RECT 4.435000  1.820000 4.685000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_hs__o221a_2
MACRO sky130_fd_sc_hs__o221a_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925000 1.350000 5.320000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.365000 1.445000 4.695000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.445000 4.195000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.445000 2.755000 1.780000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.445000 0.890000 1.780000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  1.235700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.735000 0.475000 5.985000 1.010000 ;
        RECT 5.735000 1.010000 7.065000 1.180000 ;
        RECT 5.830000 1.850000 7.115000 2.020000 ;
        RECT 5.830000 2.020000 6.160000 2.980000 ;
        RECT 6.735000 0.475000 7.065000 1.010000 ;
        RECT 6.785000 1.180000 7.065000 1.550000 ;
        RECT 6.785000 1.550000 7.555000 1.780000 ;
        RECT 6.785000 1.780000 7.115000 1.850000 ;
        RECT 6.785000 2.020000 7.115000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.680000 0.085000 ;
      RECT 0.000000  3.245000 7.680000 3.415000 ;
      RECT 0.115000  0.265000 2.305000 0.285000 ;
      RECT 0.115000  0.285000 3.170000 0.435000 ;
      RECT 0.115000  0.435000 0.365000 1.275000 ;
      RECT 0.115000  1.950000 0.365000 3.245000 ;
      RECT 0.545000  0.605000 0.795000 1.105000 ;
      RECT 0.545000  1.105000 1.230000 1.275000 ;
      RECT 0.565000  1.950000 5.660000 2.120000 ;
      RECT 0.565000  2.120000 0.895000 2.955000 ;
      RECT 0.975000  0.435000 1.305000 0.935000 ;
      RECT 1.060000  1.275000 1.230000 1.950000 ;
      RECT 1.095000  2.290000 1.345000 3.245000 ;
      RECT 1.475000  0.605000 1.805000 1.025000 ;
      RECT 1.475000  1.025000 2.740000 1.105000 ;
      RECT 1.475000  1.105000 5.055000 1.180000 ;
      RECT 1.475000  1.180000 4.115000 1.275000 ;
      RECT 1.475000  1.275000 1.805000 1.285000 ;
      RECT 1.515000  2.290000 1.845000 2.905000 ;
      RECT 1.515000  2.905000 2.745000 3.075000 ;
      RECT 1.975000  0.435000 3.170000 0.455000 ;
      RECT 1.975000  0.455000 2.305000 0.855000 ;
      RECT 2.045000  2.120000 2.215000 2.735000 ;
      RECT 2.415000  2.290000 2.745000 2.905000 ;
      RECT 2.475000  0.635000 2.670000 1.025000 ;
      RECT 2.840000  0.455000 3.170000 0.855000 ;
      RECT 2.915000  2.290000 3.630000 3.245000 ;
      RECT 3.430000  0.085000 3.760000 0.935000 ;
      RECT 3.800000  2.290000 4.130000 2.905000 ;
      RECT 3.800000  2.905000 5.130000 3.075000 ;
      RECT 3.940000  0.585000 4.115000 1.010000 ;
      RECT 3.940000  1.010000 5.055000 1.105000 ;
      RECT 4.295000  0.085000 4.625000 0.840000 ;
      RECT 4.300000  2.120000 4.630000 2.735000 ;
      RECT 4.800000  2.290000 5.130000 2.905000 ;
      RECT 4.805000  0.590000 5.055000 1.010000 ;
      RECT 5.235000  0.085000 5.565000 1.180000 ;
      RECT 5.300000  2.290000 5.630000 3.245000 ;
      RECT 5.490000  1.350000 6.615000 1.680000 ;
      RECT 5.490000  1.680000 5.660000 1.950000 ;
      RECT 6.165000  0.085000 6.565000 0.805000 ;
      RECT 6.360000  2.190000 6.610000 3.245000 ;
      RECT 7.235000  0.085000 7.565000 1.255000 ;
      RECT 7.315000  1.950000 7.565000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
  END
END sky130_fd_sc_hs__o221a_4
MACRO sky130_fd_sc_hs__o221ai_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.300000 3.715000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 1.350000 2.775000 1.680000 ;
        RECT 2.525000 1.680000 2.775000 2.890000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965000 1.350000 1.635000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.875000 1.350000 2.275000 1.780000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.300000 0.435000 1.780000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.011700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.350000 0.445000 0.960000 ;
        RECT 0.115000 0.960000 0.775000 1.130000 ;
        RECT 0.325000 1.950000 2.355000 2.120000 ;
        RECT 0.325000 2.120000 0.575000 2.980000 ;
        RECT 0.605000 1.130000 0.775000 1.950000 ;
        RECT 2.025000 2.120000 2.355000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.615000  0.350000 2.005000 0.520000 ;
      RECT 0.615000  0.520000 0.945000 0.770000 ;
      RECT 0.745000  2.290000 1.560000 3.245000 ;
      RECT 1.175000  0.800000 1.505000 1.010000 ;
      RECT 1.175000  1.010000 3.725000 1.130000 ;
      RECT 1.175000  1.130000 2.505000 1.180000 ;
      RECT 1.675000  0.520000 2.005000 0.795000 ;
      RECT 2.175000  0.350000 2.505000 0.960000 ;
      RECT 2.175000  0.960000 3.725000 1.010000 ;
      RECT 2.675000  0.085000 3.225000 0.790000 ;
      RECT 3.165000  1.950000 3.495000 3.245000 ;
      RECT 3.395000  0.350000 3.725000 0.960000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__o221ai_1
MACRO sky130_fd_sc_hs__o221ai_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.645000 1.350000 3.975000 1.950000 ;
        RECT 3.645000 1.950000 5.635000 2.120000 ;
        RECT 4.925000 1.350000 5.635000 1.950000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.345000 1.350000 4.675000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.350000 2.275000 1.950000 ;
        RECT 1.085000 1.950000 3.405000 2.120000 ;
        RECT 3.075000 1.350000 3.405000 1.950000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.520000 1.350000 2.850000 1.780000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.300000 0.435000 1.780000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.232000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.595000 0.875000 2.290000 ;
        RECT 0.605000 2.290000 4.615000 2.460000 ;
        RECT 0.605000 2.460000 0.855000 2.980000 ;
        RECT 2.365000 2.460000 2.695000 2.735000 ;
        RECT 4.365000 2.460000 4.615000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.115000  0.255000 1.305000 0.425000 ;
      RECT 0.115000  0.425000 0.365000 1.130000 ;
      RECT 0.155000  1.950000 0.405000 3.245000 ;
      RECT 1.055000  0.425000 1.305000 1.010000 ;
      RECT 1.055000  1.010000 3.280000 1.180000 ;
      RECT 1.055000  2.630000 1.695000 3.245000 ;
      RECT 1.535000  0.255000 3.710000 0.425000 ;
      RECT 1.535000  0.425000 1.865000 0.820000 ;
      RECT 1.865000  2.630000 2.195000 2.905000 ;
      RECT 1.865000  2.905000 3.195000 3.075000 ;
      RECT 2.045000  0.595000 2.215000 1.010000 ;
      RECT 2.395000  0.425000 2.725000 0.820000 ;
      RECT 2.865000  2.630000 3.195000 2.905000 ;
      RECT 2.895000  0.595000 3.280000 1.010000 ;
      RECT 3.365000  2.630000 3.695000 3.245000 ;
      RECT 3.460000  0.425000 3.710000 1.010000 ;
      RECT 3.460000  1.010000 5.645000 1.180000 ;
      RECT 3.865000  2.630000 4.195000 2.905000 ;
      RECT 3.865000  2.905000 5.145000 3.075000 ;
      RECT 3.880000  0.085000 4.210000 0.820000 ;
      RECT 4.380000  0.405000 4.710000 1.010000 ;
      RECT 4.815000  2.290000 5.145000 2.905000 ;
      RECT 4.880000  0.085000 5.210000 0.820000 ;
      RECT 5.315000  2.290000 5.645000 3.245000 ;
      RECT 5.390000  0.405000 5.645000 1.010000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_hs__o221ai_2
MACRO sky130_fd_sc_hs__o221ai_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.210000 1.260000 6.575000 1.590000 ;
        RECT 6.405000 1.090000 8.455000 1.260000 ;
        RECT 8.285000 1.260000 9.955000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.845000 1.430000 8.035000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.545000 1.350000 3.555000 1.710000 ;
        RECT 2.545000 1.710000 6.000000 1.880000 ;
        RECT 5.405000 1.350000 6.000000 1.710000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.185000 1.180000 5.195000 1.540000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.405000 1.780000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  2.514400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.595000 0.875000 1.010000 ;
        RECT 0.545000 1.010000 1.745000 1.180000 ;
        RECT 0.565000 1.950000 1.825000 2.050000 ;
        RECT 0.565000 2.050000 8.160000 2.120000 ;
        RECT 0.565000 2.120000 0.895000 2.980000 ;
        RECT 1.405000 0.595000 1.745000 1.010000 ;
        RECT 1.575000 1.180000 1.745000 1.820000 ;
        RECT 1.575000 1.820000 1.825000 1.950000 ;
        RECT 1.575000 2.120000 7.260000 2.220000 ;
        RECT 1.575000 2.220000 1.825000 2.980000 ;
        RECT 4.055000 2.220000 4.225000 2.735000 ;
        RECT 4.925000 2.220000 5.255000 2.735000 ;
        RECT 6.845000 1.950000 8.160000 2.050000 ;
        RECT 6.845000 2.220000 7.260000 2.520000 ;
        RECT 6.930000 2.520000 7.260000 2.735000 ;
        RECT 7.830000 2.120000 8.160000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.115000  0.255000  2.165000 0.425000 ;
      RECT 0.115000  0.425000  0.375000 1.180000 ;
      RECT 0.115000  1.950000  0.365000 3.245000 ;
      RECT 1.045000  0.425000  1.235000 0.840000 ;
      RECT 1.065000  2.290000  1.395000 3.245000 ;
      RECT 1.915000  0.425000  2.165000 0.770000 ;
      RECT 1.915000  0.770000  3.155000 1.010000 ;
      RECT 1.915000  1.010000  4.015000 1.180000 ;
      RECT 2.025000  2.390000  2.355000 3.245000 ;
      RECT 2.395000  0.350000  6.235000 0.600000 ;
      RECT 2.525000  2.390000  3.855000 2.560000 ;
      RECT 2.525000  2.560000  2.855000 2.980000 ;
      RECT 3.025000  2.730000  3.355000 3.245000 ;
      RECT 3.335000  0.600000  3.505000 0.840000 ;
      RECT 3.525000  2.560000  3.855000 2.905000 ;
      RECT 3.525000  2.905000  5.755000 3.075000 ;
      RECT 3.685000  0.770000  5.735000 1.010000 ;
      RECT 4.425000  2.390000  4.755000 2.905000 ;
      RECT 5.405000  1.010000  5.735000 1.050000 ;
      RECT 5.425000  2.390000  5.755000 2.905000 ;
      RECT 5.905000  0.600000  6.235000 0.750000 ;
      RECT 5.905000  0.750000  9.025000 0.920000 ;
      RECT 5.905000  0.920000  6.235000 1.090000 ;
      RECT 5.925000  2.390000  6.255000 3.245000 ;
      RECT 6.405000  0.085000  6.735000 0.580000 ;
      RECT 6.425000  2.650000  6.675000 2.730000 ;
      RECT 6.425000  2.730000  6.760000 2.905000 ;
      RECT 6.425000  2.905000  8.530000 3.075000 ;
      RECT 6.905000  0.350000  7.155000 0.750000 ;
      RECT 7.335000  0.085000  7.665000 0.580000 ;
      RECT 7.460000  2.290000  7.630000 2.905000 ;
      RECT 7.835000  0.350000  8.085000 0.750000 ;
      RECT 8.265000  0.085000  8.605000 0.580000 ;
      RECT 8.360000  1.950000  9.510000 2.120000 ;
      RECT 8.360000  2.120000  8.530000 2.905000 ;
      RECT 8.730000  2.290000  8.980000 3.245000 ;
      RECT 8.775000  0.350000  9.025000 0.750000 ;
      RECT 8.775000  0.920000  9.965000 1.090000 ;
      RECT 9.180000  2.120000  9.510000 2.980000 ;
      RECT 9.205000  0.085000  9.535000 0.750000 ;
      RECT 9.710000  1.950000  9.960000 3.245000 ;
      RECT 9.715000  0.350000  9.965000 0.920000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
  END
END sky130_fd_sc_hs__o221ai_4
MACRO sky130_fd_sc_hs__o22a_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.235000 1.470000 3.715000 1.800000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.470000 2.995000 1.800000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.335000 1.470000 2.005000 1.800000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 0.255000 2.470000 0.585000 ;
        RECT 1.085000 0.585000 1.305000 0.670000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.350000 0.365000 1.130000 ;
        RECT 0.085000 1.130000 0.255000 1.820000 ;
        RECT 0.085000 1.820000 0.445000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.425000  1.300000 1.095000 1.630000 ;
      RECT 0.545000  0.085000 0.875000 0.960000 ;
      RECT 0.615000  1.985000 1.850000 3.245000 ;
      RECT 0.925000  1.130000 2.345000 1.300000 ;
      RECT 1.475000  0.755000 2.705000 0.935000 ;
      RECT 1.905000  1.105000 2.345000 1.130000 ;
      RECT 2.175000  1.300000 2.345000 1.970000 ;
      RECT 2.175000  1.970000 2.725000 2.140000 ;
      RECT 2.395000  2.140000 2.725000 2.980000 ;
      RECT 2.535000  0.935000 2.705000 1.130000 ;
      RECT 2.535000  1.130000 3.725000 1.300000 ;
      RECT 2.885000  0.085000 3.225000 0.960000 ;
      RECT 3.385000  1.970000 3.715000 3.245000 ;
      RECT 3.395000  0.630000 3.725000 1.130000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__o22a_1
MACRO sky130_fd_sc_hs__o22a_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405000 1.300000 3.735000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.710000 1.430000 3.235000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.545000 1.430000 1.875000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.430000 2.500000 1.780000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.350000 0.790000 0.820000 ;
        RECT 0.535000 0.820000 0.865000 1.130000 ;
        RECT 0.635000 1.130000 0.805000 1.820000 ;
        RECT 0.635000 1.820000 0.965000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.105000  0.085000 0.365000 1.130000 ;
      RECT 0.135000  1.820000 0.465000 3.245000 ;
      RECT 0.965000  0.085000 1.295000 0.640000 ;
      RECT 0.975000  1.300000 1.305000 1.630000 ;
      RECT 1.135000  0.880000 2.295000 1.130000 ;
      RECT 1.135000  1.130000 1.305000 1.300000 ;
      RECT 1.135000  1.630000 1.305000 1.950000 ;
      RECT 1.135000  1.950000 2.680000 2.120000 ;
      RECT 1.135000  2.290000 1.790000 3.245000 ;
      RECT 1.505000  0.350000 2.795000 0.520000 ;
      RECT 1.505000  0.520000 1.835000 0.710000 ;
      RECT 2.005000  0.800000 2.295000 0.880000 ;
      RECT 2.350000  2.120000 2.680000 2.940000 ;
      RECT 2.465000  0.520000 2.795000 0.960000 ;
      RECT 2.465000  0.960000 3.725000 1.130000 ;
      RECT 2.965000  0.085000 3.295000 0.790000 ;
      RECT 3.400000  1.950000 3.730000 3.245000 ;
      RECT 3.475000  0.350000 3.725000 0.960000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__o22a_2
MACRO sky130_fd_sc_hs__o22a_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.845000 1.450000 2.275000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.845000 1.450000 1.515000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 0.255000 2.610000 0.570000 ;
        RECT 2.045000 0.570000 2.275000 0.670000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.450000 3.505000 1.780000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  1.125600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.600000 1.850000 6.105000 2.020000 ;
        RECT 4.600000 2.020000 4.930000 2.980000 ;
        RECT 4.980000 0.350000 5.230000 1.010000 ;
        RECT 4.980000 1.010000 6.105000 1.180000 ;
        RECT 5.775000 2.020000 6.105000 2.980000 ;
        RECT 5.920000 0.350000 6.105000 1.010000 ;
        RECT 5.935000 1.180000 6.595000 1.410000 ;
        RECT 5.935000 1.410000 6.105000 1.850000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.720000 0.085000 ;
      RECT 0.000000  3.245000 6.720000 3.415000 ;
      RECT 0.115000  0.660000 0.445000 1.110000 ;
      RECT 0.115000  1.110000 4.240000 1.280000 ;
      RECT 0.115000  1.280000 0.445000 1.340000 ;
      RECT 0.115000  1.940000 0.365000 3.245000 ;
      RECT 0.565000  1.950000 0.895000 2.905000 ;
      RECT 0.565000  2.905000 1.895000 3.075000 ;
      RECT 0.615000  0.085000 0.945000 0.940000 ;
      RECT 1.065000  1.950000 3.845000 2.120000 ;
      RECT 1.065000  2.120000 1.395000 2.735000 ;
      RECT 1.125000  0.660000 1.375000 1.110000 ;
      RECT 1.545000  0.085000 1.875000 0.940000 ;
      RECT 1.565000  2.290000 1.895000 2.905000 ;
      RECT 2.045000  0.840000 2.375000 1.090000 ;
      RECT 2.045000  1.090000 4.240000 1.110000 ;
      RECT 2.065000  2.290000 2.395000 3.245000 ;
      RECT 2.545000  0.740000 3.810000 0.750000 ;
      RECT 2.545000  0.750000 4.585000 0.920000 ;
      RECT 2.565000  2.290000 2.895000 2.905000 ;
      RECT 2.565000  2.905000 3.895000 3.075000 ;
      RECT 3.065000  2.120000 3.395000 2.735000 ;
      RECT 3.480000  0.660000 3.810000 0.740000 ;
      RECT 3.565000  2.290000 3.895000 2.905000 ;
      RECT 3.675000  1.510000 5.765000 1.680000 ;
      RECT 3.675000  1.680000 3.845000 1.950000 ;
      RECT 3.910000  1.280000 4.240000 1.340000 ;
      RECT 4.100000  1.850000 4.430000 3.245000 ;
      RECT 4.415000  0.920000 4.585000 1.350000 ;
      RECT 4.415000  1.350000 5.765000 1.510000 ;
      RECT 4.470000  0.085000 4.800000 0.580000 ;
      RECT 5.200000  2.190000 5.530000 3.245000 ;
      RECT 5.410000  0.085000 5.740000 0.790000 ;
      RECT 6.275000  0.085000 6.605000 1.010000 ;
      RECT 6.275000  1.820000 6.605000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
  END
END sky130_fd_sc_hs__o22a_4
MACRO sky130_fd_sc_hs__o22ai_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.880000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.300000 2.775000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.535000 1.350000 1.865000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 1.180000 0.445000 1.550000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965000 1.350000 1.315000 1.780000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.895900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.615000 0.655000 1.065000 1.130000 ;
        RECT 0.625000 1.130000 0.795000 1.950000 ;
        RECT 0.625000 1.950000 1.550000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.880000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.880000 0.085000 ;
      RECT 0.000000  3.245000 2.880000 3.415000 ;
      RECT 0.115000  0.315000 1.670000 0.485000 ;
      RECT 0.115000  0.485000 0.445000 1.010000 ;
      RECT 0.125000  1.820000 0.455000 3.245000 ;
      RECT 1.340000  0.485000 1.670000 0.960000 ;
      RECT 1.340000  0.960000 2.670000 1.130000 ;
      RECT 1.840000  0.085000 2.170000 0.790000 ;
      RECT 2.255000  1.950000 2.585000 3.245000 ;
      RECT 2.340000  0.350000 2.670000 0.960000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
  END
END sky130_fd_sc_hs__o22ai_1
MACRO sky130_fd_sc_hs__o22ai_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.910000 1.350000 4.675000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.665000 1.300000 3.335000 1.390000 ;
        RECT 2.665000 1.390000 3.715000 1.630000 ;
        RECT 3.485000 1.630000 3.715000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.315000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 1.350000 1.815000 1.780000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.212200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.615000 0.595000 0.945000 1.010000 ;
        RECT 0.615000 1.010000 2.275000 1.180000 ;
        RECT 1.570000 1.950000 3.310000 1.970000 ;
        RECT 1.570000 1.970000 2.275000 2.120000 ;
        RECT 1.570000 2.120000 1.800000 2.735000 ;
        RECT 1.615000 0.595000 1.945000 1.010000 ;
        RECT 2.045000 1.180000 2.275000 1.800000 ;
        RECT 2.045000 1.800000 3.310000 1.950000 ;
        RECT 3.060000 1.970000 3.310000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.115000  0.255000 2.785000 0.425000 ;
      RECT 0.115000  0.425000 0.445000 1.130000 ;
      RECT 0.120000  1.950000 1.400000 2.120000 ;
      RECT 0.120000  2.120000 0.370000 2.980000 ;
      RECT 0.570000  2.290000 0.900000 3.245000 ;
      RECT 1.070000  2.120000 1.400000 2.905000 ;
      RECT 1.070000  2.905000 2.300000 3.075000 ;
      RECT 1.115000  0.425000 1.445000 0.840000 ;
      RECT 1.970000  2.290000 2.300000 2.905000 ;
      RECT 2.115000  0.425000 2.785000 0.840000 ;
      RECT 2.455000  0.840000 2.785000 0.960000 ;
      RECT 2.455000  0.960000 3.755000 1.010000 ;
      RECT 2.455000  1.010000 4.685000 1.130000 ;
      RECT 2.530000  2.140000 2.860000 2.905000 ;
      RECT 2.530000  2.905000 3.680000 3.075000 ;
      RECT 2.955000  0.085000 3.285000 0.790000 ;
      RECT 3.505000  0.350000 3.755000 0.960000 ;
      RECT 3.505000  1.130000 4.685000 1.180000 ;
      RECT 3.510000  1.950000 4.660000 2.120000 ;
      RECT 3.510000  2.120000 3.680000 2.905000 ;
      RECT 3.880000  2.290000 4.130000 3.245000 ;
      RECT 3.925000  0.085000 4.255000 0.840000 ;
      RECT 4.330000  2.120000 4.660000 2.980000 ;
      RECT 4.435000  0.350000 4.685000 1.010000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_hs__o22ai_2
MACRO sky130_fd_sc_hs__o22ai_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.540000 1.320000 1.550000 1.650000 ;
        RECT 1.380000 1.650000 1.550000 1.720000 ;
        RECT 1.380000 1.720000 3.810000 1.890000 ;
        RECT 2.525000 1.890000 3.235000 2.150000 ;
        RECT 3.640000 1.350000 3.970000 1.680000 ;
        RECT 3.640000 1.680000 3.810000 1.720000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.885000 1.180000 3.235000 1.550000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.290000 1.300000 5.635000 1.630000 ;
        RECT 5.405000 1.090000 7.730000 1.260000 ;
        RECT 5.405000 1.260000 5.635000 1.300000 ;
        RECT 7.400000 1.260000 7.730000 1.550000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.805000 1.430000 7.155000 1.680000 ;
        RECT 6.365000 1.680000 7.155000 1.780000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  2.388000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.020000 2.060000 2.350000 2.320000 ;
        RECT 2.020000 2.320000 4.150000 2.490000 ;
        RECT 3.980000 1.850000 6.100000 1.950000 ;
        RECT 3.980000 1.950000 8.070000 2.020000 ;
        RECT 3.980000 2.020000 4.150000 2.320000 ;
        RECT 4.405000 0.750000 8.070000 0.920000 ;
        RECT 4.405000 0.920000 5.155000 1.130000 ;
        RECT 5.770000 2.020000 8.070000 2.120000 ;
        RECT 5.770000 2.120000 6.100000 2.735000 ;
        RECT 6.205000 0.595000 6.535000 0.750000 ;
        RECT 6.670000 2.120000 7.000000 2.735000 ;
        RECT 7.205000 0.595000 7.535000 0.750000 ;
        RECT 7.900000 0.920000 8.070000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.115000  0.350000 0.445000 0.980000 ;
      RECT 0.115000  0.980000 4.235000 1.010000 ;
      RECT 0.115000  1.010000 1.375000 1.150000 ;
      RECT 0.120000  1.820000 0.370000 3.245000 ;
      RECT 0.570000  1.820000 0.900000 2.060000 ;
      RECT 0.570000  2.060000 1.850000 2.230000 ;
      RECT 0.570000  2.230000 0.850000 2.980000 ;
      RECT 0.615000  0.085000 0.945000 0.810000 ;
      RECT 1.020000  2.400000 1.350000 3.245000 ;
      RECT 1.125000  0.350000 1.375000 0.840000 ;
      RECT 1.125000  0.840000 4.235000 0.980000 ;
      RECT 1.520000  2.230000 1.850000 2.660000 ;
      RECT 1.520000  2.660000 3.700000 2.980000 ;
      RECT 1.545000  0.085000 1.875000 0.670000 ;
      RECT 2.055000  0.350000 2.305000 0.840000 ;
      RECT 2.475000  0.085000 2.805000 0.670000 ;
      RECT 2.985000  0.350000 3.235000 0.840000 ;
      RECT 3.405000  0.085000 3.735000 0.670000 ;
      RECT 3.870000  2.660000 4.200000 3.245000 ;
      RECT 3.905000  0.255000 8.045000 0.425000 ;
      RECT 3.905000  0.425000 6.035000 0.580000 ;
      RECT 3.905000  0.580000 4.235000 0.840000 ;
      RECT 3.905000  1.010000 4.235000 1.130000 ;
      RECT 4.370000  2.190000 5.570000 2.360000 ;
      RECT 4.370000  2.360000 4.700000 2.980000 ;
      RECT 4.900000  2.530000 5.150000 3.245000 ;
      RECT 5.320000  2.360000 5.570000 2.905000 ;
      RECT 5.320000  2.905000 7.500000 3.075000 ;
      RECT 6.300000  2.290000 6.470000 2.905000 ;
      RECT 6.705000  0.425000 7.035000 0.580000 ;
      RECT 7.170000  2.290000 7.500000 2.905000 ;
      RECT 7.670000  2.290000 8.000000 3.245000 ;
      RECT 7.715000  0.425000 8.045000 0.580000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_hs__o22ai_4
MACRO sky130_fd_sc_hs__o2bb2a_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965000 1.420000 1.315000 1.710000 ;
        RECT 1.085000 1.710000 1.315000 1.780000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505000 1.430000 1.835000 1.780000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.885000 1.180000 4.215000 1.510000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.180000 3.715000 1.510000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.350000 0.455000 1.130000 ;
        RECT 0.085000 1.130000 0.255000 1.820000 ;
        RECT 0.085000 1.820000 0.445000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.425000  1.300000 0.795000 1.630000 ;
      RECT 0.615000  1.950000 0.945000 3.245000 ;
      RECT 0.625000  0.085000 1.120000 0.910000 ;
      RECT 0.625000  1.080000 1.460000 1.250000 ;
      RECT 0.625000  1.250000 0.795000 1.300000 ;
      RECT 1.150000  1.950000 2.380000 2.280000 ;
      RECT 1.290000  0.255000 2.815000 0.425000 ;
      RECT 1.290000  0.425000 1.460000 1.080000 ;
      RECT 1.630000  0.595000 1.880000 1.090000 ;
      RECT 1.630000  1.090000 2.380000 1.260000 ;
      RECT 1.655000  2.450000 2.820000 3.245000 ;
      RECT 2.050000  1.260000 2.380000 1.950000 ;
      RECT 2.485000  0.425000 2.815000 0.920000 ;
      RECT 2.645000  0.920000 2.815000 1.900000 ;
      RECT 2.645000  1.900000 3.320000 2.070000 ;
      RECT 2.990000  2.070000 3.320000 2.780000 ;
      RECT 2.995000  0.340000 3.245000 0.840000 ;
      RECT 2.995000  0.840000 4.205000 1.010000 ;
      RECT 3.415000  0.085000 3.745000 0.670000 ;
      RECT 3.870000  1.900000 4.200000 3.245000 ;
      RECT 3.955000  0.340000 4.205000 0.840000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__o2bb2a_1
MACRO sky130_fd_sc_hs__o2bb2a_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.475000 2.865000 1.805000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.995000 1.475000 2.325000 1.805000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.450000 0.570000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.810000 1.450000 1.285000 1.780000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.425000 1.820000 3.770000 2.980000 ;
        RECT 3.430000 0.350000 3.770000 1.130000 ;
        RECT 3.600000 1.130000 3.770000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  0.350000 0.365000 1.110000 ;
      RECT 0.115000  1.110000 1.305000 1.280000 ;
      RECT 0.120000  1.950000 0.450000 3.245000 ;
      RECT 0.545000  0.085000 0.875000 0.940000 ;
      RECT 1.050000  1.950000 1.380000 2.395000 ;
      RECT 1.050000  2.395000 3.255000 2.565000 ;
      RECT 1.050000  2.565000 1.380000 2.980000 ;
      RECT 1.055000  0.350000 1.305000 1.110000 ;
      RECT 1.455000  1.450000 1.785000 1.780000 ;
      RECT 1.475000  0.255000 2.715000 0.425000 ;
      RECT 1.475000  0.425000 1.805000 0.965000 ;
      RECT 1.585000  2.735000 1.940000 3.245000 ;
      RECT 1.615000  1.135000 2.375000 1.305000 ;
      RECT 1.615000  1.305000 1.785000 1.450000 ;
      RECT 1.615000  1.780000 1.785000 1.975000 ;
      RECT 1.615000  1.975000 2.565000 2.225000 ;
      RECT 2.045000  0.595000 2.375000 1.135000 ;
      RECT 2.545000  0.425000 2.715000 1.135000 ;
      RECT 2.545000  1.135000 3.255000 1.305000 ;
      RECT 2.770000  2.735000 3.220000 3.245000 ;
      RECT 2.885000  0.085000 3.215000 0.965000 ;
      RECT 3.085000  1.305000 3.430000 1.635000 ;
      RECT 3.085000  1.635000 3.255000 2.395000 ;
      RECT 3.940000  0.085000 4.190000 1.130000 ;
      RECT 3.955000  1.820000 4.205000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__o2bb2a_2
MACRO sky130_fd_sc_hs__o2bb2a_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.415000 1.350000 4.745000 1.780000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.845000 1.350000 4.195000 1.780000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.260000 1.115000 1.770000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.470000 1.450000 2.275000 1.780000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  1.311300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.255000 0.350000 5.585000 0.810000 ;
        RECT 5.255000 0.810000 6.585000 1.050000 ;
        RECT 5.255000 1.720000 6.585000 1.890000 ;
        RECT 5.255000 1.890000 5.585000 2.980000 ;
        RECT 6.255000 0.350000 6.585000 0.810000 ;
        RECT 6.255000 1.050000 6.585000 1.720000 ;
        RECT 6.255000 1.890000 6.585000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.200000 0.085000 ;
      RECT 0.000000  3.245000 7.200000 3.415000 ;
      RECT 0.115000  0.350000 0.445000 0.920000 ;
      RECT 0.115000  0.920000 3.335000 1.090000 ;
      RECT 0.185000  1.940000 0.515000 1.950000 ;
      RECT 0.185000  1.950000 1.415000 2.120000 ;
      RECT 0.185000  2.120000 0.515000 2.980000 ;
      RECT 0.615000  0.085000 0.945000 0.750000 ;
      RECT 0.715000  2.290000 0.885000 3.245000 ;
      RECT 1.085000  2.120000 1.415000 2.905000 ;
      RECT 1.085000  2.905000 2.315000 3.075000 ;
      RECT 1.115000  0.350000 1.445000 0.780000 ;
      RECT 1.115000  0.780000 3.335000 0.920000 ;
      RECT 1.615000  0.085000 1.945000 0.610000 ;
      RECT 1.615000  1.950000 3.335000 2.120000 ;
      RECT 1.615000  2.120000 1.785000 2.735000 ;
      RECT 1.985000  2.290000 2.315000 2.905000 ;
      RECT 2.490000  1.300000 3.675000 1.630000 ;
      RECT 2.505000  0.255000 4.370000 0.425000 ;
      RECT 2.505000  0.425000 2.835000 0.610000 ;
      RECT 2.545000  2.320000 2.875000 3.245000 ;
      RECT 2.995000  1.820000 3.335000 1.950000 ;
      RECT 2.995000  2.120000 3.335000 2.150000 ;
      RECT 3.005000  0.595000 3.335000 0.780000 ;
      RECT 3.165000  2.150000 3.335000 2.450000 ;
      RECT 3.165000  2.450000 5.085000 2.620000 ;
      RECT 3.505000  0.960000 4.030000 1.130000 ;
      RECT 3.505000  1.130000 3.675000 1.300000 ;
      RECT 3.505000  1.630000 3.675000 1.950000 ;
      RECT 3.505000  1.950000 4.465000 2.280000 ;
      RECT 3.600000  2.790000 3.930000 3.245000 ;
      RECT 3.700000  0.635000 4.030000 0.960000 ;
      RECT 4.200000  0.425000 4.370000 0.950000 ;
      RECT 4.200000  0.950000 5.085000 1.120000 ;
      RECT 4.540000  0.085000 5.080000 0.780000 ;
      RECT 4.670000  2.790000 5.000000 3.245000 ;
      RECT 4.915000  1.120000 5.085000 1.220000 ;
      RECT 4.915000  1.220000 6.065000 1.550000 ;
      RECT 4.915000  1.550000 5.085000 2.450000 ;
      RECT 5.755000  0.085000 6.085000 0.640000 ;
      RECT 5.755000  2.060000 6.085000 3.245000 ;
      RECT 6.755000  0.085000 7.085000 1.130000 ;
      RECT 6.755000  1.820000 7.085000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
  END
END sky130_fd_sc_hs__o2bb2a_4
MACRO sky130_fd_sc_hs__o2bb2ai_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.435000 1.510000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.120000 1.100000 1.450000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925000 1.300000 3.255000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.225000 1.300000 2.755000 1.780000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.546900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.610000 0.350000 1.860000 1.010000 ;
        RECT 1.610000 1.010000 2.030000 1.180000 ;
        RECT 1.860000 1.180000 2.030000 1.950000 ;
        RECT 1.860000 1.950000 2.315000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 0.950000 ;
      RECT 0.140000  1.895000 0.470000 3.245000 ;
      RECT 0.640000  1.620000 1.690000 1.790000 ;
      RECT 0.640000  1.790000 0.970000 2.775000 ;
      RECT 0.935000  0.350000 1.440000 0.950000 ;
      RECT 1.140000  1.975000 1.690000 3.245000 ;
      RECT 1.270000  0.950000 1.440000 1.350000 ;
      RECT 1.270000  1.350000 1.690000 1.620000 ;
      RECT 2.030000  0.445000 2.370000 0.840000 ;
      RECT 2.200000  0.840000 2.370000 0.960000 ;
      RECT 2.200000  0.960000 3.220000 1.130000 ;
      RECT 2.540000  0.085000 2.710000 0.790000 ;
      RECT 2.890000  0.350000 3.220000 0.960000 ;
      RECT 2.995000  1.950000 3.245000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__o2bb2ai_1
MACRO sky130_fd_sc_hs__o2bb2ai_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  0.444000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.480000 1.630000 ;
        RECT 0.125000 1.630000 0.355000 2.415000 ;
        RECT 0.125000 2.415000 0.820000 2.450000 ;
        RECT 0.125000 2.450000 2.335000 2.585000 ;
        RECT 0.650000 2.585000 2.335000 2.620000 ;
        RECT 1.965000 1.350000 2.335000 1.680000 ;
        RECT 2.165000 1.680000 2.335000 2.450000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.444000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.375000 1.445000 1.795000 1.780000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.695000 1.350000 4.025000 1.720000 ;
        RECT 3.695000 1.720000 5.495000 1.780000 ;
        RECT 3.695000 1.780000 5.095000 1.890000 ;
        RECT 4.925000 1.350000 5.495000 1.720000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.345000 1.180000 4.675000 1.550000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.896000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.000000 0.595000 3.290000 1.130000 ;
        RECT 3.005000 1.130000 3.290000 2.060000 ;
        RECT 3.005000 2.060000 4.695000 2.230000 ;
        RECT 3.005000 2.230000 3.290000 2.980000 ;
        RECT 4.465000 2.230000 4.695000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.115000  2.755000 0.445000 3.245000 ;
      RECT 0.145000  0.085000 0.475000 1.030000 ;
      RECT 0.645000  0.255000 1.910000 0.425000 ;
      RECT 0.645000  0.425000 0.975000 0.935000 ;
      RECT 0.650000  1.105000 2.675000 1.180000 ;
      RECT 0.650000  1.180000 1.405000 1.275000 ;
      RECT 0.650000  1.275000 0.980000 1.950000 ;
      RECT 0.650000  1.950000 1.995000 2.245000 ;
      RECT 1.155000  0.605000 1.405000 1.010000 ;
      RECT 1.155000  1.010000 2.675000 1.105000 ;
      RECT 1.185000  2.790000 1.515000 3.245000 ;
      RECT 1.580000  0.425000 1.910000 0.825000 ;
      RECT 1.720000  2.245000 1.995000 2.280000 ;
      RECT 2.080000  0.085000 2.340000 0.825000 ;
      RECT 2.505000  1.180000 2.675000 1.300000 ;
      RECT 2.505000  1.300000 2.835000 1.630000 ;
      RECT 2.505000  1.820000 2.835000 3.245000 ;
      RECT 2.570000  0.255000 3.790000 0.425000 ;
      RECT 2.570000  0.425000 2.820000 0.825000 ;
      RECT 3.460000  0.425000 3.790000 0.840000 ;
      RECT 3.460000  0.840000 5.645000 1.010000 ;
      RECT 3.460000  1.010000 3.790000 1.130000 ;
      RECT 3.460000  2.400000 3.790000 3.245000 ;
      RECT 3.960000  0.085000 4.290000 0.670000 ;
      RECT 3.965000  2.400000 4.295000 2.905000 ;
      RECT 3.965000  2.905000 5.195000 3.075000 ;
      RECT 4.470000  0.350000 4.690000 0.770000 ;
      RECT 4.470000  0.770000 5.645000 0.840000 ;
      RECT 4.865000  2.060000 5.195000 2.905000 ;
      RECT 4.870000  0.085000 5.215000 0.600000 ;
      RECT 5.315000  1.010000 5.645000 1.130000 ;
      RECT 5.395000  0.350000 5.645000 0.770000 ;
      RECT 5.395000  1.950000 5.645000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_hs__o2bb2ai_2
MACRO sky130_fd_sc_hs__o2bb2ai_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.935000 1.780000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.225000 1.350000 3.235000 1.780000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.150000 1.350000 9.955000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885000 1.350000 7.640000 1.780000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.758400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.155000 1.800000 5.715000 1.950000 ;
        RECT 4.155000 1.950000 7.725000 1.970000 ;
        RECT 4.155000 1.970000 4.485000 2.980000 ;
        RECT 4.695000 0.595000 5.025000 0.960000 ;
        RECT 4.695000 0.960000 5.885000 1.130000 ;
        RECT 5.055000 1.970000 7.725000 2.120000 ;
        RECT 5.055000 2.120000 5.635000 2.150000 ;
        RECT 5.055000 2.150000 5.305000 2.980000 ;
        RECT 5.545000 0.595000 5.885000 0.960000 ;
        RECT 5.545000 1.130000 5.715000 1.800000 ;
        RECT 6.495000 2.120000 6.825000 2.735000 ;
        RECT 7.395000 2.120000 7.725000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.105000  1.950000  0.355000 3.245000 ;
      RECT 0.115000  0.350000  0.365000 1.010000 ;
      RECT 0.115000  1.010000  2.095000 1.180000 ;
      RECT 0.545000  0.085000  0.875000 0.840000 ;
      RECT 0.555000  1.950000  3.585000 2.120000 ;
      RECT 0.555000  2.120000  0.885000 2.980000 ;
      RECT 1.055000  0.350000  1.235000 1.010000 ;
      RECT 1.085000  2.290000  1.255000 3.245000 ;
      RECT 1.415000  0.085000  1.745000 0.840000 ;
      RECT 1.455000  2.120000  1.785000 2.980000 ;
      RECT 1.925000  0.255000  4.035000 0.425000 ;
      RECT 1.925000  0.425000  2.095000 1.010000 ;
      RECT 1.985000  2.290000  2.155000 3.245000 ;
      RECT 2.275000  0.595000  2.605000 1.010000 ;
      RECT 2.275000  1.010000  3.605000 1.180000 ;
      RECT 2.355000  2.120000  2.685000 2.980000 ;
      RECT 2.775000  0.425000  3.105000 0.840000 ;
      RECT 2.885000  2.290000  3.055000 3.245000 ;
      RECT 3.255000  2.120000  3.585000 2.980000 ;
      RECT 3.275000  0.595000  3.605000 1.010000 ;
      RECT 3.415000  1.180000  3.605000 1.300000 ;
      RECT 3.415000  1.300000  5.375000 1.630000 ;
      RECT 3.415000  1.630000  3.585000 1.950000 ;
      RECT 3.785000  0.425000  4.035000 1.130000 ;
      RECT 3.785000  1.820000  3.955000 3.245000 ;
      RECT 4.265000  0.255000  6.235000 0.425000 ;
      RECT 4.265000  0.425000  4.515000 1.130000 ;
      RECT 4.685000  2.140000  4.855000 3.245000 ;
      RECT 5.205000  0.425000  5.375000 0.790000 ;
      RECT 5.505000  2.320000  5.835000 3.245000 ;
      RECT 6.045000  2.290000  6.310000 2.905000 ;
      RECT 6.045000  2.905000  8.110000 3.075000 ;
      RECT 6.065000  0.425000  6.235000 1.010000 ;
      RECT 6.065000  1.010000  9.965000 1.180000 ;
      RECT 6.415000  0.085000  6.745000 0.830000 ;
      RECT 6.915000  0.350000  7.165000 1.010000 ;
      RECT 7.010000  2.290000  7.210000 2.905000 ;
      RECT 7.345000  0.085000  7.675000 0.830000 ;
      RECT 7.845000  0.350000  8.095000 1.010000 ;
      RECT 7.910000  1.950000  9.975000 2.120000 ;
      RECT 7.910000  2.120000  8.110000 2.905000 ;
      RECT 8.275000  0.085000  8.605000 0.830000 ;
      RECT 8.295000  2.290000  8.560000 3.245000 ;
      RECT 8.745000  2.120000  9.075000 2.980000 ;
      RECT 8.785000  0.350000  9.035000 1.010000 ;
      RECT 9.205000  0.085000  9.535000 0.830000 ;
      RECT 9.260000  2.290000  9.465000 3.245000 ;
      RECT 9.645000  2.120000  9.975000 2.980000 ;
      RECT 9.715000  0.350000  9.965000 1.010000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
  END
END sky130_fd_sc_hs__o2bb2ai_4
MACRO sky130_fd_sc_hs__o311a_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.015000 1.120000 3.385000 1.450000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455000 1.140000 1.805000 1.470000 ;
        RECT 1.635000 1.470000 1.805000 2.320000 ;
        RECT 1.635000 2.320000 2.845000 2.490000 ;
        RECT 2.515000 1.445000 2.845000 2.320000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975000 1.120000 2.305000 2.150000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.920000 1.140000 1.285000 1.470000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.140000 0.410000 1.470000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.855000 1.960000 4.235000 2.980000 ;
        RECT 3.870000 0.350000 4.235000 1.130000 ;
        RECT 4.065000 1.130000 4.235000 1.960000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.135000  1.640000 1.465000 1.810000 ;
      RECT 0.135000  1.810000 0.465000 2.955000 ;
      RECT 0.200000  0.350000 0.530000 0.800000 ;
      RECT 0.200000  0.800000 0.750000 0.970000 ;
      RECT 0.580000  0.970000 0.750000 1.640000 ;
      RECT 0.635000  1.980000 0.965000 3.245000 ;
      RECT 1.060000  0.280000 3.180000 0.610000 ;
      RECT 1.060000  0.610000 1.390000 0.970000 ;
      RECT 1.135000  1.810000 1.465000 2.785000 ;
      RECT 1.135000  2.785000 3.185000 2.955000 ;
      RECT 1.560000  0.780000 3.690000 0.950000 ;
      RECT 3.015000  1.620000 3.895000 1.790000 ;
      RECT 3.015000  1.790000 3.185000 2.785000 ;
      RECT 3.355000  1.960000 3.685000 3.245000 ;
      RECT 3.360000  0.085000 3.690000 0.780000 ;
      RECT 3.595000  1.350000 3.895000 1.620000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__o311a_1
MACRO sky130_fd_sc_hs__o311a_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.350000 2.925000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.025000 1.350000 2.355000 2.890000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 1.350000 1.815000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945000 1.350000 1.315000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.435000 1.550000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.330000 1.720000 4.195000 1.890000 ;
        RECT 3.330000 1.890000 3.660000 2.980000 ;
        RECT 3.435000 0.350000 3.685000 0.810000 ;
        RECT 3.435000 0.810000 4.195000 1.050000 ;
        RECT 3.965000 1.050000 4.195000 1.720000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.205000  0.350000 0.775000 1.010000 ;
      RECT 0.225000  1.820000 0.775000 1.950000 ;
      RECT 0.225000  1.950000 1.665000 2.120000 ;
      RECT 0.225000  2.120000 0.605000 2.860000 ;
      RECT 0.605000  1.010000 3.265000 1.180000 ;
      RECT 0.605000  1.180000 0.775000 1.820000 ;
      RECT 0.775000  2.290000 1.105000 3.245000 ;
      RECT 1.180000  0.350000 1.510000 0.670000 ;
      RECT 1.180000  0.670000 2.660000 0.840000 ;
      RECT 1.335000  2.120000 1.665000 2.980000 ;
      RECT 1.690000  0.085000 2.150000 0.500000 ;
      RECT 2.330000  0.350000 2.660000 0.670000 ;
      RECT 2.745000  1.950000 3.075000 3.245000 ;
      RECT 2.830000  0.085000 3.160000 0.840000 ;
      RECT 3.095000  1.180000 3.265000 1.220000 ;
      RECT 3.095000  1.220000 3.510000 1.550000 ;
      RECT 3.830000  2.060000 4.160000 3.245000 ;
      RECT 3.855000  0.085000 4.205000 0.600000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__o311a_2
MACRO sky130_fd_sc_hs__o311a_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.105000 1.470000 8.035000 1.800000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.525000 1.220000 8.535000 1.300000 ;
        RECT 6.525000 1.300000 6.935000 1.550000 ;
        RECT 6.765000 1.130000 8.535000 1.220000 ;
        RECT 8.205000 1.300000 8.535000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.870000 1.420000 6.200000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505000 1.220000 4.165000 1.265000 ;
        RECT 2.505000 1.265000 2.910000 1.550000 ;
        RECT 2.740000 1.095000 4.165000 1.220000 ;
        RECT 3.995000 1.265000 4.165000 1.470000 ;
        RECT 3.995000 1.470000 5.360000 1.640000 ;
        RECT 4.925000 1.640000 5.360000 1.800000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.435000 3.825000 1.780000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  1.345400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.140000 0.945000 1.310000 ;
        RECT 0.125000 1.310000 0.355000 1.480000 ;
        RECT 0.125000 1.480000 0.895000 1.650000 ;
        RECT 0.565000 1.650000 0.895000 1.720000 ;
        RECT 0.565000 1.720000 1.895000 1.890000 ;
        RECT 0.565000 1.890000 0.895000 2.980000 ;
        RECT 0.615000 0.350000 0.945000 0.880000 ;
        RECT 0.615000 0.880000 2.070000 1.050000 ;
        RECT 0.615000 1.050000 0.945000 1.140000 ;
        RECT 1.565000 1.890000 1.895000 2.980000 ;
        RECT 1.740000 0.350000 2.070000 0.880000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
      RECT 0.000000  3.245000 8.640000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 0.970000 ;
      RECT 0.115000  1.820000 0.365000 3.245000 ;
      RECT 1.065000  2.060000 1.395000 3.245000 ;
      RECT 1.115000  0.085000 1.570000 0.680000 ;
      RECT 1.255000  1.220000 2.265000 1.550000 ;
      RECT 2.095000  1.550000 2.265000 1.720000 ;
      RECT 2.095000  1.720000 2.985000 1.890000 ;
      RECT 2.150000  2.060000 2.480000 3.245000 ;
      RECT 2.240000  0.085000 2.570000 1.050000 ;
      RECT 2.655000  1.890000 2.985000 1.950000 ;
      RECT 2.655000  1.950000 4.420000 1.970000 ;
      RECT 2.655000  1.970000 6.100000 2.120000 ;
      RECT 2.655000  2.120000 2.985000 2.980000 ;
      RECT 2.800000  0.255000 5.595000 0.425000 ;
      RECT 2.800000  0.425000 3.130000 0.925000 ;
      RECT 3.225000  2.290000 3.920000 3.245000 ;
      RECT 3.300000  0.595000 5.095000 0.765000 ;
      RECT 3.300000  0.765000 4.075000 0.925000 ;
      RECT 4.090000  1.940000 4.420000 1.950000 ;
      RECT 4.090000  2.120000 6.100000 2.140000 ;
      RECT 4.090000  2.140000 4.420000 2.980000 ;
      RECT 4.335000  0.935000 4.585000 1.130000 ;
      RECT 4.335000  1.130000 5.700000 1.300000 ;
      RECT 4.590000  2.310000 4.920000 2.370000 ;
      RECT 4.590000  2.370000 7.575000 2.395000 ;
      RECT 4.590000  2.395000 6.550000 2.540000 ;
      RECT 4.590000  2.540000 4.920000 3.245000 ;
      RECT 4.765000  0.765000 5.095000 0.960000 ;
      RECT 5.150000  2.710000 6.550000 2.905000 ;
      RECT 5.150000  2.905000 8.525000 2.960000 ;
      RECT 5.265000  0.425000 5.595000 0.790000 ;
      RECT 5.265000  0.790000 8.525000 0.960000 ;
      RECT 5.530000  1.300000 5.700000 1.950000 ;
      RECT 5.530000  1.950000 6.100000 1.970000 ;
      RECT 5.750000  2.140000 6.100000 2.200000 ;
      RECT 5.765000  0.085000 6.095000 0.620000 ;
      RECT 6.220000  2.960000 8.525000 3.075000 ;
      RECT 6.265000  0.370000 6.595000 0.790000 ;
      RECT 6.265000  0.960000 6.595000 1.050000 ;
      RECT 6.380000  1.970000 7.575000 2.370000 ;
      RECT 6.720000  2.565000 8.025000 2.735000 ;
      RECT 6.765000  0.085000 7.095000 0.620000 ;
      RECT 7.265000  0.350000 7.595000 0.790000 ;
      RECT 7.765000  0.085000 8.095000 0.620000 ;
      RECT 7.775000  1.970000 8.025000 2.565000 ;
      RECT 8.195000  1.970000 8.525000 2.905000 ;
      RECT 8.275000  0.350000 8.525000 0.790000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
  END
END sky130_fd_sc_hs__o311a_4
MACRO sky130_fd_sc_hs__o311ai_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 0.705000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945000 1.350000 1.315000 2.890000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.515000 1.180000 1.845000 1.550000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.180000 2.415000 1.550000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925000 1.180000 3.255000 1.550000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.011700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.785000 1.720000 3.235000 1.890000 ;
        RECT 1.785000 1.890000 2.115000 2.980000 ;
        RECT 2.585000 0.350000 3.110000 1.010000 ;
        RECT 2.585000 1.010000 2.755000 1.720000 ;
        RECT 2.805000 1.890000 3.235000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 1.130000 ;
      RECT 0.225000  1.950000 0.555000 3.245000 ;
      RECT 0.615000  0.350000 0.945000 0.840000 ;
      RECT 0.615000  0.840000 2.220000 1.010000 ;
      RECT 0.615000  1.010000 0.945000 1.130000 ;
      RECT 1.115000  0.085000 1.675000 0.650000 ;
      RECT 1.890000  0.330000 2.220000 0.840000 ;
      RECT 2.285000  2.060000 2.615000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__o311ai_1
MACRO sky130_fd_sc_hs__o311ai_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 0.835000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.350000 2.275000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.350000 3.235000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.350000 4.195000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925000 1.300000 5.635000 1.780000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.754600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.600000 1.950000 5.630000 2.120000 ;
        RECT 2.600000 2.120000 2.930000 2.735000 ;
        RECT 3.500000 2.120000 3.750000 2.980000 ;
        RECT 4.400000 0.595000 4.705000 0.960000 ;
        RECT 4.400000 0.960000 5.645000 1.130000 ;
        RECT 4.400000 1.130000 4.730000 1.950000 ;
        RECT 4.480000 2.120000 4.650000 2.980000 ;
        RECT 5.300000 2.120000 5.630000 2.980000 ;
        RECT 5.395000 0.350000 5.645000 0.960000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.115000  0.350000 0.365000 1.010000 ;
      RECT 0.115000  1.010000 4.225000 1.180000 ;
      RECT 0.120000  1.950000 2.370000 2.120000 ;
      RECT 0.120000  2.120000 0.450000 2.980000 ;
      RECT 0.545000  0.085000 0.875000 0.840000 ;
      RECT 0.650000  2.290000 0.900000 3.245000 ;
      RECT 1.070000  2.120000 1.400000 2.980000 ;
      RECT 1.115000  0.350000 1.365000 1.010000 ;
      RECT 1.535000  0.085000 1.865000 0.840000 ;
      RECT 1.590000  2.290000 1.920000 2.905000 ;
      RECT 1.590000  2.905000 3.300000 3.075000 ;
      RECT 2.045000  0.350000 2.295000 1.010000 ;
      RECT 2.120000  2.120000 2.370000 2.735000 ;
      RECT 2.465000  0.085000 2.795000 0.840000 ;
      RECT 2.975000  0.350000 3.225000 1.010000 ;
      RECT 3.130000  2.290000 3.300000 2.905000 ;
      RECT 3.395000  0.255000 5.215000 0.425000 ;
      RECT 3.395000  0.425000 3.725000 0.840000 ;
      RECT 3.895000  0.595000 4.225000 1.010000 ;
      RECT 3.950000  2.290000 4.280000 3.245000 ;
      RECT 4.850000  2.290000 5.100000 3.245000 ;
      RECT 4.885000  0.425000 5.215000 0.790000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_hs__o311ai_2
MACRO sky130_fd_sc_hs__o311ai_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.165000 1.350000 10.435000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.765000 1.350000 7.775000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.485000 1.430000 6.195000 1.640000 ;
        RECT 5.185000 1.640000 6.195000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.245000 1.430000 4.195000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 1.240000 1.780000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  2.271700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.770000 1.740000 1.090000 ;
        RECT 0.545000 1.090000 6.595000 1.100000 ;
        RECT 0.740000 1.950000 6.595000 2.120000 ;
        RECT 0.740000 2.120000 1.070000 2.980000 ;
        RECT 1.410000 1.100000 6.595000 1.260000 ;
        RECT 1.740000 1.820000 2.070000 1.950000 ;
        RECT 1.740000 2.120000 2.070000 2.980000 ;
        RECT 4.685000 1.820000 5.015000 1.950000 ;
        RECT 4.685000 2.120000 5.015000 2.735000 ;
        RECT 5.685000 2.120000 6.015000 2.735000 ;
        RECT 6.365000 1.260000 6.595000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.040000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 11.040000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  3.245000 11.040000 3.415000 ;
      RECT  0.115000  0.350000  2.090000 0.600000 ;
      RECT  0.115000  0.600000  0.365000 1.130000 ;
      RECT  0.115000  1.950000  0.445000 3.245000 ;
      RECT  1.240000  2.290000  1.570000 3.245000 ;
      RECT  1.920000  0.600000  2.090000 0.750000 ;
      RECT  1.920000  0.750000  3.900000 0.920000 ;
      RECT  2.240000  2.290000  3.905000 3.245000 ;
      RECT  2.270000  0.330000  4.240000 0.580000 ;
      RECT  4.070000  0.580000  4.240000 0.750000 ;
      RECT  4.070000  0.750000  7.140000 0.920000 ;
      RECT  4.185000  2.290000  4.515000 2.905000 ;
      RECT  4.185000  2.905000  8.565000 3.075000 ;
      RECT  4.410000  0.085000  4.740000 0.580000 ;
      RECT  4.920000  0.350000  5.170000 0.750000 ;
      RECT  5.185000  2.290000  5.515000 2.905000 ;
      RECT  5.350000  0.085000  5.680000 0.580000 ;
      RECT  5.860000  0.350000  6.190000 0.750000 ;
      RECT  6.285000  2.290000  6.615000 2.905000 ;
      RECT  6.370000  0.085000  6.710000 0.580000 ;
      RECT  6.785000  1.950000 10.475000 2.120000 ;
      RECT  6.785000  2.120000  7.115000 2.735000 ;
      RECT  6.890000  0.350000  7.140000 0.750000 ;
      RECT  6.890000  0.920000  7.140000 1.010000 ;
      RECT  6.890000  1.010000  8.115000 1.180000 ;
      RECT  7.285000  2.290000  7.615000 2.905000 ;
      RECT  7.320000  0.085000  7.650000 0.825000 ;
      RECT  7.785000  2.120000 10.475000 2.150000 ;
      RECT  7.785000  2.150000  8.065000 2.735000 ;
      RECT  7.945000  0.350000  8.115000 1.010000 ;
      RECT  7.945000  1.180000  8.115000 1.300000 ;
      RECT  7.945000  1.300000  8.975000 1.470000 ;
      RECT  8.235000  2.330000  8.565000 2.905000 ;
      RECT  8.295000  0.085000  8.545000 1.130000 ;
      RECT  8.725000  0.350000  8.975000 0.960000 ;
      RECT  8.725000  0.960000 10.415000 1.130000 ;
      RECT  8.725000  1.130000  8.975000 1.300000 ;
      RECT  8.795000  2.330000  9.125000 3.245000 ;
      RECT  9.155000  0.085000  9.995000 0.790000 ;
      RECT  9.295000  2.150000  9.525000 2.980000 ;
      RECT  9.695000  2.330000 10.025000 3.245000 ;
      RECT 10.165000  0.350000 10.415000 0.960000 ;
      RECT 10.195000  2.150000 10.475000 2.980000 ;
      RECT 10.595000  0.085000 10.925000 1.130000 ;
      RECT 10.675000  1.820000 10.925000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
  END
END sky130_fd_sc_hs__o311ai_4
MACRO sky130_fd_sc_hs__o31a_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965000 1.350000 1.315000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505000 1.300000 1.835000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.350000 2.375000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.545000 1.350000 2.915000 1.780000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.350000 0.445000 1.130000 ;
        RECT 0.085000 1.130000 0.255000 1.820000 ;
        RECT 0.085000 1.820000 0.455000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.425000  1.320000 0.795000 1.650000 ;
      RECT 0.615000  0.085000 0.945000 1.130000 ;
      RECT 0.625000  1.650000 0.795000 1.950000 ;
      RECT 0.625000  1.950000 3.255000 2.120000 ;
      RECT 0.625000  2.290000 1.090000 3.245000 ;
      RECT 1.125000  0.450000 1.460000 0.960000 ;
      RECT 1.125000  0.960000 2.745000 1.130000 ;
      RECT 1.765000  0.085000 2.130000 0.780000 ;
      RECT 2.195000  2.120000 2.525000 2.880000 ;
      RECT 2.415000  0.450000 2.745000 0.960000 ;
      RECT 2.735000  2.290000 3.050000 3.245000 ;
      RECT 2.915000  0.450000 3.255000 1.130000 ;
      RECT 3.085000  1.130000 3.255000 1.950000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__o31a_1
MACRO sky130_fd_sc_hs__o31a_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415000 1.350000 1.795000 2.150000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 1.470000 2.315000 2.150000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.180000 2.885000 1.550000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.395000 1.300000 3.725000 1.780000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.604800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565000 1.820000 0.950000 2.150000 ;
        RECT 0.615000 0.350000 0.945000 1.130000 ;
        RECT 0.775000 1.130000 0.945000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 1.130000 ;
      RECT 0.115000  2.660000 0.445000 3.245000 ;
      RECT 0.225000  1.320000 0.605000 1.650000 ;
      RECT 0.225000  1.650000 0.395000 2.320000 ;
      RECT 0.225000  2.320000 3.225000 2.490000 ;
      RECT 1.070000  2.660000 1.595000 3.245000 ;
      RECT 1.115000  0.085000 1.445000 1.130000 ;
      RECT 1.615000  0.350000 1.945000 0.770000 ;
      RECT 1.615000  0.770000 3.225000 0.790000 ;
      RECT 1.615000  0.790000 2.850000 0.940000 ;
      RECT 1.615000  0.940000 1.945000 1.130000 ;
      RECT 2.115000  0.085000 2.510000 0.600000 ;
      RECT 2.680000  0.460000 3.225000 0.770000 ;
      RECT 2.765000  1.940000 3.225000 2.320000 ;
      RECT 2.765000  2.490000 3.225000 2.980000 ;
      RECT 3.055000  0.960000 3.725000 1.130000 ;
      RECT 3.055000  1.130000 3.225000 1.940000 ;
      RECT 3.395000  0.350000 3.725000 0.960000 ;
      RECT 3.395000  1.950000 3.725000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__o31a_2
MACRO sky130_fd_sc_hs__o31a_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.405000 1.455000 5.875000 1.785000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.115000 1.455000 6.595000 1.785000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.455000 5.155000 1.785000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905000 1.470000 3.235000 2.150000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.575000 0.350000 0.905000 0.960000 ;
        RECT 0.575000 0.960000 1.700000 1.130000 ;
        RECT 0.575000 1.130000 0.835000 1.800000 ;
        RECT 0.575000 1.800000 1.810000 1.970000 ;
        RECT 0.575000 1.970000 0.835000 2.980000 ;
        RECT 1.450000 0.350000 1.700000 0.960000 ;
        RECT 1.480000 1.970000 1.810000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.720000 0.085000 ;
      RECT 0.000000  3.245000 6.720000 3.415000 ;
      RECT 0.130000  1.820000 0.380000 3.245000 ;
      RECT 0.145000  0.085000 0.395000 1.130000 ;
      RECT 1.005000  1.300000 2.715000 1.630000 ;
      RECT 1.030000  2.140000 1.280000 3.245000 ;
      RECT 1.085000  0.085000 1.255000 0.790000 ;
      RECT 1.880000  0.085000 2.210000 1.130000 ;
      RECT 2.010000  1.820000 2.260000 3.245000 ;
      RECT 2.440000  0.265000 3.780000 0.435000 ;
      RECT 2.440000  0.435000 2.770000 0.960000 ;
      RECT 2.465000  1.630000 2.715000 2.375000 ;
      RECT 2.465000  2.375000 4.255000 2.545000 ;
      RECT 2.465000  2.545000 2.715000 2.980000 ;
      RECT 2.545000  1.130000 3.270000 1.300000 ;
      RECT 2.915000  2.715000 3.245000 3.245000 ;
      RECT 2.940000  0.605000 3.270000 1.130000 ;
      RECT 3.450000  0.435000 3.780000 1.115000 ;
      RECT 3.450000  1.115000 6.580000 1.285000 ;
      RECT 3.475000  1.955000 6.605000 2.125000 ;
      RECT 3.475000  2.125000 4.645000 2.205000 ;
      RECT 3.925000  2.545000 4.255000 2.980000 ;
      RECT 3.960000  0.085000 4.210000 0.945000 ;
      RECT 4.390000  0.605000 4.640000 1.115000 ;
      RECT 4.435000  2.205000 4.645000 2.980000 ;
      RECT 4.820000  0.085000 5.150000 0.945000 ;
      RECT 4.825000  2.295000 6.105000 2.465000 ;
      RECT 4.825000  2.465000 5.075000 2.980000 ;
      RECT 5.275000  2.635000 5.605000 3.245000 ;
      RECT 5.320000  0.605000 5.570000 1.115000 ;
      RECT 5.750000  0.085000 6.080000 0.945000 ;
      RECT 5.775000  2.465000 6.105000 2.980000 ;
      RECT 6.250000  0.605000 6.580000 1.115000 ;
      RECT 6.275000  2.125000 6.605000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
  END
END sky130_fd_sc_hs__o31a_4
MACRO sky130_fd_sc_hs__o31ai_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.880000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.435000 1.550000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.300000 1.180000 2.890000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.690000 1.350000 2.275000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 1.300000 2.775000 1.780000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.020700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.350000 0.960000 2.765000 1.130000 ;
        RECT 1.350000 1.130000 1.520000 1.950000 ;
        RECT 1.350000 1.950000 2.230000 2.980000 ;
        RECT 2.435000 0.350000 2.765000 0.960000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.880000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.880000 0.085000 ;
      RECT 0.000000  3.245000 2.880000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 1.010000 ;
      RECT 0.130000  1.820000 0.380000 3.245000 ;
      RECT 0.625000  0.350000 0.875000 0.620000 ;
      RECT 0.625000  0.620000 2.265000 0.790000 ;
      RECT 0.625000  0.790000 0.875000 1.130000 ;
      RECT 1.055000  0.085000 1.755000 0.450000 ;
      RECT 1.935000  0.350000 2.265000 0.620000 ;
      RECT 2.410000  1.950000 2.740000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
  END
END sky130_fd_sc_hs__o31ai_1
MACRO sky130_fd_sc_hs__o31ai_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.315000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.350000 2.275000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.350000 3.445000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.685000 1.350000 4.695000 1.680000 ;
        RECT 4.365000 1.180000 4.695000 1.350000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.297000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505000 1.820000 2.835000 1.950000 ;
        RECT 2.505000 1.950000 4.685000 2.020000 ;
        RECT 2.505000 2.020000 3.785000 2.120000 ;
        RECT 2.505000 2.120000 2.755000 2.735000 ;
        RECT 2.665000 1.010000 4.180000 1.180000 ;
        RECT 2.665000 1.180000 2.835000 1.820000 ;
        RECT 3.455000 2.120000 3.785000 2.980000 ;
        RECT 3.615000 1.850000 4.685000 1.950000 ;
        RECT 3.850000 0.610000 4.180000 1.010000 ;
        RECT 4.355000 2.020000 4.685000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.115000  0.350000 0.445000 1.010000 ;
      RECT 0.115000  1.010000 2.445000 1.180000 ;
      RECT 0.120000  1.950000 2.250000 2.120000 ;
      RECT 0.120000  2.120000 0.370000 2.980000 ;
      RECT 0.570000  2.290000 0.820000 3.245000 ;
      RECT 0.615000  0.085000 0.945000 0.825000 ;
      RECT 1.020000  2.120000 1.350000 2.980000 ;
      RECT 1.115000  0.350000 1.445000 1.010000 ;
      RECT 1.550000  2.290000 1.720000 2.905000 ;
      RECT 1.550000  2.905000 3.285000 3.075000 ;
      RECT 1.615000  0.085000 1.945000 0.825000 ;
      RECT 1.920000  2.120000 2.250000 2.735000 ;
      RECT 2.115000  0.350000 2.445000 0.670000 ;
      RECT 2.115000  0.670000 3.670000 0.840000 ;
      RECT 2.115000  0.840000 2.445000 1.010000 ;
      RECT 2.625000  0.085000 3.240000 0.500000 ;
      RECT 2.955000  2.290000 3.285000 2.905000 ;
      RECT 3.420000  0.255000 4.680000 0.425000 ;
      RECT 3.420000  0.425000 3.670000 0.670000 ;
      RECT 3.985000  2.190000 4.155000 3.245000 ;
      RECT 4.350000  0.425000 4.680000 1.010000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_hs__o31ai_2
MACRO sky130_fd_sc_hs__o31ai_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.795000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.350000 3.715000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.835000 1.350000 6.115000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365000 1.350000 7.790000 1.780000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.803200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.550000 4.665000 1.950000 ;
        RECT 3.965000 1.950000 8.525000 2.120000 ;
        RECT 3.965000 2.120000 4.970000 2.150000 ;
        RECT 4.495000 1.010000 8.095000 1.180000 ;
        RECT 4.495000 1.180000 4.665000 1.550000 ;
        RECT 4.700000 2.150000 4.970000 2.735000 ;
        RECT 5.600000 2.120000 5.930000 2.735000 ;
        RECT 6.550000 2.120000 6.880000 2.980000 ;
        RECT 6.905000 0.920000 8.095000 1.010000 ;
        RECT 8.195000 1.820000 8.525000 1.950000 ;
        RECT 8.195000 2.120000 8.525000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
      RECT 0.000000  3.245000 8.640000 3.415000 ;
      RECT 0.115000  0.390000 0.445000 0.920000 ;
      RECT 0.115000  0.920000 2.305000 1.010000 ;
      RECT 0.115000  1.010000 4.325000 1.180000 ;
      RECT 0.120000  1.950000 3.300000 2.120000 ;
      RECT 0.120000  2.120000 0.370000 2.980000 ;
      RECT 0.570000  2.290000 0.900000 3.245000 ;
      RECT 0.615000  0.085000 0.945000 0.750000 ;
      RECT 1.100000  2.120000 1.270000 2.980000 ;
      RECT 1.470000  2.290000 1.800000 3.245000 ;
      RECT 1.475000  0.085000 1.805000 0.750000 ;
      RECT 1.970000  1.820000 2.300000 1.950000 ;
      RECT 1.970000  2.120000 2.300000 2.980000 ;
      RECT 1.975000  0.390000 2.305000 0.920000 ;
      RECT 2.470000  2.290000 2.800000 2.905000 ;
      RECT 2.470000  2.905000 6.380000 3.075000 ;
      RECT 2.495000  0.085000 2.960000 0.805000 ;
      RECT 2.970000  2.120000 3.300000 2.370000 ;
      RECT 2.970000  2.370000 4.470000 2.540000 ;
      RECT 2.970000  2.540000 3.300000 2.735000 ;
      RECT 3.145000  0.390000 3.475000 1.010000 ;
      RECT 3.640000  2.710000 3.970000 2.905000 ;
      RECT 3.645000  0.085000 3.975000 0.840000 ;
      RECT 4.140000  2.540000 4.470000 2.735000 ;
      RECT 4.155000  0.390000 4.325000 0.670000 ;
      RECT 4.155000  0.670000 6.805000 0.750000 ;
      RECT 4.155000  0.750000 5.775000 0.840000 ;
      RECT 4.155000  0.840000 4.325000 1.010000 ;
      RECT 4.585000  0.085000 5.265000 0.500000 ;
      RECT 5.150000  2.290000 5.400000 2.905000 ;
      RECT 5.445000  0.390000 5.775000 0.580000 ;
      RECT 5.445000  0.580000 6.805000 0.670000 ;
      RECT 5.955000  0.085000 6.295000 0.410000 ;
      RECT 6.130000  2.290000 6.380000 2.905000 ;
      RECT 6.475000  0.390000 8.525000 0.560000 ;
      RECT 6.475000  0.560000 6.805000 0.580000 ;
      RECT 7.050000  2.290000 8.025000 3.245000 ;
      RECT 7.335000  0.560000 7.665000 0.750000 ;
      RECT 8.265000  0.560000 8.525000 1.170000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
  END
END sky130_fd_sc_hs__o31ai_4
MACRO sky130_fd_sc_hs__o32a_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955000 1.350000 1.315000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.495000 1.350000 1.825000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.035000 1.350000 2.365000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.410000 1.180000 3.735000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.535000 1.350000 2.895000 1.780000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.350000 0.560000 1.130000 ;
        RECT 0.085000 1.130000 0.255000 1.820000 ;
        RECT 0.085000 1.820000 0.445000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.425000  1.320000 0.785000 1.650000 ;
      RECT 0.615000  1.650000 0.785000 1.950000 ;
      RECT 0.615000  1.950000 3.235000 2.120000 ;
      RECT 0.615000  2.290000 0.945000 3.245000 ;
      RECT 0.730000  0.085000 1.060000 1.030000 ;
      RECT 1.230000  0.350000 1.560000 1.010000 ;
      RECT 1.230000  1.010000 2.560000 1.180000 ;
      RECT 1.730000  0.085000 2.060000 0.820000 ;
      RECT 2.205000  2.120000 2.595000 2.880000 ;
      RECT 2.230000  0.340000 3.655000 0.520000 ;
      RECT 2.230000  0.520000 2.560000 1.010000 ;
      RECT 2.730000  0.700000 3.225000 1.010000 ;
      RECT 2.730000  1.010000 3.235000 1.180000 ;
      RECT 3.065000  1.180000 3.235000 1.950000 ;
      RECT 3.320000  2.290000 3.650000 3.245000 ;
      RECT 3.405000  0.520000 3.655000 1.010000 ;
      RECT 3.410000  1.970000 3.650000 2.290000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__o32a_1
MACRO sky130_fd_sc_hs__o32a_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415000 1.350000 1.795000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 1.350000 2.315000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.350000 2.855000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.355000 1.180000 4.685000 2.890000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.095000 1.350000 3.715000 1.780000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.960000 1.050000 1.130000 ;
        RECT 0.535000 1.130000 0.705000 1.820000 ;
        RECT 0.535000 1.820000 0.895000 2.980000 ;
        RECT 0.720000 0.350000 1.050000 0.960000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.115000  0.085000 0.540000 0.790000 ;
      RECT 0.115000  0.790000 0.365000 1.140000 ;
      RECT 0.115000  1.820000 0.365000 3.245000 ;
      RECT 0.875000  1.320000 1.235000 1.650000 ;
      RECT 1.065000  1.650000 1.235000 1.950000 ;
      RECT 1.065000  1.950000 4.185000 2.120000 ;
      RECT 1.065000  2.290000 1.600000 3.245000 ;
      RECT 1.220000  0.085000 1.550000 1.130000 ;
      RECT 1.720000  0.350000 2.050000 1.010000 ;
      RECT 1.720000  1.010000 3.050000 1.180000 ;
      RECT 2.220000  0.085000 2.550000 0.840000 ;
      RECT 2.675000  2.120000 3.110000 2.880000 ;
      RECT 2.720000  0.350000 4.615000 0.520000 ;
      RECT 2.720000  0.520000 3.050000 1.010000 ;
      RECT 3.220000  0.715000 4.185000 1.045000 ;
      RECT 3.815000  2.290000 4.145000 3.245000 ;
      RECT 4.015000  1.045000 4.185000 1.950000 ;
      RECT 4.355000  0.520000 4.615000 1.010000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_hs__o32a_2
MACRO sky130_fd_sc_hs__o32a_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.845000 1.120000 7.295000 1.410000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.075000 1.130000 6.405000 1.580000 ;
        RECT 6.075000 1.580000 8.035000 1.780000 ;
        RECT 6.075000 1.780000 6.405000 1.800000 ;
        RECT 7.565000 1.450000 8.035000 1.580000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.065000 1.180000 5.735000 1.510000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.450000 2.855000 1.780000 ;
        RECT 2.685000 1.780000 2.855000 2.360000 ;
        RECT 2.685000 2.360000 5.905000 2.530000 ;
        RECT 4.495000 1.450000 4.825000 1.680000 ;
        RECT 4.495000 1.680000 5.905000 1.850000 ;
        RECT 5.735000 1.850000 5.905000 2.360000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.925000 1.270000 4.255000 1.780000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  1.313300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.140000 1.015000 1.310000 ;
        RECT 0.125000 1.310000 0.355000 1.480000 ;
        RECT 0.125000 1.480000 0.895000 1.650000 ;
        RECT 0.565000 1.650000 0.895000 1.780000 ;
        RECT 0.565000 1.780000 1.895000 1.950000 ;
        RECT 0.565000 1.950000 0.895000 2.980000 ;
        RECT 0.685000 0.350000 1.015000 0.940000 ;
        RECT 0.685000 0.940000 2.015000 1.110000 ;
        RECT 0.685000 1.110000 1.015000 1.140000 ;
        RECT 1.565000 1.950000 1.895000 2.980000 ;
        RECT 1.685000 0.350000 2.015000 0.940000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.115000  1.820000 0.365000 3.245000 ;
      RECT 0.185000  0.085000 0.515000 0.970000 ;
      RECT 1.065000  2.120000 1.395000 3.245000 ;
      RECT 1.185000  0.085000 1.515000 0.770000 ;
      RECT 1.255000  1.280000 2.355000 1.610000 ;
      RECT 2.085000  1.950000 2.415000 3.245000 ;
      RECT 2.185000  1.110000 3.560000 1.280000 ;
      RECT 2.240000  0.085000 2.570000 0.940000 ;
      RECT 2.655000  2.700000 4.025000 2.960000 ;
      RECT 2.800000  0.255000 5.060000 0.425000 ;
      RECT 2.800000  0.425000 3.130000 0.940000 ;
      RECT 3.230000  1.280000 3.560000 1.920000 ;
      RECT 3.230000  1.920000 3.575000 2.020000 ;
      RECT 3.230000  2.020000 5.565000 2.190000 ;
      RECT 3.300000  0.595000 3.560000 0.930000 ;
      RECT 3.300000  0.930000 4.560000 1.100000 ;
      RECT 3.300000  1.100000 3.560000 1.110000 ;
      RECT 3.730000  0.425000 4.060000 0.760000 ;
      RECT 4.195000  2.700000 4.525000 3.245000 ;
      RECT 4.230000  0.595000 4.560000 0.930000 ;
      RECT 4.730000  0.425000 5.060000 0.790000 ;
      RECT 4.730000  0.790000 8.045000 0.950000 ;
      RECT 4.730000  0.950000 6.060000 0.960000 ;
      RECT 4.730000  0.960000 5.060000 1.010000 ;
      RECT 4.785000  2.700000 6.245000 2.980000 ;
      RECT 5.230000  0.085000 5.560000 0.620000 ;
      RECT 5.730000  0.350000 6.060000 0.780000 ;
      RECT 5.730000  0.780000 8.045000 0.790000 ;
      RECT 6.075000  2.390000 8.045000 2.560000 ;
      RECT 6.075000  2.560000 6.245000 2.700000 ;
      RECT 6.155000  1.970000 7.595000 2.200000 ;
      RECT 6.155000  2.200000 6.675000 2.220000 ;
      RECT 6.230000  0.085000 6.560000 0.610000 ;
      RECT 6.740000  0.350000 6.990000 0.780000 ;
      RECT 6.805000  2.730000 7.135000 3.245000 ;
      RECT 7.160000  0.085000 7.545000 0.600000 ;
      RECT 7.265000  1.950000 7.595000 1.970000 ;
      RECT 7.715000  0.350000 8.045000 0.780000 ;
      RECT 7.715000  0.950000 8.045000 1.030000 ;
      RECT 7.715000  2.560000 8.045000 2.980000 ;
      RECT 7.765000  1.950000 8.045000 2.390000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_hs__o32a_4
MACRO sky130_fd_sc_hs__o32ai_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.880000 1.180000 3.235000 1.550000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.350000 2.445000 2.890000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.545000 1.350000 1.875000 2.520000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 1.180000 0.445000 1.550000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.975000 1.350000 1.315000 1.780000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.992900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.615000 0.720000 1.140000 1.130000 ;
        RECT 0.635000 1.130000 0.805000 1.950000 ;
        RECT 0.635000 1.950000 1.375000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.115000  0.350000 1.680000 0.520000 ;
      RECT 0.115000  0.520000 0.445000 1.010000 ;
      RECT 0.135000  1.820000 0.465000 3.245000 ;
      RECT 1.350000  0.520000 1.680000 1.010000 ;
      RECT 1.350000  1.010000 2.710000 1.180000 ;
      RECT 1.850000  0.085000 2.180000 0.810000 ;
      RECT 2.380000  0.350000 2.710000 1.010000 ;
      RECT 2.835000  1.820000 3.165000 3.245000 ;
      RECT 2.880000  0.085000 3.140000 1.010000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__o32ai_1
MACRO sky130_fd_sc_hs__o32ai_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.350000 6.115000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.350000 4.195000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.350000 2.755000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 1.350000 1.815000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.315000 1.780000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.138200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.610000 0.875000 1.010000 ;
        RECT 0.545000 1.010000 3.095000 1.180000 ;
        RECT 0.565000 1.950000 3.255000 2.120000 ;
        RECT 0.565000 2.120000 0.895000 2.735000 ;
        RECT 1.545000 0.610000 1.875000 1.010000 ;
        RECT 2.925000 1.180000 3.095000 1.820000 ;
        RECT 2.925000 1.820000 3.255000 1.950000 ;
        RECT 2.925000 2.120000 3.255000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.240000 0.085000 ;
      RECT 0.000000  3.245000 6.240000 3.415000 ;
      RECT 0.115000  0.255000 2.375000 0.425000 ;
      RECT 0.115000  0.425000 0.365000 1.130000 ;
      RECT 0.115000  1.950000 0.365000 2.905000 ;
      RECT 0.115000  2.905000 1.265000 3.075000 ;
      RECT 1.045000  0.425000 1.375000 0.825000 ;
      RECT 1.095000  2.290000 2.245000 2.460000 ;
      RECT 1.095000  2.460000 1.265000 2.905000 ;
      RECT 1.465000  2.630000 1.715000 3.245000 ;
      RECT 1.915000  2.460000 2.245000 2.980000 ;
      RECT 2.045000  0.425000 2.375000 0.670000 ;
      RECT 2.045000  0.670000 3.635000 0.840000 ;
      RECT 2.475000  2.290000 2.725000 2.905000 ;
      RECT 2.475000  2.905000 4.605000 3.075000 ;
      RECT 2.555000  0.085000 3.125000 0.500000 ;
      RECT 3.305000  0.350000 3.635000 0.670000 ;
      RECT 3.305000  0.840000 3.635000 1.010000 ;
      RECT 3.305000  1.010000 6.125000 1.180000 ;
      RECT 3.455000  1.950000 3.625000 2.905000 ;
      RECT 3.805000  0.085000 4.135000 0.800000 ;
      RECT 3.825000  1.950000 5.670000 2.120000 ;
      RECT 3.825000  2.120000 4.075000 2.735000 ;
      RECT 4.275000  2.290000 4.605000 2.905000 ;
      RECT 4.305000  0.350000 4.635000 1.010000 ;
      RECT 4.805000  0.085000 5.625000 0.805000 ;
      RECT 4.835000  2.290000 5.165000 3.245000 ;
      RECT 5.335000  2.120000 5.670000 2.980000 ;
      RECT 5.795000  0.350000 6.125000 1.010000 ;
      RECT 5.870000  1.950000 6.120000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
  END
END sky130_fd_sc_hs__o32ai_2
MACRO sky130_fd_sc_hs__o32ai_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.765000 1.350000 10.915000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365000 1.350000 8.515000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.430000 5.635000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.430000 4.195000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.430000 1.795000 1.780000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  2.287500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.595000 0.875000 1.090000 ;
        RECT 0.545000 1.090000 5.975000 1.260000 ;
        RECT 0.645000 1.950000 5.975000 2.120000 ;
        RECT 0.645000 2.120000 0.815000 2.735000 ;
        RECT 1.465000 2.120000 1.795000 2.735000 ;
        RECT 1.555000 0.595000 1.805000 1.090000 ;
        RECT 2.475000 0.595000 2.805000 1.090000 ;
        RECT 3.475000 0.595000 3.805000 1.090000 ;
        RECT 4.735000 2.120000 5.065000 2.735000 ;
        RECT 5.635000 2.120000 5.965000 2.735000 ;
        RECT 5.805000 1.260000 5.975000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.040000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 11.040000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  3.245000 11.040000 3.415000 ;
      RECT  0.115000  0.255000  4.305000 0.425000 ;
      RECT  0.115000  0.425000  0.365000 1.130000 ;
      RECT  0.115000  1.950000  0.445000 2.905000 ;
      RECT  0.115000  2.905000  2.245000 3.075000 ;
      RECT  1.015000  2.290000  1.265000 2.905000 ;
      RECT  1.045000  0.425000  1.375000 0.920000 ;
      RECT  1.975000  0.425000  2.305000 0.920000 ;
      RECT  1.995000  2.290000  4.055000 2.460000 ;
      RECT  1.995000  2.460000  2.245000 2.905000 ;
      RECT  2.445000  2.630000  2.615000 3.245000 ;
      RECT  2.815000  2.460000  3.145000 2.980000 ;
      RECT  2.975000  0.425000  3.305000 0.920000 ;
      RECT  3.345000  2.630000  3.515000 3.245000 ;
      RECT  3.725000  2.460000  4.055000 2.980000 ;
      RECT  3.975000  0.425000  4.305000 0.750000 ;
      RECT  3.975000  0.750000  6.670000 0.920000 ;
      RECT  4.285000  2.290000  4.535000 2.905000 ;
      RECT  4.285000  2.905000  8.465000 3.075000 ;
      RECT  4.485000  0.085000  4.815000 0.580000 ;
      RECT  4.995000  0.330000  5.325000 0.750000 ;
      RECT  5.265000  2.290000  5.435000 2.905000 ;
      RECT  5.495000  0.085000  5.825000 0.580000 ;
      RECT  5.995000  0.330000  6.670000 0.750000 ;
      RECT  6.145000  1.950000  6.465000 2.905000 ;
      RECT  6.330000  0.920000  6.670000 1.010000 ;
      RECT  6.330000  1.010000 10.670000 1.180000 ;
      RECT  6.635000  1.950000 10.475000 2.120000 ;
      RECT  6.635000  2.120000  6.965000 2.735000 ;
      RECT  6.840000  0.085000  7.170000 0.840000 ;
      RECT  7.135000  2.290000  7.465000 2.905000 ;
      RECT  7.340000  0.350000  7.670000 1.010000 ;
      RECT  7.635000  2.120000  7.965000 2.735000 ;
      RECT  7.840000  0.085000  8.170000 0.840000 ;
      RECT  8.135000  2.290000  8.465000 2.905000 ;
      RECT  8.340000  0.350000  8.670000 1.010000 ;
      RECT  8.695000  2.290000  8.945000 3.245000 ;
      RECT  8.840000  0.085000  9.170000 0.840000 ;
      RECT  9.145000  2.120000  9.475000 2.980000 ;
      RECT  9.340000  0.350000  9.670000 1.010000 ;
      RECT  9.645000  2.290000  9.975000 3.245000 ;
      RECT  9.840000  0.085000 10.170000 0.840000 ;
      RECT 10.145000  2.120000 10.475000 2.980000 ;
      RECT 10.340000  0.350000 10.670000 1.010000 ;
      RECT 10.675000  1.950000 10.925000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
  END
END sky130_fd_sc_hs__o32ai_4
MACRO sky130_fd_sc_hs__o41a_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.264000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.610000 1.350000 4.195000 2.150000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.264000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.300000 3.370000 2.890000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.264000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.470000 1.220000 2.800000 2.890000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.264000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.870000 1.190000 2.275000 1.780000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.450000 1.580000 1.780000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.350000 0.375000 1.130000 ;
        RECT 0.115000 1.130000 0.285000 2.290000 ;
        RECT 0.115000 2.290000 0.445000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.455000  1.350000 0.785000 1.950000 ;
      RECT 0.455000  1.950000 2.080000 2.120000 ;
      RECT 0.545000  0.085000 0.945000 0.940000 ;
      RECT 0.615000  1.110000 1.505000 1.280000 ;
      RECT 0.615000  1.280000 0.785000 1.350000 ;
      RECT 0.615000  2.290000 1.540000 3.245000 ;
      RECT 1.175000  0.350000 1.505000 1.110000 ;
      RECT 1.675000  0.350000 2.005000 0.850000 ;
      RECT 1.675000  0.850000 4.205000 1.020000 ;
      RECT 1.750000  2.120000 2.080000 2.845000 ;
      RECT 2.175000  0.085000 2.505000 0.680000 ;
      RECT 2.675000  0.350000 3.005000 0.850000 ;
      RECT 3.175000  0.085000 3.705000 0.680000 ;
      RECT 3.760000  2.320000 4.205000 3.245000 ;
      RECT 3.875000  0.350000 4.205000 0.850000 ;
      RECT 3.875000  1.020000 4.205000 1.030000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__o41a_1
MACRO sky130_fd_sc_hs__o41a_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 0.595000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.835000 1.350000 1.165000 1.920000 ;
        RECT 0.835000 1.920000 1.315000 2.890000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.405000 1.350000 1.795000 1.680000 ;
        RECT 1.565000 1.680000 1.795000 2.890000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975000 1.350000 2.305000 1.780000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.350000 3.235000 1.780000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.855000 0.350000 4.185000 1.130000 ;
        RECT 3.950000 1.130000 4.185000 1.180000 ;
        RECT 3.950000 1.180000 4.195000 1.410000 ;
        RECT 3.950000 1.410000 4.155000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.115000  0.350000 0.445000 1.010000 ;
      RECT 0.115000  1.010000 2.625000 1.180000 ;
      RECT 0.115000  1.950000 0.445000 3.245000 ;
      RECT 0.615000  0.085000 0.945000 0.840000 ;
      RECT 1.115000  0.350000 1.445000 1.010000 ;
      RECT 1.615000  0.085000 2.125000 0.815000 ;
      RECT 2.125000  1.950000 3.735000 2.120000 ;
      RECT 2.125000  2.120000 2.455000 2.980000 ;
      RECT 2.295000  0.350000 2.625000 1.010000 ;
      RECT 2.695000  2.290000 3.780000 3.245000 ;
      RECT 2.795000  0.350000 3.125000 1.010000 ;
      RECT 2.795000  1.010000 3.575000 1.180000 ;
      RECT 3.355000  0.085000 3.685000 0.820000 ;
      RECT 3.405000  1.180000 3.575000 1.300000 ;
      RECT 3.405000  1.300000 3.735000 1.950000 ;
      RECT 4.355000  0.085000 4.615000 1.010000 ;
      RECT 4.355000  1.820000 4.685000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_hs__o41a_2
MACRO sky130_fd_sc_hs__o41a_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.528000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.330000 1.420000 7.075000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.528000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.305000 0.255000 7.635000 0.335000 ;
        RECT 7.305000 0.335000 8.035000 0.505000 ;
        RECT 7.805000 0.505000 8.035000 0.670000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.528000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.875000 0.255000 4.205000 0.670000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.528000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.425000 5.180000 1.780000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.444000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.280000 1.440000 4.195000 1.780000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.930000 1.855000 1.100000 ;
        RECT 0.125000 1.100000 0.295000 1.770000 ;
        RECT 0.125000 1.770000 2.125000 1.940000 ;
        RECT 0.125000 1.940000 0.355000 2.890000 ;
        RECT 0.675000 0.350000 0.925000 0.930000 ;
        RECT 0.895000 1.940000 1.225000 2.980000 ;
        RECT 1.605000 0.350000 1.855000 0.930000 ;
        RECT 1.795000 1.940000 2.125000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.175000  0.085000 0.505000 0.760000 ;
      RECT 0.525000  2.110000 0.695000 3.245000 ;
      RECT 0.585000  1.270000 3.110000 1.600000 ;
      RECT 1.105000  0.085000 1.435000 0.760000 ;
      RECT 1.425000  2.110000 1.595000 3.245000 ;
      RECT 2.035000  0.085000 2.365000 1.100000 ;
      RECT 2.325000  1.910000 2.575000 3.245000 ;
      RECT 2.595000  0.260000 3.705000 0.430000 ;
      RECT 2.595000  0.430000 2.925000 0.930000 ;
      RECT 2.780000  1.600000 3.110000 1.950000 ;
      RECT 2.780000  1.950000 5.030000 2.120000 ;
      RECT 2.780000  2.120000 3.110000 2.790000 ;
      RECT 2.940000  1.100000 3.275000 1.270000 ;
      RECT 3.105000  0.600000 3.275000 1.100000 ;
      RECT 3.310000  2.290000 3.560000 3.245000 ;
      RECT 3.455000  0.430000 3.705000 1.085000 ;
      RECT 3.455000  1.085000 7.635000 1.250000 ;
      RECT 3.455000  1.250000 5.845000 1.255000 ;
      RECT 3.455000  1.255000 3.705000 1.270000 ;
      RECT 3.790000  2.290000 5.850000 2.460000 ;
      RECT 3.790000  2.460000 4.040000 2.980000 ;
      RECT 4.240000  2.630000 5.480000 2.980000 ;
      RECT 4.375000  0.085000 4.545000 0.915000 ;
      RECT 4.725000  0.580000 4.975000 1.085000 ;
      RECT 5.155000  0.085000 5.485000 0.915000 ;
      RECT 5.665000  0.580000 5.845000 1.080000 ;
      RECT 5.665000  1.080000 7.635000 1.085000 ;
      RECT 5.680000  1.820000 5.850000 1.950000 ;
      RECT 5.680000  1.950000 7.870000 2.120000 ;
      RECT 5.680000  2.120000 5.850000 2.290000 ;
      RECT 5.680000  2.460000 5.850000 2.980000 ;
      RECT 6.025000  0.085000 6.275000 0.910000 ;
      RECT 6.050000  2.290000 7.370000 2.460000 ;
      RECT 6.050000  2.460000 6.380000 2.980000 ;
      RECT 6.455000  0.580000 6.705000 1.080000 ;
      RECT 6.580000  2.650000 6.870000 3.245000 ;
      RECT 6.885000  0.085000 7.135000 0.910000 ;
      RECT 7.040000  2.460000 7.370000 2.980000 ;
      RECT 7.385000  0.675000 7.635000 1.080000 ;
      RECT 7.385000  1.250000 7.635000 1.275000 ;
      RECT 7.540000  1.820000 7.870000 1.950000 ;
      RECT 7.540000  2.120000 7.870000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_hs__o41a_4
MACRO sky130_fd_sc_hs__o41ai_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.810000 1.350000 3.235000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.920000 2.295000 2.890000 ;
        RECT 2.125000 1.350000 2.525000 1.680000 ;
        RECT 2.125000 1.680000 2.295000 1.920000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.350000 1.955000 1.680000 ;
        RECT 1.565000 1.680000 1.795000 2.890000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055000 1.350000 1.385000 1.780000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.435000 1.550000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.602900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.350000 0.775000 1.010000 ;
        RECT 0.605000 1.010000 0.775000 1.350000 ;
        RECT 0.605000 1.350000 0.885000 1.520000 ;
        RECT 0.715000 1.520000 0.885000 1.950000 ;
        RECT 0.715000 1.950000 1.165000 2.120000 ;
        RECT 0.835000 2.120000 1.165000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.115000  1.820000 0.545000 2.650000 ;
      RECT 0.115000  2.650000 0.665000 3.245000 ;
      RECT 0.955000  0.350000 1.205000 1.010000 ;
      RECT 0.955000  1.010000 3.220000 1.180000 ;
      RECT 1.375000  0.085000 1.705000 0.840000 ;
      RECT 1.890000  0.350000 2.220000 1.010000 ;
      RECT 2.390000  0.085000 2.720000 0.840000 ;
      RECT 2.890000  0.350000 3.220000 1.010000 ;
      RECT 2.995000  1.950000 3.245000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__o41ai_1
MACRO sky130_fd_sc_hs__o41ai_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.350000 1.350000 6.115000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.765000 1.350000 5.155000 1.680000 ;
        RECT 4.925000 1.680000 5.155000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.350000 3.455000 1.780000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405000 1.350000 2.755000 1.780000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.280000 0.455000 1.180000 ;
        RECT 0.125000 1.180000 0.900000 1.550000 ;
        RECT 0.125000 1.550000 0.455000 1.630000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.879200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.635000 1.720000 2.235000 1.890000 ;
        RECT 0.635000 1.890000 0.805000 2.980000 ;
        RECT 1.070000 0.645000 1.400000 1.550000 ;
        RECT 1.070000 1.550000 2.235000 1.720000 ;
        RECT 2.035000 1.890000 2.235000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.240000 0.085000 ;
      RECT 0.000000  3.245000 6.240000 3.415000 ;
      RECT 0.105000  1.820000 0.435000 3.245000 ;
      RECT 0.640000  0.255000 1.900000 0.425000 ;
      RECT 0.640000  0.425000 0.890000 1.010000 ;
      RECT 1.005000  2.060000 1.335000 3.245000 ;
      RECT 1.535000  2.060000 1.865000 2.905000 ;
      RECT 1.535000  2.905000 2.765000 3.075000 ;
      RECT 1.570000  0.425000 1.900000 1.010000 ;
      RECT 1.570000  1.010000 5.790000 1.180000 ;
      RECT 2.070000  0.085000 2.400000 0.795000 ;
      RECT 2.435000  1.950000 3.800000 2.120000 ;
      RECT 2.435000  2.120000 2.765000 2.905000 ;
      RECT 2.580000  0.350000 2.830000 1.010000 ;
      RECT 3.000000  0.085000 3.330000 0.795000 ;
      RECT 3.020000  2.290000 3.270000 2.905000 ;
      RECT 3.020000  2.905000 4.705000 3.075000 ;
      RECT 3.470000  2.120000 3.800000 2.735000 ;
      RECT 3.510000  0.350000 3.790000 1.010000 ;
      RECT 3.960000  0.085000 4.290000 0.795000 ;
      RECT 4.005000  1.850000 4.335000 1.950000 ;
      RECT 4.005000  1.950000 6.135000 2.120000 ;
      RECT 4.005000  2.120000 4.335000 2.735000 ;
      RECT 4.460000  0.350000 4.790000 1.010000 ;
      RECT 4.535000  2.290000 4.705000 2.905000 ;
      RECT 4.905000  2.120000 5.235000 2.980000 ;
      RECT 4.960000  0.085000 5.290000 0.795000 ;
      RECT 5.435000  2.290000 5.605000 3.245000 ;
      RECT 5.460000  0.350000 5.790000 1.010000 ;
      RECT 5.805000  2.120000 6.135000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
  END
END sky130_fd_sc_hs__o41ai_2
MACRO sky130_fd_sc_hs__o41ai_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAPARTIALMETALSIDEAREA  0.136000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.285000 1.180000 9.955000 1.550000 ;
    END
  END A1
  PIN A2
    ANTENNAPARTIALMETALSIDEAREA  0.136000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365000 1.180000 8.035000 1.550000 ;
    END
  END A2
  PIN A3
    ANTENNAPARTIALMETALSIDEAREA  0.146000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.395000 1.180000 6.115000 1.550000 ;
    END
  END A3
  PIN A4
    ANTENNAPARTIALMETALSIDEAREA  0.161000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.180000 3.160000 1.550000 ;
    END
  END A4
  PIN B1
    ANTENNAPARTIALMETALSIDEAREA  0.142000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 1.145000 1.550000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.586200 ;
    ANTENNAPARTIALMETALSIDEAREA  1.389000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.615000 1.720000 3.330000 1.890000 ;
        RECT 0.615000 1.890000 0.945000 2.980000 ;
        RECT 0.625000 0.595000 0.795000 0.840000 ;
        RECT 0.625000 0.840000 1.805000 1.010000 ;
        RECT 1.475000 0.595000 1.805000 0.840000 ;
        RECT 1.475000 1.010000 1.805000 1.720000 ;
        RECT 2.150000 1.890000 3.330000 2.150000 ;
        RECT 2.150000 2.150000 2.430000 2.735000 ;
        RECT 3.050000 2.150000 3.330000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.115000  0.255000  2.305000 0.425000 ;
      RECT 0.115000  0.425000  0.445000 1.010000 ;
      RECT 0.115000  1.820000  0.445000 3.245000 ;
      RECT 0.975000  0.425000  1.305000 0.670000 ;
      RECT 1.115000  2.060000  1.445000 3.245000 ;
      RECT 1.675000  2.060000  1.980000 2.905000 ;
      RECT 1.675000  2.905000  5.705000 3.075000 ;
      RECT 1.975000  0.425000  2.305000 0.840000 ;
      RECT 1.975000  0.840000  3.500000 1.010000 ;
      RECT 2.475000  0.085000  2.990000 0.600000 ;
      RECT 2.600000  2.320000  2.880000 2.905000 ;
      RECT 3.160000  0.350000  3.500000 0.840000 ;
      RECT 3.330000  1.010000  3.500000 1.300000 ;
      RECT 3.330000  1.300000  4.190000 1.470000 ;
      RECT 3.500000  1.800000  3.805000 2.905000 ;
      RECT 3.670000  0.085000  3.840000 1.130000 ;
      RECT 3.975000  1.720000  7.565000 1.890000 ;
      RECT 3.975000  1.890000  4.305000 2.735000 ;
      RECT 4.020000  0.350000  4.350000 0.840000 ;
      RECT 4.020000  0.840000  9.965000 1.010000 ;
      RECT 4.020000  1.010000  4.190000 1.300000 ;
      RECT 4.475000  2.060000  4.805000 2.905000 ;
      RECT 4.520000  0.085000  4.850000 0.670000 ;
      RECT 4.975000  1.890000  5.205000 2.735000 ;
      RECT 5.030000  0.350000  5.280000 0.840000 ;
      RECT 5.375000  2.060000  5.705000 2.905000 ;
      RECT 5.450000  0.085000  5.780000 0.670000 ;
      RECT 5.935000  2.060000  6.265000 2.890000 ;
      RECT 5.935000  2.890000  7.165000 2.905000 ;
      RECT 5.935000  2.905000  8.015000 3.075000 ;
      RECT 5.960000  0.350000  6.210000 0.840000 ;
      RECT 6.380000  0.085000  6.710000 0.670000 ;
      RECT 6.435000  1.890000  6.665000 2.720000 ;
      RECT 6.835000  2.060000  7.165000 2.890000 ;
      RECT 6.890000  0.350000  7.060000 0.840000 ;
      RECT 7.240000  0.085000  7.570000 0.670000 ;
      RECT 7.335000  1.890000  7.565000 2.735000 ;
      RECT 7.735000  1.720000  9.965000 1.890000 ;
      RECT 7.735000  1.890000  8.015000 2.905000 ;
      RECT 7.785000  0.350000  8.035000 0.840000 ;
      RECT 8.185000  2.060000  8.515000 3.245000 ;
      RECT 8.205000  0.085000  8.535000 0.670000 ;
      RECT 8.685000  1.890000  9.015000 3.000000 ;
      RECT 8.705000  0.350000  9.035000 0.840000 ;
      RECT 9.185000  2.060000  9.515000 3.245000 ;
      RECT 9.205000  0.085000  9.535000 0.670000 ;
      RECT 9.685000  1.890000  9.965000 3.000000 ;
      RECT 9.715000  0.350000  9.965000 0.840000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
  END
END sky130_fd_sc_hs__o41ai_4
MACRO sky130_fd_sc_hs__or2_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.400000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045000 1.350000 1.375000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.775000 1.550000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.955000 0.350000 2.310000 1.130000 ;
        RECT 1.955000 1.820000 2.310000 2.980000 ;
        RECT 2.140000 1.130000 2.310000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.400000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.400000 0.085000 ;
      RECT 0.000000  3.245000 2.400000 3.415000 ;
      RECT 0.295000  0.085000 0.650000 0.995000 ;
      RECT 0.295000  1.820000 0.625000 1.950000 ;
      RECT 0.295000  1.950000 1.785000 2.120000 ;
      RECT 0.295000  2.120000 0.625000 2.700000 ;
      RECT 0.945000  0.540000 1.240000 1.010000 ;
      RECT 0.945000  1.010000 1.785000 1.180000 ;
      RECT 1.165000  2.290000 1.785000 3.245000 ;
      RECT 1.455000  0.085000 1.785000 0.840000 ;
      RECT 1.615000  1.180000 1.785000 1.300000 ;
      RECT 1.615000  1.300000 1.970000 1.630000 ;
      RECT 1.615000  1.630000 1.785000 1.950000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
  END
END sky130_fd_sc_hs__or2_1
MACRO sky130_fd_sc_hs__or2_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.400000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.350000 1.045000 2.150000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.435000 1.550000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.565600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.555000 0.350000 1.795000 1.820000 ;
        RECT 1.555000 1.820000 1.835000 2.150000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.400000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.400000 0.085000 ;
      RECT 0.000000  3.245000 2.400000 3.415000 ;
      RECT 0.105000  1.820000 0.435000 2.320000 ;
      RECT 0.105000  2.320000 2.295000 2.490000 ;
      RECT 0.105000  2.490000 0.435000 2.860000 ;
      RECT 0.110000  0.085000 0.440000 1.000000 ;
      RECT 0.620000  0.450000 0.870000 1.010000 ;
      RECT 0.620000  1.010000 1.385000 1.180000 ;
      RECT 1.035000  2.660000 1.365000 3.245000 ;
      RECT 1.045000  0.085000 1.375000 0.825000 ;
      RECT 1.215000  1.180000 1.385000 2.320000 ;
      RECT 1.955000  2.660000 2.285000 3.245000 ;
      RECT 1.965000  1.300000 2.295000 1.630000 ;
      RECT 1.970000  0.085000 2.300000 1.130000 ;
      RECT 2.125000  1.630000 2.295000 2.320000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
  END
END sky130_fd_sc_hs__or2_2
MACRO sky130_fd_sc_hs__or2_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.210000 1.350000 2.755000 1.950000 ;
        RECT 2.520000 1.950000 3.895000 2.120000 ;
        RECT 3.590000 1.450000 3.895000 1.950000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925000 1.450000 3.255000 1.780000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  1.149300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.960000 1.700000 1.130000 ;
        RECT 0.125000 1.130000 0.355000 1.800000 ;
        RECT 0.125000 1.800000 1.795000 1.970000 ;
        RECT 0.545000 0.350000 0.795000 0.960000 ;
        RECT 0.565000 1.970000 0.895000 2.980000 ;
        RECT 1.405000 0.350000 1.700000 0.960000 ;
        RECT 1.465000 1.970000 1.795000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  0.085000 0.365000 0.790000 ;
      RECT 0.115000  2.140000 0.365000 3.245000 ;
      RECT 0.595000  1.300000 2.040000 1.630000 ;
      RECT 0.975000  0.085000 1.225000 0.790000 ;
      RECT 1.095000  2.140000 1.265000 3.245000 ;
      RECT 1.870000  1.010000 4.235000 1.180000 ;
      RECT 1.870000  1.180000 2.040000 1.300000 ;
      RECT 1.920000  0.085000 2.250000 0.840000 ;
      RECT 1.995000  2.120000 2.245000 3.245000 ;
      RECT 2.420000  0.350000 2.750000 1.010000 ;
      RECT 2.450000  2.290000 2.780000 2.905000 ;
      RECT 2.450000  2.905000 3.730000 3.075000 ;
      RECT 2.920000  0.085000 4.205000 0.840000 ;
      RECT 2.980000  2.290000 4.235000 2.460000 ;
      RECT 2.980000  2.460000 3.230000 2.735000 ;
      RECT 3.400000  2.630000 3.730000 2.905000 ;
      RECT 3.930000  2.630000 4.205000 3.245000 ;
      RECT 4.065000  1.180000 4.235000 2.290000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__or2_4
MACRO sky130_fd_sc_hs__or2b_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.233000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.035000 1.350000 2.365000 1.780000 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 0.455000 1.550000 ;
    END
  END B_N
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.755000 1.820000 3.275000 2.980000 ;
        RECT 2.875000 0.350000 3.275000 1.130000 ;
        RECT 3.105000 1.130000 3.275000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.115000  0.680000 0.830000 1.010000 ;
      RECT 0.115000  1.760000 0.830000 1.930000 ;
      RECT 0.115000  1.930000 0.445000 2.980000 ;
      RECT 0.615000  2.100000 0.945000 3.245000 ;
      RECT 0.660000  1.010000 0.830000 1.300000 ;
      RECT 0.660000  1.300000 1.525000 1.630000 ;
      RECT 0.660000  1.630000 0.830000 1.760000 ;
      RECT 1.000000  0.085000 1.525000 1.130000 ;
      RECT 1.300000  1.820000 1.865000 1.990000 ;
      RECT 1.300000  1.990000 1.630000 2.860000 ;
      RECT 1.695000  0.540000 2.045000 1.010000 ;
      RECT 1.695000  1.010000 2.705000 1.180000 ;
      RECT 1.695000  1.180000 1.865000 1.820000 ;
      RECT 2.255000  1.950000 2.585000 3.245000 ;
      RECT 2.265000  0.085000 2.680000 0.840000 ;
      RECT 2.535000  1.180000 2.705000 1.300000 ;
      RECT 2.535000  1.300000 2.935000 1.630000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__or2b_1
MACRO sky130_fd_sc_hs__or2b_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.035000 1.350000 2.365000 1.780000 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 0.550000 1.780000 ;
    END
  END B_N
  PIN X
    ANTENNADIFFAREA  0.787700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.060000 0.350000 1.390000 1.130000 ;
        RECT 1.060000 1.130000 1.230000 1.820000 ;
        RECT 1.060000 1.820000 1.645000 2.070000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.115000  1.950000 0.890000 2.240000 ;
      RECT 0.115000  2.240000 2.705000 2.410000 ;
      RECT 0.115000  2.410000 0.445000 2.700000 ;
      RECT 0.120000  0.540000 0.450000 1.010000 ;
      RECT 0.120000  1.010000 0.890000 1.180000 ;
      RECT 0.630000  0.085000 0.880000 0.840000 ;
      RECT 0.650000  2.580000 0.980000 3.245000 ;
      RECT 0.720000  1.180000 0.890000 1.950000 ;
      RECT 1.465000  1.300000 1.795000 1.630000 ;
      RECT 1.560000  0.085000 2.235000 0.810000 ;
      RECT 1.625000  0.980000 3.275000 1.150000 ;
      RECT 1.625000  1.150000 1.795000 1.300000 ;
      RECT 1.765000  2.580000 2.095000 3.245000 ;
      RECT 2.405000  0.350000 2.735000 0.980000 ;
      RECT 2.535000  1.320000 2.935000 1.650000 ;
      RECT 2.535000  1.650000 2.705000 2.240000 ;
      RECT 2.875000  1.820000 3.275000 2.860000 ;
      RECT 2.915000  0.085000 3.245000 0.810000 ;
      RECT 3.105000  1.150000 3.275000 1.820000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__or2b_2
MACRO sky130_fd_sc_hs__or2b_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.450000 3.235000 1.780000 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.905000 1.120000 5.235000 1.790000 ;
    END
  END B_N
  PIN X
    ANTENNADIFFAREA  1.104900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 0.775000 1.410000 ;
        RECT 0.545000 0.350000 0.795000 0.960000 ;
        RECT 0.545000 0.960000 1.805000 1.130000 ;
        RECT 0.545000 1.130000 0.775000 1.180000 ;
        RECT 0.605000 1.410000 0.775000 1.800000 ;
        RECT 0.605000 1.800000 1.785000 1.970000 ;
        RECT 0.605000 1.970000 0.805000 2.980000 ;
        RECT 1.455000 1.970000 1.785000 2.980000 ;
        RECT 1.475000 0.350000 1.805000 0.960000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.105000  1.820000 0.435000 3.245000 ;
      RECT 0.115000  0.085000 0.365000 1.010000 ;
      RECT 0.945000  1.300000 2.145000 1.630000 ;
      RECT 0.975000  0.085000 1.305000 0.765000 ;
      RECT 1.005000  2.140000 1.255000 3.245000 ;
      RECT 1.975000  0.085000 2.305000 0.940000 ;
      RECT 1.975000  1.110000 3.755000 1.280000 ;
      RECT 1.975000  1.280000 2.145000 1.300000 ;
      RECT 1.985000  1.940000 2.235000 3.245000 ;
      RECT 2.430000  1.950000 3.675000 2.120000 ;
      RECT 2.430000  2.120000 2.760000 2.980000 ;
      RECT 2.475000  0.350000 2.805000 1.110000 ;
      RECT 2.960000  2.290000 3.210000 3.245000 ;
      RECT 3.005000  0.085000 3.335000 0.940000 ;
      RECT 3.425000  1.915000 3.675000 1.950000 ;
      RECT 3.425000  2.120000 3.675000 2.905000 ;
      RECT 3.425000  2.905000 4.655000 3.075000 ;
      RECT 3.505000  0.350000 3.755000 1.110000 ;
      RECT 3.505000  1.280000 4.125000 1.450000 ;
      RECT 3.875000  1.450000 4.125000 2.735000 ;
      RECT 3.935000  0.085000 4.265000 1.030000 ;
      RECT 4.295000  1.445000 4.625000 1.775000 ;
      RECT 4.325000  1.945000 4.655000 2.905000 ;
      RECT 4.435000  0.350000 5.655000 0.950000 ;
      RECT 4.435000  0.950000 4.625000 1.445000 ;
      RECT 4.875000  1.960000 5.205000 3.245000 ;
      RECT 5.405000  0.950000 5.655000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_hs__or2b_4
MACRO sky130_fd_sc_hs__or3_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.880000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.233000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 1.350000 1.815000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.233000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.835000 1.350000 1.315000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.233000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 0.570000 1.780000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.430000 0.350000 2.795000 1.130000 ;
        RECT 2.515000 1.820000 2.795000 2.980000 ;
        RECT 2.625000 1.130000 2.795000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.880000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.880000 0.085000 ;
      RECT 0.000000  3.245000 2.880000 3.415000 ;
      RECT 0.115000  0.350000 0.365000 1.010000 ;
      RECT 0.115000  1.010000 2.260000 1.180000 ;
      RECT 0.115000  1.950000 2.260000 2.120000 ;
      RECT 0.115000  2.120000 0.445000 2.860000 ;
      RECT 0.545000  0.085000 0.875000 0.810000 ;
      RECT 1.045000  0.455000 1.760000 1.010000 ;
      RECT 1.555000  2.290000 2.315000 3.245000 ;
      RECT 1.930000  0.085000 2.260000 0.810000 ;
      RECT 2.090000  1.180000 2.260000 1.300000 ;
      RECT 2.090000  1.300000 2.455000 1.630000 ;
      RECT 2.090000  1.630000 2.260000 1.950000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
  END
END sky130_fd_sc_hs__or3_1
MACRO sky130_fd_sc_hs__or3_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.180000 1.905000 1.550000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.130000 1.335000 2.890000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.435000 1.120000 0.835000 1.790000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.335000 1.800000 3.235000 1.970000 ;
        RECT 2.335000 1.970000 2.665000 2.980000 ;
        RECT 2.415000 0.350000 2.745000 0.960000 ;
        RECT 2.415000 0.960000 3.235000 1.130000 ;
        RECT 3.005000 1.130000 3.235000 1.800000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.095000  0.350000 0.445000 0.780000 ;
      RECT 0.095000  0.780000 1.530000 0.790000 ;
      RECT 0.095000  0.790000 2.245000 0.950000 ;
      RECT 0.095000  0.950000 0.265000 1.960000 ;
      RECT 0.095000  1.960000 0.615000 2.130000 ;
      RECT 0.285000  2.130000 0.615000 2.980000 ;
      RECT 0.615000  0.085000 1.030000 0.600000 ;
      RECT 1.200000  0.350000 1.530000 0.780000 ;
      RECT 1.200000  0.950000 2.245000 0.960000 ;
      RECT 1.700000  0.085000 2.245000 0.600000 ;
      RECT 1.725000  1.940000 2.055000 3.245000 ;
      RECT 2.075000  0.960000 2.245000 1.300000 ;
      RECT 2.075000  1.300000 2.815000 1.630000 ;
      RECT 2.835000  2.140000 3.165000 3.245000 ;
      RECT 2.915000  0.085000 3.245000 0.790000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__or3_2
MACRO sky130_fd_sc_hs__or3_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.280000 0.435000 1.110000 ;
        RECT 0.105000 1.110000 3.055000 1.280000 ;
        RECT 0.105000 1.280000 0.435000 1.630000 ;
        RECT 2.755000 1.280000 3.055000 1.550000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.450000 2.545000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.050000 0.270000 1.380000 0.940000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  1.090100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.565000 0.350000 3.735000 0.960000 ;
        RECT 3.565000 0.960000 5.155000 1.130000 ;
        RECT 3.565000 1.800000 5.155000 1.970000 ;
        RECT 3.565000 1.970000 3.735000 2.980000 ;
        RECT 4.385000 1.970000 4.715000 2.980000 ;
        RECT 4.405000 0.350000 4.655000 0.960000 ;
        RECT 4.925000 1.130000 5.155000 1.800000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.280000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.245000 5.280000 3.415000 ;
      RECT 0.115000  1.920000 0.365000 3.245000 ;
      RECT 0.565000  1.950000 0.815000 2.370000 ;
      RECT 0.565000  2.370000 2.830000 2.540000 ;
      RECT 0.565000  2.540000 0.815000 2.960000 ;
      RECT 1.015000  2.710000 2.330000 2.960000 ;
      RECT 1.495000  1.950000 3.395000 2.120000 ;
      RECT 1.495000  2.120000 1.825000 2.200000 ;
      RECT 1.550000  0.350000 1.880000 0.770000 ;
      RECT 1.550000  0.770000 3.395000 0.940000 ;
      RECT 2.050000  0.085000 2.380000 0.600000 ;
      RECT 2.500000  2.290000 2.830000 2.370000 ;
      RECT 2.500000  2.540000 2.830000 2.960000 ;
      RECT 2.550000  0.350000 2.880000 0.770000 ;
      RECT 3.035000  2.290000 3.365000 3.245000 ;
      RECT 3.050000  0.085000 3.380000 0.600000 ;
      RECT 3.225000  0.940000 3.395000 1.300000 ;
      RECT 3.225000  1.300000 4.685000 1.630000 ;
      RECT 3.225000  1.630000 3.395000 1.950000 ;
      RECT 3.915000  0.085000 4.165000 0.790000 ;
      RECT 3.935000  2.140000 4.185000 3.245000 ;
      RECT 4.835000  0.085000 5.165000 0.790000 ;
      RECT 4.915000  2.140000 5.165000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
  END
END sky130_fd_sc_hs__or3_4
MACRO sky130_fd_sc_hs__or3b_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.233000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.515000 1.300000 2.845000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.233000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.915000 1.190000 2.275000 2.890000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.110000 0.605000 1.780000 ;
    END
  END C_N
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.250000 1.820000 3.755000 2.980000 ;
        RECT 3.395000 0.350000 3.755000 1.130000 ;
        RECT 3.585000 1.130000 3.755000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 0.940000 ;
      RECT 0.115000  2.100000 0.445000 3.245000 ;
      RECT 0.615000  0.350000 0.945000 0.940000 ;
      RECT 0.615000  2.100000 0.945000 2.980000 ;
      RECT 0.775000  0.940000 0.945000 1.210000 ;
      RECT 0.775000  1.210000 1.205000 1.880000 ;
      RECT 0.775000  1.880000 0.945000 2.100000 ;
      RECT 1.175000  0.350000 1.505000 0.850000 ;
      RECT 1.175000  0.850000 3.225000 1.020000 ;
      RECT 1.375000  1.020000 1.705000 2.975000 ;
      RECT 1.675000  0.085000 2.005000 0.680000 ;
      RECT 2.175000  0.350000 2.505000 0.850000 ;
      RECT 2.675000  0.085000 3.225000 0.680000 ;
      RECT 2.750000  1.950000 3.080000 3.245000 ;
      RECT 3.055000  1.020000 3.225000 1.300000 ;
      RECT 3.055000  1.300000 3.415000 1.630000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__or3b_1
MACRO sky130_fd_sc_hs__or3b_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975000 1.350000 2.305000 2.150000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.515000 1.350000 2.845000 1.780000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.300000 0.435000 1.780000 ;
    END
  END C_N
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 0.960000 1.455000 1.130000 ;
        RECT 1.065000 1.130000 1.235000 1.820000 ;
        RECT 1.065000 1.820000 1.795000 2.150000 ;
        RECT 1.125000 0.350000 1.455000 0.960000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.115000  1.950000 0.775000 2.320000 ;
      RECT 0.115000  2.320000 2.645000 2.490000 ;
      RECT 0.115000  2.490000 0.445000 2.700000 ;
      RECT 0.185000  0.540000 0.605000 0.960000 ;
      RECT 0.185000  0.960000 0.775000 1.130000 ;
      RECT 0.605000  1.130000 0.775000 1.950000 ;
      RECT 0.650000  2.660000 0.980000 3.245000 ;
      RECT 0.775000  0.085000 0.945000 0.790000 ;
      RECT 1.405000  1.300000 1.795000 1.630000 ;
      RECT 1.625000  0.085000 2.135000 0.780000 ;
      RECT 1.625000  1.010000 3.755000 1.180000 ;
      RECT 1.625000  1.180000 1.795000 1.300000 ;
      RECT 1.635000  2.660000 2.070000 3.245000 ;
      RECT 2.350000  0.450000 2.680000 1.010000 ;
      RECT 2.475000  1.950000 3.415000 2.120000 ;
      RECT 2.475000  2.120000 2.645000 2.320000 ;
      RECT 2.850000  0.085000 3.180000 0.840000 ;
      RECT 3.085000  1.350000 3.415000 1.950000 ;
      RECT 3.235000  2.290000 3.755000 2.860000 ;
      RECT 3.350000  0.450000 3.755000 1.010000 ;
      RECT 3.585000  1.180000 3.755000 2.290000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__or3b_2
MACRO sky130_fd_sc_hs__or3b_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.800000 1.150000 3.545000 1.320000 ;
        RECT 0.800000 1.320000 1.130000 1.760000 ;
        RECT 3.005000 1.320000 3.545000 1.380000 ;
        RECT 3.285000 1.380000 3.545000 1.550000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.340000 1.490000 1.670000 1.550000 ;
        RECT 1.340000 1.550000 3.075000 1.800000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.255000 0.775000 0.640000 ;
    END
  END C_N
  PIN X
    ANTENNADIFFAREA  1.104900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.055000 0.350000 4.225000 0.960000 ;
        RECT 4.055000 0.960000 5.635000 1.130000 ;
        RECT 4.055000 1.800000 5.635000 1.970000 ;
        RECT 4.055000 1.970000 4.225000 2.980000 ;
        RECT 4.875000 1.970000 5.205000 2.980000 ;
        RECT 4.885000 0.350000 5.135000 0.960000 ;
        RECT 5.405000 1.130000 5.635000 1.800000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.110000  0.810000 1.910000 0.980000 ;
      RECT 0.110000  0.980000 0.465000 1.340000 ;
      RECT 0.110000  1.340000 0.360000 2.980000 ;
      RECT 0.560000  1.940000 0.890000 3.245000 ;
      RECT 0.945000  0.085000 1.410000 0.640000 ;
      RECT 1.070000  1.970000 1.400000 2.360000 ;
      RECT 1.070000  2.360000 3.335000 2.530000 ;
      RECT 1.070000  2.530000 1.400000 2.980000 ;
      RECT 1.580000  0.310000 1.910000 0.810000 ;
      RECT 1.580000  2.700000 2.835000 2.980000 ;
      RECT 2.030000  1.970000 3.885000 2.140000 ;
      RECT 2.030000  2.140000 2.385000 2.190000 ;
      RECT 2.080000  0.350000 2.410000 0.810000 ;
      RECT 2.080000  0.810000 3.885000 0.980000 ;
      RECT 2.580000  0.085000 2.910000 0.640000 ;
      RECT 3.005000  2.310000 3.335000 2.360000 ;
      RECT 3.005000  2.530000 3.335000 2.980000 ;
      RECT 3.090000  0.350000 3.340000 0.810000 ;
      RECT 3.505000  2.310000 3.835000 3.245000 ;
      RECT 3.510000  0.085000 3.850000 0.600000 ;
      RECT 3.715000  0.980000 3.885000 1.300000 ;
      RECT 3.715000  1.300000 5.175000 1.630000 ;
      RECT 3.715000  1.630000 3.885000 1.970000 ;
      RECT 4.405000  0.085000 4.655000 0.790000 ;
      RECT 4.425000  2.140000 4.675000 3.245000 ;
      RECT 5.315000  0.085000 5.645000 0.790000 ;
      RECT 5.405000  2.140000 5.655000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_hs__or3b_4
MACRO sky130_fd_sc_hs__or4_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.233000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.350000 2.390000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.233000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.490000 1.420000 1.820000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.233000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.920000 1.420000 1.295000 1.780000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.233000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.420000 0.650000 1.780000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.900000 1.820000 3.275000 2.980000 ;
        RECT 2.960000 0.350000 3.275000 1.130000 ;
        RECT 3.105000 1.130000 3.275000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 1.130000 ;
      RECT 0.200000  1.950000 2.730000 2.120000 ;
      RECT 0.200000  2.120000 0.530000 2.980000 ;
      RECT 0.615000  0.540000 0.945000 1.010000 ;
      RECT 0.615000  1.010000 2.730000 1.180000 ;
      RECT 1.125000  0.085000 1.600000 0.840000 ;
      RECT 1.860000  0.540000 2.190000 1.010000 ;
      RECT 2.150000  2.290000 2.565000 3.245000 ;
      RECT 2.450000  0.085000 2.780000 0.840000 ;
      RECT 2.560000  1.180000 2.730000 1.300000 ;
      RECT 2.560000  1.300000 2.935000 1.630000 ;
      RECT 2.560000  1.630000 2.730000 1.950000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__or4_1
MACRO sky130_fd_sc_hs__or4_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.350000 2.455000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.545000 1.350000 1.875000 2.890000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.165000 1.335000 2.890000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.180000 0.835000 1.770000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.860000 1.800000 3.715000 1.970000 ;
        RECT 2.860000 1.970000 3.190000 2.980000 ;
        RECT 2.965000 0.350000 3.215000 0.960000 ;
        RECT 2.965000 0.960000 3.715000 1.130000 ;
        RECT 3.485000 1.130000 3.715000 1.800000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.085000  0.825000 2.190000 0.995000 ;
      RECT 0.085000  0.995000 0.255000 1.940000 ;
      RECT 0.085000  1.940000 0.735000 2.110000 ;
      RECT 0.115000  0.085000 0.510000 0.655000 ;
      RECT 0.405000  2.110000 0.735000 2.980000 ;
      RECT 0.690000  0.350000 1.020000 0.825000 ;
      RECT 1.200000  0.085000 1.680000 0.655000 ;
      RECT 1.860000  0.350000 2.190000 0.825000 ;
      RECT 1.860000  0.995000 2.190000 1.010000 ;
      RECT 1.860000  1.010000 2.795000 1.180000 ;
      RECT 2.360000  0.085000 2.795000 0.825000 ;
      RECT 2.360000  1.950000 2.690000 3.245000 ;
      RECT 2.625000  1.180000 2.795000 1.300000 ;
      RECT 2.625000  1.300000 3.040000 1.630000 ;
      RECT 3.360000  2.140000 3.690000 3.245000 ;
      RECT 3.395000  0.085000 3.725000 0.775000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__or4_2
MACRO sky130_fd_sc_hs__or4_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405000 1.470000 3.735000 1.800000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.130000 4.395000 1.300000 ;
        RECT 2.525000 1.300000 3.235000 1.410000 ;
        RECT 2.615000 1.410000 3.235000 1.550000 ;
        RECT 4.065000 1.300000 4.395000 1.550000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.605000 1.365000 6.285000 1.770000 ;
        RECT 4.925000 1.770000 6.285000 1.780000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.285000 0.255000 6.615000 0.855000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  1.326900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.945000 1.820000 ;
        RECT 0.125000 1.820000 2.275000 2.150000 ;
        RECT 0.615000 0.350000 0.945000 0.980000 ;
        RECT 0.615000 0.980000 1.945000 1.150000 ;
        RECT 0.615000 1.150000 0.945000 1.300000 ;
        RECT 0.615000 2.150000 0.845000 2.980000 ;
        RECT 1.515000 2.150000 1.745000 2.980000 ;
        RECT 1.615000 0.350000 1.945000 0.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.720000 0.085000 ;
      RECT 0.000000  3.245000 6.720000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 1.130000 ;
      RECT 0.115000  2.320000 0.445000 3.245000 ;
      RECT 1.015000  2.320000 1.345000 3.245000 ;
      RECT 1.115000  0.085000 1.445000 0.810000 ;
      RECT 1.315000  1.320000 2.325000 1.650000 ;
      RECT 1.915000  2.320000 2.245000 3.245000 ;
      RECT 2.155000  0.790000 5.100000 0.960000 ;
      RECT 2.155000  0.960000 2.325000 1.320000 ;
      RECT 2.380000  0.085000 2.740000 0.620000 ;
      RECT 2.475000  1.940000 2.805000 1.970000 ;
      RECT 2.475000  1.970000 4.675000 2.140000 ;
      RECT 2.475000  2.140000 2.805000 2.190000 ;
      RECT 2.475000  2.190000 2.755000 2.980000 ;
      RECT 2.920000  0.350000 3.250000 0.790000 ;
      RECT 2.925000  2.360000 4.175000 2.560000 ;
      RECT 2.925000  2.560000 3.205000 2.980000 ;
      RECT 3.375000  2.730000 3.705000 3.245000 ;
      RECT 3.430000  0.085000 4.590000 0.620000 ;
      RECT 3.825000  2.310000 4.175000 2.360000 ;
      RECT 3.895000  2.560000 4.175000 2.980000 ;
      RECT 4.345000  1.940000 4.675000 1.970000 ;
      RECT 4.345000  2.140000 4.675000 2.360000 ;
      RECT 4.345000  2.360000 6.575000 2.530000 ;
      RECT 4.345000  2.530000 4.675000 2.980000 ;
      RECT 4.770000  0.350000 5.100000 0.790000 ;
      RECT 4.770000  0.960000 5.100000 1.025000 ;
      RECT 4.770000  1.025000 6.635000 1.195000 ;
      RECT 4.845000  2.700000 6.075000 2.980000 ;
      RECT 5.270000  0.085000 6.115000 0.680000 ;
      RECT 5.295000  1.950000 6.635000 2.120000 ;
      RECT 5.295000  2.120000 5.625000 2.190000 ;
      RECT 6.245000  2.290000 6.575000 2.360000 ;
      RECT 6.245000  2.530000 6.575000 2.980000 ;
      RECT 6.465000  1.195000 6.635000 1.950000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
  END
END sky130_fd_sc_hs__or4_4
MACRO sky130_fd_sc_hs__or4b_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.233000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.995000 1.350000 3.325000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.233000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.455000 1.180000 2.785000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.233000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.885000 1.045000 2.275000 1.780000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.450000 0.570000 1.780000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.835000 0.350000 4.235000 1.130000 ;
        RECT 3.835000 1.820000 4.235000 2.980000 ;
        RECT 4.065000 1.130000 4.235000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  0.350000 0.445000 1.110000 ;
      RECT 0.115000  1.110000 0.980000 1.280000 ;
      RECT 0.120000  1.950000 0.980000 2.120000 ;
      RECT 0.120000  2.120000 0.450000 2.980000 ;
      RECT 0.615000  0.085000 0.945000 0.940000 ;
      RECT 0.620000  2.290000 0.950000 3.245000 ;
      RECT 0.810000  1.280000 0.980000 1.580000 ;
      RECT 0.810000  1.580000 1.140000 1.910000 ;
      RECT 0.810000  1.910000 0.980000 1.950000 ;
      RECT 1.115000  0.545000 2.090000 0.875000 ;
      RECT 1.315000  0.875000 1.645000 1.950000 ;
      RECT 1.315000  1.950000 3.665000 2.120000 ;
      RECT 1.315000  2.120000 1.645000 2.860000 ;
      RECT 2.260000  0.085000 2.590000 0.875000 ;
      RECT 2.760000  0.350000 3.125000 0.940000 ;
      RECT 2.955000  0.940000 3.125000 1.010000 ;
      RECT 2.955000  1.010000 3.665000 1.180000 ;
      RECT 3.295000  0.085000 3.625000 0.840000 ;
      RECT 3.335000  2.290000 3.665000 3.245000 ;
      RECT 3.495000  1.180000 3.665000 1.300000 ;
      RECT 3.495000  1.300000 3.895000 1.630000 ;
      RECT 3.495000  1.630000 3.665000 1.950000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__or4b_1
MACRO sky130_fd_sc_hs__or4b_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945000 1.350000 2.275000 2.150000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.485000 1.470000 2.815000 2.150000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.470000 3.355000 2.520000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 0.550000 1.780000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.060000 0.350000 1.405000 1.130000 ;
        RECT 1.060000 1.130000 1.230000 1.820000 ;
        RECT 1.060000 1.820000 1.430000 2.150000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  1.950000 0.890000 2.320000 ;
      RECT 0.115000  2.320000 2.465000 2.490000 ;
      RECT 0.115000  2.490000 0.445000 2.700000 ;
      RECT 0.130000  0.540000 0.460000 1.010000 ;
      RECT 0.130000  1.010000 0.890000 1.180000 ;
      RECT 0.640000  0.085000 0.890000 0.840000 ;
      RECT 0.650000  2.660000 0.980000 3.245000 ;
      RECT 0.720000  1.180000 0.890000 1.950000 ;
      RECT 1.400000  1.300000 1.745000 1.630000 ;
      RECT 1.550000  2.730000 2.125000 3.245000 ;
      RECT 1.575000  0.085000 1.995000 0.780000 ;
      RECT 1.575000  0.960000 3.705000 1.100000 ;
      RECT 1.575000  1.100000 4.235000 1.130000 ;
      RECT 1.575000  1.130000 1.745000 1.300000 ;
      RECT 2.175000  0.450000 2.505000 0.960000 ;
      RECT 2.295000  2.490000 2.465000 2.690000 ;
      RECT 2.295000  2.690000 3.695000 2.860000 ;
      RECT 2.685000  0.085000 3.205000 0.780000 ;
      RECT 3.375000  0.450000 3.705000 0.960000 ;
      RECT 3.375000  1.130000 4.235000 1.270000 ;
      RECT 3.525000  1.440000 3.895000 1.770000 ;
      RECT 3.525000  1.770000 3.695000 2.690000 ;
      RECT 3.865000  1.940000 4.235000 2.980000 ;
      RECT 3.875000  0.085000 4.205000 0.930000 ;
      RECT 4.065000  1.270000 4.235000 1.940000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__or4b_2
MACRO sky130_fd_sc_hs__or4b_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.450000 1.335000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.110000 2.035000 1.280000 ;
        RECT 0.125000 1.280000 0.835000 1.550000 ;
        RECT 1.705000 1.280000 2.035000 1.550000 ;
    END
  END B
  PIN C
    ANTENNAPARTIALMETALSIDEAREA  1.197000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2.495000 1.180000 2.785000 1.225000 ;
        RECT 2.495000 1.225000 4.225000 1.365000 ;
        RECT 2.495000 1.365000 2.785000 1.410000 ;
        RECT 3.935000 1.180000 4.225000 1.225000 ;
        RECT 3.935000 1.365000 4.225000 1.410000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.180000 4.815000 1.550000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  1.178900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.325000 0.350000 5.655000 0.980000 ;
        RECT 5.325000 0.980000 6.575000 1.150000 ;
        RECT 5.410000 1.820000 7.075000 2.150000 ;
        RECT 5.410000 2.150000 5.690000 2.980000 ;
        RECT 6.325000 0.350000 6.575000 0.980000 ;
        RECT 6.325000 1.150000 6.575000 1.300000 ;
        RECT 6.325000 1.300000 6.655000 1.470000 ;
        RECT 6.360000 2.150000 6.590000 2.980000 ;
        RECT 6.365000 1.470000 6.655000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.200000 0.085000 ;
      RECT 0.000000  3.245000 7.200000 3.415000 ;
      RECT 0.115000  0.350000 0.445000 0.770000 ;
      RECT 0.115000  0.770000 3.270000 0.840000 ;
      RECT 0.115000  0.840000 5.155000 0.940000 ;
      RECT 0.115000  1.940000 0.445000 1.950000 ;
      RECT 0.115000  1.950000 2.345000 2.120000 ;
      RECT 0.115000  2.120000 0.445000 2.980000 ;
      RECT 0.615000  0.085000 0.945000 0.600000 ;
      RECT 0.645000  2.290000 1.845000 2.460000 ;
      RECT 0.645000  2.460000 0.815000 2.980000 ;
      RECT 1.015000  2.630000 1.345000 3.245000 ;
      RECT 1.115000  0.350000 2.200000 0.770000 ;
      RECT 1.515000  2.460000 1.845000 2.980000 ;
      RECT 2.015000  2.120000 2.345000 2.360000 ;
      RECT 2.015000  2.360000 4.195000 2.530000 ;
      RECT 2.015000  2.530000 2.345000 2.980000 ;
      RECT 2.245000  1.180000 2.725000 1.780000 ;
      RECT 2.370000  0.085000 2.725000 0.600000 ;
      RECT 2.515000  2.700000 3.745000 2.980000 ;
      RECT 2.895000  0.350000 3.270000 0.770000 ;
      RECT 2.895000  0.940000 5.155000 1.010000 ;
      RECT 2.895000  1.010000 3.270000 1.130000 ;
      RECT 2.895000  1.130000 3.065000 2.020000 ;
      RECT 2.895000  2.020000 3.295000 2.190000 ;
      RECT 3.235000  1.470000 3.635000 1.720000 ;
      RECT 3.235000  1.720000 4.755000 1.800000 ;
      RECT 3.440000  0.340000 4.565000 0.670000 ;
      RECT 3.465000  1.800000 4.755000 1.890000 ;
      RECT 3.865000  1.180000 4.195000 1.510000 ;
      RECT 3.945000  2.060000 4.195000 2.360000 ;
      RECT 3.945000  2.530000 4.195000 2.980000 ;
      RECT 4.425000  1.890000 4.755000 2.860000 ;
      RECT 4.825000  0.085000 5.155000 0.670000 ;
      RECT 4.960000  1.820000 5.210000 3.245000 ;
      RECT 4.985000  1.010000 5.155000 1.320000 ;
      RECT 4.985000  1.320000 6.155000 1.650000 ;
      RECT 5.825000  0.085000 6.155000 0.810000 ;
      RECT 5.860000  2.320000 6.190000 3.245000 ;
      RECT 6.755000  0.085000 7.085000 1.130000 ;
      RECT 6.760000  2.320000 7.090000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  1.210000 2.725000 1.380000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  1.210000 4.165000 1.380000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
  END
END sky130_fd_sc_hs__or4b_4
MACRO sky130_fd_sc_hs__or4bb_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.233000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.350000 3.835000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.233000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.965000 1.350000 3.295000 2.890000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.455000 1.780000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965000 1.050000 1.315000 1.720000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.240000 1.820000 4.715000 2.980000 ;
        RECT 4.345000 0.350000 4.715000 1.130000 ;
        RECT 4.545000 1.130000 4.715000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.115000  2.100000 0.795000 2.310000 ;
      RECT 0.115000  2.310000 1.285000 2.480000 ;
      RECT 0.115000  2.480000 0.445000 2.980000 ;
      RECT 0.140000  0.350000 0.470000 0.960000 ;
      RECT 0.140000  0.960000 0.795000 1.130000 ;
      RECT 0.615000  2.650000 0.945000 3.245000 ;
      RECT 0.625000  1.130000 0.795000 2.100000 ;
      RECT 0.640000  0.085000 0.970000 0.790000 ;
      RECT 1.115000  2.480000 1.285000 2.905000 ;
      RECT 1.115000  2.905000 2.755000 3.075000 ;
      RECT 1.140000  0.350000 1.655000 0.880000 ;
      RECT 1.150000  1.890000 1.655000 2.140000 ;
      RECT 1.485000  0.880000 1.655000 1.030000 ;
      RECT 1.485000  1.030000 1.905000 1.700000 ;
      RECT 1.485000  1.700000 1.655000 1.890000 ;
      RECT 1.825000  0.085000 2.075000 0.680000 ;
      RECT 1.845000  1.870000 2.245000 2.735000 ;
      RECT 2.075000  0.850000 3.640000 1.010000 ;
      RECT 2.075000  1.010000 4.175000 1.020000 ;
      RECT 2.075000  1.020000 2.245000 1.870000 ;
      RECT 2.245000  0.350000 2.575000 0.850000 ;
      RECT 2.425000  1.190000 2.755000 2.905000 ;
      RECT 2.745000  0.085000 3.140000 0.680000 ;
      RECT 3.310000  0.350000 3.640000 0.850000 ;
      RECT 3.310000  1.020000 4.175000 1.180000 ;
      RECT 3.740000  1.950000 4.070000 3.245000 ;
      RECT 3.810000  0.085000 4.140000 0.840000 ;
      RECT 4.005000  1.180000 4.175000 1.300000 ;
      RECT 4.005000  1.300000 4.375000 1.630000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_hs__or4bb_1
MACRO sky130_fd_sc_hs__or4bb_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.470000 3.925000 1.800000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.150000 0.255000 3.715000 0.570000 ;
        RECT 3.485000 0.570000 3.715000 0.670000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.435000 1.300000 4.695000 1.780000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 0.550000 1.780000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.060000 0.440000 1.315000 1.180000 ;
        RECT 1.060000 1.180000 1.230000 1.850000 ;
        RECT 1.060000 1.850000 1.390000 2.100000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.105000  2.100000 0.890000 2.270000 ;
      RECT 0.105000  2.270000 2.265000 2.440000 ;
      RECT 0.105000  2.440000 0.435000 2.980000 ;
      RECT 0.120000  0.670000 0.450000 1.010000 ;
      RECT 0.120000  1.010000 0.890000 1.180000 ;
      RECT 0.605000  2.610000 0.935000 3.245000 ;
      RECT 0.630000  0.085000 0.880000 0.840000 ;
      RECT 0.720000  1.180000 0.890000 2.100000 ;
      RECT 1.400000  1.350000 1.730000 1.680000 ;
      RECT 1.510000  2.610000 1.840000 3.245000 ;
      RECT 1.560000  1.130000 3.735000 1.300000 ;
      RECT 1.560000  1.300000 1.730000 1.350000 ;
      RECT 1.575000  0.085000 2.035000 0.910000 ;
      RECT 1.970000  1.470000 2.265000 2.270000 ;
      RECT 2.050000  2.610000 2.605000 2.780000 ;
      RECT 2.050000  2.780000 2.380000 2.980000 ;
      RECT 2.310000  0.580000 2.640000 1.130000 ;
      RECT 2.435000  1.300000 2.605000 2.610000 ;
      RECT 2.775000  1.470000 3.070000 1.970000 ;
      RECT 2.775000  1.970000 4.690000 2.140000 ;
      RECT 2.810000  0.085000 2.980000 0.740000 ;
      RECT 2.810000  0.740000 3.195000 0.960000 ;
      RECT 3.405000  0.840000 3.735000 1.130000 ;
      RECT 3.820000  2.310000 4.150000 3.245000 ;
      RECT 3.925000  0.085000 4.255000 0.790000 ;
      RECT 4.095000  0.960000 4.685000 1.130000 ;
      RECT 4.095000  1.130000 4.265000 1.950000 ;
      RECT 4.095000  1.950000 4.690000 1.970000 ;
      RECT 4.360000  2.140000 4.690000 2.820000 ;
      RECT 4.435000  0.435000 4.685000 0.960000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_hs__or4bb_2
MACRO sky130_fd_sc_hs__or4bb_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.525000 1.180000 8.535000 1.550000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365000 1.450000 7.075000 1.780000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.375000 1.350000 3.715000 1.780000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.350000 0.835000 1.780000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  1.677500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.180000 1.450000 2.050000 ;
        RECT 1.085000 2.050000 2.525000 2.220000 ;
        RECT 1.120000 0.350000 1.450000 0.580000 ;
        RECT 1.120000 0.580000 2.775000 0.750000 ;
        RECT 1.120000 0.750000 1.450000 1.180000 ;
        RECT 2.140000 0.420000 2.775000 0.580000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
      RECT 0.000000  3.245000 8.640000 3.415000 ;
      RECT 0.085000  0.450000 0.445000 1.130000 ;
      RECT 0.085000  1.130000 0.255000 1.950000 ;
      RECT 0.085000  1.950000 0.445000 2.390000 ;
      RECT 0.085000  2.390000 2.865000 2.560000 ;
      RECT 0.085000  2.560000 0.445000 2.860000 ;
      RECT 0.615000  0.085000 0.915000 1.130000 ;
      RECT 0.650000  2.730000 0.995000 3.245000 ;
      RECT 1.565000  2.730000 1.990000 3.245000 ;
      RECT 1.620000  0.920000 4.275000 1.090000 ;
      RECT 1.620000  1.090000 1.790000 1.710000 ;
      RECT 1.620000  1.710000 2.865000 1.880000 ;
      RECT 1.630000  0.085000 1.960000 0.410000 ;
      RECT 1.960000  1.260000 3.205000 1.540000 ;
      RECT 2.695000  1.880000 2.865000 2.390000 ;
      RECT 2.840000  2.730000 3.170000 3.245000 ;
      RECT 2.945000  0.085000 3.275000 0.750000 ;
      RECT 3.035000  1.540000 3.205000 2.290000 ;
      RECT 3.035000  2.290000 4.715000 2.460000 ;
      RECT 3.375000  1.950000 4.055000 2.120000 ;
      RECT 3.455000  0.450000 3.785000 0.580000 ;
      RECT 3.455000  0.580000 4.615000 0.750000 ;
      RECT 3.885000  1.420000 5.805000 1.590000 ;
      RECT 3.885000  1.590000 4.055000 1.950000 ;
      RECT 3.935000  2.630000 5.165000 2.905000 ;
      RECT 3.935000  2.905000 6.115000 2.980000 ;
      RECT 3.945000  1.090000 4.275000 1.250000 ;
      RECT 4.015000  0.085000 4.605000 0.410000 ;
      RECT 4.385000  1.760000 6.145000 1.930000 ;
      RECT 4.385000  1.930000 4.715000 2.290000 ;
      RECT 4.445000  0.750000 4.615000 1.260000 ;
      RECT 4.445000  1.260000 5.805000 1.420000 ;
      RECT 4.785000  0.350000 6.280000 1.090000 ;
      RECT 4.835000  2.980000 6.115000 3.075000 ;
      RECT 5.335000  2.100000 7.045000 2.270000 ;
      RECT 5.335000  2.270000 5.665000 2.735000 ;
      RECT 5.865000  2.440000 6.115000 2.905000 ;
      RECT 5.975000  1.090000 7.355000 1.260000 ;
      RECT 5.975000  1.260000 6.145000 1.760000 ;
      RECT 6.345000  2.440000 6.675000 2.905000 ;
      RECT 6.345000  2.905000 7.575000 3.075000 ;
      RECT 6.450000  0.085000 6.780000 0.920000 ;
      RECT 6.575000  1.950000 7.045000 2.100000 ;
      RECT 6.875000  2.270000 7.045000 2.735000 ;
      RECT 7.025000  0.350000 7.355000 1.090000 ;
      RECT 7.245000  1.950000 8.525000 2.240000 ;
      RECT 7.245000  2.240000 7.575000 2.905000 ;
      RECT 7.640000  0.085000 8.310000 0.985000 ;
      RECT 7.745000  2.410000 8.075000 3.245000 ;
      RECT 8.195000  1.940000 8.525000 1.950000 ;
      RECT 8.250000  2.240000 8.525000 2.990000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
  END
END sky130_fd_sc_hs__or4bb_4
MACRO sky130_fd_sc_hs__sdfbbn_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  16.80000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 1.480000 1.815000 1.810000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.335000 0.350000 16.715000 1.050000 ;
        RECT 16.355000 1.820000 16.715000 2.980000 ;
        RECT 16.545000 1.050000 16.715000 1.820000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.890000 1.820000 15.275000 2.980000 ;
        RECT 14.915000 0.350000 15.275000 1.130000 ;
        RECT 15.105000 1.130000 15.275000 1.820000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.075000 1.190000 14.380000 1.550000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.205000 0.550000 1.875000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.805000 1.205000 1.315000 1.875000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAPARTIALMETALSIDEAREA  2.541000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  8.255000 1.920000  8.545000 1.965000 ;
        RECT  8.255000 1.965000 11.905000 2.105000 ;
        RECT  8.255000 2.105000  8.545000 2.150000 ;
        RECT 11.615000 1.920000 11.905000 1.965000 ;
        RECT 11.615000 2.105000 11.905000 2.150000 ;
    END
  END SET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.470000 1.350000 3.800000 1.780000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 16.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 16.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 16.800000 0.085000 ;
      RECT  0.000000  3.245000 16.800000 3.415000 ;
      RECT  0.115000  2.045000  1.235000 2.215000 ;
      RECT  0.115000  2.215000  0.395000 2.980000 ;
      RECT  0.140000  0.085000  0.470000 1.035000 ;
      RECT  0.565000  2.385000  0.895000 3.245000 ;
      RECT  0.960000  0.575000  1.290000 0.865000 ;
      RECT  0.960000  0.865000  1.655000 1.035000 ;
      RECT  1.065000  2.215000  1.235000 2.905000 ;
      RECT  1.065000  2.905000  2.245000 3.075000 ;
      RECT  1.465000  2.300000  1.715000 2.735000 ;
      RECT  1.485000  1.035000  1.655000 1.140000 ;
      RECT  1.485000  1.140000  2.560000 1.310000 ;
      RECT  1.545000  1.980000  2.155000 2.150000 ;
      RECT  1.545000  2.150000  1.715000 2.300000 ;
      RECT  1.890000  0.085000  2.220000 0.970000 ;
      RECT  1.915000  2.320000  2.245000 2.905000 ;
      RECT  1.985000  1.310000  2.155000 1.980000 ;
      RECT  2.390000  0.255000  3.400000 0.425000 ;
      RECT  2.390000  0.425000  2.560000 1.140000 ;
      RECT  2.470000  2.300000  2.720000 3.245000 ;
      RECT  2.510000  1.480000  3.060000 1.810000 ;
      RECT  2.730000  0.595000  3.060000 1.480000 ;
      RECT  2.890000  1.810000  3.060000 2.300000 ;
      RECT  2.890000  2.300000  3.250000 2.980000 ;
      RECT  3.230000  0.425000  3.400000 0.580000 ;
      RECT  3.230000  0.580000  5.130000 0.750000 ;
      RECT  3.290000  0.920000  4.140000 1.170000 ;
      RECT  3.480000  1.950000  4.140000 2.120000 ;
      RECT  3.480000  2.120000  3.730000 2.980000 ;
      RECT  3.800000  0.085000  4.130000 0.410000 ;
      RECT  3.930000  2.290000  4.180000 3.245000 ;
      RECT  3.970000  1.170000  4.140000 1.340000 ;
      RECT  3.970000  1.340000  4.440000 1.670000 ;
      RECT  3.970000  1.670000  4.140000 1.950000 ;
      RECT  4.310000  0.920000  4.790000 1.170000 ;
      RECT  4.380000  1.840000  4.780000 2.980000 ;
      RECT  4.610000  1.170000  4.790000 1.550000 ;
      RECT  4.610000  1.550000  6.710000 1.720000 ;
      RECT  4.610000  1.720000  4.780000 1.840000 ;
      RECT  4.950000  1.965000  5.215000 2.125000 ;
      RECT  4.950000  2.125000  5.610000 2.295000 ;
      RECT  4.960000  0.750000  5.130000 1.205000 ;
      RECT  4.960000  1.205000  5.970000 1.375000 ;
      RECT  5.020000  2.465000  5.270000 3.245000 ;
      RECT  5.300000  0.085000  5.630000 1.035000 ;
      RECT  5.405000  1.720000  6.710000 1.800000 ;
      RECT  5.405000  1.800000  5.755000 1.905000 ;
      RECT  5.440000  2.295000  5.610000 2.905000 ;
      RECT  5.440000  2.905000  7.505000 3.075000 ;
      RECT  5.800000  0.255000  6.925000 0.425000 ;
      RECT  5.800000  0.425000  5.970000 1.205000 ;
      RECT  5.865000  2.245000  6.195000 2.735000 ;
      RECT  6.025000  1.970000  7.250000 2.140000 ;
      RECT  6.025000  2.140000  6.195000 2.245000 ;
      RECT  6.170000  0.595000  6.420000 1.130000 ;
      RECT  6.170000  1.130000  7.250000 1.300000 ;
      RECT  6.365000  2.310000  7.590000 2.480000 ;
      RECT  6.365000  2.480000  6.695000 2.735000 ;
      RECT  6.380000  1.470000  6.710000 1.550000 ;
      RECT  6.595000  0.425000  6.925000 0.790000 ;
      RECT  6.595000  0.790000  7.590000 0.960000 ;
      RECT  6.920000  1.300000  7.250000 1.970000 ;
      RECT  6.925000  2.650000  7.930000 2.820000 ;
      RECT  6.925000  2.820000  7.505000 2.905000 ;
      RECT  7.150000  0.255000  8.590000 0.425000 ;
      RECT  7.150000  0.425000  7.480000 0.620000 ;
      RECT  7.420000  0.960000  7.590000 2.310000 ;
      RECT  7.760000  0.595000  8.090000 1.080000 ;
      RECT  7.760000  1.080000  7.930000 2.310000 ;
      RECT  7.760000  2.310000  8.830000 2.480000 ;
      RECT  7.760000  2.480000  7.930000 2.650000 ;
      RECT  8.100000  1.290000  9.555000 1.460000 ;
      RECT  8.100000  1.460000  8.430000 1.620000 ;
      RECT  8.125000  2.650000  8.295000 3.245000 ;
      RECT  8.260000  0.425000  8.590000 1.080000 ;
      RECT  8.285000  1.790000  8.990000 1.960000 ;
      RECT  8.285000  1.960000  8.490000 2.140000 ;
      RECT  8.495000  2.480000  8.830000 2.980000 ;
      RECT  8.660000  1.630000  8.990000 1.790000 ;
      RECT  8.660000  2.130000  9.530000 2.300000 ;
      RECT  8.660000  2.300000  8.830000 2.310000 ;
      RECT  8.795000  0.085000  9.125000 1.080000 ;
      RECT  9.050000  2.470000  9.380000 3.245000 ;
      RECT  9.200000  1.630000  9.530000 2.130000 ;
      RECT  9.385000  0.365000 10.920000 0.535000 ;
      RECT  9.385000  0.535000  9.555000 1.290000 ;
      RECT  9.725000  1.260000 11.000000 1.555000 ;
      RECT  9.725000  1.555000 10.070000 1.940000 ;
      RECT  9.745000  0.705000 10.580000 0.920000 ;
      RECT  9.745000  0.920000 11.340000 1.090000 ;
      RECT  9.890000  2.110000 10.410000 2.280000 ;
      RECT  9.890000  2.280000 10.220000 2.980000 ;
      RECT 10.240000  1.725000 11.340000 1.895000 ;
      RECT 10.240000  1.895000 10.410000 2.110000 ;
      RECT 10.665000  2.065000 10.995000 2.630000 ;
      RECT 10.665000  2.630000 13.280000 2.800000 ;
      RECT 10.750000  0.535000 10.920000 0.580000 ;
      RECT 10.750000  0.580000 11.680000 0.750000 ;
      RECT 10.900000  2.970000 11.230000 3.245000 ;
      RECT 11.170000  1.090000 11.340000 1.725000 ;
      RECT 11.170000  1.895000 11.340000 2.290000 ;
      RECT 11.170000  2.290000 12.780000 2.460000 ;
      RECT 11.415000  0.085000 11.755000 0.410000 ;
      RECT 11.460000  2.800000 11.790000 2.980000 ;
      RECT 11.510000  0.750000 11.680000 1.130000 ;
      RECT 11.510000  1.130000 13.905000 1.300000 ;
      RECT 11.630000  1.470000 11.960000 2.120000 ;
      RECT 11.935000  0.255000 13.225000 0.425000 ;
      RECT 11.935000  0.425000 12.265000 0.960000 ;
      RECT 11.995000  2.970000 12.325000 3.245000 ;
      RECT 12.200000  1.300000 12.530000 1.550000 ;
      RECT 12.465000  0.595000 12.795000 0.790000 ;
      RECT 12.465000  0.790000 13.565000 0.960000 ;
      RECT 12.610000  1.720000 13.440000 1.890000 ;
      RECT 12.610000  1.890000 12.780000 2.290000 ;
      RECT 12.770000  1.470000 13.440000 1.720000 ;
      RECT 12.950000  2.060000 13.280000 2.210000 ;
      RECT 12.950000  2.210000 14.720000 2.380000 ;
      RECT 12.950000  2.380000 13.280000 2.630000 ;
      RECT 12.950000  2.800000 13.280000 2.980000 ;
      RECT 12.975000  0.425000 13.225000 0.620000 ;
      RECT 13.395000  0.330000 14.245000 0.500000 ;
      RECT 13.395000  0.500000 13.565000 0.790000 ;
      RECT 13.610000  1.300000 13.780000 1.790000 ;
      RECT 13.610000  1.790000 14.130000 2.040000 ;
      RECT 13.735000  0.670000 13.905000 1.130000 ;
      RECT 14.000000  2.550000 14.690000 3.245000 ;
      RECT 14.075000  0.500000 14.245000 0.850000 ;
      RECT 14.075000  0.850000 14.720000 1.020000 ;
      RECT 14.415000  0.085000 14.735000 0.680000 ;
      RECT 14.550000  1.020000 14.720000 1.300000 ;
      RECT 14.550000  1.300000 14.935000 1.630000 ;
      RECT 14.550000  1.630000 14.720000 2.210000 ;
      RECT 15.450000  0.350000 15.725000 1.220000 ;
      RECT 15.450000  1.220000 16.375000 1.550000 ;
      RECT 15.450000  1.550000 15.700000 2.780000 ;
      RECT 15.905000  0.085000 16.155000 1.050000 ;
      RECT 15.905000  1.900000 16.155000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  1.580000  5.605000 1.750000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  1.950000  8.485000 2.120000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  1.580000  9.925000 1.750000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  1.950000 11.845000 2.120000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.245000 15.205000 3.415000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.245000 15.685000 3.415000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.245000 16.165000 3.415000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  3.245000 16.645000 3.415000 ;
    LAYER met1 ;
      RECT 5.375000 1.550000 5.665000 1.595000 ;
      RECT 5.375000 1.595000 9.985000 1.735000 ;
      RECT 5.375000 1.735000 5.665000 1.780000 ;
      RECT 9.695000 1.550000 9.985000 1.595000 ;
      RECT 9.695000 1.735000 9.985000 1.780000 ;
  END
END sky130_fd_sc_hs__sdfbbn_1
MACRO sky130_fd_sc_hs__sdfbbn_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  18.24000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 1.460000 1.815000 1.790000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 17.370000 0.350000 17.705000 1.050000 ;
        RECT 17.395000 1.820000 17.705000 2.980000 ;
        RECT 17.535000 1.050000 17.705000 1.820000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.280000 0.350000 15.610000 1.220000 ;
        RECT 15.375000 1.220000 15.610000 1.550000 ;
        RECT 15.375000 1.550000 15.715000 1.780000 ;
        RECT 15.375000 1.780000 15.625000 2.980000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.945000 1.505000 14.275000 1.835000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.125000 0.550000 2.135000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.805000 1.125000 1.315000 1.795000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAPARTIALMETALSIDEAREA  2.205000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  9.215000 1.550000  9.505000 1.595000 ;
        RECT  9.215000 1.595000 12.385000 1.735000 ;
        RECT  9.215000 1.735000  9.505000 1.780000 ;
        RECT 12.095000 1.550000 12.385000 1.595000 ;
        RECT 12.095000 1.735000 12.385000 1.780000 ;
    END
  END SET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.350000 3.895000 1.780000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 18.240000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 18.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 18.240000 0.085000 ;
      RECT  0.000000  3.245000 18.240000 3.415000 ;
      RECT  0.115000  2.305000  1.235000 2.475000 ;
      RECT  0.115000  2.475000  0.365000 2.980000 ;
      RECT  0.140000  0.085000  0.470000 0.955000 ;
      RECT  0.565000  2.645000  0.895000 3.245000 ;
      RECT  0.960000  0.625000  1.690000 0.955000 ;
      RECT  1.065000  2.475000  1.235000 2.905000 ;
      RECT  1.065000  2.905000  2.185000 3.075000 ;
      RECT  1.405000  2.300000  1.655000 2.735000 ;
      RECT  1.485000  0.955000  1.690000 1.120000 ;
      RECT  1.485000  1.120000  2.770000 1.290000 ;
      RECT  1.485000  1.960000  2.155000 2.130000 ;
      RECT  1.485000  2.130000  1.655000 2.300000 ;
      RECT  1.855000  2.300000  2.185000 2.905000 ;
      RECT  1.985000  1.290000  2.155000 1.960000 ;
      RECT  2.180000  0.085000  2.430000 0.950000 ;
      RECT  2.415000  2.300000  2.745000 3.245000 ;
      RECT  2.600000  0.255000  3.535000 0.425000 ;
      RECT  2.600000  0.425000  2.770000 1.120000 ;
      RECT  2.605000  1.480000  3.195000 1.810000 ;
      RECT  2.940000  0.595000  3.195000 1.480000 ;
      RECT  2.945000  1.810000  3.195000 2.980000 ;
      RECT  3.365000  0.425000  3.535000 0.660000 ;
      RECT  3.365000  0.660000  4.520000 0.830000 ;
      RECT  3.420000  1.000000  4.235000 1.170000 ;
      RECT  3.425000  1.950000  4.235000 2.120000 ;
      RECT  3.425000  2.120000  3.675000 2.980000 ;
      RECT  3.875000  2.290000  4.205000 3.245000 ;
      RECT  3.930000  0.085000  4.180000 0.490000 ;
      RECT  4.065000  1.170000  4.235000 1.340000 ;
      RECT  4.065000  1.340000  4.445000 1.670000 ;
      RECT  4.065000  1.670000  4.235000 1.950000 ;
      RECT  4.350000  0.255000  5.280000 0.425000 ;
      RECT  4.350000  0.425000  4.520000 0.660000 ;
      RECT  4.405000  1.840000  4.785000 2.980000 ;
      RECT  4.615000  1.180000  6.115000 1.350000 ;
      RECT  4.615000  1.350000  4.785000 1.840000 ;
      RECT  4.690000  0.595000  4.940000 1.180000 ;
      RECT  4.965000  2.350000  5.215000 3.245000 ;
      RECT  5.035000  1.830000  5.365000 2.010000 ;
      RECT  5.035000  2.010000  5.555000 2.180000 ;
      RECT  5.110000  0.425000  5.280000 0.840000 ;
      RECT  5.110000  0.840000  6.115000 1.010000 ;
      RECT  5.385000  2.180000  5.555000 2.905000 ;
      RECT  5.385000  2.905000  7.825000 3.075000 ;
      RECT  5.450000  0.085000  5.720000 0.670000 ;
      RECT  5.595000  1.350000  6.115000 1.525000 ;
      RECT  5.595000  1.525000  6.825000 1.840000 ;
      RECT  5.840000  2.040000  7.365000 2.210000 ;
      RECT  5.840000  2.210000  6.170000 2.735000 ;
      RECT  5.945000  0.265000  7.115000 0.435000 ;
      RECT  5.945000  0.435000  6.115000 0.840000 ;
      RECT  6.285000  0.605000  6.615000 1.185000 ;
      RECT  6.285000  1.185000  7.365000 1.355000 ;
      RECT  6.340000  2.380000  7.705000 2.550000 ;
      RECT  6.340000  2.550000  6.670000 2.735000 ;
      RECT  6.495000  1.840000  6.825000 1.855000 ;
      RECT  6.785000  0.435000  7.115000 0.845000 ;
      RECT  6.785000  0.845000  7.705000 1.015000 ;
      RECT  6.900000  2.730000  8.045000 2.900000 ;
      RECT  6.900000  2.900000  7.825000 2.905000 ;
      RECT  7.035000  1.355000  7.365000 2.040000 ;
      RECT  7.345000  0.265000  8.620000 0.435000 ;
      RECT  7.345000  0.435000  7.770000 0.675000 ;
      RECT  7.535000  1.015000  7.705000 2.380000 ;
      RECT  7.875000  0.945000  8.280000 1.115000 ;
      RECT  7.875000  1.115000  8.045000 2.125000 ;
      RECT  7.875000  2.125000  9.235000 2.295000 ;
      RECT  7.875000  2.295000  8.045000 2.730000 ;
      RECT  7.950000  0.605000  8.280000 0.945000 ;
      RECT  8.215000  1.285000  8.620000 1.955000 ;
      RECT  8.365000  2.465000  8.695000 3.245000 ;
      RECT  8.450000  0.435000  8.620000 0.605000 ;
      RECT  8.450000  0.605000  8.885000 0.935000 ;
      RECT  8.450000  1.110000  9.725000 1.280000 ;
      RECT  8.450000  1.280000  8.620000 1.285000 ;
      RECT  8.790000  1.450000  9.445000 1.780000 ;
      RECT  8.905000  1.950000  9.945000 2.120000 ;
      RECT  8.905000  2.120000  9.235000 2.125000 ;
      RECT  8.905000  2.295000  9.235000 2.980000 ;
      RECT  9.055000  0.085000  9.385000 0.940000 ;
      RECT  9.465000  2.290000  9.795000 3.245000 ;
      RECT  9.555000  0.260000 11.510000 0.430000 ;
      RECT  9.555000  0.430000  9.725000 1.110000 ;
      RECT  9.615000  1.580000  9.945000 1.950000 ;
      RECT  9.960000  0.600000 11.110000 0.850000 ;
      RECT 10.155000  1.180000 10.485000 1.280000 ;
      RECT 10.155000  1.280000 11.385000 1.580000 ;
      RECT 10.155000  1.580000 10.485000 1.755000 ;
      RECT 10.305000  2.100000 10.910000 2.270000 ;
      RECT 10.305000  2.270000 10.635000 2.980000 ;
      RECT 10.740000  1.750000 11.750000 1.920000 ;
      RECT 10.740000  1.920000 10.910000 2.100000 ;
      RECT 10.940000  0.850000 11.110000 0.940000 ;
      RECT 10.940000  0.940000 11.725000 1.110000 ;
      RECT 11.080000  2.090000 11.410000 2.260000 ;
      RECT 11.080000  2.260000 13.435000 2.430000 ;
      RECT 11.230000  2.600000 11.560000 3.245000 ;
      RECT 11.340000  0.430000 11.510000 0.600000 ;
      RECT 11.340000  0.600000 12.065000 0.770000 ;
      RECT 11.555000  1.110000 11.725000 1.750000 ;
      RECT 11.580000  1.920000 12.665000 2.090000 ;
      RECT 11.680000  0.085000 12.055000 0.430000 ;
      RECT 11.805000  2.430000 12.135000 2.980000 ;
      RECT 11.895000  0.770000 12.665000 0.940000 ;
      RECT 11.955000  1.180000 12.325000 1.750000 ;
      RECT 12.235000  0.255000 13.595000 0.425000 ;
      RECT 12.235000  0.425000 12.655000 0.600000 ;
      RECT 12.305000  2.600000 12.635000 3.245000 ;
      RECT 12.495000  0.940000 12.665000 1.130000 ;
      RECT 12.495000  1.130000 14.150000 1.300000 ;
      RECT 12.495000  1.300000 12.825000 1.550000 ;
      RECT 12.495000  1.720000 13.365000 1.890000 ;
      RECT 12.495000  1.890000 12.665000 1.920000 ;
      RECT 12.835000  0.595000 13.085000 0.665000 ;
      RECT 12.835000  0.665000 14.490000 0.835000 ;
      RECT 12.835000  0.835000 13.085000 0.960000 ;
      RECT 13.035000  1.470000 13.365000 1.720000 ;
      RECT 13.185000  2.060000 13.435000 2.260000 ;
      RECT 13.185000  2.430000 13.435000 2.505000 ;
      RECT 13.185000  2.505000 14.655000 2.675000 ;
      RECT 13.185000  2.675000 13.435000 2.980000 ;
      RECT 13.265000  0.425000 13.595000 0.495000 ;
      RECT 13.605000  1.005000 14.150000 1.130000 ;
      RECT 13.605000  1.300000 14.150000 1.335000 ;
      RECT 13.605000  1.335000 13.775000 2.005000 ;
      RECT 13.605000  2.005000 14.075000 2.335000 ;
      RECT 14.280000  2.845000 15.170000 3.245000 ;
      RECT 14.320000  0.835000 14.655000 1.005000 ;
      RECT 14.485000  1.005000 14.655000 1.430000 ;
      RECT 14.485000  1.430000 14.815000 1.760000 ;
      RECT 14.485000  1.760000 14.655000 2.505000 ;
      RECT 14.825000  0.085000 15.110000 1.130000 ;
      RECT 14.825000  1.950000 15.170000 2.845000 ;
      RECT 15.780000  0.085000 16.110000 1.130000 ;
      RECT 15.825000  1.950000 16.155000 3.245000 ;
      RECT 16.340000  0.540000 16.670000 1.220000 ;
      RECT 16.340000  1.220000 17.365000 1.550000 ;
      RECT 16.340000  1.550000 16.700000 2.940000 ;
      RECT 16.870000  0.085000 17.200000 1.050000 ;
      RECT 16.895000  1.820000 17.225000 3.245000 ;
      RECT 17.875000  1.820000 18.125000 3.245000 ;
      RECT 17.880000  0.085000 18.130000 1.130000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  1.210000  6.085000 1.380000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  1.580000  9.445000 1.750000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  1.210000 10.405000 1.380000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  1.580000 12.325000 1.750000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.245000 15.205000 3.415000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.245000 15.685000 3.415000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.245000 16.165000 3.415000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  3.245000 16.645000 3.415000 ;
      RECT 16.955000 -0.085000 17.125000 0.085000 ;
      RECT 16.955000  3.245000 17.125000 3.415000 ;
      RECT 17.435000 -0.085000 17.605000 0.085000 ;
      RECT 17.435000  3.245000 17.605000 3.415000 ;
      RECT 17.915000 -0.085000 18.085000 0.085000 ;
      RECT 17.915000  3.245000 18.085000 3.415000 ;
    LAYER met1 ;
      RECT  5.855000 1.180000  6.145000 1.225000 ;
      RECT  5.855000 1.225000 10.465000 1.365000 ;
      RECT  5.855000 1.365000  6.145000 1.410000 ;
      RECT 10.175000 1.180000 10.465000 1.225000 ;
      RECT 10.175000 1.365000 10.465000 1.410000 ;
  END
END sky130_fd_sc_hs__sdfbbn_2
MACRO sky130_fd_sc_hs__sdfbbp_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  15.84000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455000 1.525000 1.765000 1.855000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.530100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.395000 0.350000 15.735000 2.980000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.518900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.770000 0.350000 14.275000 1.050000 ;
        RECT 13.870000 1.720000 14.275000 2.890000 ;
        RECT 14.105000 1.050000 14.275000 1.720000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.065000 1.180000 13.360000 1.550000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.125000 0.550000 2.135000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.805000 1.550000 1.285000 2.095000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.470000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  7.045000 1.410000  7.375000 1.655000 ;
        RECT  7.095000 1.655000  7.265000 2.905000 ;
        RECT  7.095000 2.905000  8.105000 3.075000 ;
        RECT  7.935000 2.165000  9.025000 2.335000 ;
        RECT  7.935000 2.335000  8.105000 2.905000 ;
        RECT  8.855000 2.335000  9.025000 2.905000 ;
        RECT  8.855000 2.905000 10.265000 3.075000 ;
        RECT 10.095000 2.015000 10.295000 2.185000 ;
        RECT 10.095000 2.185000 10.265000 2.905000 ;
        RECT 10.125000 1.690000 11.385000 1.800000 ;
        RECT 10.125000 1.800000 11.365000 1.860000 ;
        RECT 10.125000 1.860000 10.295000 2.015000 ;
        RECT 11.055000 1.520000 11.385000 1.690000 ;
        RECT 11.055000 1.860000 11.365000 2.150000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.430000 1.180000 3.760000 1.670000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 15.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 15.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 15.840000 0.085000 ;
      RECT  0.000000  3.245000 15.840000 3.415000 ;
      RECT  0.115000  2.305000  1.285000 2.475000 ;
      RECT  0.115000  2.475000  0.445000 2.980000 ;
      RECT  0.140000  0.085000  0.470000 0.955000 ;
      RECT  0.615000  2.645000  0.945000 3.245000 ;
      RECT  1.040000  0.575000  1.370000 1.185000 ;
      RECT  1.040000  1.185000  2.420000 1.355000 ;
      RECT  1.115000  2.475000  1.285000 2.905000 ;
      RECT  1.115000  2.905000  2.275000 3.075000 ;
      RECT  1.495000  2.025000  2.105000 2.195000 ;
      RECT  1.495000  2.195000  1.745000 2.735000 ;
      RECT  1.830000  0.085000  2.080000 1.015000 ;
      RECT  1.935000  1.355000  2.105000 2.025000 ;
      RECT  1.945000  2.520000  2.275000 2.905000 ;
      RECT  2.250000  0.255000  3.680000 0.425000 ;
      RECT  2.250000  0.425000  2.420000 1.185000 ;
      RECT  2.275000  1.830000  2.780000 2.180000 ;
      RECT  2.275000  2.180000  3.285000 2.350000 ;
      RECT  2.505000  2.520000  2.755000 3.245000 ;
      RECT  2.610000  0.595000  2.860000 1.035000 ;
      RECT  2.610000  1.035000  2.780000 1.830000 ;
      RECT  2.955000  2.350000  3.285000 2.980000 ;
      RECT  3.090000  0.595000  3.340000 1.010000 ;
      RECT  3.090000  1.010000  3.260000 1.840000 ;
      RECT  3.090000  1.840000  4.245000 2.010000 ;
      RECT  3.510000  0.425000  3.680000 0.660000 ;
      RECT  3.510000  0.660000  5.335000 0.830000 ;
      RECT  3.515000  2.010000  3.845000 2.980000 ;
      RECT  3.850000  0.085000  4.180000 0.490000 ;
      RECT  4.045000  2.180000  4.215000 3.245000 ;
      RECT  4.075000  1.340000  4.565000 1.670000 ;
      RECT  4.075000  1.670000  4.245000 1.840000 ;
      RECT  4.360000  1.000000  4.905000 1.170000 ;
      RECT  4.415000  1.840000  4.905000 2.980000 ;
      RECT  4.735000  1.170000  4.905000 1.365000 ;
      RECT  4.735000  1.365000  5.445000 1.695000 ;
      RECT  4.735000  1.695000  4.905000 1.840000 ;
      RECT  5.005000  0.460000  5.335000 0.660000 ;
      RECT  5.075000  1.865000  5.785000 2.035000 ;
      RECT  5.075000  2.035000  5.405000 2.755000 ;
      RECT  5.165000  0.830000  5.335000 1.025000 ;
      RECT  5.165000  1.025000  5.785000 1.195000 ;
      RECT  5.505000  0.460000  5.835000 0.685000 ;
      RECT  5.505000  0.685000  6.125000 0.855000 ;
      RECT  5.575000  2.205000  6.125000 2.535000 ;
      RECT  5.615000  1.195000  5.785000 1.865000 ;
      RECT  5.955000  0.855000  6.125000 1.655000 ;
      RECT  5.955000  1.655000  6.875000 1.825000 ;
      RECT  5.955000  1.825000  6.125000 2.205000 ;
      RECT  6.295000  0.730000  8.855000 0.900000 ;
      RECT  6.295000  0.900000  6.535000 1.485000 ;
      RECT  6.490000  0.085000  6.885000 0.560000 ;
      RECT  6.595000  2.075000  6.925000 3.245000 ;
      RECT  6.705000  1.070000  7.915000 1.240000 ;
      RECT  6.705000  1.240000  6.875000 1.655000 ;
      RECT  7.145000  0.310000  8.715000 0.480000 ;
      RECT  7.145000  0.480000  7.640000 0.560000 ;
      RECT  7.435000  1.825000  9.015000 1.995000 ;
      RECT  7.435000  1.995000  7.765000 2.735000 ;
      RECT  7.585000  1.240000  7.915000 1.585000 ;
      RECT  7.820000  0.655000  8.150000 0.730000 ;
      RECT  8.125000  1.180000  8.515000 1.585000 ;
      RECT  8.315000  2.505000  8.685000 3.245000 ;
      RECT  8.330000  0.480000  8.715000 0.560000 ;
      RECT  8.685000  0.900000  8.855000 1.335000 ;
      RECT  8.685000  1.335000  9.015000 1.825000 ;
      RECT  9.025000  0.085000  9.275000 1.050000 ;
      RECT  9.255000  1.335000  9.615000 1.505000 ;
      RECT  9.255000  1.505000  9.585000 1.940000 ;
      RECT  9.375000  2.110000  9.925000 2.735000 ;
      RECT  9.445000  0.255000 10.485000 0.425000 ;
      RECT  9.445000  0.425000  9.615000 1.335000 ;
      RECT  9.755000  1.675000  9.955000 1.845000 ;
      RECT  9.755000  1.845000  9.925000 2.110000 ;
      RECT  9.785000  0.595000  9.985000 1.350000 ;
      RECT  9.785000  1.350000 10.885000 1.520000 ;
      RECT  9.785000  1.520000  9.955000 1.675000 ;
      RECT 10.155000  0.425000 10.485000 1.180000 ;
      RECT 10.435000  2.660000 11.150000 3.245000 ;
      RECT 10.465000  2.030000 10.795000 2.320000 ;
      RECT 10.465000  2.320000 11.785000 2.490000 ;
      RECT 10.715000  1.180000 11.875000 1.350000 ;
      RECT 10.900000  0.085000 11.150000 1.010000 ;
      RECT 11.330000  0.255000 12.555000 0.425000 ;
      RECT 11.330000  0.425000 11.660000 1.010000 ;
      RECT 11.535000  1.970000 12.215000 2.140000 ;
      RECT 11.535000  2.140000 13.700000 2.310000 ;
      RECT 11.535000  2.310000 11.785000 2.320000 ;
      RECT 11.535000  2.490000 11.785000 2.980000 ;
      RECT 11.595000  1.350000 11.875000 1.550000 ;
      RECT 11.870000  0.595000 12.215000 1.010000 ;
      RECT 12.045000  1.010000 12.215000 1.970000 ;
      RECT 12.295000  2.480000 12.625000 3.245000 ;
      RECT 12.385000  0.425000 12.555000 1.010000 ;
      RECT 12.445000  1.180000 12.895000 1.720000 ;
      RECT 12.725000  0.670000 13.115000 1.010000 ;
      RECT 12.725000  1.010000 12.895000 1.180000 ;
      RECT 12.725000  1.720000 13.155000 1.970000 ;
      RECT 13.295000  0.085000 13.590000 1.000000 ;
      RECT 13.340000  2.480000 13.670000 3.245000 ;
      RECT 13.530000  1.220000 13.915000 1.550000 ;
      RECT 13.530000  1.550000 13.700000 2.140000 ;
      RECT 14.445000  0.350000 14.715000 1.355000 ;
      RECT 14.445000  1.355000 14.845000 1.685000 ;
      RECT 14.445000  1.685000 14.775000 2.980000 ;
      RECT 14.895000  0.085000 15.225000 0.940000 ;
      RECT 14.945000  2.115000 15.205000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  1.210000  8.485000 1.380000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  1.210000 12.805000 1.380000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.245000 15.205000 3.415000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.245000 15.685000 3.415000 ;
    LAYER met1 ;
      RECT  8.255000 1.180000  8.545000 1.225000 ;
      RECT  8.255000 1.225000 12.865000 1.365000 ;
      RECT  8.255000 1.365000  8.545000 1.410000 ;
      RECT 12.575000 1.180000 12.865000 1.225000 ;
      RECT 12.575000 1.365000 12.865000 1.410000 ;
  END
END sky130_fd_sc_hs__sdfbbp_1
MACRO sky130_fd_sc_hs__sdfrbp_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.92000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 0.810000 2.100000 1.310000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.518900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.470000 0.350000 13.835000 1.130000 ;
        RECT 13.555000 1.820000 13.835000 2.980000 ;
        RECT 13.665000 1.130000 13.835000 1.820000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.537600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.015000 0.350000 12.345000 2.980000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  3.935000 1.920000  4.225000 1.965000 ;
        RECT  3.935000 1.965000 10.945000 2.105000 ;
        RECT  3.935000 2.105000  4.225000 2.150000 ;
        RECT  7.775000 1.920000  8.065000 1.965000 ;
        RECT  7.775000 2.105000  8.065000 2.150000 ;
        RECT 10.655000 1.920000 10.945000 1.965000 ;
        RECT 10.655000 2.105000 10.945000 2.150000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.935000 1.440000 3.265000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.490000 2.725000 1.660000 ;
        RECT 0.605000 1.660000 1.795000 1.880000 ;
        RECT 2.395000 1.260000 2.725000 1.490000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.785000 0.920000 4.060000 1.180000 ;
        RECT 3.785000 1.180000 4.645000 1.630000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 13.920000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 13.920000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.920000 0.085000 ;
      RECT  0.000000  3.245000 13.920000 3.415000 ;
      RECT  0.115000  0.350000  0.365000 0.980000 ;
      RECT  0.115000  0.980000  1.395000 1.310000 ;
      RECT  0.115000  1.310000  0.285000 2.050000 ;
      RECT  0.115000  2.050000  2.695000 2.220000 ;
      RECT  0.115000  2.220000  1.055000 2.975000 ;
      RECT  0.545000  0.085000  0.875000 0.810000 ;
      RECT  1.105000  0.255000  3.410000 0.425000 ;
      RECT  1.105000  0.425000  1.355000 0.810000 ;
      RECT  1.225000  2.390000  1.555000 3.245000 ;
      RECT  2.095000  2.390000  4.230000 2.400000 ;
      RECT  2.095000  2.400000  4.250000 2.420000 ;
      RECT  2.095000  2.420000  6.075000 2.560000 ;
      RECT  2.095000  2.560000  2.945000 2.600000 ;
      RECT  2.095000  2.600000  2.555000 2.980000 ;
      RECT  2.270000  0.595000  2.600000 0.920000 ;
      RECT  2.270000  0.920000  3.615000 1.090000 ;
      RECT  2.365000  1.830000  2.695000 2.050000 ;
      RECT  3.060000  0.425000  3.410000 0.750000 ;
      RECT  3.095000  2.730000  3.425000 3.245000 ;
      RECT  3.445000  1.090000  3.615000 2.330000 ;
      RECT  3.445000  2.330000  3.785000 2.385000 ;
      RECT  3.445000  2.385000  4.230000 2.390000 ;
      RECT  3.590000  0.085000  3.880000 0.750000 ;
      RECT  3.665000  2.560000  6.075000 2.580000 ;
      RECT  3.665000  2.580000  4.645000 2.585000 ;
      RECT  3.665000  2.585000  4.630000 2.590000 ;
      RECT  3.665000  2.590000  4.610000 2.600000 ;
      RECT  3.665000  2.600000  4.580000 2.620000 ;
      RECT  3.665000  2.620000  3.995000 2.980000 ;
      RECT  3.785000  1.830000  4.165000 2.160000 ;
      RECT  3.920000  2.160000  4.165000 2.190000 ;
      RECT  4.135000  0.500000  4.535000 0.750000 ;
      RECT  4.230000  0.750000  4.535000 0.840000 ;
      RECT  4.230000  0.840000  5.045000 1.010000 ;
      RECT  4.335000  1.800000  4.985000 2.195000 ;
      RECT  4.335000  2.195000  4.505000 2.250000 ;
      RECT  4.555000  2.415000  6.075000 2.420000 ;
      RECT  4.570000  2.410000  6.075000 2.415000 ;
      RECT  4.590000  2.400000  6.075000 2.410000 ;
      RECT  4.615000  2.385000  6.075000 2.400000 ;
      RECT  4.705000  0.085000  5.035000 0.670000 ;
      RECT  4.705000  2.750000  5.035000 3.245000 ;
      RECT  4.815000  1.010000  5.045000 1.455000 ;
      RECT  4.815000  1.455000  5.280000 1.775000 ;
      RECT  4.815000  1.775000  4.985000 1.800000 ;
      RECT  5.155000  1.955000  5.630000 2.215000 ;
      RECT  5.215000  0.255000  7.220000 0.425000 ;
      RECT  5.215000  0.425000  5.620000 1.070000 ;
      RECT  5.215000  1.070000  5.630000 1.285000 ;
      RECT  5.450000  1.285000  5.630000 1.545000 ;
      RECT  5.450000  1.545000  6.175000 1.875000 ;
      RECT  5.450000  1.875000  5.630000 1.955000 ;
      RECT  5.795000  0.595000  5.975000 0.995000 ;
      RECT  5.800000  0.995000  5.975000 1.200000 ;
      RECT  5.800000  1.200000  6.515000 1.370000 ;
      RECT  5.825000  2.045000  6.515000 2.215000 ;
      RECT  5.825000  2.215000  6.075000 2.385000 ;
      RECT  5.825000  2.580000  6.075000 2.725000 ;
      RECT  6.145000  0.595000  6.470000 0.860000 ;
      RECT  6.145000  0.860000  6.855000 1.030000 ;
      RECT  6.250000  2.385000  6.855000 2.725000 ;
      RECT  6.345000  1.370000  6.515000 2.045000 ;
      RECT  6.685000  1.030000  6.855000 1.985000 ;
      RECT  6.685000  1.985000  7.605000 2.165000 ;
      RECT  6.685000  2.165000  6.855000 2.385000 ;
      RECT  7.025000  0.920000  8.655000 1.090000 ;
      RECT  7.025000  1.090000  7.265000 1.805000 ;
      RECT  7.025000  2.345000  7.265000 3.245000 ;
      RECT  7.050000  0.425000  7.220000 0.580000 ;
      RECT  7.050000  0.580000  8.100000 0.750000 ;
      RECT  7.430000  0.085000  7.760000 0.410000 ;
      RECT  7.435000  1.260000  8.315000 1.545000 ;
      RECT  7.435000  1.545000  7.605000 1.985000 ;
      RECT  7.435000  2.165000  7.605000 2.320000 ;
      RECT  7.435000  2.320000  7.765000 2.745000 ;
      RECT  7.775000  1.795000  8.035000 2.150000 ;
      RECT  7.930000  0.255000  8.995000 0.425000 ;
      RECT  7.930000  0.425000  8.100000 0.580000 ;
      RECT  8.235000  1.715000  8.485000 3.245000 ;
      RECT  8.270000  0.595000  8.655000 0.920000 ;
      RECT  8.485000  1.090000  8.655000 1.245000 ;
      RECT  8.485000  1.245000  8.935000 1.415000 ;
      RECT  8.685000  1.415000  8.935000 2.755000 ;
      RECT  8.825000  0.425000  8.995000 0.905000 ;
      RECT  8.825000  0.905000  9.435000 1.075000 ;
      RECT  9.105000  1.075000  9.435000 1.345000 ;
      RECT  9.105000  1.345000  9.755000 1.575000 ;
      RECT  9.105000  1.755000  9.325000 2.425000 ;
      RECT  9.105000  2.425000 10.095000 2.755000 ;
      RECT  9.165000  0.405000  9.775000 0.735000 ;
      RECT  9.505000  1.575000  9.755000 2.230000 ;
      RECT  9.605000  0.735000  9.775000 1.005000 ;
      RECT  9.605000  1.005000 11.425000 1.175000 ;
      RECT  9.925000  1.175000 11.425000 1.435000 ;
      RECT  9.925000  1.435000 10.095000 2.425000 ;
      RECT 10.165000  0.085000 10.495000 0.760000 ;
      RECT 10.265000  1.650000 10.525000 2.320000 ;
      RECT 10.265000  2.320000 11.405000 2.490000 ;
      RECT 10.305000  2.660000 10.650000 3.245000 ;
      RECT 10.695000  1.685000 11.065000 2.150000 ;
      RECT 10.855000  2.490000 11.185000 2.885000 ;
      RECT 10.955000  0.350000 11.285000 0.580000 ;
      RECT 10.955000  0.580000 11.845000 0.750000 ;
      RECT 11.235000  1.630000 11.845000 1.800000 ;
      RECT 11.235000  1.800000 11.405000 2.320000 ;
      RECT 11.370000  2.695000 11.815000 3.245000 ;
      RECT 11.510000  0.085000 11.840000 0.410000 ;
      RECT 11.585000  1.970000 11.815000 2.695000 ;
      RECT 11.675000  0.750000 11.845000 1.630000 ;
      RECT 12.570000  0.455000 12.855000 1.300000 ;
      RECT 12.570000  1.300000 13.485000 1.630000 ;
      RECT 12.570000  1.630000 12.855000 2.980000 ;
      RECT 13.045000  1.820000 13.325000 3.245000 ;
      RECT 13.120000  0.085000 13.290000 1.130000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  1.950000  4.165000 2.120000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  1.950000  8.005000 2.120000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  1.950000 10.885000 2.120000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
  END
END sky130_fd_sc_hs__sdfrbp_1
MACRO sky130_fd_sc_hs__sdfrbp_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.88000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 0.810000 2.090000 1.190000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.055000 0.350000 14.325000 2.980000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.030000 0.915000 12.465000 1.085000 ;
        RECT 12.030000 1.085000 12.360000 2.980000 ;
        RECT 12.135000 0.350000 12.465000 0.915000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  3.935000 1.920000  4.225000 1.965000 ;
        RECT  3.935000 1.965000 10.945000 2.105000 ;
        RECT  3.935000 2.105000  4.225000 2.150000 ;
        RECT  7.775000 1.920000  8.065000 1.965000 ;
        RECT  7.775000 2.105000  8.065000 2.150000 ;
        RECT 10.655000 1.920000 10.945000 1.965000 ;
        RECT 10.655000 2.105000 10.945000 2.150000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.945000 1.440000 3.275000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.540000 1.820000 1.795000 2.150000 ;
        RECT 1.625000 1.360000 2.735000 1.620000 ;
        RECT 1.625000 1.620000 1.795000 1.820000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.905000 1.180000 4.235000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 14.880000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 14.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.880000 0.085000 ;
      RECT  0.000000  3.245000 14.880000 3.415000 ;
      RECT  0.115000  0.375000  0.365000 1.250000 ;
      RECT  0.115000  1.250000  1.395000 1.580000 ;
      RECT  0.115000  1.580000  0.285000 2.320000 ;
      RECT  0.115000  2.320000  2.605000 2.490000 ;
      RECT  0.115000  2.490000  0.445000 2.980000 ;
      RECT  0.545000  0.085000  0.875000 0.835000 ;
      RECT  0.615000  2.730000  1.400000 3.245000 ;
      RECT  1.095000  0.255000  3.430000 0.425000 ;
      RECT  1.095000  0.425000  1.345000 0.835000 ;
      RECT  1.940000  2.660000  2.945000 2.910000 ;
      RECT  2.260000  0.595000  2.610000 1.005000 ;
      RECT  2.260000  1.005000  3.615000 1.175000 ;
      RECT  2.275000  1.830000  2.605000 2.320000 ;
      RECT  2.775000  2.320000  3.995000 2.420000 ;
      RECT  2.775000  2.420000  5.985000 2.490000 ;
      RECT  2.775000  2.490000  2.945000 2.660000 ;
      RECT  3.100000  0.425000  3.430000 0.835000 ;
      RECT  3.115000  2.660000  3.445000 3.245000 ;
      RECT  3.445000  1.175000  3.615000 2.320000 ;
      RECT  3.615000  2.490000  5.985000 2.580000 ;
      RECT  3.615000  2.580000  4.645000 2.590000 ;
      RECT  3.615000  2.590000  3.995000 2.980000 ;
      RECT  3.640000  0.085000  3.970000 0.835000 ;
      RECT  3.785000  1.820000  4.165000 2.150000 ;
      RECT  4.240000  0.595000  4.575000 1.010000 ;
      RECT  4.335000  1.820000  4.985000 1.990000 ;
      RECT  4.335000  1.990000  4.505000 2.250000 ;
      RECT  4.405000  1.010000  4.575000 1.445000 ;
      RECT  4.405000  1.445000  5.305000 1.775000 ;
      RECT  4.405000  1.775000  4.985000 1.820000 ;
      RECT  4.570000  2.410000  5.985000 2.420000 ;
      RECT  4.705000  2.750000  5.035000 3.245000 ;
      RECT  4.750000  0.085000  4.920000 1.130000 ;
      RECT  5.100000  0.310000  7.170000 0.480000 ;
      RECT  5.100000  0.480000  5.430000 0.990000 ;
      RECT  5.100000  0.990000  5.645000 1.275000 ;
      RECT  5.155000  1.945000  6.150000 1.985000 ;
      RECT  5.155000  1.985000  5.675000 2.030000 ;
      RECT  5.155000  2.030000  5.630000 2.240000 ;
      RECT  5.430000  1.900000  6.150000 1.945000 ;
      RECT  5.475000  1.275000  5.645000 1.500000 ;
      RECT  5.475000  1.500000  6.150000 1.900000 ;
      RECT  5.660000  0.650000  5.990000 0.820000 ;
      RECT  5.710000  2.580000  5.985000 2.725000 ;
      RECT  5.800000  2.155000  6.490000 2.325000 ;
      RECT  5.800000  2.325000  5.985000 2.410000 ;
      RECT  5.820000  0.820000  5.990000 1.120000 ;
      RECT  5.820000  1.120000  6.490000 1.290000 ;
      RECT  6.160000  0.650000  6.830000 0.950000 ;
      RECT  6.160000  2.495000  7.915000 2.510000 ;
      RECT  6.160000  2.510000  6.900000 2.725000 ;
      RECT  6.320000  1.290000  6.490000 2.155000 ;
      RECT  6.660000  0.950000  6.830000 2.340000 ;
      RECT  6.660000  2.340000  7.915000 2.495000 ;
      RECT  7.000000  0.480000  7.170000 0.580000 ;
      RECT  7.000000  0.580000  8.325000 0.750000 ;
      RECT  7.000000  0.920000  8.930000 1.090000 ;
      RECT  7.000000  1.090000  7.210000 1.780000 ;
      RECT  7.070000  2.680000  7.320000 3.245000 ;
      RECT  7.380000  1.260000  8.590000 1.575000 ;
      RECT  7.380000  1.575000  7.550000 2.320000 ;
      RECT  7.380000  2.320000  7.915000 2.340000 ;
      RECT  7.450000  0.085000  7.985000 0.410000 ;
      RECT  7.550000  2.510000  7.915000 2.725000 ;
      RECT  7.720000  1.795000  8.020000 2.150000 ;
      RECT  8.155000  0.255000  9.270000 0.425000 ;
      RECT  8.155000  0.425000  8.325000 0.580000 ;
      RECT  8.190000  1.745000  8.440000 3.245000 ;
      RECT  8.495000  0.595000  8.930000 0.920000 ;
      RECT  8.640000  1.745000  8.930000 2.755000 ;
      RECT  8.760000  1.090000  8.930000 1.745000 ;
      RECT  9.100000  0.425000  9.270000 0.905000 ;
      RECT  9.100000  0.905000  9.640000 1.235000 ;
      RECT  9.100000  2.365000 10.095000 2.695000 ;
      RECT  9.310000  1.235000  9.640000 1.865000 ;
      RECT  9.310000  1.865000  9.755000 2.195000 ;
      RECT  9.440000  0.405000 10.095000 0.735000 ;
      RECT  9.925000  0.735000 10.095000 1.045000 ;
      RECT  9.925000  1.045000 11.520000 1.310000 ;
      RECT  9.925000  1.310000 10.095000 2.365000 ;
      RECT 10.265000  1.480000 11.860000 1.650000 ;
      RECT 10.265000  1.650000 10.545000 2.320000 ;
      RECT 10.265000  2.320000 11.395000 2.490000 ;
      RECT 10.265000  2.660000 10.860000 3.245000 ;
      RECT 10.335000  0.085000 10.665000 0.810000 ;
      RECT 10.715000  1.820000 11.395000 2.150000 ;
      RECT 11.065000  2.490000 11.395000 2.795000 ;
      RECT 11.125000  0.350000 11.455000 0.705000 ;
      RECT 11.125000  0.705000 11.860000 0.875000 ;
      RECT 11.600000  1.820000 11.850000 3.245000 ;
      RECT 11.645000  0.085000 11.895000 0.535000 ;
      RECT 11.690000  0.875000 11.860000 1.480000 ;
      RECT 12.540000  1.920000 12.830000 3.245000 ;
      RECT 12.635000  0.085000 12.895000 1.050000 ;
      RECT 13.065000  0.350000 13.325000 1.300000 ;
      RECT 13.065000  1.300000 13.885000 1.630000 ;
      RECT 13.065000  1.630000 13.325000 2.980000 ;
      RECT 13.545000  1.820000 13.875000 3.245000 ;
      RECT 13.670000  0.085000 13.840000 1.130000 ;
      RECT 14.495000  0.085000 14.780000 1.130000 ;
      RECT 14.495000  1.820000 14.775000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  1.950000  4.165000 2.120000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  1.950000  8.005000 2.120000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  1.950000 10.885000 2.120000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
  END
END sky130_fd_sc_hs__sdfrbp_2
MACRO sky130_fd_sc_hs__sdfrtn_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.92000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.780000 1.980000 2.120000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.546900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.475000 0.350000 13.805000 2.980000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  3.455000 1.550000  3.745000 1.595000 ;
        RECT  3.455000 1.595000 11.425000 1.735000 ;
        RECT  3.455000 1.735000  3.745000 1.780000 ;
        RECT  7.775000 1.550000  8.065000 1.595000 ;
        RECT  7.775000 1.735000  8.065000 1.780000 ;
        RECT 11.135000 1.550000 11.425000 1.595000 ;
        RECT 11.135000 1.735000 11.425000 1.780000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.800000 1.525000 3.235000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 1.410000 2.045000 1.580000 ;
        RECT 0.535000 1.580000 0.865000 2.080000 ;
        RECT 1.875000 0.955000 2.550000 1.410000 ;
    END
  END SCE
  PIN CLK_N
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.275000 1.210000 4.675000 1.550000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 13.920000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 13.920000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.920000 0.085000 ;
      RECT  0.000000  3.245000 13.920000 3.415000 ;
      RECT  0.115000  0.420000  0.445000 1.050000 ;
      RECT  0.115000  1.050000  1.620000 1.240000 ;
      RECT  0.115000  1.240000  0.365000 2.290000 ;
      RECT  0.115000  2.290000  2.545000 2.460000 ;
      RECT  0.115000  2.460000  0.365000 2.980000 ;
      RECT  0.565000  2.630000  0.895000 3.245000 ;
      RECT  0.615000  0.085000  0.945000 0.880000 ;
      RECT  1.165000  0.255000  3.390000 0.425000 ;
      RECT  1.165000  0.425000  1.495000 0.765000 ;
      RECT  1.290000  0.935000  1.620000 1.050000 ;
      RECT  1.405000  2.630000  3.680000 2.800000 ;
      RECT  1.405000  2.800000  2.220000 2.960000 ;
      RECT  1.955000  0.595000  2.890000 0.765000 ;
      RECT  2.215000  1.580000  2.545000 2.290000 ;
      RECT  2.720000  0.765000  2.890000 1.015000 ;
      RECT  2.720000  1.015000  4.075000 1.185000 ;
      RECT  2.815000  2.970000  3.145000 3.245000 ;
      RECT  3.060000  0.425000  3.390000 0.845000 ;
      RECT  3.405000  1.355000  3.735000 2.025000 ;
      RECT  3.430000  2.195000  6.115000 2.330000 ;
      RECT  3.430000  2.330000  4.720000 2.340000 ;
      RECT  3.430000  2.340000  4.700000 2.350000 ;
      RECT  3.430000  2.350000  4.645000 2.395000 ;
      RECT  3.430000  2.395000  3.680000 2.630000 ;
      RECT  3.430000  2.800000  3.680000 2.980000 ;
      RECT  3.575000  0.085000  4.065000 0.360000 ;
      RECT  3.905000  0.530000  6.155000 0.700000 ;
      RECT  3.905000  0.700000  4.075000 1.015000 ;
      RECT  3.905000  1.185000  4.075000 2.170000 ;
      RECT  3.905000  2.170000  6.115000 2.195000 ;
      RECT  4.245000  0.870000  5.165000 1.040000 ;
      RECT  4.255000  1.820000  5.030000 1.990000 ;
      RECT  4.255000  1.990000  4.600000 2.000000 ;
      RECT  4.660000  2.160000  6.115000 2.170000 ;
      RECT  4.780000  2.500000  5.110000 3.245000 ;
      RECT  4.805000  0.085000  5.165000 0.360000 ;
      RECT  4.845000  1.040000  5.165000 1.235000 ;
      RECT  4.845000  1.235000  5.255000 1.605000 ;
      RECT  4.845000  1.605000  5.030000 1.820000 ;
      RECT  5.230000  1.775000  6.715000 1.990000 ;
      RECT  5.345000  0.870000  5.675000 1.085000 ;
      RECT  5.425000  1.085000  5.675000 1.265000 ;
      RECT  5.425000  1.265000  6.495000 1.465000 ;
      RECT  5.425000  1.465000  5.675000 1.735000 ;
      RECT  5.425000  1.735000  6.715000 1.775000 ;
      RECT  5.855000  2.330000  6.115000 2.735000 ;
      RECT  5.905000  0.700000  6.155000 1.095000 ;
      RECT  6.285000  2.235000  7.055000 2.445000 ;
      RECT  6.285000  2.445000  6.570000 2.735000 ;
      RECT  6.325000  0.255000  7.720000 0.545000 ;
      RECT  6.325000  0.545000  6.495000 1.265000 ;
      RECT  6.495000  1.990000  6.715000 2.065000 ;
      RECT  6.665000  0.725000  7.055000 1.095000 ;
      RECT  6.885000  1.095000  7.055000 2.040000 ;
      RECT  6.885000  2.040000  8.520000 2.140000 ;
      RECT  6.885000  2.140000  7.950000 2.210000 ;
      RECT  6.885000  2.210000  7.055000 2.235000 ;
      RECT  7.225000  1.130000  9.010000 1.300000 ;
      RECT  7.225000  1.300000  7.475000 1.870000 ;
      RECT  7.225000  2.380000  7.395000 3.245000 ;
      RECT  7.495000  0.545000  7.720000 0.790000 ;
      RECT  7.495000  0.790000  9.825000 0.960000 ;
      RECT  7.575000  2.210000  7.950000 2.735000 ;
      RECT  7.645000  1.970000  8.520000 2.040000 ;
      RECT  7.685000  1.470000  8.035000 1.800000 ;
      RECT  7.890000  0.085000  8.220000 0.620000 ;
      RECT  8.225000  1.470000  8.520000 1.970000 ;
      RECT  8.295000  2.310000  8.625000 3.245000 ;
      RECT  8.690000  1.300000  8.860000 1.970000 ;
      RECT  8.690000  1.970000  9.565000 2.140000 ;
      RECT  8.795000  2.140000  9.565000 2.980000 ;
      RECT  9.030000  1.470000 10.395000 1.540000 ;
      RECT  9.030000  1.540000  9.350000 1.800000 ;
      RECT  9.180000  1.370000 10.395000 1.470000 ;
      RECT  9.190000  0.290000 10.165000 0.620000 ;
      RECT  9.495000  0.960000  9.825000 1.200000 ;
      RECT  9.735000  1.710000 11.025000 1.880000 ;
      RECT  9.735000  1.880000 10.065000 2.980000 ;
      RECT  9.995000  0.620000 10.165000 0.870000 ;
      RECT  9.995000  0.870000 11.895000 1.040000 ;
      RECT 10.065000  1.225000 10.395000 1.370000 ;
      RECT 10.435000  2.050000 10.685000 2.290000 ;
      RECT 10.435000  2.290000 12.235000 2.460000 ;
      RECT 10.605000  2.650000 11.210000 3.245000 ;
      RECT 10.730000  0.085000 11.200000 0.680000 ;
      RECT 10.855000  1.880000 11.025000 1.950000 ;
      RECT 10.855000  1.950000 11.895000 2.120000 ;
      RECT 10.995000  1.210000 11.395000 1.540000 ;
      RECT 11.195000  1.540000 11.395000 1.780000 ;
      RECT 11.380000  2.460000 11.710000 2.980000 ;
      RECT 11.565000  1.040000 11.895000 1.950000 ;
      RECT 11.690000  0.450000 12.235000 0.700000 ;
      RECT 11.880000  2.630000 12.210000 3.245000 ;
      RECT 12.065000  0.700000 12.235000 2.290000 ;
      RECT 12.440000  0.350000 12.795000 1.355000 ;
      RECT 12.440000  1.355000 12.810000 1.685000 ;
      RECT 12.440000  1.685000 12.795000 2.980000 ;
      RECT 12.975000  0.085000 13.305000 1.130000 ;
      RECT 12.975000  1.820000 13.305000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  1.580000  3.685000 1.750000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  1.580000  8.005000 1.750000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  1.580000 11.365000 1.750000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
  END
END sky130_fd_sc_hs__sdfrtn_1
MACRO sky130_fd_sc_hs__sdfrtp_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.44000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 0.810000 2.100000 1.265000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.995000 0.350000 13.325000 1.130000 ;
        RECT 13.070000 1.130000 13.325000 2.980000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  3.935000 1.920000  4.225000 1.965000 ;
        RECT  3.935000 1.965000 10.945000 2.105000 ;
        RECT  3.935000 2.105000  4.225000 2.150000 ;
        RECT  7.775000 1.920000  8.065000 1.965000 ;
        RECT  7.775000 2.105000  8.065000 2.150000 ;
        RECT 10.655000 1.920000 10.945000 1.965000 ;
        RECT 10.655000 2.105000 10.945000 2.150000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.945000 1.440000 3.275000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455000 1.490000 2.725000 1.660000 ;
        RECT 0.455000 1.660000 1.795000 1.835000 ;
        RECT 2.345000 1.260000 2.725000 1.490000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.785000 0.920000 4.195000 1.260000 ;
        RECT 3.785000 1.260000 4.640000 1.650000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 13.440000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 13.440000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.440000 0.085000 ;
      RECT  0.000000  3.245000 13.440000 3.415000 ;
      RECT  0.115000  0.420000  0.365000 1.050000 ;
      RECT  0.115000  1.050000  1.375000 1.265000 ;
      RECT  0.115000  1.265000  0.285000 2.005000 ;
      RECT  0.115000  2.005000  2.705000 2.175000 ;
      RECT  0.115000  2.175000  0.445000 2.980000 ;
      RECT  0.545000  0.085000  0.875000 0.880000 ;
      RECT  0.615000  2.345000  0.945000 3.245000 ;
      RECT  1.045000  0.935000  1.375000 1.050000 ;
      RECT  1.105000  0.255000  3.410000 0.425000 ;
      RECT  1.105000  0.425000  1.435000 0.640000 ;
      RECT  1.485000  2.345000  3.785000 2.385000 ;
      RECT  1.485000  2.385000  4.230000 2.400000 ;
      RECT  1.485000  2.400000  4.250000 2.420000 ;
      RECT  1.485000  2.420000  6.075000 2.515000 ;
      RECT  1.485000  2.515000  2.555000 2.980000 ;
      RECT  2.035000  1.830000  2.705000 2.005000 ;
      RECT  2.270000  0.595000  2.600000 0.920000 ;
      RECT  2.270000  0.920000  3.615000 1.090000 ;
      RECT  3.060000  0.425000  3.410000 0.750000 ;
      RECT  3.095000  2.685000  3.425000 3.245000 ;
      RECT  3.445000  1.090000  3.615000 2.330000 ;
      RECT  3.445000  2.330000  3.785000 2.345000 ;
      RECT  3.590000  0.085000  3.880000 0.750000 ;
      RECT  3.665000  2.515000  6.075000 2.580000 ;
      RECT  3.665000  2.580000  4.645000 2.585000 ;
      RECT  3.665000  2.585000  4.630000 2.590000 ;
      RECT  3.665000  2.590000  4.610000 2.600000 ;
      RECT  3.665000  2.600000  4.580000 2.620000 ;
      RECT  3.665000  2.620000  3.995000 2.980000 ;
      RECT  3.785000  1.830000  4.165000 2.160000 ;
      RECT  3.920000  2.160000  4.165000 2.190000 ;
      RECT  4.135000  0.500000  4.535000 0.750000 ;
      RECT  4.335000  1.820000  4.980000 2.195000 ;
      RECT  4.335000  2.195000  4.505000 2.250000 ;
      RECT  4.365000  0.750000  4.535000 0.920000 ;
      RECT  4.365000  0.920000  5.045000 1.090000 ;
      RECT  4.555000  2.415000  6.075000 2.420000 ;
      RECT  4.570000  2.410000  6.075000 2.415000 ;
      RECT  4.590000  2.400000  6.075000 2.410000 ;
      RECT  4.615000  2.385000  6.075000 2.400000 ;
      RECT  4.705000  0.085000  5.035000 0.750000 ;
      RECT  4.705000  2.750000  5.035000 3.245000 ;
      RECT  4.810000  1.090000  5.045000 1.455000 ;
      RECT  4.810000  1.455000  5.280000 1.775000 ;
      RECT  4.810000  1.775000  4.980000 1.820000 ;
      RECT  5.155000  1.955000  5.630000 2.215000 ;
      RECT  5.215000  0.255000  7.220000 0.425000 ;
      RECT  5.215000  0.425000  5.620000 1.070000 ;
      RECT  5.215000  1.070000  5.630000 1.285000 ;
      RECT  5.450000  1.285000  5.630000 1.545000 ;
      RECT  5.450000  1.545000  6.200000 1.875000 ;
      RECT  5.450000  1.875000  5.630000 1.955000 ;
      RECT  5.795000  0.595000  5.975000 0.995000 ;
      RECT  5.800000  0.995000  5.975000 1.200000 ;
      RECT  5.800000  1.200000  6.540000 1.370000 ;
      RECT  5.825000  2.045000  6.540000 2.215000 ;
      RECT  5.825000  2.215000  6.075000 2.385000 ;
      RECT  5.825000  2.580000  6.075000 2.725000 ;
      RECT  6.145000  0.595000  6.470000 0.860000 ;
      RECT  6.145000  0.860000  6.880000 1.030000 ;
      RECT  6.250000  2.385000  8.075000 2.490000 ;
      RECT  6.250000  2.490000  6.880000 2.725000 ;
      RECT  6.370000  1.370000  6.540000 2.045000 ;
      RECT  6.710000  1.030000  6.880000 2.320000 ;
      RECT  6.710000  2.320000  8.075000 2.385000 ;
      RECT  7.050000  0.425000  7.220000 0.580000 ;
      RECT  7.050000  0.580000  8.100000 0.750000 ;
      RECT  7.050000  0.920000  8.895000 1.090000 ;
      RECT  7.050000  1.090000  7.325000 1.805000 ;
      RECT  7.205000  2.660000  7.540000 3.245000 ;
      RECT  7.430000  0.085000  7.760000 0.410000 ;
      RECT  7.495000  1.260000  8.315000 1.575000 ;
      RECT  7.495000  1.575000  7.665000 2.320000 ;
      RECT  7.745000  2.490000  8.075000 2.745000 ;
      RECT  7.835000  1.815000  8.165000 2.150000 ;
      RECT  7.930000  0.255000  9.235000 0.425000 ;
      RECT  7.930000  0.425000  8.100000 0.580000 ;
      RECT  8.270000  0.595000  8.655000 0.920000 ;
      RECT  8.385000  1.745000  8.555000 3.245000 ;
      RECT  8.725000  1.090000  8.895000 1.715000 ;
      RECT  8.725000  1.715000  9.005000 2.755000 ;
      RECT  9.065000  0.425000  9.235000 0.940000 ;
      RECT  9.065000  0.940000  9.415000 1.270000 ;
      RECT  9.245000  1.270000  9.415000 2.125000 ;
      RECT  9.245000  2.125000  9.975000 2.380000 ;
      RECT  9.290000  2.550000 10.315000 2.880000 ;
      RECT  9.405000  0.350000  9.755000 0.770000 ;
      RECT  9.585000  0.770000  9.755000 1.095000 ;
      RECT  9.585000  1.095000 11.395000 1.265000 ;
      RECT  9.585000  1.265000  9.755000 1.785000 ;
      RECT  9.585000  1.785000 10.315000 1.955000 ;
      RECT  9.985000  1.435000 10.315000 1.445000 ;
      RECT  9.985000  1.445000 11.735000 1.615000 ;
      RECT 10.145000  1.955000 10.315000 2.550000 ;
      RECT 10.195000  0.085000 10.525000 0.810000 ;
      RECT 10.485000  2.520000 10.735000 3.245000 ;
      RECT 10.640000  1.820000 10.970000 2.150000 ;
      RECT 10.945000  2.520000 11.310000 2.980000 ;
      RECT 11.010000  0.350000 11.340000 0.755000 ;
      RECT 11.010000  0.755000 11.735000 0.925000 ;
      RECT 11.065000  1.265000 11.395000 1.275000 ;
      RECT 11.140000  1.615000 11.310000 2.520000 ;
      RECT 11.480000  2.100000 11.810000 3.245000 ;
      RECT 11.565000  0.925000 11.735000 1.445000 ;
      RECT 11.570000  0.085000 11.905000 0.585000 ;
      RECT 11.980000  2.100000 12.310000 2.980000 ;
      RECT 12.085000  0.350000 12.335000 1.300000 ;
      RECT 12.085000  1.300000 12.870000 1.630000 ;
      RECT 12.085000  1.630000 12.310000 2.100000 ;
      RECT 12.540000  1.820000 12.870000 3.245000 ;
      RECT 12.565000  0.085000 12.815000 1.130000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  1.950000  4.165000 2.120000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  1.950000  8.005000 2.120000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  1.950000 10.885000 2.120000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
  END
END sky130_fd_sc_hs__sdfrtp_1
MACRO sky130_fd_sc_hs__sdfrtp_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.40000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 0.810000 2.100000 1.265000 ;
        RECT 1.605000 0.595000 2.100000 0.810000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.525000 0.350000 13.855000 1.410000 ;
        RECT 13.525000 1.410000 13.785000 2.980000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  3.935000 1.920000  4.225000 1.965000 ;
        RECT  3.935000 1.965000 11.425000 2.105000 ;
        RECT  3.935000 2.105000  4.225000 2.150000 ;
        RECT  8.255000 1.920000  8.545000 1.965000 ;
        RECT  8.255000 2.105000  8.545000 2.150000 ;
        RECT 11.135000 1.920000 11.425000 1.965000 ;
        RECT 11.135000 2.105000 11.425000 2.150000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.875000 2.000000 3.275000 2.175000 ;
        RECT 2.945000 1.440000 3.275000 2.000000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455000 1.490000 2.705000 1.660000 ;
        RECT 0.455000 1.660000 2.205000 1.835000 ;
        RECT 2.375000 1.260000 2.705000 1.490000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.785000 0.920000 4.060000 1.180000 ;
        RECT 3.785000 1.180000 4.195000 1.260000 ;
        RECT 3.785000 1.260000 4.645000 1.630000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 14.400000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 14.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.400000 0.085000 ;
      RECT  0.000000  3.245000 14.400000 3.415000 ;
      RECT  0.115000  0.350000  0.365000 0.935000 ;
      RECT  0.115000  0.935000  1.140000 1.265000 ;
      RECT  0.115000  1.265000  0.285000 2.005000 ;
      RECT  0.115000  2.005000  2.705000 2.175000 ;
      RECT  0.115000  2.175000  0.445000 2.980000 ;
      RECT  0.545000  0.085000  0.875000 0.765000 ;
      RECT  0.615000  2.345000  1.565000 3.245000 ;
      RECT  1.105000  0.255000  3.430000 0.425000 ;
      RECT  1.105000  0.425000  1.435000 0.640000 ;
      RECT  2.095000  2.345000  3.785000 2.385000 ;
      RECT  2.095000  2.385000  4.230000 2.400000 ;
      RECT  2.095000  2.400000  4.250000 2.420000 ;
      RECT  2.095000  2.420000  6.075000 2.515000 ;
      RECT  2.095000  2.515000  2.425000 2.980000 ;
      RECT  2.270000  0.595000  3.020000 0.810000 ;
      RECT  2.270000  0.810000  3.040000 0.835000 ;
      RECT  2.270000  0.835000  3.055000 0.845000 ;
      RECT  2.375000  1.830000  2.705000 2.005000 ;
      RECT  2.785000  0.845000  3.055000 0.855000 ;
      RECT  2.785000  0.855000  3.065000 0.865000 ;
      RECT  2.810000  0.865000  3.085000 0.880000 ;
      RECT  2.830000  0.880000  3.110000 0.890000 ;
      RECT  2.840000  0.890000  3.110000 0.900000 ;
      RECT  2.840000  0.900000  3.615000 0.910000 ;
      RECT  2.855000  0.910000  3.615000 0.935000 ;
      RECT  2.875000  0.935000  3.615000 1.270000 ;
      RECT  3.095000  2.685000  3.425000 3.245000 ;
      RECT  3.190000  0.425000  3.430000 0.730000 ;
      RECT  3.445000  1.270000  3.615000 2.330000 ;
      RECT  3.445000  2.330000  3.785000 2.345000 ;
      RECT  3.610000  0.085000  3.880000 0.730000 ;
      RECT  3.615000  2.515000  6.075000 2.580000 ;
      RECT  3.615000  2.580000  4.645000 2.585000 ;
      RECT  3.615000  2.585000  4.630000 2.590000 ;
      RECT  3.615000  2.590000  4.610000 2.600000 ;
      RECT  3.615000  2.600000  4.580000 2.620000 ;
      RECT  3.615000  2.620000  3.995000 2.980000 ;
      RECT  3.785000  1.830000  4.165000 2.160000 ;
      RECT  3.920000  2.160000  4.165000 2.190000 ;
      RECT  4.135000  0.500000  4.535000 0.750000 ;
      RECT  4.230000  0.750000  4.535000 0.790000 ;
      RECT  4.230000  0.790000  4.555000 0.815000 ;
      RECT  4.230000  0.815000  4.570000 0.835000 ;
      RECT  4.230000  0.835000  4.580000 0.845000 ;
      RECT  4.300000  0.845000  4.600000 0.860000 ;
      RECT  4.300000  0.860000  4.625000 0.865000 ;
      RECT  4.325000  0.865000  4.625000 0.880000 ;
      RECT  4.335000  1.820000  4.985000 2.195000 ;
      RECT  4.335000  2.195000  4.505000 2.250000 ;
      RECT  4.345000  0.880000  5.045000 0.890000 ;
      RECT  4.355000  0.890000  5.045000 0.910000 ;
      RECT  4.370000  0.910000  5.045000 0.935000 ;
      RECT  4.390000  0.935000  5.045000 1.080000 ;
      RECT  4.555000  2.415000  6.075000 2.420000 ;
      RECT  4.570000  2.410000  6.075000 2.415000 ;
      RECT  4.590000  2.400000  6.075000 2.410000 ;
      RECT  4.615000  2.385000  6.075000 2.400000 ;
      RECT  4.705000  0.085000  5.035000 0.710000 ;
      RECT  4.705000  2.750000  5.035000 3.245000 ;
      RECT  4.815000  1.080000  5.045000 1.455000 ;
      RECT  4.815000  1.455000  5.280000 1.775000 ;
      RECT  4.815000  1.775000  4.985000 1.820000 ;
      RECT  5.155000  1.955000  5.630000 2.215000 ;
      RECT  5.215000  0.255000  7.220000 0.425000 ;
      RECT  5.215000  0.425000  5.620000 1.070000 ;
      RECT  5.215000  1.070000  5.630000 1.285000 ;
      RECT  5.450000  1.285000  5.630000 1.545000 ;
      RECT  5.450000  1.545000  6.175000 1.875000 ;
      RECT  5.450000  1.875000  5.630000 1.955000 ;
      RECT  5.795000  0.595000  5.975000 0.995000 ;
      RECT  5.800000  0.995000  5.975000 1.200000 ;
      RECT  5.800000  1.200000  6.515000 1.370000 ;
      RECT  5.825000  2.045000  6.515000 2.215000 ;
      RECT  5.825000  2.215000  6.075000 2.385000 ;
      RECT  5.825000  2.580000  6.075000 2.725000 ;
      RECT  6.145000  0.595000  6.470000 0.860000 ;
      RECT  6.145000  0.860000  6.855000 1.030000 ;
      RECT  6.250000  2.385000  6.855000 2.725000 ;
      RECT  6.345000  1.370000  6.515000 2.045000 ;
      RECT  6.685000  1.030000  6.855000 1.985000 ;
      RECT  6.685000  1.985000  7.605000 2.165000 ;
      RECT  6.685000  2.165000  6.855000 2.385000 ;
      RECT  7.025000  0.920000  8.920000 1.090000 ;
      RECT  7.025000  1.090000  7.265000 1.805000 ;
      RECT  7.025000  2.345000  7.265000 3.245000 ;
      RECT  7.050000  0.425000  7.220000 0.580000 ;
      RECT  7.050000  0.580000  8.100000 0.750000 ;
      RECT  7.430000  0.085000  7.760000 0.410000 ;
      RECT  7.435000  1.260000  8.485000 1.545000 ;
      RECT  7.435000  1.545000  7.605000 1.985000 ;
      RECT  7.435000  2.165000  7.605000 2.320000 ;
      RECT  7.435000  2.320000  7.765000 2.745000 ;
      RECT  7.775000  1.795000  8.570000 2.150000 ;
      RECT  7.930000  0.255000  9.260000 0.425000 ;
      RECT  7.930000  0.425000  8.100000 0.580000 ;
      RECT  8.245000  2.330000  8.580000 3.245000 ;
      RECT  8.270000  0.595000  8.920000 0.920000 ;
      RECT  8.750000  1.090000  8.920000 1.715000 ;
      RECT  8.750000  1.715000  9.115000 2.755000 ;
      RECT  9.090000  0.425000  9.260000 1.005000 ;
      RECT  9.090000  1.005000 10.050000 1.335000 ;
      RECT  9.320000  1.840000  9.600000 2.520000 ;
      RECT  9.320000  2.520000 10.390000 2.850000 ;
      RECT  9.430000  0.480000 10.390000 0.810000 ;
      RECT  9.785000  1.335000 10.050000 2.330000 ;
      RECT 10.220000  0.810000 10.390000 1.030000 ;
      RECT 10.220000  1.030000 11.190000 1.110000 ;
      RECT 10.220000  1.110000 11.890000 1.200000 ;
      RECT 10.220000  1.200000 10.390000 2.520000 ;
      RECT 10.560000  1.370000 10.850000 1.580000 ;
      RECT 10.560000  1.580000 12.230000 1.750000 ;
      RECT 10.560000  1.750000 10.850000 2.390000 ;
      RECT 10.560000  2.390000 11.740000 2.560000 ;
      RECT 10.560000  2.730000 11.240000 3.245000 ;
      RECT 10.755000  0.085000 11.085000 0.810000 ;
      RECT 11.020000  1.200000 11.890000 1.410000 ;
      RECT 11.110000  1.920000 11.440000 2.220000 ;
      RECT 11.410000  2.560000 11.740000 2.980000 ;
      RECT 11.545000  0.350000 11.875000 0.770000 ;
      RECT 11.545000  0.770000 12.230000 0.940000 ;
      RECT 11.945000  1.940000 12.275000 3.245000 ;
      RECT 12.060000  0.940000 12.230000 1.580000 ;
      RECT 12.105000  0.085000 12.435000 0.600000 ;
      RECT 12.445000  1.940000 12.775000 2.980000 ;
      RECT 12.605000  0.350000 12.865000 1.300000 ;
      RECT 12.605000  1.300000 13.355000 1.630000 ;
      RECT 12.605000  1.630000 12.775000 1.940000 ;
      RECT 13.005000  1.820000 13.335000 3.245000 ;
      RECT 13.095000  0.085000 13.345000 1.130000 ;
      RECT 13.955000  1.820000 14.285000 3.245000 ;
      RECT 14.035000  0.085000 14.285000 1.130000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  1.950000  4.165000 2.120000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  1.950000  8.485000 2.120000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  1.950000 11.365000 2.120000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
  END
END sky130_fd_sc_hs__sdfrtp_2
MACRO sky130_fd_sc_hs__sdfrtp_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.88000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 0.810000 2.100000 1.265000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.535000 0.350000 12.865000 0.930000 ;
        RECT 12.535000 0.930000 14.255000 1.100000 ;
        RECT 13.085000 1.770000 14.755000 1.940000 ;
        RECT 13.085000 1.940000 13.415000 2.980000 ;
        RECT 14.065000 1.940000 14.280000 2.980000 ;
        RECT 14.085000 0.350000 14.255000 0.930000 ;
        RECT 14.085000 1.100000 14.255000 1.300000 ;
        RECT 14.085000 1.300000 14.755000 1.770000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  3.935000 1.920000  4.225000 1.965000 ;
        RECT  3.935000 1.965000 10.945000 2.105000 ;
        RECT  3.935000 2.105000  4.225000 2.150000 ;
        RECT  7.775000 1.920000  8.065000 1.965000 ;
        RECT  7.775000 2.105000  8.065000 2.150000 ;
        RECT 10.655000 1.920000 10.945000 1.965000 ;
        RECT 10.655000 2.105000 10.945000 2.150000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.945000 1.440000 3.275000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.490000 2.735000 1.660000 ;
        RECT 0.605000 1.660000 1.795000 1.835000 ;
        RECT 2.405000 1.260000 2.735000 1.490000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.840000 1.180000 4.195000 1.260000 ;
        RECT 3.840000 1.260000 4.635000 1.590000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 14.880000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 14.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.880000 0.085000 ;
      RECT  0.000000  3.245000 14.880000 3.415000 ;
      RECT  0.115000  0.350000  0.365000 0.935000 ;
      RECT  0.115000  0.935000  1.140000 1.265000 ;
      RECT  0.115000  1.265000  0.285000 2.005000 ;
      RECT  0.115000  2.005000  2.705000 2.175000 ;
      RECT  0.115000  2.175000  0.445000 2.980000 ;
      RECT  0.545000  0.085000  0.875000 0.765000 ;
      RECT  0.615000  2.345000  1.565000 3.245000 ;
      RECT  1.105000  0.255000  3.500000 0.425000 ;
      RECT  1.105000  0.425000  1.435000 0.640000 ;
      RECT  2.105000  2.345000  3.995000 2.420000 ;
      RECT  2.105000  2.420000  6.075000 2.515000 ;
      RECT  2.105000  2.515000  2.435000 2.980000 ;
      RECT  2.270000  0.595000  2.735000 0.845000 ;
      RECT  2.375000  1.830000  2.705000 2.005000 ;
      RECT  2.565000  0.845000  2.735000 0.920000 ;
      RECT  2.565000  0.920000  3.615000 1.090000 ;
      RECT  3.095000  2.685000  3.425000 3.245000 ;
      RECT  3.225000  0.425000  3.500000 0.750000 ;
      RECT  3.445000  1.090000  3.615000 2.330000 ;
      RECT  3.445000  2.330000  3.995000 2.345000 ;
      RECT  3.615000  2.515000  6.075000 2.580000 ;
      RECT  3.615000  2.580000  4.645000 2.590000 ;
      RECT  3.615000  2.590000  3.995000 2.980000 ;
      RECT  3.670000  0.085000  3.995000 0.750000 ;
      RECT  3.785000  1.830000  4.165000 2.160000 ;
      RECT  4.165000  0.550000  4.535000 0.750000 ;
      RECT  4.335000  1.820000  4.975000 1.990000 ;
      RECT  4.335000  1.990000  4.515000 2.250000 ;
      RECT  4.365000  0.750000  4.535000 0.920000 ;
      RECT  4.365000  0.920000  4.975000 1.090000 ;
      RECT  4.580000  2.410000  6.075000 2.420000 ;
      RECT  4.705000  2.750000  5.035000 3.245000 ;
      RECT  4.715000  0.085000  5.045000 0.750000 ;
      RECT  4.805000  1.090000  4.975000 1.410000 ;
      RECT  4.805000  1.410000  5.280000 1.740000 ;
      RECT  4.805000  1.740000  4.975000 1.820000 ;
      RECT  5.155000  1.910000  6.205000 1.915000 ;
      RECT  5.155000  1.915000  5.655000 2.240000 ;
      RECT  5.195000  0.920000  5.620000 1.240000 ;
      RECT  5.215000  0.330000  7.225000 0.500000 ;
      RECT  5.215000  0.500000  5.620000 0.920000 ;
      RECT  5.450000  1.240000  5.620000 1.585000 ;
      RECT  5.450000  1.585000  6.205000 1.910000 ;
      RECT  5.745000  2.580000  6.075000 2.755000 ;
      RECT  5.790000  0.670000  5.990000 1.245000 ;
      RECT  5.790000  1.245000  6.545000 1.415000 ;
      RECT  5.825000  2.085000  6.545000 2.255000 ;
      RECT  5.825000  2.255000  6.075000 2.410000 ;
      RECT  6.160000  0.670000  6.470000 0.905000 ;
      RECT  6.160000  0.905000  6.885000 1.075000 ;
      RECT  6.245000  2.425000  8.055000 2.490000 ;
      RECT  6.245000  2.490000  6.885000 2.755000 ;
      RECT  6.375000  1.415000  6.545000 2.085000 ;
      RECT  6.715000  1.075000  6.885000 2.320000 ;
      RECT  6.715000  2.320000  8.055000 2.425000 ;
      RECT  7.055000  0.500000  7.225000 0.580000 ;
      RECT  7.055000  0.580000  8.100000 0.750000 ;
      RECT  7.055000  0.920000  8.655000 1.090000 ;
      RECT  7.055000  1.090000  7.325000 1.945000 ;
      RECT  7.170000  2.660000  7.520000 3.245000 ;
      RECT  7.430000  0.085000  7.760000 0.410000 ;
      RECT  7.495000  1.260000  8.315000 1.575000 ;
      RECT  7.495000  1.575000  7.665000 2.320000 ;
      RECT  7.725000  2.490000  8.055000 2.755000 ;
      RECT  7.835000  1.820000  8.145000 2.150000 ;
      RECT  7.930000  0.255000  8.995000 0.425000 ;
      RECT  7.930000  0.425000  8.100000 0.580000 ;
      RECT  8.270000  0.595000  8.655000 0.920000 ;
      RECT  8.365000  1.745000  8.535000 3.245000 ;
      RECT  8.485000  1.090000  8.655000 1.405000 ;
      RECT  8.485000  1.405000  9.065000 1.575000 ;
      RECT  8.735000  1.575000  9.065000 2.755000 ;
      RECT  8.825000  0.425000  8.995000 0.905000 ;
      RECT  8.825000  0.905000  9.415000 1.235000 ;
      RECT  9.165000  0.405000  9.755000 0.735000 ;
      RECT  9.245000  1.235000  9.415000 2.065000 ;
      RECT  9.245000  2.065000  9.955000 2.380000 ;
      RECT  9.270000  2.550000 10.295000 2.880000 ;
      RECT  9.585000  0.735000  9.755000 0.885000 ;
      RECT  9.585000  0.885000 11.245000 1.055000 ;
      RECT  9.585000  1.055000  9.755000 1.725000 ;
      RECT  9.585000  1.725000 10.295000 1.895000 ;
      RECT 10.015000  1.225000 10.345000 1.385000 ;
      RECT 10.015000  1.385000 11.585000 1.555000 ;
      RECT 10.125000  1.895000 10.295000 2.550000 ;
      RECT 10.140000  0.085000 10.580000 0.680000 ;
      RECT 10.465000  2.520000 10.795000 3.245000 ;
      RECT 10.585000  1.820000 10.915000 2.150000 ;
      RECT 10.915000  1.055000 11.245000 1.215000 ;
      RECT 11.000000  2.520000 11.330000 2.980000 ;
      RECT 11.040000  0.385000 11.585000 0.715000 ;
      RECT 11.160000  1.555000 11.330000 2.520000 ;
      RECT 11.415000  0.715000 11.585000 1.385000 ;
      RECT 11.650000  1.820000 11.900000 3.245000 ;
      RECT 11.755000  0.350000 11.925000 1.270000 ;
      RECT 11.755000  1.270000 13.850000 1.600000 ;
      RECT 12.100000  1.600000 12.430000 2.700000 ;
      RECT 12.105000  0.085000 12.365000 1.100000 ;
      RECT 12.635000  1.820000 12.885000 3.245000 ;
      RECT 13.035000  0.085000 13.905000 0.760000 ;
      RECT 13.615000  2.110000 13.865000 3.245000 ;
      RECT 14.435000  0.085000 14.765000 1.130000 ;
      RECT 14.470000  2.110000 14.765000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  1.950000  4.165000 2.120000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  1.950000  8.005000 2.120000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  1.950000 10.885000 2.120000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
  END
END sky130_fd_sc_hs__sdfrtp_4
MACRO sky130_fd_sc_hs__sdfsbp_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.40000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.790000 1.585000 2.120000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.535700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.955000 0.350000 14.290000 2.980000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.535700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.125000 0.350000 12.620000 1.130000 ;
        RECT 12.450000 1.130000 12.620000 1.820000 ;
        RECT 12.450000 1.820000 12.705000 2.980000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555000 1.140000 2.765000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.505000 1.450000 2.045000 1.620000 ;
        RECT 0.505000 1.620000 0.835000 1.850000 ;
        RECT 1.795000 1.260000 2.045000 1.450000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAPARTIALMETALSIDEAREA  1.869000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 7.295000 1.550000 7.585000 1.595000 ;
        RECT 7.295000 1.595000 9.985000 1.735000 ;
        RECT 7.295000 1.735000 7.585000 1.780000 ;
        RECT 9.695000 1.550000 9.985000 1.595000 ;
        RECT 9.695000 1.735000 9.985000 1.780000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.275000 1.180000 3.715000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 14.400000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 14.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.400000 0.085000 ;
      RECT  0.000000  3.245000 14.400000 3.415000 ;
      RECT  0.115000  0.350000  0.445000 0.950000 ;
      RECT  0.115000  0.950000  1.140000 1.280000 ;
      RECT  0.115000  1.280000  0.335000 2.290000 ;
      RECT  0.115000  2.290000  2.045000 2.460000 ;
      RECT  0.115000  2.460000  0.365000 2.980000 ;
      RECT  0.565000  2.630000  0.895000 3.245000 ;
      RECT  0.615000  0.085000  0.945000 0.780000 ;
      RECT  1.435000  2.630000  2.385000 2.800000 ;
      RECT  1.435000  2.800000  1.945000 2.960000 ;
      RECT  1.505000  0.350000  1.835000 0.920000 ;
      RECT  1.505000  0.920000  2.385000 1.090000 ;
      RECT  1.795000  1.830000  2.045000 2.290000 ;
      RECT  2.215000  1.090000  2.385000 2.320000 ;
      RECT  2.215000  2.320000  4.925000 2.380000 ;
      RECT  2.215000  2.380000  3.795000 2.490000 ;
      RECT  2.215000  2.490000  2.385000 2.630000 ;
      RECT  2.325000  0.085000  2.655000 0.750000 ;
      RECT  2.555000  2.660000  2.820000 3.245000 ;
      RECT  2.935000  0.340000  3.200000 1.010000 ;
      RECT  2.935000  1.010000  3.105000 1.820000 ;
      RECT  2.935000  1.820000  4.215000 1.990000 ;
      RECT  2.935000  1.990000  3.455000 2.150000 ;
      RECT  3.380000  0.085000  3.710000 1.010000 ;
      RECT  3.575000  2.660000  3.905000 3.245000 ;
      RECT  3.625000  2.210000  4.925000 2.320000 ;
      RECT  3.880000  0.255000  5.030000 0.425000 ;
      RECT  3.880000  0.425000  4.210000 1.010000 ;
      RECT  3.885000  1.220000  4.215000 1.820000 ;
      RECT  4.105000  2.550000  4.355000 2.905000 ;
      RECT  4.105000  2.905000  5.810000 3.075000 ;
      RECT  4.420000  0.595000  4.690000 0.925000 ;
      RECT  4.420000  0.925000  4.590000 2.210000 ;
      RECT  4.590000  2.380000  4.925000 2.735000 ;
      RECT  4.760000  1.370000  5.030000 2.040000 ;
      RECT  4.860000  0.425000  5.030000 1.370000 ;
      RECT  5.120000  2.370000  5.450000 2.735000 ;
      RECT  5.200000  0.350000  5.450000 1.350000 ;
      RECT  5.200000  1.350000  7.110000 1.520000 ;
      RECT  5.200000  1.520000  5.370000 2.370000 ;
      RECT  5.540000  1.690000  5.810000 2.020000 ;
      RECT  5.640000  2.020000  5.810000 2.085000 ;
      RECT  5.640000  2.085000  6.765000 2.255000 ;
      RECT  5.640000  2.255000  5.810000 2.905000 ;
      RECT  5.815000  0.735000  6.770000 0.905000 ;
      RECT  5.815000  0.905000  6.485000 1.180000 ;
      RECT  6.020000  0.085000  6.370000 0.565000 ;
      RECT  6.050000  1.690000  7.105000 1.915000 ;
      RECT  6.175000  2.425000  6.425000 3.245000 ;
      RECT  6.595000  2.255000  6.765000 2.905000 ;
      RECT  6.595000  2.905000  7.445000 3.075000 ;
      RECT  6.600000  0.350000  6.930000 0.735000 ;
      RECT  6.725000  1.190000  7.110000 1.350000 ;
      RECT  6.935000  1.915000  7.105000 2.735000 ;
      RECT  6.940000  0.905000  8.165000 1.075000 ;
      RECT  6.940000  1.075000  7.110000 1.190000 ;
      RECT  7.275000  1.950000  8.830000 2.120000 ;
      RECT  7.275000  2.120000  7.445000 2.905000 ;
      RECT  7.295000  1.245000  7.625000 1.780000 ;
      RECT  7.500000  0.085000  8.295000 0.735000 ;
      RECT  7.615000  2.295000  7.785000 3.245000 ;
      RECT  7.835000  1.075000  8.165000 1.450000 ;
      RECT  7.985000  2.290000  8.315000 2.350000 ;
      RECT  7.985000  2.350000  9.830000 2.520000 ;
      RECT  7.985000  2.520000  8.315000 2.755000 ;
      RECT  8.530000  2.690000  8.860000 2.905000 ;
      RECT  8.530000  2.905000 10.380000 3.075000 ;
      RECT  8.660000  1.350000  8.990000 1.680000 ;
      RECT  8.660000  1.680000  8.830000 1.950000 ;
      RECT  8.785000  0.350000  9.380000 1.050000 ;
      RECT  9.045000  1.850000  9.380000 1.950000 ;
      RECT  9.045000  1.950000 10.170000 2.095000 ;
      RECT  9.045000  2.095000 11.280000 2.120000 ;
      RECT  9.045000  2.120000  9.380000 2.180000 ;
      RECT  9.210000  1.050000  9.380000 1.850000 ;
      RECT  9.580000  2.290000  9.830000 2.350000 ;
      RECT  9.580000  2.520000  9.830000 2.735000 ;
      RECT  9.620000  0.900000 11.395000 1.070000 ;
      RECT  9.620000  1.070000  9.950000 1.230000 ;
      RECT  9.725000  1.550000 10.915000 1.780000 ;
      RECT 10.000000  2.120000 11.280000 2.265000 ;
      RECT 10.050000  2.520000 10.380000 2.905000 ;
      RECT 10.285000  0.085000 10.895000 0.680000 ;
      RECT 10.580000  2.520000 10.750000 3.245000 ;
      RECT 10.585000  1.255000 10.915000 1.550000 ;
      RECT 10.585000  1.780000 10.915000 1.925000 ;
      RECT 10.950000  2.520000 11.280000 2.980000 ;
      RECT 11.065000  0.350000 11.395000 0.900000 ;
      RECT 11.110000  1.640000 11.895000 1.970000 ;
      RECT 11.110000  1.970000 11.280000 2.095000 ;
      RECT 11.110000  2.265000 11.280000 2.520000 ;
      RECT 11.225000  1.070000 11.395000 1.300000 ;
      RECT 11.225000  1.300000 12.235000 1.470000 ;
      RECT 11.500000  2.180000 12.235000 2.350000 ;
      RECT 11.500000  2.350000 11.750000 2.980000 ;
      RECT 11.625000  0.085000 11.955000 1.130000 ;
      RECT 11.950000  2.520000 12.280000 3.245000 ;
      RECT 12.065000  1.470000 12.235000 2.180000 ;
      RECT 12.840000  0.540000 13.255000 1.130000 ;
      RECT 13.005000  1.130000 13.255000 1.220000 ;
      RECT 13.005000  1.220000 13.785000 1.550000 ;
      RECT 13.005000  1.550000 13.255000 2.875000 ;
      RECT 13.455000  0.085000 13.785000 1.050000 ;
      RECT 13.455000  1.995000 13.785000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  1.580000  7.525000 1.750000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  1.580000  9.925000 1.750000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
  END
END sky130_fd_sc_hs__sdfsbp_1
MACRO sky130_fd_sc_hs__sdfsbp_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  17.76000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.385000 0.440000 1.795000 1.230000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.865000 1.820000 17.225000 2.980000 ;
        RECT 16.885000 0.350000 17.225000 1.130000 ;
        RECT 17.055000 1.130000 17.225000 1.820000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.558000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.850000 0.350000 15.235000 1.410000 ;
        RECT 14.850000 1.410000 15.105000 2.980000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.805000 0.950000 3.205000 1.620000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.400000 2.295000 1.570000 ;
        RECT 0.425000 1.570000 1.085000 1.800000 ;
        RECT 1.965000 0.900000 2.295000 1.400000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAPARTIALMETALSIDEAREA  3.885000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  7.775000 1.550000  8.065000 1.595000 ;
        RECT  7.775000 1.595000 13.345000 1.735000 ;
        RECT  7.775000 1.735000  8.065000 1.780000 ;
        RECT 13.055000 1.550000 13.345000 1.595000 ;
        RECT 13.055000 1.735000 13.345000 1.780000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.715000 1.180000 4.195000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 17.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 17.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 17.760000 0.085000 ;
      RECT  0.000000  3.245000 17.760000 3.415000 ;
      RECT  0.085000  0.350000  0.445000 0.900000 ;
      RECT  0.085000  0.900000  1.145000 1.230000 ;
      RECT  0.085000  1.230000  0.255000 1.970000 ;
      RECT  0.085000  1.970000  2.105000 2.140000 ;
      RECT  0.085000  2.140000  0.465000 2.980000 ;
      RECT  0.615000  0.085000  1.020000 0.680000 ;
      RECT  0.635000  2.310000  0.965000 3.245000 ;
      RECT  1.505000  2.310000  3.885000 2.480000 ;
      RECT  1.505000  2.480000  1.955000 2.980000 ;
      RECT  1.775000  1.810000  2.105000 1.970000 ;
      RECT  1.965000  0.400000  2.350000 0.560000 ;
      RECT  1.965000  0.560000  2.635000 0.730000 ;
      RECT  2.465000  0.730000  2.635000 2.310000 ;
      RECT  2.495000  2.650000  2.845000 3.245000 ;
      RECT  2.840000  0.085000  3.170000 0.780000 ;
      RECT  3.075000  1.790000  4.720000 1.960000 ;
      RECT  3.075000  1.960000  3.545000 2.140000 ;
      RECT  3.375000  0.340000  3.650000 1.010000 ;
      RECT  3.375000  1.010000  3.545000 1.790000 ;
      RECT  3.525000  2.650000  4.220000 3.245000 ;
      RECT  3.715000  2.130000  5.370000 2.300000 ;
      RECT  3.715000  2.300000  3.885000 2.310000 ;
      RECT  3.830000  0.085000  4.160000 1.010000 ;
      RECT  4.330000  0.255000  5.560000 0.425000 ;
      RECT  4.330000  0.425000  4.660000 1.010000 ;
      RECT  4.390000  1.350000  4.720000 1.790000 ;
      RECT  4.390000  2.470000  4.720000 2.905000 ;
      RECT  4.390000  2.905000  6.240000 3.075000 ;
      RECT  4.890000  0.595000  5.220000 0.845000 ;
      RECT  4.890000  0.845000  5.060000 2.130000 ;
      RECT  4.890000  2.300000  5.370000 2.735000 ;
      RECT  5.230000  1.290000  5.560000 1.960000 ;
      RECT  5.390000  0.425000  5.560000 1.290000 ;
      RECT  5.540000  2.295000  5.900000 2.735000 ;
      RECT  5.730000  0.470000  6.645000 0.800000 ;
      RECT  5.730000  0.800000  5.900000 2.295000 ;
      RECT  6.070000  0.970000  6.305000 2.165000 ;
      RECT  6.070000  2.165000  7.325000 2.335000 ;
      RECT  6.070000  2.335000  6.240000 2.905000 ;
      RECT  6.410000  2.505000  6.985000 3.245000 ;
      RECT  6.475000  0.800000  6.645000 1.395000 ;
      RECT  6.475000  1.395000  7.665000 1.565000 ;
      RECT  6.635000  1.735000  7.665000 1.995000 ;
      RECT  6.815000  0.085000  7.150000 0.700000 ;
      RECT  6.815000  0.870000  7.710000 1.040000 ;
      RECT  6.815000  1.040000  7.145000 1.225000 ;
      RECT  7.155000  2.335000  7.325000 2.905000 ;
      RECT  7.155000  2.905000  8.165000 3.075000 ;
      RECT  7.355000  1.210000  8.050000 1.380000 ;
      RECT  7.355000  1.380000  7.665000 1.395000 ;
      RECT  7.380000  0.350000  7.710000 0.870000 ;
      RECT  7.495000  1.995000  7.665000 2.295000 ;
      RECT  7.495000  2.295000  7.825000 2.735000 ;
      RECT  7.835000  1.550000  8.225000 1.880000 ;
      RECT  7.880000  0.900000  8.860000 1.175000 ;
      RECT  7.880000  1.175000  8.050000 1.210000 ;
      RECT  7.995000  2.050000  8.565000 2.220000 ;
      RECT  7.995000  2.220000  8.165000 2.905000 ;
      RECT  8.200000  0.085000  8.530000 0.680000 ;
      RECT  8.335000  2.390000  8.665000 3.245000 ;
      RECT  8.395000  1.345000 11.390000 1.515000 ;
      RECT  8.395000  1.515000  8.565000 2.050000 ;
      RECT  8.735000  1.685000  9.065000 1.700000 ;
      RECT  8.735000  1.700000 12.050000 1.870000 ;
      RECT  8.735000  1.870000  9.065000 1.960000 ;
      RECT  8.925000  2.130000 10.125000 2.300000 ;
      RECT  8.925000  2.300000  9.255000 2.980000 ;
      RECT  9.030000  0.350000  9.280000 1.005000 ;
      RECT  9.030000  1.005000 10.210000 1.175000 ;
      RECT  9.425000  2.470000  9.675000 3.245000 ;
      RECT  9.450000  0.085000  9.780000 0.835000 ;
      RECT  9.875000  2.100000 10.125000 2.130000 ;
      RECT  9.875000  2.300000 10.125000 2.905000 ;
      RECT  9.875000  2.905000 11.105000 3.075000 ;
      RECT  9.960000  0.255000 11.210000 0.425000 ;
      RECT  9.960000  0.425000 10.210000 1.005000 ;
      RECT 10.325000  2.040000 12.390000 2.140000 ;
      RECT 10.325000  2.140000 13.975000 2.210000 ;
      RECT 10.325000  2.210000 10.575000 2.700000 ;
      RECT 10.380000  0.595000 10.710000 0.860000 ;
      RECT 10.380000  0.860000 11.550000 1.030000 ;
      RECT 10.380000  1.200000 11.390000 1.345000 ;
      RECT 10.380000  1.515000 11.390000 1.530000 ;
      RECT 10.775000  2.380000 11.105000 2.905000 ;
      RECT 10.880000  0.425000 11.210000 0.690000 ;
      RECT 11.365000  2.385000 11.620000 2.885000 ;
      RECT 11.365000  2.885000 12.740000 3.055000 ;
      RECT 11.380000  0.400000 12.390000 0.730000 ;
      RECT 11.380000  0.730000 11.550000 0.860000 ;
      RECT 11.720000  0.900000 12.050000 1.700000 ;
      RECT 11.820000  2.210000 13.975000 2.310000 ;
      RECT 11.820000  2.310000 12.220000 2.715000 ;
      RECT 12.220000  0.730000 12.390000 2.040000 ;
      RECT 12.410000  2.520000 12.740000 2.885000 ;
      RECT 12.565000  0.960000 14.315000 1.130000 ;
      RECT 12.565000  1.130000 12.895000 1.960000 ;
      RECT 12.940000  2.520000 13.110000 3.245000 ;
      RECT 13.085000  1.300000 13.435000 1.970000 ;
      RECT 13.260000  0.085000 13.590000 0.790000 ;
      RECT 13.310000  2.310000 13.640000 2.980000 ;
      RECT 13.645000  1.300000 13.975000 2.140000 ;
      RECT 13.770000  0.350000 14.100000 0.960000 ;
      RECT 13.870000  2.480000 14.315000 2.910000 ;
      RECT 14.145000  1.130000 14.315000 2.480000 ;
      RECT 14.350000  0.085000 14.680000 0.790000 ;
      RECT 14.485000  1.820000 14.655000 3.245000 ;
      RECT 15.305000  1.820000 15.635000 3.245000 ;
      RECT 15.405000  0.085000 15.655000 1.130000 ;
      RECT 15.865000  0.450000 16.220000 1.300000 ;
      RECT 15.865000  1.300000 16.885000 1.630000 ;
      RECT 15.865000  1.630000 16.195000 2.860000 ;
      RECT 16.415000  1.820000 16.665000 3.245000 ;
      RECT 16.455000  0.085000 16.705000 1.130000 ;
      RECT 17.395000  0.085000 17.645000 1.130000 ;
      RECT 17.395000  1.820000 17.645000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  1.580000  8.005000 1.750000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  1.580000 13.285000 1.750000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.245000 15.205000 3.415000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.245000 15.685000 3.415000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.245000 16.165000 3.415000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  3.245000 16.645000 3.415000 ;
      RECT 16.955000 -0.085000 17.125000 0.085000 ;
      RECT 16.955000  3.245000 17.125000 3.415000 ;
      RECT 17.435000 -0.085000 17.605000 0.085000 ;
      RECT 17.435000  3.245000 17.605000 3.415000 ;
  END
END sky130_fd_sc_hs__sdfsbp_2
MACRO sky130_fd_sc_hs__sdfstp_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.92000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.820000 1.580000 2.150000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.530100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.380000 0.350000 13.815000 1.050000 ;
        RECT 13.565000 1.050000 13.815000 2.980000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555000 1.140000 2.805000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.280000 0.680000 1.440000 ;
        RECT 0.425000 1.440000 2.045000 1.610000 ;
        RECT 0.425000 1.610000 0.835000 1.950000 ;
        RECT 1.790000 1.260000 2.045000 1.440000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAPARTIALMETALSIDEAREA  2.541000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  7.295000 1.550000  7.585000 1.595000 ;
        RECT  7.295000 1.595000 10.945000 1.735000 ;
        RECT  7.295000 1.735000  7.585000 1.780000 ;
        RECT 10.655000 1.550000 10.945000 1.595000 ;
        RECT 10.655000 1.735000 10.945000 1.780000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.315000 1.180000 3.715000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 13.920000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 13.920000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.920000 0.085000 ;
      RECT  0.000000  3.245000 13.920000 3.415000 ;
      RECT  0.085000  0.350000  0.525000 0.940000 ;
      RECT  0.085000  0.940000  1.220000 1.110000 ;
      RECT  0.085000  1.110000  0.255000 2.300000 ;
      RECT  0.085000  2.300000  0.360000 2.320000 ;
      RECT  0.085000  2.320000  2.045000 2.490000 ;
      RECT  0.085000  2.490000  0.360000 2.980000 ;
      RECT  0.560000  2.660000  0.890000 3.245000 ;
      RECT  0.695000  0.085000  1.025000 0.770000 ;
      RECT  0.890000  1.110000  1.220000 1.270000 ;
      RECT  1.430000  2.660000  2.385000 2.910000 ;
      RECT  1.555000  0.350000  1.885000 0.920000 ;
      RECT  1.555000  0.920000  2.385000 1.090000 ;
      RECT  1.790000  1.830000  2.045000 2.320000 ;
      RECT  2.215000  1.090000  2.385000 2.490000 ;
      RECT  2.215000  2.490000  3.405000 2.660000 ;
      RECT  2.375000  0.085000  2.705000 0.750000 ;
      RECT  2.565000  2.830000  2.895000 3.245000 ;
      RECT  2.975000  0.350000  3.305000 1.010000 ;
      RECT  2.975000  1.010000  3.145000 1.820000 ;
      RECT  2.975000  1.820000  4.215000 2.070000 ;
      RECT  3.235000  2.240000  5.005000 2.410000 ;
      RECT  3.235000  2.410000  3.405000 2.490000 ;
      RECT  3.475000  0.085000  3.805000 1.010000 ;
      RECT  3.575000  2.580000  3.905000 3.245000 ;
      RECT  3.885000  1.350000  4.215000 1.820000 ;
      RECT  3.975000  0.255000  5.205000 0.425000 ;
      RECT  3.975000  0.425000  4.225000 1.130000 ;
      RECT  4.105000  2.580000  4.275000 2.895000 ;
      RECT  4.105000  2.895000  5.845000 3.065000 ;
      RECT  4.445000  0.595000  4.865000 0.765000 ;
      RECT  4.445000  0.765000  4.615000 2.240000 ;
      RECT  4.445000  2.410000  5.005000 2.725000 ;
      RECT  4.785000  0.935000  5.205000 1.105000 ;
      RECT  4.785000  1.105000  5.005000 2.070000 ;
      RECT  5.035000  0.425000  5.205000 0.935000 ;
      RECT  5.175000  1.275000  6.070000 1.435000 ;
      RECT  5.175000  1.435000  6.935000 1.445000 ;
      RECT  5.175000  1.445000  5.345000 2.265000 ;
      RECT  5.175000  2.265000  5.505000 2.725000 ;
      RECT  5.375000  0.385000  5.625000 1.275000 ;
      RECT  5.515000  1.615000  5.730000 1.775000 ;
      RECT  5.515000  1.775000  5.845000 1.945000 ;
      RECT  5.675000  1.945000  5.845000 2.345000 ;
      RECT  5.675000  2.345000  6.815000 2.515000 ;
      RECT  5.675000  2.515000  5.845000 2.895000 ;
      RECT  5.900000  1.445000  6.935000 1.605000 ;
      RECT  6.015000  1.795000  6.345000 2.005000 ;
      RECT  6.015000  2.005000  7.155000 2.175000 ;
      RECT  6.115000  0.085000  6.445000 0.690000 ;
      RECT  6.225000  2.685000  6.475000 3.245000 ;
      RECT  6.240000  0.860000  7.005000 1.030000 ;
      RECT  6.240000  1.030000  6.480000 1.265000 ;
      RECT  6.645000  2.515000  6.815000 2.895000 ;
      RECT  6.645000  2.895000  7.495000 3.065000 ;
      RECT  6.650000  1.200000  8.430000 1.370000 ;
      RECT  6.650000  1.370000  6.935000 1.435000 ;
      RECT  6.650000  1.605000  6.935000 1.835000 ;
      RECT  6.675000  0.570000  7.005000 0.860000 ;
      RECT  6.985000  2.175000  7.155000 2.725000 ;
      RECT  7.145000  1.540000  7.555000 1.800000 ;
      RECT  7.325000  1.970000  7.945000 2.140000 ;
      RECT  7.325000  2.140000  7.495000 2.895000 ;
      RECT  7.455000  0.085000  8.305000 0.940000 ;
      RECT  7.665000  2.310000  7.915000 3.245000 ;
      RECT  7.760000  1.120000  8.430000 1.200000 ;
      RECT  7.760000  1.370000  8.430000 1.410000 ;
      RECT  7.775000  1.580000  8.840000 1.750000 ;
      RECT  7.775000  1.750000  7.945000 1.970000 ;
      RECT  8.115000  1.920000  8.365000 2.350000 ;
      RECT  8.115000  2.350000  9.895000 2.520000 ;
      RECT  8.115000  2.520000  8.365000 2.725000 ;
      RECT  8.585000  2.690000  8.915000 2.905000 ;
      RECT  8.585000  2.905000 10.430000 3.075000 ;
      RECT  8.670000  1.120000  9.000000 1.450000 ;
      RECT  8.670000  1.450000  8.840000 1.580000 ;
      RECT  8.795000  0.350000  9.365000 0.940000 ;
      RECT  9.090000  1.620000 10.235000 1.790000 ;
      RECT  9.090000  1.790000  9.365000 2.180000 ;
      RECT  9.195000  0.940000  9.365000 1.620000 ;
      RECT  9.565000  1.960000  9.895000 2.350000 ;
      RECT  9.565000  2.520000  9.895000 2.735000 ;
      RECT  9.790000  0.980000 11.770000 1.040000 ;
      RECT  9.790000  1.040000 11.940000 1.210000 ;
      RECT  9.790000  1.210000 10.460000 1.310000 ;
      RECT 10.065000  1.790000 10.235000 2.220000 ;
      RECT 10.065000  2.220000 11.370000 2.390000 ;
      RECT 10.100000  2.560000 10.430000 2.905000 ;
      RECT 10.630000  2.560000 10.800000 3.245000 ;
      RECT 10.685000  1.380000 11.030000 2.050000 ;
      RECT 10.825000  0.085000 11.155000 0.810000 ;
      RECT 11.000000  2.390000 11.370000 2.980000 ;
      RECT 11.200000  1.380000 11.600000 2.050000 ;
      RECT 11.200000  2.050000 11.370000 2.220000 ;
      RECT 11.395000  0.350000 11.770000 0.980000 ;
      RECT 11.540000  2.220000 11.940000 2.390000 ;
      RECT 11.540000  2.390000 11.870000 2.980000 ;
      RECT 11.770000  1.210000 11.940000 2.220000 ;
      RECT 11.955000  0.540000 12.700000 0.870000 ;
      RECT 12.070000  2.560000 12.320000 3.245000 ;
      RECT 12.370000  0.870000 12.700000 1.005000 ;
      RECT 12.530000  1.005000 12.700000 1.220000 ;
      RECT 12.530000  1.220000 13.395000 1.550000 ;
      RECT 12.530000  1.550000 12.700000 1.995000 ;
      RECT 12.530000  1.995000 12.860000 2.875000 ;
      RECT 12.880000  0.085000 13.210000 1.050000 ;
      RECT 13.030000  1.995000 13.360000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  1.580000  7.525000 1.750000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  1.580000 10.885000 1.750000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
  END
END sky130_fd_sc_hs__sdfstp_1
MACRO sky130_fd_sc_hs__sdfstp_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.88000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.820000 1.585000 2.150000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.990000 0.370000 14.345000 1.150000 ;
        RECT 13.995000 1.820000 14.755000 2.150000 ;
        RECT 13.995000 2.150000 14.275000 2.980000 ;
        RECT 14.175000 1.150000 14.345000 1.320000 ;
        RECT 14.175000 1.320000 14.755000 1.490000 ;
        RECT 14.325000 1.490000 14.755000 1.820000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555000 1.140000 2.780000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.475000 1.410000 2.045000 1.580000 ;
        RECT 0.475000 1.580000 0.805000 2.140000 ;
        RECT 1.795000 1.250000 2.045000 1.410000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAPARTIALMETALSIDEAREA  3.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  7.295000 1.180000  7.585000 1.225000 ;
        RECT  7.295000 1.225000 11.905000 1.365000 ;
        RECT  7.295000 1.365000  7.585000 1.410000 ;
        RECT 11.615000 1.180000 11.905000 1.225000 ;
        RECT 11.615000 1.365000 11.905000 1.410000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.300000 1.180000 3.715000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 14.880000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 14.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.880000 0.085000 ;
      RECT  0.000000  3.245000 14.880000 3.415000 ;
      RECT  0.115000  0.350000  0.445000 0.900000 ;
      RECT  0.115000  0.900000  1.225000 1.230000 ;
      RECT  0.115000  1.230000  0.285000 2.310000 ;
      RECT  0.115000  2.310000  0.365000 2.320000 ;
      RECT  0.115000  2.320000  2.045000 2.490000 ;
      RECT  0.115000  2.490000  0.365000 2.980000 ;
      RECT  0.565000  2.660000  0.895000 3.245000 ;
      RECT  0.615000  0.085000  1.070000 0.680000 ;
      RECT  1.435000  2.660000  2.385000 2.910000 ;
      RECT  1.560000  0.350000  1.890000 0.910000 ;
      RECT  1.560000  0.910000  2.385000 1.080000 ;
      RECT  1.795000  1.830000  2.045000 2.320000 ;
      RECT  2.215000  1.080000  2.385000 2.490000 ;
      RECT  2.215000  2.490000  3.120000 2.660000 ;
      RECT  2.460000  0.085000  2.790000 0.740000 ;
      RECT  2.560000  2.830000  2.890000 3.245000 ;
      RECT  2.950000  2.240000  4.915000 2.410000 ;
      RECT  2.950000  2.410000  3.120000 2.490000 ;
      RECT  2.960000  0.350000  3.350000 1.010000 ;
      RECT  2.960000  1.010000  3.130000 1.820000 ;
      RECT  2.960000  1.820000  4.215000 2.070000 ;
      RECT  3.520000  0.085000  3.850000 1.010000 ;
      RECT  3.545000  2.580000  3.875000 3.245000 ;
      RECT  3.885000  1.350000  4.215000 1.820000 ;
      RECT  4.030000  0.255000  5.170000 0.425000 ;
      RECT  4.030000  0.425000  4.200000 1.130000 ;
      RECT  4.075000  2.580000  4.325000 2.895000 ;
      RECT  4.075000  2.895000  5.730000 3.065000 ;
      RECT  4.420000  0.595000  4.830000 0.845000 ;
      RECT  4.420000  0.845000  4.590000 1.900000 ;
      RECT  4.420000  1.900000  4.915000 2.070000 ;
      RECT  4.585000  2.070000  4.915000 2.240000 ;
      RECT  4.585000  2.410000  4.915000 2.725000 ;
      RECT  4.760000  1.015000  5.170000 1.185000 ;
      RECT  4.760000  1.185000  4.965000 1.730000 ;
      RECT  5.000000  0.425000  5.170000 1.015000 ;
      RECT  5.115000  2.265000  5.365000 2.725000 ;
      RECT  5.135000  1.375000  6.880000 1.545000 ;
      RECT  5.135000  1.545000  5.305000 2.265000 ;
      RECT  5.340000  0.385000  5.590000 1.375000 ;
      RECT  5.475000  1.715000  5.730000 2.045000 ;
      RECT  5.560000  2.045000  5.730000 2.085000 ;
      RECT  5.560000  2.085000  6.685000 2.255000 ;
      RECT  5.560000  2.255000  5.730000 2.895000 ;
      RECT  5.940000  1.715000  6.270000 1.745000 ;
      RECT  5.940000  1.745000  7.025000 1.915000 ;
      RECT  5.980000  0.530000  7.020000 0.700000 ;
      RECT  5.980000  0.700000  6.310000 1.205000 ;
      RECT  6.095000  2.425000  6.345000 3.245000 ;
      RECT  6.130000  0.085000  6.460000 0.360000 ;
      RECT  6.515000  2.255000  6.685000 2.905000 ;
      RECT  6.515000  2.905000  7.365000 3.075000 ;
      RECT  6.550000  0.870000  7.925000 1.040000 ;
      RECT  6.550000  1.040000  6.880000 1.375000 ;
      RECT  6.550000  1.545000  6.880000 1.570000 ;
      RECT  6.690000  0.350000  7.020000 0.530000 ;
      RECT  6.855000  1.915000  7.025000 2.735000 ;
      RECT  7.195000  1.725000 10.170000 1.805000 ;
      RECT  7.195000  1.805000  8.425000 1.895000 ;
      RECT  7.195000  1.895000  7.365000 2.905000 ;
      RECT  7.205000  1.210000  7.555000 1.555000 ;
      RECT  7.510000  0.085000  8.010000 0.680000 ;
      RECT  7.535000  2.065000  7.705000 3.245000 ;
      RECT  7.755000  1.040000  7.925000 1.225000 ;
      RECT  7.755000  1.225000  8.085000 1.555000 ;
      RECT  7.905000  2.065000  9.830000 2.145000 ;
      RECT  7.905000  2.145000  8.765000 2.235000 ;
      RECT  7.905000  2.235000  8.235000 2.755000 ;
      RECT  8.180000  0.350000  8.510000 0.885000 ;
      RECT  8.180000  0.885000 10.080000 1.055000 ;
      RECT  8.255000  1.475000 10.170000 1.725000 ;
      RECT  8.435000  2.405000  8.685000 3.245000 ;
      RECT  8.595000  1.975000  9.830000 2.065000 ;
      RECT  8.690000  0.085000  9.020000 0.715000 ;
      RECT  9.000000  2.315000  9.330000 2.905000 ;
      RECT  9.000000  2.905000 10.435000 3.075000 ;
      RECT  9.250000  0.255000 10.580000 0.425000 ;
      RECT  9.250000  0.425000  9.580000 0.715000 ;
      RECT  9.500000  2.145000  9.830000 2.735000 ;
      RECT  9.750000  0.595000 10.080000 0.885000 ;
      RECT 10.000000  1.805000 10.720000 2.135000 ;
      RECT 10.105000  2.305000 11.860000 2.475000 ;
      RECT 10.105000  2.475000 10.435000 2.905000 ;
      RECT 10.250000  0.425000 10.580000 0.810000 ;
      RECT 10.410000  0.810000 10.580000 1.400000 ;
      RECT 10.410000  1.400000 11.060000 1.570000 ;
      RECT 10.890000  1.570000 11.060000 1.970000 ;
      RECT 10.890000  1.970000 12.465000 2.140000 ;
      RECT 10.890000  2.140000 11.860000 2.305000 ;
      RECT 10.945000  0.790000 12.805000 0.960000 ;
      RECT 10.945000  0.960000 11.275000 1.230000 ;
      RECT 11.080000  2.645000 11.330000 3.245000 ;
      RECT 11.445000  1.180000 11.875000 1.800000 ;
      RECT 11.530000  2.475000 11.860000 2.980000 ;
      RECT 11.640000  0.085000 12.330000 0.600000 ;
      RECT 12.060000  2.310000 12.805000 2.480000 ;
      RECT 12.060000  2.480000 12.310000 2.980000 ;
      RECT 12.135000  1.130000 12.465000 1.970000 ;
      RECT 12.500000  0.350000 12.805000 0.790000 ;
      RECT 12.510000  2.650000 12.840000 3.245000 ;
      RECT 12.635000  0.960000 12.805000 2.310000 ;
      RECT 13.035000  0.470000 13.365000 1.320000 ;
      RECT 13.035000  1.320000 14.005000 1.650000 ;
      RECT 13.035000  1.650000 13.370000 2.980000 ;
      RECT 13.540000  1.820000 13.825000 3.245000 ;
      RECT 13.555000  0.085000 13.805000 1.150000 ;
      RECT 14.445000  2.320000 14.775000 3.245000 ;
      RECT 14.515000  0.085000 14.765000 1.150000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  1.210000  7.525000 1.380000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  1.210000 11.845000 1.380000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
  END
END sky130_fd_sc_hs__sdfstp_2
MACRO sky130_fd_sc_hs__sdfstp_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  15.84000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.105000 1.820000 1.575000 2.150000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.201100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.895000 0.350000 14.225000 0.980000 ;
        RECT 13.895000 0.980000 15.225000 1.150000 ;
        RECT 14.045000 1.820000 15.195000 2.150000 ;
        RECT 14.045000 2.150000 14.325000 2.980000 ;
        RECT 14.895000 0.350000 15.225000 0.980000 ;
        RECT 14.895000 1.150000 15.225000 1.270000 ;
        RECT 14.895000 1.270000 15.715000 1.440000 ;
        RECT 15.025000 1.610000 15.715000 1.780000 ;
        RECT 15.025000 1.780000 15.195000 1.820000 ;
        RECT 15.025000 2.150000 15.195000 2.980000 ;
        RECT 15.485000 1.440000 15.715000 1.610000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555000 1.100000 2.835000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525000 1.410000 2.045000 1.580000 ;
        RECT 0.525000 1.580000 0.855000 2.150000 ;
        RECT 1.715000 1.250000 2.045000 1.410000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAPARTIALMETALSIDEAREA  3.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  7.295000 1.550000  7.585000 1.595000 ;
        RECT  7.295000 1.595000 11.905000 1.735000 ;
        RECT  7.295000 1.735000  7.585000 1.780000 ;
        RECT 11.615000 1.550000 11.905000 1.595000 ;
        RECT 11.615000 1.735000 11.905000 1.780000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.345000 1.180000 3.715000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 15.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 15.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 15.840000 0.085000 ;
      RECT  0.000000  3.245000 15.840000 3.415000 ;
      RECT  0.105000  0.350000  0.445000 0.910000 ;
      RECT  0.105000  0.910000  1.140000 1.240000 ;
      RECT  0.105000  1.240000  0.355000 2.320000 ;
      RECT  0.105000  2.320000  2.045000 2.490000 ;
      RECT  0.105000  2.490000  0.355000 2.980000 ;
      RECT  0.555000  2.660000  0.885000 3.245000 ;
      RECT  0.615000  0.085000  0.945000 0.740000 ;
      RECT  1.425000  2.660000  2.385000 2.910000 ;
      RECT  1.475000  0.410000  1.960000 0.740000 ;
      RECT  1.785000  1.830000  2.045000 2.320000 ;
      RECT  1.790000  0.740000  1.960000 0.910000 ;
      RECT  1.790000  0.910000  2.385000 1.080000 ;
      RECT  2.215000  1.080000  2.385000 2.490000 ;
      RECT  2.215000  2.490000  3.175000 2.660000 ;
      RECT  2.450000  0.085000  2.780000 0.740000 ;
      RECT  2.560000  2.830000  2.890000 3.245000 ;
      RECT  3.005000  0.350000  3.390000 1.010000 ;
      RECT  3.005000  1.010000  3.175000 1.820000 ;
      RECT  3.005000  1.820000  4.215000 2.070000 ;
      RECT  3.005000  2.240000  5.030000 2.410000 ;
      RECT  3.005000  2.410000  3.175000 2.490000 ;
      RECT  3.560000  0.085000  3.890000 1.010000 ;
      RECT  3.570000  2.580000  3.900000 3.245000 ;
      RECT  3.885000  1.350000  4.215000 1.820000 ;
      RECT  4.070000  0.255000  5.140000 0.425000 ;
      RECT  4.070000  0.425000  4.240000 1.130000 ;
      RECT  4.070000  2.580000  4.400000 2.895000 ;
      RECT  4.070000  2.895000  5.830000 3.065000 ;
      RECT  4.410000  0.595000  4.800000 0.925000 ;
      RECT  4.410000  0.925000  4.580000 1.900000 ;
      RECT  4.410000  1.900000  5.030000 2.240000 ;
      RECT  4.700000  2.410000  5.030000 2.725000 ;
      RECT  4.750000  1.095000  5.140000 1.265000 ;
      RECT  4.750000  1.265000  5.030000 1.730000 ;
      RECT  4.970000  0.425000  5.140000 1.095000 ;
      RECT  5.200000  1.435000  6.955000 1.605000 ;
      RECT  5.200000  1.605000  5.370000 2.275000 ;
      RECT  5.200000  2.275000  5.480000 2.725000 ;
      RECT  5.310000  0.385000  5.640000 1.435000 ;
      RECT  5.540000  1.775000  5.830000 2.105000 ;
      RECT  5.660000  2.105000  5.830000 2.290000 ;
      RECT  5.660000  2.290000  6.865000 2.460000 ;
      RECT  5.660000  2.460000  5.830000 2.895000 ;
      RECT  6.005000  0.770000  7.100000 0.940000 ;
      RECT  6.005000  0.940000  6.335000 1.265000 ;
      RECT  6.040000  1.780000  6.370000 1.950000 ;
      RECT  6.040000  1.950000  7.205000 2.120000 ;
      RECT  6.210000  0.085000  6.540000 0.600000 ;
      RECT  6.275000  2.630000  6.525000 3.245000 ;
      RECT  6.625000  1.110000  8.265000 1.280000 ;
      RECT  6.625000  1.280000  6.955000 1.435000 ;
      RECT  6.625000  1.605000  6.955000 1.780000 ;
      RECT  6.695000  2.460000  6.865000 2.895000 ;
      RECT  6.695000  2.895000  7.545000 3.065000 ;
      RECT  6.770000  0.350000  7.100000 0.770000 ;
      RECT  7.035000  2.120000  7.205000 2.725000 ;
      RECT  7.195000  1.450000  7.555000 1.780000 ;
      RECT  7.375000  1.950000  7.895000 2.120000 ;
      RECT  7.375000  2.120000  7.545000 2.895000 ;
      RECT  7.590000  0.085000  8.260000 0.930000 ;
      RECT  7.715000  2.290000  7.885000 3.245000 ;
      RECT  7.725000  1.780000 10.765000 1.930000 ;
      RECT  7.725000  1.930000  9.375000 1.950000 ;
      RECT  7.935000  1.280000  8.265000 1.450000 ;
      RECT  8.085000  2.120000  9.875000 2.290000 ;
      RECT  8.085000  2.290000  8.365000 2.715000 ;
      RECT  8.440000  0.350000  8.610000 1.110000 ;
      RECT  8.440000  1.110000 10.030000 1.280000 ;
      RECT  8.535000  2.460000  8.865000 3.245000 ;
      RECT  8.790000  0.085000  9.120000 0.940000 ;
      RECT  9.045000  1.450000  9.375000 1.760000 ;
      RECT  9.045000  1.760000 10.765000 1.780000 ;
      RECT  9.095000  2.600000  9.375000 2.860000 ;
      RECT  9.095000  2.860000 10.375000 3.075000 ;
      RECT  9.350000  0.255000 10.540000 0.425000 ;
      RECT  9.350000  0.425000  9.680000 0.940000 ;
      RECT  9.545000  2.100000  9.875000 2.120000 ;
      RECT  9.545000  2.290000  9.875000 2.690000 ;
      RECT  9.860000  0.595000 10.030000 1.110000 ;
      RECT 10.045000  2.310000 12.210000 2.480000 ;
      RECT 10.045000  2.480000 10.375000 2.860000 ;
      RECT 10.210000  0.425000 10.540000 1.400000 ;
      RECT 10.210000  1.400000 11.105000 1.570000 ;
      RECT 10.435000  1.930000 10.765000 2.135000 ;
      RECT 10.545000  2.650000 10.955000 2.980000 ;
      RECT 10.935000  1.570000 11.105000 2.310000 ;
      RECT 10.955000  0.900000 12.710000 1.070000 ;
      RECT 10.955000  1.070000 11.285000 1.230000 ;
      RECT 11.125000  2.650000 11.375000 3.245000 ;
      RECT 11.470000  1.470000 11.870000 2.140000 ;
      RECT 11.575000  2.480000 11.905000 2.980000 ;
      RECT 11.650000  0.085000 12.150000 0.680000 ;
      RECT 12.040000  1.340000 12.370000 2.010000 ;
      RECT 12.040000  2.010000 12.210000 2.310000 ;
      RECT 12.135000  2.650000 12.550000 2.980000 ;
      RECT 12.320000  0.350000 12.710000 0.900000 ;
      RECT 12.380000  2.180000 12.710000 2.350000 ;
      RECT 12.380000  2.350000 12.550000 2.650000 ;
      RECT 12.540000  1.070000 12.710000 2.180000 ;
      RECT 12.720000  2.520000 12.970000 3.245000 ;
      RECT 12.880000  0.350000 13.210000 1.320000 ;
      RECT 12.880000  1.320000 14.695000 1.490000 ;
      RECT 13.170000  1.490000 14.695000 1.650000 ;
      RECT 13.170000  1.650000 13.340000 2.980000 ;
      RECT 13.380000  0.085000 13.710000 1.130000 ;
      RECT 13.540000  2.100000 13.870000 3.245000 ;
      RECT 14.395000  0.085000 14.725000 0.810000 ;
      RECT 14.495000  2.320000 14.825000 3.245000 ;
      RECT 15.395000  0.085000 15.725000 1.100000 ;
      RECT 15.395000  1.950000 15.725000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  1.580000  7.525000 1.750000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  1.580000 11.845000 1.750000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.245000 15.205000 3.415000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.245000 15.685000 3.415000 ;
  END
END sky130_fd_sc_hs__sdfstp_4
MACRO sky130_fd_sc_hs__sdfxbp_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.48000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.455000 1.630000 1.785000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.518900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.500000 0.350000 10.915000 1.130000 ;
        RECT 10.650000 1.820000 10.915000 2.980000 ;
        RECT 10.745000 1.130000 10.915000 1.820000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.530100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.035000 0.350000 12.375000 1.050000 ;
        RECT 12.045000 1.820000 12.375000 2.980000 ;
        RECT 12.155000 1.050000 12.375000 1.820000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.380000 1.550000 2.725000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.955000 2.050000 1.285000 ;
        RECT 1.565000 0.810000 2.050000 0.955000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.235000 1.180000 3.685000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.480000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 12.480000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.480000 0.085000 ;
      RECT  0.000000  3.245000 12.480000 3.415000 ;
      RECT  0.085000  0.350000  0.465000 0.785000 ;
      RECT  0.085000  0.785000  0.255000 1.525000 ;
      RECT  0.085000  1.525000  0.915000 1.855000 ;
      RECT  0.085000  1.855000  0.530000 2.980000 ;
      RECT  0.635000  0.085000  0.965000 0.730000 ;
      RECT  0.700000  2.300000  1.030000 3.245000 ;
      RECT  0.745000  1.855000  0.915000 1.955000 ;
      RECT  0.745000  1.955000  2.170000 2.125000 ;
      RECT  1.455000  0.390000  2.390000 0.640000 ;
      RECT  1.570000  2.300000  1.900000 2.390000 ;
      RECT  1.570000  2.390000  4.675000 2.460000 ;
      RECT  1.570000  2.460000  5.235000 2.560000 ;
      RECT  1.570000  2.560000  1.900000 2.980000 ;
      RECT  1.840000  1.795000  2.170000 1.955000 ;
      RECT  2.220000  0.640000  2.390000 1.180000 ;
      RECT  2.220000  1.180000  3.065000 1.350000 ;
      RECT  2.560000  2.730000  3.150000 3.245000 ;
      RECT  2.615000  0.085000  2.865000 0.810000 ;
      RECT  2.895000  1.350000  3.065000 2.390000 ;
      RECT  3.035000  0.350000  3.365000 0.840000 ;
      RECT  3.035000  0.840000  4.025000 1.010000 ;
      RECT  3.270000  1.820000  4.025000 1.990000 ;
      RECT  3.270000  1.990000  3.600000 2.220000 ;
      RECT  3.595000  0.085000  3.935000 0.670000 ;
      RECT  3.830000  2.730000  4.335000 3.245000 ;
      RECT  3.855000  1.010000  4.025000 1.820000 ;
      RECT  4.195000  0.255000  6.035000 0.425000 ;
      RECT  4.195000  0.425000  4.445000 1.130000 ;
      RECT  4.195000  1.480000  4.900000 1.650000 ;
      RECT  4.195000  1.650000  4.365000 2.390000 ;
      RECT  4.505000  2.560000  5.235000 2.630000 ;
      RECT  4.535000  1.820000  5.240000 2.220000 ;
      RECT  4.650000  0.595000  4.900000 1.480000 ;
      RECT  4.910000  2.220000  5.240000 2.280000 ;
      RECT  4.985000  2.630000  5.235000 2.920000 ;
      RECT  5.070000  0.425000  5.240000 1.820000 ;
      RECT  5.410000  0.595000  5.580000 1.530000 ;
      RECT  5.410000  1.530000  7.020000 1.700000 ;
      RECT  5.410000  1.700000  5.580000 2.460000 ;
      RECT  5.410000  2.460000  5.765000 2.920000 ;
      RECT  5.750000  0.425000  6.035000 0.690000 ;
      RECT  5.750000  0.690000  7.020000 0.860000 ;
      RECT  5.750000  0.860000  6.035000 1.360000 ;
      RECT  5.750000  1.870000  6.105000 2.200000 ;
      RECT  5.935000  2.200000  6.105000 2.520000 ;
      RECT  5.935000  2.520000  7.735000 2.690000 ;
      RECT  6.245000  1.030000  7.360000 1.360000 ;
      RECT  6.430000  0.085000  6.680000 0.520000 ;
      RECT  6.450000  2.860000  6.780000 3.245000 ;
      RECT  6.690000  1.700000  7.020000 1.930000 ;
      RECT  6.850000  0.255000  7.860000 0.425000 ;
      RECT  6.850000  0.425000  7.020000 0.690000 ;
      RECT  6.985000  2.100000  7.395000 2.350000 ;
      RECT  7.190000  0.595000  7.520000 0.920000 ;
      RECT  7.190000  0.920000  7.360000 1.030000 ;
      RECT  7.190000  1.360000  7.360000 2.100000 ;
      RECT  7.530000  1.090000  7.860000 1.250000 ;
      RECT  7.530000  1.250000  8.220000 1.355000 ;
      RECT  7.530000  1.355000  8.680000 1.420000 ;
      RECT  7.565000  1.630000  7.880000 1.960000 ;
      RECT  7.565000  1.960000  7.735000 2.520000 ;
      RECT  7.690000  0.425000  7.860000 1.090000 ;
      RECT  7.905000  2.130000  8.235000 2.980000 ;
      RECT  8.030000  0.350000  8.560000 0.810000 ;
      RECT  8.050000  1.420000  8.680000 1.610000 ;
      RECT  8.065000  1.780000  9.020000 1.950000 ;
      RECT  8.065000  1.950000  8.235000 2.130000 ;
      RECT  8.390000  0.810000  8.560000 0.980000 ;
      RECT  8.390000  0.980000  9.020000 1.100000 ;
      RECT  8.390000  1.100000  9.610000 1.150000 ;
      RECT  8.710000  2.120000  9.950000 2.350000 ;
      RECT  8.740000  0.085000  9.410000 0.810000 ;
      RECT  8.850000  1.150000  9.610000 1.270000 ;
      RECT  8.850000  1.270000  9.020000 1.780000 ;
      RECT  8.860000  2.650000  9.430000 3.245000 ;
      RECT  9.280000  1.270000  9.610000 1.770000 ;
      RECT  9.590000  0.350000  9.950000 0.930000 ;
      RECT  9.600000  1.940000  9.950000 2.120000 ;
      RECT  9.600000  2.350000  9.950000 2.980000 ;
      RECT  9.780000  0.930000  9.950000 1.320000 ;
      RECT  9.780000  1.320000 10.575000 1.650000 ;
      RECT  9.780000  1.650000  9.950000 1.940000 ;
      RECT 10.120000  1.820000 10.450000 3.245000 ;
      RECT 10.150000  0.085000 10.320000 1.130000 ;
      RECT 11.090000  0.540000 11.310000 1.220000 ;
      RECT 11.090000  1.220000 11.985000 1.550000 ;
      RECT 11.090000  1.550000 11.340000 2.875000 ;
      RECT 11.490000  0.085000 11.865000 1.020000 ;
      RECT 11.540000  1.995000 11.870000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
  END
END sky130_fd_sc_hs__sdfxbp_1
MACRO sky130_fd_sc_hs__sdfxbp_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.44000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.470000 1.655000 1.800000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.590000 1.800000 10.950000 1.970000 ;
        RECT 10.590000 1.970000 10.840000 2.980000 ;
        RECT 10.620000 0.350000 10.950000 1.130000 ;
        RECT 10.780000 1.130000 10.950000 1.800000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.554300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.550000 0.900000 13.315000 1.150000 ;
        RECT 12.555000 1.820000 13.315000 2.150000 ;
        RECT 12.555000 2.150000 12.835000 2.980000 ;
        RECT 13.075000 1.150000 13.315000 1.820000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405000 1.775000 2.755000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.900000 2.075000 1.230000 ;
        RECT 1.565000 0.810000 2.075000 0.900000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.265000 1.350000 3.685000 1.780000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 13.440000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 13.440000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.440000 0.085000 ;
      RECT  0.000000  3.245000 13.440000 3.415000 ;
      RECT  0.085000  0.350000  0.490000 0.730000 ;
      RECT  0.085000  0.730000  0.255000 1.470000 ;
      RECT  0.085000  1.470000  0.915000 1.800000 ;
      RECT  0.085000  1.800000  0.520000 2.925000 ;
      RECT  0.660000  0.085000  0.990000 0.730000 ;
      RECT  0.725000  2.310000  1.055000 3.245000 ;
      RECT  0.745000  1.800000  0.915000 1.970000 ;
      RECT  0.745000  1.970000  2.195000 2.140000 ;
      RECT  1.480000  0.390000  2.415000 0.640000 ;
      RECT  1.650000  2.310000  1.980000 2.370000 ;
      RECT  1.650000  2.370000  4.745000 2.495000 ;
      RECT  1.650000  2.495000  5.335000 2.540000 ;
      RECT  1.650000  2.540000  1.980000 2.925000 ;
      RECT  1.865000  1.725000  2.195000 1.970000 ;
      RECT  2.245000  0.640000  2.415000 1.350000 ;
      RECT  2.245000  1.350000  3.095000 1.520000 ;
      RECT  2.670000  2.710000  3.090000 3.245000 ;
      RECT  2.695000  0.085000  2.945000 1.130000 ;
      RECT  2.925000  1.520000  3.095000 2.370000 ;
      RECT  3.125000  0.350000  3.455000 1.010000 ;
      RECT  3.125000  1.010000  4.025000 1.180000 ;
      RECT  3.295000  1.950000  4.095000 2.200000 ;
      RECT  3.685000  0.085000  4.015000 0.840000 ;
      RECT  3.855000  1.180000  4.025000 1.350000 ;
      RECT  3.855000  1.350000  4.095000 1.950000 ;
      RECT  4.075000  2.710000  4.405000 3.245000 ;
      RECT  4.195000  0.255000  6.080000 0.425000 ;
      RECT  4.195000  0.425000  4.445000 1.130000 ;
      RECT  4.265000  1.480000  4.900000 1.650000 ;
      RECT  4.265000  1.650000  4.435000 2.370000 ;
      RECT  4.575000  2.540000  5.335000 2.665000 ;
      RECT  4.605000  1.820000  4.855000 2.005000 ;
      RECT  4.605000  2.005000  5.335000 2.200000 ;
      RECT  4.650000  0.595000  4.900000 1.480000 ;
      RECT  5.005000  2.200000  5.335000 2.325000 ;
      RECT  5.070000  0.425000  5.240000 2.005000 ;
      RECT  5.085000  2.665000  5.335000 2.935000 ;
      RECT  5.410000  0.595000  5.740000 0.875000 ;
      RECT  5.410000  0.875000  5.580000 1.575000 ;
      RECT  5.410000  1.575000  7.010000 1.745000 ;
      RECT  5.505000  1.745000  5.675000 2.475000 ;
      RECT  5.505000  2.475000  5.865000 2.935000 ;
      RECT  5.750000  1.045000  6.080000 1.375000 ;
      RECT  5.845000  1.915000  6.205000 2.245000 ;
      RECT  5.910000  0.425000  6.080000 0.770000 ;
      RECT  5.910000  0.770000  7.010000 0.940000 ;
      RECT  5.910000  0.940000  6.080000 1.045000 ;
      RECT  6.035000  2.245000  6.205000 2.615000 ;
      RECT  6.035000  2.615000  7.735000 2.785000 ;
      RECT  6.250000  1.110000  7.350000 1.405000 ;
      RECT  6.340000  0.085000  6.670000 0.600000 ;
      RECT  6.575000  2.955000  6.905000 3.245000 ;
      RECT  6.730000  1.745000  7.010000 1.945000 ;
      RECT  6.840000  0.255000  7.690000 0.425000 ;
      RECT  6.840000  0.425000  7.010000 0.770000 ;
      RECT  7.110000  2.115000  7.395000 2.445000 ;
      RECT  7.180000  0.595000  7.350000 1.110000 ;
      RECT  7.180000  1.405000  7.350000 2.115000 ;
      RECT  7.520000  0.425000  7.690000 1.030000 ;
      RECT  7.520000  1.030000  7.780000 1.225000 ;
      RECT  7.520000  1.225000  8.680000 1.395000 ;
      RECT  7.565000  1.600000  7.895000 1.930000 ;
      RECT  7.565000  1.930000  7.735000 2.615000 ;
      RECT  7.860000  0.350000  8.190000 0.810000 ;
      RECT  7.905000  2.100000  8.235000 2.980000 ;
      RECT  8.020000  0.810000  8.190000 0.885000 ;
      RECT  8.020000  0.885000  9.020000 1.055000 ;
      RECT  8.065000  1.720000  9.020000 1.890000 ;
      RECT  8.065000  1.890000  8.235000 2.100000 ;
      RECT  8.350000  1.395000  8.680000 1.550000 ;
      RECT  8.680000  0.085000  9.390000 0.715000 ;
      RECT  8.710000  2.060000  9.950000 2.380000 ;
      RECT  8.850000  1.055000  9.610000 1.225000 ;
      RECT  8.850000  1.225000  9.020000 1.720000 ;
      RECT  8.860000  2.650000  9.430000 3.245000 ;
      RECT  9.280000  1.225000  9.610000 1.550000 ;
      RECT  9.560000  0.350000  9.950000 0.885000 ;
      RECT  9.600000  1.940000  9.950000 2.060000 ;
      RECT  9.600000  2.380000  9.950000 2.980000 ;
      RECT  9.780000  0.885000  9.950000 1.300000 ;
      RECT  9.780000  1.300000 10.610000 1.630000 ;
      RECT  9.780000  1.630000  9.950000 1.940000 ;
      RECT 10.120000  0.085000 10.450000 1.130000 ;
      RECT 10.140000  1.820000 10.390000 3.245000 ;
      RECT 11.040000  2.140000 11.370000 3.245000 ;
      RECT 11.120000  1.820000 11.370000 2.140000 ;
      RECT 11.130000  0.085000 11.380000 1.130000 ;
      RECT 11.580000  0.560000 11.940000 1.320000 ;
      RECT 11.580000  1.320000 12.735000 1.650000 ;
      RECT 11.580000  1.650000 11.910000 2.860000 ;
      RECT 12.105000  1.820000 12.355000 3.245000 ;
      RECT 12.120000  0.085000 12.450000 0.730000 ;
      RECT 12.120000  0.730000 12.380000 1.150000 ;
      RECT 12.995000  0.085000 13.325000 0.730000 ;
      RECT 13.005000  2.320000 13.335000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
  END
END sky130_fd_sc_hs__sdfxbp_2
MACRO sky130_fd_sc_hs__sdfxtp_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.455000 1.655000 1.785000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.528300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.600000 0.370000 10.935000 2.980000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405000 1.470000 2.740000 2.140000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.955000 2.250000 1.285000 ;
        RECT 1.085000 0.810000 1.315000 0.900000 ;
        RECT 1.085000 0.900000 2.250000 0.955000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.250000 1.180000 3.685000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.040000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 11.040000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  3.245000 11.040000 3.415000 ;
      RECT  0.085000  0.350000  0.405000 0.785000 ;
      RECT  0.085000  0.785000  0.255000 1.525000 ;
      RECT  0.085000  1.525000  0.825000 1.955000 ;
      RECT  0.085000  1.955000  2.195000 2.125000 ;
      RECT  0.085000  2.125000  0.555000 2.980000 ;
      RECT  0.585000  0.085000  0.915000 0.785000 ;
      RECT  0.725000  2.300000  1.055000 3.245000 ;
      RECT  1.485000  0.400000  2.590000 0.730000 ;
      RECT  1.595000  2.310000  4.395000 2.390000 ;
      RECT  1.595000  2.390000  4.705000 2.480000 ;
      RECT  1.595000  2.480000  1.925000 2.980000 ;
      RECT  1.865000  1.470000  2.195000 1.955000 ;
      RECT  1.865000  2.125000  2.195000 2.140000 ;
      RECT  2.420000  0.730000  2.590000 1.130000 ;
      RECT  2.420000  1.130000  3.080000 1.300000 ;
      RECT  2.670000  2.650000  3.175000 3.245000 ;
      RECT  2.775000  0.085000  2.945000 0.790000 ;
      RECT  2.910000  1.300000  3.080000 2.310000 ;
      RECT  3.125000  0.350000  3.455000 0.790000 ;
      RECT  3.125000  0.790000  4.025000 0.960000 ;
      RECT  3.295000  1.820000  4.055000 2.140000 ;
      RECT  3.345000  2.480000  4.705000 2.560000 ;
      RECT  3.685000  0.085000  4.015000 0.620000 ;
      RECT  3.855000  0.960000  4.025000 1.300000 ;
      RECT  3.855000  1.300000  4.055000 1.820000 ;
      RECT  3.855000  2.730000  4.365000 3.245000 ;
      RECT  4.195000  0.255000  5.905000 0.425000 ;
      RECT  4.195000  0.425000  4.445000 1.130000 ;
      RECT  4.225000  1.480000  4.785000 1.650000 ;
      RECT  4.225000  1.650000  4.395000 2.310000 ;
      RECT  4.535000  2.560000  4.705000 2.710000 ;
      RECT  4.535000  2.710000  5.375000 2.980000 ;
      RECT  4.565000  1.820000  4.815000 2.050000 ;
      RECT  4.565000  2.050000  5.225000 2.220000 ;
      RECT  4.615000  0.595000  4.885000 0.940000 ;
      RECT  4.615000  0.940000  4.785000 1.480000 ;
      RECT  4.955000  2.220000  5.225000 2.380000 ;
      RECT  5.055000  0.425000  5.225000 2.050000 ;
      RECT  5.395000  0.595000  5.565000 1.530000 ;
      RECT  5.395000  1.530000  6.975000 1.700000 ;
      RECT  5.395000  1.700000  5.565000 2.370000 ;
      RECT  5.395000  2.370000  5.875000 2.540000 ;
      RECT  5.545000  2.540000  5.875000 2.980000 ;
      RECT  5.735000  0.425000  5.905000 0.690000 ;
      RECT  5.735000  0.690000  6.975000 0.860000 ;
      RECT  5.735000  0.860000  5.985000 1.360000 ;
      RECT  5.735000  1.870000  6.215000 2.200000 ;
      RECT  6.045000  2.200000  6.215000 2.520000 ;
      RECT  6.045000  2.520000  7.715000 2.690000 ;
      RECT  6.195000  1.030000  7.315000 1.360000 ;
      RECT  6.385000  0.085000  6.635000 0.520000 ;
      RECT  6.480000  2.860000  6.810000 3.245000 ;
      RECT  6.645000  1.700000  6.975000 1.930000 ;
      RECT  6.805000  0.255000  7.815000 0.425000 ;
      RECT  6.805000  0.425000  6.975000 0.690000 ;
      RECT  7.015000  2.100000  7.375000 2.350000 ;
      RECT  7.145000  0.595000  7.475000 0.860000 ;
      RECT  7.145000  0.860000  7.315000 1.030000 ;
      RECT  7.145000  1.360000  7.315000 2.100000 ;
      RECT  7.485000  1.030000  7.815000 1.190000 ;
      RECT  7.485000  1.190000  8.240000 1.320000 ;
      RECT  7.485000  1.320000  8.555000 1.360000 ;
      RECT  7.545000  1.600000  7.900000 1.930000 ;
      RECT  7.545000  1.930000  7.715000 2.520000 ;
      RECT  7.645000  0.425000  7.815000 1.030000 ;
      RECT  7.885000  2.100000  8.135000 2.245000 ;
      RECT  7.885000  2.245000  8.895000 2.415000 ;
      RECT  7.885000  2.415000  8.135000 2.980000 ;
      RECT  7.985000  0.480000  8.315000 0.770000 ;
      RECT  7.985000  0.770000  8.580000 0.940000 ;
      RECT  8.070000  1.360000  8.555000 1.490000 ;
      RECT  8.305000  1.490000  8.555000 2.075000 ;
      RECT  8.410000  0.940000  8.580000 0.980000 ;
      RECT  8.410000  0.980000  8.895000 1.150000 ;
      RECT  8.725000  1.150000  8.895000 1.600000 ;
      RECT  8.725000  1.600000  9.595000 1.930000 ;
      RECT  8.725000  1.930000  8.895000 2.245000 ;
      RECT  8.805000  0.085000  9.480000 0.810000 ;
      RECT  8.845000  2.650000  9.420000 3.245000 ;
      RECT  9.065000  1.030000  9.980000 1.320000 ;
      RECT  9.065000  1.320000 10.245000 1.360000 ;
      RECT  9.590000  2.100000  9.935000 2.980000 ;
      RECT  9.650000  0.350000  9.980000 1.030000 ;
      RECT  9.765000  1.360000 10.245000 1.650000 ;
      RECT  9.765000  1.650000  9.935000 2.100000 ;
      RECT 10.150000  1.820000 10.400000 3.245000 ;
      RECT 10.175000  0.085000 10.425000 1.150000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
  END
END sky130_fd_sc_hs__sdfxtp_1
MACRO sky130_fd_sc_hs__sdfxtp_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.190000 1.665000 1.845000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.576500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.055000 0.350000 11.385000 1.050000 ;
        RECT 11.105000 1.820000 11.435000 2.980000 ;
        RECT 11.215000 1.050000 11.385000 1.820000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.450000 1.435000 2.780000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.810000 0.835000 0.850000 ;
        RECT 0.425000 0.850000 2.205000 1.020000 ;
        RECT 0.425000 1.020000 0.835000 1.230000 ;
        RECT 1.875000 1.020000 2.205000 1.230000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.290000 1.350000 3.685000 1.780000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.000000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 12.000000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.000000 0.085000 ;
      RECT  0.000000  3.245000 12.000000 3.415000 ;
      RECT  0.085000  0.390000  0.490000 0.640000 ;
      RECT  0.085000  0.640000  0.255000 1.470000 ;
      RECT  0.085000  1.470000  0.915000 2.015000 ;
      RECT  0.085000  2.015000  2.210000 2.185000 ;
      RECT  0.085000  2.185000  0.445000 2.925000 ;
      RECT  0.615000  2.355000  0.945000 3.245000 ;
      RECT  0.660000  0.085000  0.990000 0.640000 ;
      RECT  1.480000  0.350000  2.545000 0.680000 ;
      RECT  1.485000  2.355000  3.120000 2.450000 ;
      RECT  1.485000  2.450000  5.385000 2.620000 ;
      RECT  1.485000  2.620000  2.060000 2.945000 ;
      RECT  1.880000  1.775000  2.210000 2.015000 ;
      RECT  2.375000  0.680000  2.545000 1.095000 ;
      RECT  2.375000  1.095000  3.120000 1.265000 ;
      RECT  2.685000  2.790000  3.135000 3.245000 ;
      RECT  2.715000  0.085000  2.975000 0.810000 ;
      RECT  2.950000  1.265000  3.120000 2.355000 ;
      RECT  3.145000  0.330000  3.475000 0.920000 ;
      RECT  3.305000  0.920000  3.475000 1.010000 ;
      RECT  3.305000  1.010000  4.025000 1.180000 ;
      RECT  3.340000  1.950000  4.145000 2.280000 ;
      RECT  3.705000  0.085000  4.035000 0.840000 ;
      RECT  3.855000  1.180000  4.025000 1.300000 ;
      RECT  3.855000  1.300000  4.145000 1.950000 ;
      RECT  3.900000  2.790000  4.370000 3.245000 ;
      RECT  4.205000  0.255000  6.115000 0.425000 ;
      RECT  4.205000  0.425000  4.535000 1.130000 ;
      RECT  4.315000  1.300000  4.875000 1.470000 ;
      RECT  4.315000  1.470000  4.485000 2.450000 ;
      RECT  4.655000  1.820000  5.375000 2.280000 ;
      RECT  4.705000  0.595000  5.015000 0.940000 ;
      RECT  4.705000  0.940000  4.875000 1.300000 ;
      RECT  5.045000  1.610000  5.375000 1.820000 ;
      RECT  5.135000  2.620000  5.385000 2.980000 ;
      RECT  5.185000  0.425000  5.355000 1.610000 ;
      RECT  5.525000  0.595000  5.775000 0.940000 ;
      RECT  5.555000  0.940000  5.775000 1.630000 ;
      RECT  5.555000  1.630000  7.175000 1.800000 ;
      RECT  5.555000  1.800000  5.725000 2.520000 ;
      RECT  5.555000  2.520000  5.915000 2.980000 ;
      RECT  5.895000  1.970000  6.225000 2.130000 ;
      RECT  5.895000  2.130000  7.175000 2.300000 ;
      RECT  5.945000  0.425000  6.115000 0.720000 ;
      RECT  5.945000  0.720000  7.390000 0.890000 ;
      RECT  5.945000  0.890000  6.275000 1.360000 ;
      RECT  6.485000  1.060000  7.890000 1.230000 ;
      RECT  6.485000  1.230000  7.515000 1.390000 ;
      RECT  6.585000  2.520000  6.835000 3.245000 ;
      RECT  6.720000  0.085000  7.050000 0.550000 ;
      RECT  6.845000  1.800000  7.175000 1.960000 ;
      RECT  7.005000  2.300000  7.175000 2.905000 ;
      RECT  7.005000  2.905000  7.855000 3.075000 ;
      RECT  7.220000  0.255000  8.230000 0.425000 ;
      RECT  7.220000  0.425000  7.390000 0.720000 ;
      RECT  7.345000  1.390000  7.515000 2.610000 ;
      RECT  7.560000  0.595000  7.890000 1.060000 ;
      RECT  7.685000  1.600000  8.115000 1.930000 ;
      RECT  7.685000  1.930000  7.855000 2.905000 ;
      RECT  8.025000  2.490000  9.060000 2.660000 ;
      RECT  8.025000  2.660000  8.275000 2.920000 ;
      RECT  8.060000  0.425000  8.230000 1.030000 ;
      RECT  8.060000  1.030000  8.455000 1.360000 ;
      RECT  8.285000  1.360000  8.455000 1.990000 ;
      RECT  8.285000  1.990000  8.720000 2.320000 ;
      RECT  8.400000  0.350000  8.795000 0.640000 ;
      RECT  8.400000  0.640000  9.060000 0.810000 ;
      RECT  8.890000  0.810000  9.060000 2.075000 ;
      RECT  8.890000  2.075000 10.105000 2.245000 ;
      RECT  8.890000  2.245000  9.060000 2.490000 ;
      RECT  9.230000  1.070000 10.445000 1.220000 ;
      RECT  9.230000  1.220000 11.045000 1.240000 ;
      RECT  9.230000  1.240000  9.535000 1.905000 ;
      RECT  9.295000  2.590000  9.925000 3.245000 ;
      RECT  9.300000  0.085000  9.630000 0.810000 ;
      RECT  9.775000  1.410000 10.105000 2.075000 ;
      RECT  9.800000  0.350000 10.130000 1.070000 ;
      RECT 10.095000  2.415000 10.445000 2.920000 ;
      RECT 10.275000  1.240000 11.045000 1.550000 ;
      RECT 10.275000  1.550000 10.445000 2.415000 ;
      RECT 10.615000  0.085000 10.885000 1.050000 ;
      RECT 10.655000  1.820000 10.905000 3.245000 ;
      RECT 11.555000  0.085000 11.885000 1.130000 ;
      RECT 11.635000  1.820000 11.885000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
  END
END sky130_fd_sc_hs__sdfxtp_2
MACRO sky130_fd_sc_hs__sdfxtp_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.48000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.455000 1.655000 1.785000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.149300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.685000 1.800000 12.355000 1.970000 ;
        RECT 10.685000 1.970000 11.015000 2.980000 ;
        RECT 10.745000 0.350000 10.995000 0.880000 ;
        RECT 10.745000 0.880000 12.355000 1.130000 ;
        RECT 11.665000 1.970000 12.355000 2.015000 ;
        RECT 11.665000 2.015000 11.855000 2.980000 ;
        RECT 11.675000 0.350000 11.865000 0.880000 ;
        RECT 11.760000 1.130000 12.355000 1.800000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.435000 1.550000 2.765000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.955000 2.195000 1.285000 ;
        RECT 1.565000 0.810000 2.195000 0.955000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.275000 1.180000 3.685000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.480000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 12.480000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.480000 0.085000 ;
      RECT  0.000000  3.245000 12.480000 3.415000 ;
      RECT  0.085000  0.350000  0.490000 0.785000 ;
      RECT  0.085000  0.785000  0.255000 1.525000 ;
      RECT  0.085000  1.525000  0.915000 1.955000 ;
      RECT  0.085000  1.955000  2.195000 2.125000 ;
      RECT  0.085000  2.125000  0.555000 2.980000 ;
      RECT  0.660000  0.085000  0.990000 0.785000 ;
      RECT  0.725000  2.300000  1.055000 3.245000 ;
      RECT  1.480000  0.390000  2.535000 0.640000 ;
      RECT  1.595000  2.310000  1.925000 2.390000 ;
      RECT  1.595000  2.390000  4.815000 2.540000 ;
      RECT  1.595000  2.540000  5.405000 2.560000 ;
      RECT  1.595000  2.560000  1.925000 2.980000 ;
      RECT  1.865000  1.470000  2.195000 1.955000 ;
      RECT  1.865000  2.125000  2.195000 2.140000 ;
      RECT  2.365000  0.640000  2.535000 1.180000 ;
      RECT  2.365000  1.180000  3.105000 1.350000 ;
      RECT  2.585000  2.730000  3.205000 3.245000 ;
      RECT  2.705000  0.085000  2.955000 0.810000 ;
      RECT  2.935000  1.350000  3.105000 2.390000 ;
      RECT  3.125000  0.350000  3.455000 0.840000 ;
      RECT  3.125000  0.840000  4.025000 1.010000 ;
      RECT  3.325000  1.820000  4.165000 1.990000 ;
      RECT  3.325000  1.990000  3.655000 2.220000 ;
      RECT  3.685000  0.085000  4.015000 0.670000 ;
      RECT  3.855000  1.010000  4.025000 1.300000 ;
      RECT  3.855000  1.300000  4.165000 1.820000 ;
      RECT  3.885000  2.730000  4.475000 3.245000 ;
      RECT  4.195000  0.255000  5.945000 0.425000 ;
      RECT  4.195000  0.425000  4.445000 1.130000 ;
      RECT  4.335000  1.480000  4.925000 1.650000 ;
      RECT  4.335000  1.650000  4.505000 2.390000 ;
      RECT  4.645000  2.560000  5.405000 2.710000 ;
      RECT  4.675000  0.595000  4.925000 1.480000 ;
      RECT  4.675000  1.820000  4.925000 2.040000 ;
      RECT  4.675000  2.040000  5.405000 2.220000 ;
      RECT  5.075000  2.220000  5.405000 2.370000 ;
      RECT  5.095000  0.425000  5.265000 2.040000 ;
      RECT  5.155000  2.710000  5.405000 2.970000 ;
      RECT  5.435000  0.595000  5.605000 1.610000 ;
      RECT  5.435000  1.610000  7.160000 1.780000 ;
      RECT  5.575000  1.780000  5.745000 2.510000 ;
      RECT  5.575000  2.510000  5.935000 2.970000 ;
      RECT  5.775000  0.425000  5.945000 0.770000 ;
      RECT  5.775000  0.770000  7.160000 0.940000 ;
      RECT  5.775000  0.940000  6.075000 1.360000 ;
      RECT  5.915000  1.950000  6.275000 2.280000 ;
      RECT  6.105000  2.280000  6.275000 2.515000 ;
      RECT  6.105000  2.515000  8.100000 2.685000 ;
      RECT  6.295000  1.110000  7.500000 1.440000 ;
      RECT  6.490000  0.085000  6.820000 0.600000 ;
      RECT  6.680000  2.855000  7.010000 3.245000 ;
      RECT  6.835000  1.780000  7.160000 1.940000 ;
      RECT  6.990000  0.295000  8.125000 0.465000 ;
      RECT  6.990000  0.465000  7.160000 0.770000 ;
      RECT  7.215000  2.175000  7.760000 2.345000 ;
      RECT  7.330000  0.635000  7.785000 0.885000 ;
      RECT  7.330000  0.885000  7.500000 1.110000 ;
      RECT  7.330000  1.440000  7.500000 2.175000 ;
      RECT  7.670000  1.055000  8.125000 1.240000 ;
      RECT  7.670000  1.240000  8.845000 1.410000 ;
      RECT  7.770000  1.625000  8.100000 1.955000 ;
      RECT  7.930000  1.955000  8.100000 2.515000 ;
      RECT  7.955000  0.465000  8.125000 1.055000 ;
      RECT  8.270000  2.020000  9.185000 2.190000 ;
      RECT  8.270000  2.190000  8.600000 2.820000 ;
      RECT  8.295000  0.350000  8.625000 0.900000 ;
      RECT  8.295000  0.900000  9.185000 1.070000 ;
      RECT  8.535000  1.410000  8.845000 1.715000 ;
      RECT  9.015000  1.070000  9.185000 1.470000 ;
      RECT  9.015000  1.470000  9.795000 1.800000 ;
      RECT  9.015000  1.800000  9.185000 2.020000 ;
      RECT  9.195000  0.085000  9.525000 0.730000 ;
      RECT  9.225000  2.360000  9.555000 3.245000 ;
      RECT  9.355000  0.900000  9.665000 1.130000 ;
      RECT  9.355000  1.130000 10.135000 1.300000 ;
      RECT  9.730000  1.970000 10.135000 2.820000 ;
      RECT  9.835000  0.350000 10.005000 1.130000 ;
      RECT  9.965000  1.300000 11.545000 1.630000 ;
      RECT  9.965000  1.630000 10.135000 1.970000 ;
      RECT 10.185000  0.085000 10.515000 0.960000 ;
      RECT 10.305000  1.940000 10.475000 3.245000 ;
      RECT 11.175000  0.085000 11.505000 0.710000 ;
      RECT 11.215000  2.140000 11.465000 3.245000 ;
      RECT 12.035000  0.085000 12.365000 0.710000 ;
      RECT 12.035000  2.185000 12.365000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
  END
END sky130_fd_sc_hs__sdfxtp_4
MACRO sky130_fd_sc_hs__sdlclkp_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN GATE
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.805000 1.630000 1.285000 2.150000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.632800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.235000 1.820000 7.585000 2.980000 ;
        RECT 7.240000 0.350000 7.585000 1.130000 ;
        RECT 7.415000 1.130000 7.585000 1.820000 ;
    END
  END GCLK
  PIN SCE
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.290000 0.545000 1.960000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.459000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 5.330000 1.355000 5.660000 1.780000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.680000 0.085000 ;
      RECT 0.000000  3.245000 7.680000 3.415000 ;
      RECT 0.115000  0.085000 0.365000 1.120000 ;
      RECT 0.115000  2.130000 0.445000 3.245000 ;
      RECT 0.545000  0.540000 2.375000 0.710000 ;
      RECT 0.545000  0.710000 0.885000 1.120000 ;
      RECT 0.715000  1.120000 0.885000 1.290000 ;
      RECT 0.715000  1.290000 1.625000 1.460000 ;
      RECT 0.955000  2.320000 2.860000 2.490000 ;
      RECT 0.955000  2.490000 1.285000 2.980000 ;
      RECT 1.055000  0.085000 1.385000 0.370000 ;
      RECT 1.455000  1.460000 1.625000 2.320000 ;
      RECT 1.515000  2.660000 1.845000 3.245000 ;
      RECT 1.565000  0.880000 1.895000 0.950000 ;
      RECT 1.565000  0.950000 1.965000 1.120000 ;
      RECT 1.795000  1.120000 1.965000 1.545000 ;
      RECT 1.795000  1.545000 2.900000 1.715000 ;
      RECT 1.795000  1.715000 2.380000 2.150000 ;
      RECT 2.125000  0.350000 2.375000 0.540000 ;
      RECT 2.125000  0.710000 2.375000 0.780000 ;
      RECT 2.135000  1.030000 2.715000 1.200000 ;
      RECT 2.135000  1.200000 2.415000 1.360000 ;
      RECT 2.545000  0.255000 3.580000 0.425000 ;
      RECT 2.545000  0.425000 2.715000 1.030000 ;
      RECT 2.610000  1.885000 2.860000 2.320000 ;
      RECT 2.610000  2.490000 2.860000 2.755000 ;
      RECT 2.625000  1.385000 2.900000 1.545000 ;
      RECT 2.885000  0.595000 3.240000 0.925000 ;
      RECT 3.060000  2.425000 3.390000 2.755000 ;
      RECT 3.070000  0.925000 3.240000 1.220000 ;
      RECT 3.070000  1.220000 4.320000 1.550000 ;
      RECT 3.070000  1.550000 3.390000 2.425000 ;
      RECT 3.410000  0.425000 3.580000 0.880000 ;
      RECT 3.410000  0.880000 4.260000 1.050000 ;
      RECT 3.600000  1.740000 4.820000 2.120000 ;
      RECT 3.750000  0.085000 3.920000 0.710000 ;
      RECT 3.985000  2.440000 4.315000 3.245000 ;
      RECT 4.090000  0.255000 5.230000 0.425000 ;
      RECT 4.090000  0.425000 4.260000 0.880000 ;
      RECT 4.430000  0.595000 4.680000 1.050000 ;
      RECT 4.490000  1.050000 4.680000 1.740000 ;
      RECT 4.490000  2.120000 4.820000 2.495000 ;
      RECT 4.490000  2.495000 6.000000 2.665000 ;
      RECT 4.490000  2.665000 4.820000 2.900000 ;
      RECT 4.900000  0.425000 5.230000 1.130000 ;
      RECT 4.990000  1.130000 5.160000 1.995000 ;
      RECT 4.990000  1.995000 5.380000 2.325000 ;
      RECT 5.410000  0.085000 5.660000 1.130000 ;
      RECT 5.585000  2.835000 5.990000 3.245000 ;
      RECT 5.830000  1.220000 6.305000 1.550000 ;
      RECT 5.830000  1.550000 6.000000 2.495000 ;
      RECT 6.165000  0.450000 6.645000 1.050000 ;
      RECT 6.195000  1.720000 6.645000 1.890000 ;
      RECT 6.195000  1.890000 6.525000 2.875000 ;
      RECT 6.475000  1.050000 6.645000 1.300000 ;
      RECT 6.475000  1.300000 7.245000 1.630000 ;
      RECT 6.475000  1.630000 6.645000 1.720000 ;
      RECT 6.695000  2.060000 7.025000 3.245000 ;
      RECT 6.815000  0.085000 7.065000 1.130000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
  END
END sky130_fd_sc_hs__sdlclkp_1
MACRO sky130_fd_sc_hs__sdlclkp_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN GATE
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.795000 1.630000 1.300000 2.150000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.210000 1.820000 7.565000 2.980000 ;
        RECT 7.295000 0.350000 7.625000 1.130000 ;
        RECT 7.395000 1.130000 7.565000 1.820000 ;
    END
  END GCLK
  PIN SCE
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.290000 0.550000 1.960000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.498000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 5.335000 1.180000 5.665000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.105000  2.130000 0.435000 3.245000 ;
      RECT 0.115000  0.085000 0.365000 1.120000 ;
      RECT 0.545000  0.540000 2.375000 0.710000 ;
      RECT 0.545000  0.710000 0.890000 1.120000 ;
      RECT 0.720000  1.120000 0.890000 1.220000 ;
      RECT 0.720000  1.220000 1.640000 1.390000 ;
      RECT 0.945000  2.320000 2.800000 2.490000 ;
      RECT 0.945000  2.490000 1.275000 2.980000 ;
      RECT 1.055000  0.085000 1.385000 0.370000 ;
      RECT 1.470000  1.390000 1.640000 2.320000 ;
      RECT 1.485000  2.660000 1.815000 3.245000 ;
      RECT 1.565000  0.880000 1.980000 1.050000 ;
      RECT 1.810000  1.050000 1.980000 1.545000 ;
      RECT 1.810000  1.545000 3.020000 1.715000 ;
      RECT 1.810000  1.715000 2.340000 2.150000 ;
      RECT 2.125000  0.350000 2.375000 0.540000 ;
      RECT 2.150000  1.030000 2.715000 1.200000 ;
      RECT 2.150000  1.200000 2.480000 1.360000 ;
      RECT 2.545000  0.255000 3.700000 0.425000 ;
      RECT 2.545000  0.425000 2.715000 1.030000 ;
      RECT 2.550000  1.885000 2.800000 2.320000 ;
      RECT 2.550000  2.490000 2.800000 2.755000 ;
      RECT 2.690000  1.385000 3.020000 1.545000 ;
      RECT 2.885000  0.595000 3.360000 0.845000 ;
      RECT 3.000000  2.235000 3.360000 2.695000 ;
      RECT 3.190000  0.845000 3.360000 1.245000 ;
      RECT 3.190000  1.245000 4.485000 1.415000 ;
      RECT 3.190000  1.415000 3.360000 2.235000 ;
      RECT 3.530000  0.425000 3.700000 0.905000 ;
      RECT 3.530000  0.905000 4.380000 1.075000 ;
      RECT 3.530000  1.585000 3.860000 1.755000 ;
      RECT 3.530000  1.755000 4.825000 1.925000 ;
      RECT 3.870000  0.085000 4.040000 0.735000 ;
      RECT 3.990000  2.095000 4.240000 3.245000 ;
      RECT 4.155000  1.415000 4.485000 1.585000 ;
      RECT 4.210000  0.255000 5.360000 0.425000 ;
      RECT 4.210000  0.425000 4.380000 0.905000 ;
      RECT 4.440000  1.925000 4.825000 2.220000 ;
      RECT 4.440000  2.220000 6.005000 2.390000 ;
      RECT 4.440000  2.390000 4.825000 2.920000 ;
      RECT 4.550000  0.595000 4.825000 1.075000 ;
      RECT 4.655000  1.075000 4.825000 1.755000 ;
      RECT 4.995000  0.425000 5.360000 1.010000 ;
      RECT 4.995000  1.010000 5.165000 1.720000 ;
      RECT 4.995000  1.720000 5.310000 2.050000 ;
      RECT 5.510000  2.560000 5.840000 3.245000 ;
      RECT 5.530000  0.085000 5.860000 1.010000 ;
      RECT 5.835000  1.300000 6.530000 1.630000 ;
      RECT 5.835000  1.630000 6.005000 2.220000 ;
      RECT 6.175000  1.800000 7.040000 1.970000 ;
      RECT 6.175000  1.970000 6.505000 2.890000 ;
      RECT 6.325000  0.350000 6.655000 0.960000 ;
      RECT 6.325000  0.960000 7.040000 1.130000 ;
      RECT 6.710000  2.140000 7.040000 3.245000 ;
      RECT 6.865000  0.085000 7.115000 0.790000 ;
      RECT 6.870000  1.130000 7.040000 1.300000 ;
      RECT 6.870000  1.300000 7.225000 1.630000 ;
      RECT 6.870000  1.630000 7.040000 1.800000 ;
      RECT 7.740000  1.820000 7.990000 3.245000 ;
      RECT 7.805000  0.085000 8.055000 1.130000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_hs__sdlclkp_2
MACRO sky130_fd_sc_hs__sdlclkp_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.600000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN GATE
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.835000 1.455000 1.315000 1.785000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  1.319400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.705000 1.800000 8.985000 1.970000 ;
        RECT 7.705000 1.970000 8.035000 2.980000 ;
        RECT 7.865000 0.350000 8.115000 0.960000 ;
        RECT 7.865000 0.960000 9.055000 1.130000 ;
        RECT 8.655000 1.970000 8.985000 2.980000 ;
        RECT 8.725000 0.350000 9.055000 0.960000 ;
        RECT 8.725000 1.130000 9.055000 1.410000 ;
        RECT 8.725000 1.410000 8.985000 1.800000 ;
    END
  END GCLK
  PIN SCE
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.455000 0.550000 1.785000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.516000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 5.785000 1.180000 6.115000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.600000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.600000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.600000 0.085000 ;
      RECT 0.000000  3.245000 9.600000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 1.285000 ;
      RECT 0.115000  1.955000 0.445000 3.245000 ;
      RECT 0.615000  0.615000 2.635000 0.785000 ;
      RECT 0.615000  0.785000 0.945000 1.285000 ;
      RECT 0.985000  1.955000 1.655000 2.310000 ;
      RECT 0.985000  2.310000 3.255000 2.480000 ;
      RECT 0.985000  2.480000 1.315000 2.835000 ;
      RECT 1.125000  0.085000 1.565000 0.445000 ;
      RECT 1.485000  0.785000 1.655000 1.955000 ;
      RECT 1.545000  2.650000 2.160000 3.245000 ;
      RECT 1.825000  0.955000 2.075000 1.565000 ;
      RECT 1.825000  1.565000 3.255000 1.735000 ;
      RECT 2.245000  1.065000 2.975000 1.235000 ;
      RECT 2.245000  1.235000 2.575000 1.395000 ;
      RECT 2.305000  0.350000 2.635000 0.615000 ;
      RECT 2.305000  0.785000 2.635000 0.895000 ;
      RECT 2.365000  1.735000 2.695000 2.140000 ;
      RECT 2.805000  0.270000 3.935000 0.440000 ;
      RECT 2.805000  0.440000 2.975000 1.065000 ;
      RECT 2.925000  1.405000 3.255000 1.565000 ;
      RECT 2.925000  1.905000 3.255000 2.310000 ;
      RECT 2.925000  2.480000 3.255000 2.755000 ;
      RECT 3.145000  0.610000 3.595000 0.940000 ;
      RECT 3.425000  0.940000 3.595000 1.235000 ;
      RECT 3.425000  1.235000 4.930000 1.405000 ;
      RECT 3.425000  1.405000 3.705000 2.755000 ;
      RECT 3.765000  0.440000 3.935000 0.895000 ;
      RECT 3.765000  0.895000 4.775000 1.065000 ;
      RECT 3.960000  1.575000 4.290000 1.735000 ;
      RECT 3.960000  1.735000 5.270000 1.905000 ;
      RECT 4.105000  0.085000 4.435000 0.725000 ;
      RECT 4.430000  2.075000 4.680000 3.245000 ;
      RECT 4.600000  1.405000 4.930000 1.565000 ;
      RECT 4.605000  0.255000 5.835000 0.425000 ;
      RECT 4.605000  0.425000 4.775000 0.895000 ;
      RECT 4.880000  1.905000 5.270000 2.240000 ;
      RECT 4.880000  2.240000 6.455000 2.410000 ;
      RECT 4.880000  2.410000 5.270000 2.895000 ;
      RECT 4.945000  0.595000 5.275000 1.065000 ;
      RECT 5.100000  1.065000 5.270000 1.735000 ;
      RECT 5.440000  1.820000 5.775000 2.070000 ;
      RECT 5.445000  0.425000 5.835000 1.010000 ;
      RECT 5.445000  1.010000 5.615000 1.820000 ;
      RECT 5.980000  2.580000 6.310000 3.245000 ;
      RECT 6.005000  0.085000 6.335000 1.010000 ;
      RECT 6.285000  1.300000 7.030000 1.630000 ;
      RECT 6.285000  1.630000 6.455000 2.240000 ;
      RECT 6.625000  1.800000 7.535000 1.970000 ;
      RECT 6.625000  1.970000 6.955000 2.980000 ;
      RECT 6.825000  0.350000 7.155000 0.960000 ;
      RECT 6.825000  0.960000 7.535000 1.130000 ;
      RECT 7.125000  2.140000 7.455000 3.245000 ;
      RECT 7.365000  1.130000 7.535000 1.300000 ;
      RECT 7.365000  1.300000 8.435000 1.630000 ;
      RECT 7.365000  1.630000 7.535000 1.800000 ;
      RECT 7.385000  0.085000 7.635000 0.790000 ;
      RECT 8.235000  2.140000 8.485000 3.245000 ;
      RECT 8.295000  0.085000 8.545000 0.790000 ;
      RECT 9.155000  1.820000 9.485000 3.245000 ;
      RECT 9.235000  0.085000 9.485000 1.130000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
  END
END sky130_fd_sc_hs__sdlclkp_4
MACRO sky130_fd_sc_hs__sedfxbp_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  16.32000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455000 1.060000 0.835000 1.780000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.450000 2.085000 1.780000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.845000 0.620000 15.015000 1.820000 ;
        RECT 14.845000 1.820000 15.240000 2.980000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.860000 1.820000 16.235000 2.980000 ;
        RECT 15.875000 0.370000 16.235000 1.150000 ;
        RECT 16.065000 1.150000 16.235000 1.820000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.075000 1.180000 5.635000 1.510000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.475000 1.450000 4.865000 1.780000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.575000 1.180000 7.075000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 16.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 16.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 16.320000 0.085000 ;
      RECT  0.000000  3.245000 16.320000 3.415000 ;
      RECT  0.115000  0.480000  0.660000 0.810000 ;
      RECT  0.115000  0.810000  0.285000 2.290000 ;
      RECT  0.115000  2.290000  1.545000 2.460000 ;
      RECT  0.115000  2.460000  0.445000 2.980000 ;
      RECT  0.955000  2.630000  1.205000 3.245000 ;
      RECT  1.025000  1.110000  2.040000 1.280000 ;
      RECT  1.025000  1.280000  1.355000 1.950000 ;
      RECT  1.025000  1.950000  2.665000 2.120000 ;
      RECT  1.150000  0.085000  1.480000 0.890000 ;
      RECT  1.375000  2.460000  1.545000 2.905000 ;
      RECT  1.375000  2.905000  2.225000 3.075000 ;
      RECT  1.710000  0.545000  2.040000 1.110000 ;
      RECT  1.715000  2.120000  1.885000 2.735000 ;
      RECT  2.055000  2.310000  3.545000 2.480000 ;
      RECT  2.055000  2.480000  2.225000 2.905000 ;
      RECT  2.210000  0.085000  2.540000 1.005000 ;
      RECT  2.335000  1.525000  2.665000 1.950000 ;
      RECT  2.395000  2.650000  2.645000 3.245000 ;
      RECT  2.875000  1.525000  3.205000 2.140000 ;
      RECT  3.030000  0.545000  3.360000 1.175000 ;
      RECT  3.030000  1.175000  3.545000 1.345000 ;
      RECT  3.185000  2.480000  3.545000 2.980000 ;
      RECT  3.375000  1.345000  3.545000 2.310000 ;
      RECT  3.530000  0.545000  3.885000 1.005000 ;
      RECT  3.715000  1.005000  3.885000 2.300000 ;
      RECT  3.715000  2.300000  3.965000 2.905000 ;
      RECT  3.715000  2.905000  4.785000 3.075000 ;
      RECT  4.055000  0.410000  4.305000 0.605000 ;
      RECT  4.055000  0.605000  4.740000 1.065000 ;
      RECT  4.055000  1.065000  4.305000 1.950000 ;
      RECT  4.055000  1.950000  5.870000 2.120000 ;
      RECT  4.135000  2.120000  4.305000 2.290000 ;
      RECT  4.135000  2.290000  4.445000 2.735000 ;
      RECT  4.615000  2.290000  6.210000 2.310000 ;
      RECT  4.615000  2.310000  8.335000 2.460000 ;
      RECT  4.615000  2.460000  4.785000 2.905000 ;
      RECT  4.910000  0.085000  5.240000 1.010000 ;
      RECT  4.955000  2.630000  5.205000 3.245000 ;
      RECT  5.565000  1.790000  5.870000 1.950000 ;
      RECT  5.715000  2.460000  8.335000 2.480000 ;
      RECT  5.715000  2.480000  6.045000 2.970000 ;
      RECT  5.740000  0.605000  6.210000 1.010000 ;
      RECT  6.040000  1.010000  6.210000 2.290000 ;
      RECT  6.275000  2.650000  6.605000 3.245000 ;
      RECT  6.380000  0.085000  6.550000 1.010000 ;
      RECT  6.725000  1.820000  7.525000 2.140000 ;
      RECT  6.730000  0.350000  7.060000 0.840000 ;
      RECT  6.730000  0.840000  7.525000 1.010000 ;
      RECT  7.055000  1.810000  7.525000 1.820000 ;
      RECT  7.290000  0.085000  7.620000 0.670000 ;
      RECT  7.355000  1.010000  7.525000 1.810000 ;
      RECT  7.665000  2.650000  7.995000 3.245000 ;
      RECT  7.775000  1.480000  8.530000 1.650000 ;
      RECT  7.775000  1.650000  7.945000 2.310000 ;
      RECT  7.800000  0.255000  9.690000 0.425000 ;
      RECT  7.800000  0.425000  8.050000 1.130000 ;
      RECT  8.115000  1.820000  8.870000 2.140000 ;
      RECT  8.165000  2.480000  8.335000 2.730000 ;
      RECT  8.165000  2.730000  9.020000 2.980000 ;
      RECT  8.280000  0.595000  8.530000 1.480000 ;
      RECT  8.585000  2.140000  8.870000 2.380000 ;
      RECT  8.700000  0.425000  8.870000 1.820000 ;
      RECT  9.040000  0.620000  9.320000 0.950000 ;
      RECT  9.040000  0.950000  9.210000 1.620000 ;
      RECT  9.040000  1.620000 10.730000 1.790000 ;
      RECT  9.040000  1.790000  9.210000 2.390000 ;
      RECT  9.040000  2.390000  9.520000 2.560000 ;
      RECT  9.190000  2.560000  9.520000 2.980000 ;
      RECT  9.380000  1.120000  9.690000 1.450000 ;
      RECT  9.380000  1.960000  9.860000 2.220000 ;
      RECT  9.490000  0.425000  9.690000 0.850000 ;
      RECT  9.490000  0.850000 10.730000 1.020000 ;
      RECT  9.490000  1.020000  9.690000 1.120000 ;
      RECT  9.690000  2.220000  9.860000 2.390000 ;
      RECT  9.690000  2.390000 12.595000 2.560000 ;
      RECT  9.860000  1.190000 11.740000 1.360000 ;
      RECT  9.860000  1.360000 10.190000 1.450000 ;
      RECT 10.065000  0.085000 10.390000 0.680000 ;
      RECT 10.080000  2.730000 10.410000 3.245000 ;
      RECT 10.400000  1.530000 10.730000 1.620000 ;
      RECT 10.400000  1.790000 10.730000 1.830000 ;
      RECT 10.560000  0.255000 11.410000 0.425000 ;
      RECT 10.560000  0.425000 10.730000 0.850000 ;
      RECT 10.615000  2.050000 11.070000 2.220000 ;
      RECT 10.900000  0.595000 11.070000 1.190000 ;
      RECT 10.900000  1.360000 11.740000 1.520000 ;
      RECT 10.900000  1.520000 11.070000 2.050000 ;
      RECT 11.175000  2.730000 11.505000 3.245000 ;
      RECT 11.240000  0.425000 11.410000 0.850000 ;
      RECT 11.240000  0.850000 12.120000 1.020000 ;
      RECT 11.580000  0.085000 11.830000 0.680000 ;
      RECT 11.950000  1.020000 12.120000 1.130000 ;
      RECT 11.950000  1.130000 13.395000 1.300000 ;
      RECT 11.950000  1.300000 12.255000 1.800000 ;
      RECT 12.290000  0.350000 12.620000 0.770000 ;
      RECT 12.290000  0.770000 13.875000 0.940000 ;
      RECT 12.425000  1.470000 12.855000 1.800000 ;
      RECT 12.425000  1.800000 12.595000 2.390000 ;
      RECT 12.765000  2.520000 13.195000 2.980000 ;
      RECT 13.025000  1.715000 13.875000 1.885000 ;
      RECT 13.025000  1.885000 13.195000 2.520000 ;
      RECT 13.065000  1.300000 13.395000 1.545000 ;
      RECT 13.190000  0.085000 14.035000 0.600000 ;
      RECT 13.460000  2.055000 14.600000 2.380000 ;
      RECT 13.640000  2.650000 14.230000 3.245000 ;
      RECT 13.705000  0.940000 13.875000 1.200000 ;
      RECT 13.705000  1.200000 14.260000 1.530000 ;
      RECT 13.705000  1.530000 13.875000 1.715000 ;
      RECT 14.045000  1.920000 14.600000 2.055000 ;
      RECT 14.205000  0.255000 15.355000 0.425000 ;
      RECT 14.205000  0.425000 14.600000 1.030000 ;
      RECT 14.430000  1.030000 14.600000 1.920000 ;
      RECT 14.430000  2.380000 14.600000 2.980000 ;
      RECT 15.185000  0.425000 15.355000 1.320000 ;
      RECT 15.185000  1.320000 15.895000 1.650000 ;
      RECT 15.440000  1.820000 15.690000 3.245000 ;
      RECT 15.525000  0.085000 15.695000 1.150000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  1.950000  3.205000 2.120000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  1.950000 14.245000 2.120000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.245000 15.205000 3.415000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.245000 15.685000 3.415000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.245000 16.165000 3.415000 ;
    LAYER met1 ;
      RECT  2.975000 1.920000  3.265000 1.965000 ;
      RECT  2.975000 1.965000 14.305000 2.105000 ;
      RECT  2.975000 2.105000  3.265000 2.150000 ;
      RECT 14.015000 1.920000 14.305000 1.965000 ;
      RECT 14.015000 2.105000 14.305000 2.150000 ;
  END
END sky130_fd_sc_hs__sedfxbp_1
MACRO sky130_fd_sc_hs__sedfxbp_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  17.28000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.980000 0.835000 1.990000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.450000 1.905000 1.780000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.485000 0.350000 15.825000 2.150000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.355000 0.350000 16.685000 0.960000 ;
        RECT 16.355000 0.960000 17.165000 1.130000 ;
        RECT 16.435000 1.805000 17.165000 1.975000 ;
        RECT 16.435000 1.975000 16.665000 3.010000 ;
        RECT 16.700000 1.130000 17.165000 1.805000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.125000 1.180000 5.635000 1.510000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.475000 1.180000 4.915000 1.510000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.705000 1.180000 7.045000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 17.280000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 17.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 17.280000 0.085000 ;
      RECT  0.000000  3.245000 17.280000 3.415000 ;
      RECT  0.085000  0.420000  0.580000 0.730000 ;
      RECT  0.085000  0.730000  0.255000 2.290000 ;
      RECT  0.085000  2.290000  1.655000 2.460000 ;
      RECT  0.085000  2.460000  0.525000 2.980000 ;
      RECT  1.005000  1.110000  2.010000 1.280000 ;
      RECT  1.005000  1.280000  1.335000 1.950000 ;
      RECT  1.005000  1.950000  2.635000 2.120000 ;
      RECT  1.065000  2.630000  1.315000 3.245000 ;
      RECT  1.070000  0.085000  1.400000 0.810000 ;
      RECT  1.485000  2.460000  1.655000 2.905000 ;
      RECT  1.485000  2.905000  2.335000 3.075000 ;
      RECT  1.680000  0.545000  2.010000 1.110000 ;
      RECT  1.825000  2.120000  1.995000 2.735000 ;
      RECT  2.165000  2.290000  3.545000 2.460000 ;
      RECT  2.165000  2.460000  2.335000 2.905000 ;
      RECT  2.180000  0.085000  2.510000 1.005000 ;
      RECT  2.305000  1.515000  2.635000 1.950000 ;
      RECT  2.505000  2.630000  2.755000 3.245000 ;
      RECT  2.875000  1.515000  3.205000 1.845000 ;
      RECT  3.000000  0.545000  3.330000 1.175000 ;
      RECT  3.000000  1.175000  3.545000 1.345000 ;
      RECT  3.265000  2.460000  3.545000 2.970000 ;
      RECT  3.375000  1.345000  3.545000 2.290000 ;
      RECT  3.500000  0.545000  3.885000 1.005000 ;
      RECT  3.715000  1.005000  3.885000 2.290000 ;
      RECT  3.715000  2.290000  3.965000 2.905000 ;
      RECT  3.715000  2.905000  4.865000 3.075000 ;
      RECT  4.055000  0.365000  4.305000 0.605000 ;
      RECT  4.055000  0.605000  4.790000 1.010000 ;
      RECT  4.055000  1.010000  4.305000 1.680000 ;
      RECT  4.055000  1.680000  6.135000 1.850000 ;
      RECT  4.055000  1.850000  4.305000 2.055000 ;
      RECT  4.135000  2.055000  4.305000 2.245000 ;
      RECT  4.135000  2.245000  4.525000 2.735000 ;
      RECT  4.695000  2.255000  6.475000 2.310000 ;
      RECT  4.695000  2.310000  8.465000 2.425000 ;
      RECT  4.695000  2.425000  4.865000 2.905000 ;
      RECT  4.960000  0.085000  5.290000 1.010000 ;
      RECT  5.035000  2.595000  5.305000 3.245000 ;
      RECT  5.805000  1.430000  6.135000 1.680000 ;
      RECT  5.805000  1.850000  6.135000 2.085000 ;
      RECT  5.820000  0.605000  6.150000 1.090000 ;
      RECT  5.820000  1.090000  6.475000 1.260000 ;
      RECT  5.845000  2.425000  8.465000 2.480000 ;
      RECT  5.845000  2.480000  6.305000 2.925000 ;
      RECT  6.305000  1.260000  6.475000 2.255000 ;
      RECT  6.415000  0.085000  6.745000 0.920000 ;
      RECT  6.485000  2.650000  6.735000 3.245000 ;
      RECT  6.855000  1.820000  7.655000 2.140000 ;
      RECT  6.915000  0.350000  7.385000 1.010000 ;
      RECT  7.215000  1.010000  7.385000 1.470000 ;
      RECT  7.215000  1.470000  7.655000 1.820000 ;
      RECT  7.555000  0.085000  7.725000 1.130000 ;
      RECT  7.795000  2.650000  8.125000 3.245000 ;
      RECT  7.905000  0.255000  9.735000 0.425000 ;
      RECT  7.905000  0.425000  8.235000 1.130000 ;
      RECT  7.905000  1.480000  8.715000 1.650000 ;
      RECT  7.905000  1.650000  8.075000 2.310000 ;
      RECT  8.245000  1.820000  9.055000 2.140000 ;
      RECT  8.295000  2.480000  9.055000 2.650000 ;
      RECT  8.465000  0.595000  8.715000 1.480000 ;
      RECT  8.725000  2.140000  9.055000 2.305000 ;
      RECT  8.805000  2.650000  9.055000 2.980000 ;
      RECT  8.885000  0.425000  9.055000 1.820000 ;
      RECT  9.225000  0.595000  9.395000 1.690000 ;
      RECT  9.225000  1.690000 10.940000 1.860000 ;
      RECT  9.225000  1.860000  9.395000 2.530000 ;
      RECT  9.225000  2.530000  9.585000 2.980000 ;
      RECT  9.565000  0.425000  9.735000 0.850000 ;
      RECT  9.565000  0.850000 10.860000 1.020000 ;
      RECT  9.565000  1.020000  9.855000 1.345000 ;
      RECT  9.565000  2.030000  9.925000 2.360000 ;
      RECT  9.755000  2.360000  9.925000 2.390000 ;
      RECT  9.755000  2.390000 12.720000 2.560000 ;
      RECT 10.065000  1.190000 11.885000 1.360000 ;
      RECT 10.065000  1.360000 10.395000 1.520000 ;
      RECT 10.225000  2.730000 10.555000 3.245000 ;
      RECT 10.270000  0.085000 10.520000 0.680000 ;
      RECT 10.610000  1.530000 10.940000 1.690000 ;
      RECT 10.690000  0.255000 11.540000 0.425000 ;
      RECT 10.690000  0.425000 10.860000 0.850000 ;
      RECT 10.760000  2.050000 11.385000 2.220000 ;
      RECT 11.030000  0.595000 11.200000 1.190000 ;
      RECT 11.215000  1.360000 11.885000 1.520000 ;
      RECT 11.215000  1.520000 11.385000 2.050000 ;
      RECT 11.320000  2.730000 11.650000 3.245000 ;
      RECT 11.370000  0.425000 11.540000 0.850000 ;
      RECT 11.370000  0.850000 12.250000 1.020000 ;
      RECT 11.710000  0.085000 11.960000 0.680000 ;
      RECT 12.080000  1.020000 12.250000 1.130000 ;
      RECT 12.080000  1.130000 13.525000 1.300000 ;
      RECT 12.080000  1.300000 12.380000 1.800000 ;
      RECT 12.420000  0.350000 12.750000 0.770000 ;
      RECT 12.420000  0.770000 13.865000 0.940000 ;
      RECT 12.550000  1.470000 12.985000 1.800000 ;
      RECT 12.550000  1.800000 12.720000 2.390000 ;
      RECT 12.890000  2.520000 13.325000 2.980000 ;
      RECT 13.155000  1.715000 13.865000 1.885000 ;
      RECT 13.155000  1.885000 13.325000 2.520000 ;
      RECT 13.195000  1.300000 13.525000 1.545000 ;
      RECT 13.320000  0.085000 14.335000 0.600000 ;
      RECT 13.585000  2.055000 15.235000 2.320000 ;
      RECT 13.585000  2.320000 16.185000 2.380000 ;
      RECT 13.695000  0.940000 13.865000 1.300000 ;
      RECT 13.695000  1.300000 14.495000 1.630000 ;
      RECT 13.695000  1.630000 13.865000 1.715000 ;
      RECT 13.765000  2.650000 14.305000 3.245000 ;
      RECT 14.065000  0.600000 14.335000 1.120000 ;
      RECT 14.475000  1.800000 15.235000 2.055000 ;
      RECT 14.475000  2.380000 16.185000 2.490000 ;
      RECT 14.475000  2.490000 14.835000 2.980000 ;
      RECT 14.505000  0.350000 14.835000 1.130000 ;
      RECT 14.665000  1.130000 14.835000 1.550000 ;
      RECT 14.665000  1.550000 15.235000 1.800000 ;
      RECT 15.035000  2.660000 15.365000 3.245000 ;
      RECT 15.065000  0.085000 15.315000 1.130000 ;
      RECT 15.935000  2.660000 16.265000 3.245000 ;
      RECT 15.995000  1.300000 16.510000 1.635000 ;
      RECT 15.995000  1.635000 16.185000 2.320000 ;
      RECT 16.005000  0.085000 16.175000 1.130000 ;
      RECT 16.835000  2.145000 17.165000 3.245000 ;
      RECT 16.855000  0.085000 17.115000 0.790000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  1.580000  3.205000 1.750000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  1.580000 15.205000 1.750000 ;
      RECT 15.035000  3.245000 15.205000 3.415000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.245000 15.685000 3.415000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.245000 16.165000 3.415000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  3.245000 16.645000 3.415000 ;
      RECT 16.955000 -0.085000 17.125000 0.085000 ;
      RECT 16.955000  3.245000 17.125000 3.415000 ;
    LAYER met1 ;
      RECT  2.975000 1.550000  3.265000 1.595000 ;
      RECT  2.975000 1.595000 15.265000 1.735000 ;
      RECT  2.975000 1.735000  3.265000 1.780000 ;
      RECT 14.975000 1.550000 15.265000 1.595000 ;
      RECT 14.975000 1.735000 15.265000 1.780000 ;
  END
END sky130_fd_sc_hs__sedfxbp_2
MACRO sky130_fd_sc_hs__sedfxtp_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  15.36000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.110000 0.805000 1.780000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.515000 1.320000 1.845000 1.780000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.518900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.475000 0.350000 14.815000 2.980000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925000 1.180000 5.280000 1.745000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.400000 1.180000 4.730000 1.510000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.330000 1.180000 6.660000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 15.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 15.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 15.360000 0.085000 ;
      RECT  0.000000  3.245000 15.360000 3.415000 ;
      RECT  0.085000  0.480000  0.590000 0.810000 ;
      RECT  0.085000  0.810000  0.255000 2.290000 ;
      RECT  0.085000  2.290000  1.535000 2.460000 ;
      RECT  0.085000  2.460000  0.435000 2.980000 ;
      RECT  0.945000  2.630000  1.195000 3.245000 ;
      RECT  0.975000  0.980000  1.890000 0.995000 ;
      RECT  0.975000  0.995000  1.810000 1.150000 ;
      RECT  0.975000  1.150000  1.305000 1.950000 ;
      RECT  0.975000  1.950000  2.385000 2.120000 ;
      RECT  1.080000  0.085000  1.410000 0.810000 ;
      RECT  1.365000  2.460000  1.535000 2.905000 ;
      RECT  1.365000  2.905000  2.215000 3.075000 ;
      RECT  1.640000  0.535000  1.890000 0.980000 ;
      RECT  1.705000  2.120000  1.875000 2.735000 ;
      RECT  2.045000  2.290000  3.395000 2.460000 ;
      RECT  2.045000  2.460000  2.215000 2.905000 ;
      RECT  2.055000  1.520000  2.385000 1.950000 ;
      RECT  2.070000  0.085000  2.400000 0.995000 ;
      RECT  2.385000  2.630000  2.635000 3.245000 ;
      RECT  2.555000  1.505000  3.055000 1.835000 ;
      RECT  2.890000  0.535000  3.220000 1.165000 ;
      RECT  2.890000  1.165000  3.395000 1.335000 ;
      RECT  3.145000  2.460000  3.395000 2.975000 ;
      RECT  3.225000  1.335000  3.395000 2.290000 ;
      RECT  3.390000  0.535000  3.735000 0.995000 ;
      RECT  3.565000  0.995000  3.735000 2.295000 ;
      RECT  3.565000  2.295000  3.845000 2.905000 ;
      RECT  3.565000  2.905000  4.710000 3.075000 ;
      RECT  3.905000  0.255000  4.185000 0.605000 ;
      RECT  3.905000  0.605000  4.575000 1.010000 ;
      RECT  3.905000  1.010000  4.185000 1.915000 ;
      RECT  3.905000  1.915000  5.820000 2.085000 ;
      RECT  4.015000  2.085000  4.185000 2.255000 ;
      RECT  4.015000  2.255000  4.370000 2.735000 ;
      RECT  4.540000  2.255000  6.160000 2.330000 ;
      RECT  4.540000  2.330000  8.180000 2.425000 ;
      RECT  4.540000  2.425000  4.710000 2.905000 ;
      RECT  4.755000  0.085000  5.005000 1.010000 ;
      RECT  4.880000  2.595000  5.130000 3.245000 ;
      RECT  5.465000  0.605000  5.795000 1.075000 ;
      RECT  5.465000  1.075000  6.160000 1.245000 ;
      RECT  5.490000  1.415000  5.820000 1.915000 ;
      RECT  5.640000  2.425000  8.180000 2.500000 ;
      RECT  5.640000  2.500000  5.990000 2.935000 ;
      RECT  5.990000  1.245000  6.160000 2.255000 ;
      RECT  6.020000  0.085000  6.280000 0.905000 ;
      RECT  6.160000  2.670000  6.490000 3.245000 ;
      RECT  6.450000  0.350000  6.780000 0.840000 ;
      RECT  6.450000  0.840000  7.000000 1.010000 ;
      RECT  6.610000  1.760000  7.000000 1.830000 ;
      RECT  6.610000  1.830000  7.390000 2.160000 ;
      RECT  6.830000  1.010000  7.000000 1.760000 ;
      RECT  7.005000  0.085000  7.335000 0.670000 ;
      RECT  7.510000  2.670000  7.840000 3.245000 ;
      RECT  7.515000  0.255000  9.255000 0.425000 ;
      RECT  7.515000  0.425000  7.765000 1.130000 ;
      RECT  7.620000  1.480000  8.235000 1.650000 ;
      RECT  7.620000  1.650000  7.790000 2.330000 ;
      RECT  7.960000  1.820000  8.575000 1.990000 ;
      RECT  7.960000  1.990000  8.665000 2.160000 ;
      RECT  7.985000  0.595000  8.235000 1.480000 ;
      RECT  8.010000  2.500000  8.180000 2.730000 ;
      RECT  8.010000  2.730000  8.815000 2.980000 ;
      RECT  8.405000  0.425000  8.575000 1.820000 ;
      RECT  8.405000  2.160000  8.665000 2.335000 ;
      RECT  8.745000  0.595000  8.915000 1.620000 ;
      RECT  8.745000  1.620000 10.465000 1.790000 ;
      RECT  8.835000  1.790000  9.005000 2.390000 ;
      RECT  8.835000  2.390000  9.315000 2.560000 ;
      RECT  8.985000  2.560000  9.315000 2.980000 ;
      RECT  9.085000  0.425000  9.255000 0.850000 ;
      RECT  9.085000  0.850000 10.340000 1.020000 ;
      RECT  9.085000  1.020000  9.340000 1.345000 ;
      RECT  9.175000  1.960000  9.655000 2.220000 ;
      RECT  9.485000  2.220000  9.655000 2.390000 ;
      RECT  9.485000  2.390000 12.200000 2.560000 ;
      RECT  9.565000  1.190000  9.895000 1.195000 ;
      RECT  9.565000  1.195000 11.385000 1.365000 ;
      RECT  9.565000  1.365000  9.895000 1.450000 ;
      RECT  9.750000  0.085000 10.000000 0.680000 ;
      RECT  9.865000  2.730000 10.195000 3.245000 ;
      RECT 10.135000  1.535000 10.465000 1.620000 ;
      RECT 10.135000  1.790000 10.465000 1.795000 ;
      RECT 10.170000  0.255000 11.020000 0.425000 ;
      RECT 10.170000  0.425000 10.340000 0.850000 ;
      RECT 10.385000  1.970000 10.805000 2.220000 ;
      RECT 10.510000  0.595000 10.680000 1.195000 ;
      RECT 10.635000  1.365000 11.385000 1.525000 ;
      RECT 10.635000  1.525000 10.805000 1.970000 ;
      RECT 10.850000  0.425000 11.020000 0.855000 ;
      RECT 10.850000  0.855000 11.730000 1.025000 ;
      RECT 10.905000  2.730000 11.235000 3.245000 ;
      RECT 11.190000  0.085000 11.440000 0.685000 ;
      RECT 11.560000  1.025000 11.730000 1.110000 ;
      RECT 11.560000  1.110000 13.005000 1.280000 ;
      RECT 11.560000  1.280000 11.860000 1.800000 ;
      RECT 11.900000  0.350000 12.230000 0.770000 ;
      RECT 11.900000  0.770000 13.345000 0.940000 ;
      RECT 12.030000  1.450000 12.465000 1.735000 ;
      RECT 12.030000  1.735000 12.200000 2.390000 ;
      RECT 12.370000  1.940000 12.805000 2.980000 ;
      RECT 12.635000  1.735000 13.785000 1.905000 ;
      RECT 12.635000  1.905000 12.805000 1.940000 ;
      RECT 12.675000  1.280000 13.005000 1.555000 ;
      RECT 12.800000  0.085000 13.755000 0.600000 ;
      RECT 13.065000  2.075000 14.285000 2.380000 ;
      RECT 13.175000  0.940000 13.345000 1.735000 ;
      RECT 13.330000  2.650000 13.785000 3.245000 ;
      RECT 13.615000  1.050000 13.945000 1.380000 ;
      RECT 13.615000  1.380000 13.785000 1.735000 ;
      RECT 13.925000  0.350000 14.285000 0.810000 ;
      RECT 13.955000  2.380000 14.285000 2.980000 ;
      RECT 14.045000  1.550000 14.285000 2.075000 ;
      RECT 14.115000  0.810000 14.285000 1.550000 ;
      RECT 14.995000  0.085000 15.245000 1.130000 ;
      RECT 15.005000  1.820000 15.255000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  1.580000  2.725000 1.750000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  1.580000 14.245000 1.750000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.245000 15.205000 3.415000 ;
    LAYER met1 ;
      RECT  2.495000 1.550000  2.785000 1.595000 ;
      RECT  2.495000 1.595000 14.305000 1.735000 ;
      RECT  2.495000 1.735000  2.785000 1.780000 ;
      RECT 14.015000 1.550000 14.305000 1.595000 ;
      RECT 14.015000 1.735000 14.305000 1.780000 ;
  END
END sky130_fd_sc_hs__sedfxtp_1
MACRO sky130_fd_sc_hs__sedfxtp_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  16.32000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.980000 0.805000 1.990000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.515000 1.320000 1.845000 1.780000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.560000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.375000 0.350000 15.705000 1.130000 ;
        RECT 15.460000 1.130000 15.705000 1.550000 ;
        RECT 15.460000 1.550000 16.195000 2.150000 ;
        RECT 15.460000 2.150000 15.705000 2.980000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.955000 1.180000 5.410000 1.745000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.465000 1.180000 4.785000 1.510000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.395000 1.180000 6.725000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 16.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 16.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 16.320000 0.085000 ;
      RECT  0.000000  3.245000 16.320000 3.415000 ;
      RECT  0.085000  0.350000  0.565000 0.810000 ;
      RECT  0.085000  0.810000  0.255000 2.290000 ;
      RECT  0.085000  2.290000  1.640000 2.460000 ;
      RECT  0.085000  2.460000  0.510000 2.980000 ;
      RECT  0.975000  0.980000  1.865000 1.150000 ;
      RECT  0.975000  1.150000  1.305000 1.950000 ;
      RECT  0.975000  1.950000  2.385000 2.120000 ;
      RECT  1.050000  2.630000  1.300000 3.245000 ;
      RECT  1.055000  0.085000  1.385000 0.810000 ;
      RECT  1.470000  2.460000  1.640000 2.905000 ;
      RECT  1.470000  2.905000  2.320000 3.075000 ;
      RECT  1.615000  0.545000  1.865000 0.980000 ;
      RECT  1.810000  2.120000  1.980000 2.735000 ;
      RECT  2.045000  0.085000  2.375000 1.005000 ;
      RECT  2.055000  1.520000  2.385000 1.950000 ;
      RECT  2.150000  2.290000  3.500000 2.460000 ;
      RECT  2.150000  2.460000  2.320000 2.905000 ;
      RECT  2.490000  2.630000  2.740000 3.245000 ;
      RECT  2.555000  1.515000  3.070000 1.845000 ;
      RECT  2.865000  0.675000  3.340000 1.005000 ;
      RECT  3.170000  1.005000  3.340000 1.175000 ;
      RECT  3.170000  1.175000  3.500000 1.345000 ;
      RECT  3.250000  2.460000  3.500000 2.975000 ;
      RECT  3.330000  1.345000  3.500000 2.290000 ;
      RECT  3.510000  0.545000  3.840000 1.005000 ;
      RECT  3.670000  1.005000  3.840000 2.295000 ;
      RECT  3.670000  2.295000  3.950000 2.905000 ;
      RECT  3.670000  2.905000  4.840000 3.075000 ;
      RECT  4.010000  0.255000  4.295000 0.605000 ;
      RECT  4.010000  0.605000  4.715000 1.010000 ;
      RECT  4.010000  1.010000  4.295000 1.915000 ;
      RECT  4.010000  1.915000  5.885000 2.085000 ;
      RECT  4.125000  2.085000  4.295000 2.255000 ;
      RECT  4.125000  2.255000  4.500000 2.735000 ;
      RECT  4.670000  2.255000  6.225000 2.370000 ;
      RECT  4.670000  2.370000  8.425000 2.425000 ;
      RECT  4.670000  2.425000  4.840000 2.905000 ;
      RECT  4.885000  0.085000  5.215000 1.010000 ;
      RECT  5.010000  2.595000  5.260000 3.245000 ;
      RECT  5.620000  1.415000  5.885000 1.915000 ;
      RECT  5.675000  0.605000  6.005000 0.895000 ;
      RECT  5.675000  0.895000  6.225000 1.065000 ;
      RECT  5.800000  2.425000  8.425000 2.520000 ;
      RECT  5.800000  2.520000  9.015000 2.540000 ;
      RECT  5.800000  2.540000  6.130000 2.935000 ;
      RECT  6.055000  1.065000  6.225000 2.255000 ;
      RECT  6.235000  0.085000  6.495000 0.680000 ;
      RECT  6.360000  2.710000  6.695000 3.245000 ;
      RECT  6.675000  0.350000  7.065000 1.010000 ;
      RECT  6.895000  1.010000  7.065000 1.530000 ;
      RECT  6.895000  1.530000  7.615000 2.200000 ;
      RECT  7.235000  0.085000  7.485000 1.130000 ;
      RECT  7.665000  0.255000  9.495000 0.425000 ;
      RECT  7.665000  0.425000  7.995000 1.130000 ;
      RECT  7.755000  2.710000  8.085000 3.245000 ;
      RECT  7.865000  1.480000  8.475000 1.650000 ;
      RECT  7.865000  1.650000  8.035000 2.370000 ;
      RECT  8.205000  1.820000  8.815000 2.020000 ;
      RECT  8.205000  2.020000  9.005000 2.200000 ;
      RECT  8.225000  0.595000  8.475000 1.480000 ;
      RECT  8.255000  2.540000  9.015000 2.690000 ;
      RECT  8.645000  0.425000  8.815000 1.820000 ;
      RECT  8.645000  2.200000  9.005000 2.350000 ;
      RECT  8.765000  2.690000  9.015000 2.980000 ;
      RECT  8.985000  0.595000  9.155000 1.660000 ;
      RECT  8.985000  1.660000 10.785000 1.830000 ;
      RECT  9.185000  1.830000  9.355000 2.520000 ;
      RECT  9.185000  2.520000  9.545000 2.980000 ;
      RECT  9.325000  0.425000  9.495000 0.850000 ;
      RECT  9.325000  0.850000 10.705000 1.020000 ;
      RECT  9.325000  1.020000  9.655000 1.345000 ;
      RECT  9.525000  2.020000  9.885000 2.350000 ;
      RECT  9.715000  2.350000  9.885000 2.390000 ;
      RECT  9.715000  2.390000 12.730000 2.560000 ;
      RECT  9.915000  1.190000 11.800000 1.360000 ;
      RECT  9.915000  1.360000 10.245000 1.490000 ;
      RECT 10.100000  0.085000 10.365000 0.680000 ;
      RECT 10.215000  2.730000 10.545000 3.245000 ;
      RECT 10.455000  1.530000 10.785000 1.660000 ;
      RECT 10.535000  0.255000 11.465000 0.425000 ;
      RECT 10.535000  0.425000 10.705000 0.850000 ;
      RECT 10.750000  2.050000 11.125000 2.220000 ;
      RECT 10.875000  0.595000 11.125000 1.190000 ;
      RECT 10.955000  1.360000 11.800000 1.520000 ;
      RECT 10.955000  1.520000 11.125000 2.050000 ;
      RECT 11.295000  0.425000 11.465000 0.850000 ;
      RECT 11.295000  0.850000 12.210000 1.020000 ;
      RECT 11.310000  2.730000 11.650000 3.245000 ;
      RECT 11.635000  0.085000 11.885000 0.680000 ;
      RECT 12.040000  1.020000 12.210000 1.190000 ;
      RECT 12.040000  1.190000 13.450000 1.360000 ;
      RECT 12.040000  1.360000 12.370000 1.800000 ;
      RECT 12.390000  0.350000 12.720000 0.850000 ;
      RECT 12.390000  0.850000 13.790000 1.020000 ;
      RECT 12.560000  1.530000 12.910000 1.755000 ;
      RECT 12.560000  1.755000 12.730000 2.390000 ;
      RECT 12.900000  1.925000 13.250000 2.980000 ;
      RECT 13.080000  1.755000 14.410000 1.925000 ;
      RECT 13.120000  1.360000 13.450000 1.585000 ;
      RECT 13.210000  0.085000 14.145000 0.680000 ;
      RECT 13.510000  2.095000 13.840000 2.300000 ;
      RECT 13.510000  2.300000 14.750000 2.470000 ;
      RECT 13.620000  1.020000 13.790000 1.755000 ;
      RECT 13.690000  2.650000 14.230000 3.245000 ;
      RECT 14.080000  1.460000 14.410000 1.755000 ;
      RECT 14.080000  1.925000 14.410000 2.130000 ;
      RECT 14.315000  0.350000 14.645000 1.120000 ;
      RECT 14.315000  1.120000 14.750000 1.290000 ;
      RECT 14.400000  2.470000 14.750000 2.980000 ;
      RECT 14.580000  1.290000 14.750000 1.550000 ;
      RECT 14.580000  1.550000 15.235000 1.780000 ;
      RECT 14.580000  1.780000 14.750000 2.300000 ;
      RECT 14.875000  0.085000 15.205000 0.950000 ;
      RECT 14.960000  1.950000 15.290000 3.245000 ;
      RECT 15.875000  0.085000 16.205000 1.130000 ;
      RECT 15.875000  2.320000 16.205000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  1.580000  2.725000 1.750000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  1.580000 15.205000 1.750000 ;
      RECT 15.035000  3.245000 15.205000 3.415000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.245000 15.685000 3.415000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.245000 16.165000 3.415000 ;
    LAYER met1 ;
      RECT  2.495000 1.550000  2.785000 1.595000 ;
      RECT  2.495000 1.595000 15.265000 1.735000 ;
      RECT  2.495000 1.735000  2.785000 1.780000 ;
      RECT 14.975000 1.550000 15.265000 1.595000 ;
      RECT 14.975000 1.735000 15.265000 1.780000 ;
  END
END sky130_fd_sc_hs__sedfxtp_2
MACRO sky130_fd_sc_hs__sedfxtp_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  16.80000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.980000 0.825000 1.990000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.535000 1.320000 1.865000 1.780000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  1.097500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.065000 1.820000 16.675000 2.150000 ;
        RECT 15.065000 2.150000 15.285000 2.980000 ;
        RECT 15.075000 0.560000 15.325000 1.090000 ;
        RECT 15.075000 1.090000 16.675000 1.340000 ;
        RECT 15.165000 1.340000 16.675000 1.820000 ;
        RECT 15.970000 2.150000 16.185000 2.980000 ;
        RECT 15.995000 0.575000 16.200000 1.090000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.955000 1.180000 5.370000 1.745000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.180000 4.785000 1.510000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.455000 1.180000 7.075000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 16.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 16.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 16.800000 0.085000 ;
      RECT  0.000000  3.245000 16.800000 3.415000 ;
      RECT  0.085000  0.340000  0.550000 0.810000 ;
      RECT  0.085000  0.810000  0.255000 2.290000 ;
      RECT  0.085000  2.290000  1.625000 2.460000 ;
      RECT  0.085000  2.460000  0.495000 2.980000 ;
      RECT  0.995000  0.980000  1.850000 1.150000 ;
      RECT  0.995000  1.150000  1.325000 1.950000 ;
      RECT  0.995000  1.950000  2.365000 2.120000 ;
      RECT  1.035000  2.630000  1.285000 3.245000 ;
      RECT  1.040000  0.085000  1.370000 0.810000 ;
      RECT  1.455000  2.460000  1.625000 2.905000 ;
      RECT  1.455000  2.905000  2.305000 3.075000 ;
      RECT  1.600000  0.545000  1.850000 0.980000 ;
      RECT  1.795000  2.120000  1.965000 2.735000 ;
      RECT  2.030000  0.085000  2.360000 1.005000 ;
      RECT  2.115000  1.520000  2.365000 1.950000 ;
      RECT  2.135000  2.290000  3.485000 2.460000 ;
      RECT  2.135000  2.460000  2.305000 2.905000 ;
      RECT  2.475000  2.630000  2.725000 3.245000 ;
      RECT  2.535000  1.520000  3.055000 1.850000 ;
      RECT  2.850000  0.545000  3.180000 1.175000 ;
      RECT  2.850000  1.175000  3.485000 1.345000 ;
      RECT  3.235000  2.460000  3.485000 2.975000 ;
      RECT  3.315000  1.345000  3.485000 2.290000 ;
      RECT  3.350000  0.675000  3.825000 1.005000 ;
      RECT  3.655000  1.005000  3.825000 2.295000 ;
      RECT  3.655000  2.295000  3.935000 2.905000 ;
      RECT  3.655000  2.905000  4.800000 3.075000 ;
      RECT  3.995000  0.255000  4.275000 0.605000 ;
      RECT  3.995000  0.605000  4.585000 1.010000 ;
      RECT  3.995000  1.010000  4.275000 1.915000 ;
      RECT  3.995000  1.915000  5.860000 2.085000 ;
      RECT  4.105000  2.085000  4.275000 2.255000 ;
      RECT  4.105000  2.255000  4.460000 2.735000 ;
      RECT  4.630000  2.255000  6.200000 2.335000 ;
      RECT  4.630000  2.335000  8.325000 2.425000 ;
      RECT  4.630000  2.425000  4.800000 2.905000 ;
      RECT  4.765000  0.085000  5.095000 1.010000 ;
      RECT  4.970000  2.595000  5.220000 3.245000 ;
      RECT  5.555000  0.605000  5.885000 1.075000 ;
      RECT  5.555000  1.075000  6.200000 1.245000 ;
      RECT  5.580000  1.415000  5.860000 1.915000 ;
      RECT  5.730000  2.425000  8.325000 2.505000 ;
      RECT  5.730000  2.505000  6.060000 2.935000 ;
      RECT  6.030000  1.245000  6.200000 2.255000 ;
      RECT  6.110000  0.085000  6.360000 0.905000 ;
      RECT  6.260000  2.675000  6.590000 3.245000 ;
      RECT  6.540000  0.350000  6.870000 0.840000 ;
      RECT  6.540000  0.840000  7.415000 1.010000 ;
      RECT  6.710000  1.785000  7.490000 2.165000 ;
      RECT  7.095000  0.085000  7.425000 0.670000 ;
      RECT  7.245000  1.010000  7.415000 1.785000 ;
      RECT  7.605000  0.255000  9.505000 0.425000 ;
      RECT  7.605000  0.425000  7.855000 1.130000 ;
      RECT  7.610000  2.675000  7.940000 3.245000 ;
      RECT  7.720000  1.480000  8.325000 1.650000 ;
      RECT  7.720000  1.650000  7.890000 2.335000 ;
      RECT  8.060000  1.820000  8.665000 1.995000 ;
      RECT  8.060000  1.995000  8.830000 2.165000 ;
      RECT  8.075000  0.595000  8.325000 1.480000 ;
      RECT  8.155000  2.505000  8.830000 2.980000 ;
      RECT  8.495000  0.425000  8.665000 1.820000 ;
      RECT  8.495000  2.165000  8.830000 2.335000 ;
      RECT  8.835000  0.595000  9.005000 1.630000 ;
      RECT  8.835000  1.630000 10.585000 1.800000 ;
      RECT  9.000000  1.800000  9.170000 2.520000 ;
      RECT  9.000000  2.520000  9.360000 2.980000 ;
      RECT  9.175000  0.425000  9.505000 0.860000 ;
      RECT  9.175000  0.860000 10.430000 1.030000 ;
      RECT  9.175000  1.030000  9.505000 1.255000 ;
      RECT  9.340000  2.000000  9.700000 2.330000 ;
      RECT  9.530000  2.330000  9.700000 2.390000 ;
      RECT  9.530000  2.390000 12.295000 2.560000 ;
      RECT  9.715000  1.200000 11.475000 1.370000 ;
      RECT  9.715000  1.370000 10.045000 1.405000 ;
      RECT  9.840000  0.085000 10.090000 0.690000 ;
      RECT  9.960000  2.730000 10.290000 3.245000 ;
      RECT 10.255000  1.540000 10.585000 1.630000 ;
      RECT 10.260000  0.255000 11.110000 0.425000 ;
      RECT 10.260000  0.425000 10.430000 0.860000 ;
      RECT 10.475000  1.970000 10.925000 2.220000 ;
      RECT 10.600000  0.595000 10.770000 1.200000 ;
      RECT 10.755000  1.370000 11.475000 1.530000 ;
      RECT 10.755000  1.530000 10.925000 1.970000 ;
      RECT 10.940000  0.425000 11.110000 0.860000 ;
      RECT 10.940000  0.860000 11.855000 1.030000 ;
      RECT 10.995000  2.730000 11.325000 3.245000 ;
      RECT 11.280000  0.085000 11.530000 0.690000 ;
      RECT 11.685000  1.030000 11.855000 1.190000 ;
      RECT 11.685000  1.190000 13.095000 1.360000 ;
      RECT 11.685000  1.360000 11.955000 1.800000 ;
      RECT 12.035000  0.350000 12.365000 0.850000 ;
      RECT 12.035000  0.850000 13.435000 0.990000 ;
      RECT 12.035000  0.990000 14.055000 1.020000 ;
      RECT 12.125000  1.530000 12.555000 1.755000 ;
      RECT 12.125000  1.755000 12.295000 2.390000 ;
      RECT 12.465000  1.925000 12.895000 2.980000 ;
      RECT 12.725000  1.755000 14.055000 1.925000 ;
      RECT 12.765000  1.360000 13.095000 1.585000 ;
      RECT 12.855000  0.085000 13.835000 0.680000 ;
      RECT 13.155000  2.095000 13.485000 2.180000 ;
      RECT 13.155000  2.180000 14.395000 2.350000 ;
      RECT 13.265000  1.020000 14.055000 1.755000 ;
      RECT 13.335000  2.650000 13.875000 3.245000 ;
      RECT 13.725000  0.980000 14.055000 0.990000 ;
      RECT 13.725000  1.925000 14.055000 1.990000 ;
      RECT 14.005000  0.350000 14.395000 0.810000 ;
      RECT 14.045000  2.350000 14.395000 2.980000 ;
      RECT 14.225000  0.810000 14.395000 1.550000 ;
      RECT 14.225000  1.550000 14.755000 1.780000 ;
      RECT 14.225000  1.780000 14.395000 2.180000 ;
      RECT 14.565000  0.085000 14.895000 1.340000 ;
      RECT 14.565000  1.950000 14.895000 3.245000 ;
      RECT 15.465000  2.320000 15.795000 3.245000 ;
      RECT 15.495000  0.085000 15.825000 0.920000 ;
      RECT 16.365000  2.320000 16.695000 3.245000 ;
      RECT 16.370000  0.085000 16.700000 0.920000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  1.580000  2.725000 1.750000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  1.580000 14.725000 1.750000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.245000 15.205000 3.415000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.245000 15.685000 3.415000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.245000 16.165000 3.415000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  3.245000 16.645000 3.415000 ;
    LAYER met1 ;
      RECT  2.495000 1.550000  2.785000 1.595000 ;
      RECT  2.495000 1.595000 14.785000 1.735000 ;
      RECT  2.495000 1.735000  2.785000 1.780000 ;
      RECT 14.495000 1.550000 14.785000 1.595000 ;
      RECT 14.495000 1.735000 14.785000 1.780000 ;
  END
END sky130_fd_sc_hs__sedfxtp_4
MACRO sky130_fd_sc_hs__tap_1
  CLASS CORE WELLTAP ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.480000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 0.480000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.265000 0.390000 1.440000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.890000 0.390000 3.065000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 0.480000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.480000 0.085000 ;
      RECT 0.000000  3.245000 0.480000 3.415000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
  END
END sky130_fd_sc_hs__tap_1
MACRO sky130_fd_sc_hs__tap_2
  CLASS CORE WELLTAP ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.960000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 0.960000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.265000 0.870000 1.440000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.890000 0.870000 3.065000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 0.960000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.960000 0.085000 ;
      RECT 0.000000  3.245000 0.960000 3.415000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
  END
END sky130_fd_sc_hs__tap_2
MACRO sky130_fd_sc_hs__tapmet1_2
  CLASS CORE WELLTAP ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.960000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 0.960000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.080000 0.425000 0.400000 0.685000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.560000 2.645000 0.880000 2.905000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 0.960000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.960000 0.085000 ;
      RECT 0.000000  3.245000 0.960000 3.415000 ;
      RECT 0.090000  0.265000 0.870000 1.105000 ;
      RECT 0.090000  2.210000 0.870000 3.065000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  0.470000 0.325000 0.640000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  2.690000 0.805000 2.860000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
  END
END sky130_fd_sc_hs__tapmet1_2
MACRO sky130_fd_sc_hs__tapvgnd_1
  CLASS CORE WELLTAP ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.480000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 0.480000 0.245000 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.080000 2.645000 0.400000 2.905000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 0.480000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.480000 0.085000 ;
      RECT 0.000000  3.245000 0.480000 3.415000 ;
      RECT 0.090000  0.085000 0.390000 1.440000 ;
      RECT 0.090000  1.890000 0.390000 3.065000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  2.690000 0.325000 2.860000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
  END
END sky130_fd_sc_hs__tapvgnd_1
MACRO sky130_fd_sc_hs__tapvgnd2_1
  CLASS CORE WELLTAP ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.480000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 0.480000 0.245000 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.080000 2.275000 0.400000 2.535000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 0.480000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.480000 0.085000 ;
      RECT 0.000000  3.245000 0.480000 3.415000 ;
      RECT 0.090000  0.085000 0.390000 1.440000 ;
      RECT 0.090000  1.890000 0.390000 3.065000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  2.320000 0.325000 2.490000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
  END
END sky130_fd_sc_hs__tapvgnd2_1
MACRO sky130_fd_sc_hs__tapvpwrvgnd_1
  CLASS CORE WELLTAP ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.480000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 0.480000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 0.480000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.480000 0.085000 ;
      RECT 0.000000  3.245000 0.480000 3.415000 ;
      RECT 0.090000  0.085000 0.390000 1.105000 ;
      RECT 0.090000  2.205000 0.390000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
  END
END sky130_fd_sc_hs__tapvpwrvgnd_1
MACRO sky130_fd_sc_hs__xnor2_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.501000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.515000 1.350000 1.845000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.501000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945000 1.435000 1.345000 1.780000 ;
        RECT 1.175000 1.780000 1.345000 1.950000 ;
        RECT 1.175000 1.950000 2.185000 2.120000 ;
        RECT 2.015000 1.350000 2.465000 1.680000 ;
        RECT 2.015000 1.680000 2.185000 1.950000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.699800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 2.290000 2.685000 2.980000 ;
        RECT 2.355000 1.850000 3.275000 2.020000 ;
        RECT 2.355000 2.020000 2.685000 2.290000 ;
        RECT 2.975000 0.350000 3.275000 1.130000 ;
        RECT 3.105000 1.130000 3.275000 1.850000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.105000  0.085000 0.435000 1.255000 ;
      RECT 0.175000  1.905000 0.425000 2.290000 ;
      RECT 0.175000  2.290000 0.505000 3.245000 ;
      RECT 0.605000  1.085000 2.805000 1.180000 ;
      RECT 0.605000  1.180000 1.225000 1.255000 ;
      RECT 0.605000  1.255000 0.775000 1.950000 ;
      RECT 0.605000  1.950000 1.005000 2.120000 ;
      RECT 0.675000  2.120000 1.005000 2.785000 ;
      RECT 0.895000  0.575000 1.225000 1.010000 ;
      RECT 0.895000  1.010000 2.805000 1.085000 ;
      RECT 1.415000  2.290000 1.745000 3.245000 ;
      RECT 1.435000  0.510000 1.765000 0.670000 ;
      RECT 1.435000  0.670000 2.770000 0.840000 ;
      RECT 1.935000  0.085000 2.265000 0.500000 ;
      RECT 2.440000  0.510000 2.770000 0.670000 ;
      RECT 2.635000  1.180000 2.805000 1.300000 ;
      RECT 2.635000  1.300000 2.935000 1.630000 ;
      RECT 2.855000  2.190000 3.185000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__xnor2_1
MACRO sky130_fd_sc_hs__xnor2_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAPARTIALMETALSIDEAREA  2.107000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.180000 3.355000 1.550000 ;
        RECT 3.025000 1.550000 3.355000 1.720000 ;
        RECT 3.025000 1.720000 4.675000 1.890000 ;
        RECT 4.445000 1.350000 4.855000 1.680000 ;
        RECT 4.445000 1.680000 4.675000 1.720000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.819000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.345000 1.350000 1.675000 1.720000 ;
        RECT 1.345000 1.720000 2.775000 1.890000 ;
        RECT 2.605000 1.890000 2.775000 2.060000 ;
        RECT 2.605000 2.060000 5.195000 2.230000 ;
        RECT 3.925000 1.010000 5.195000 1.180000 ;
        RECT 3.925000 1.180000 4.255000 1.550000 ;
        RECT 5.025000 1.180000 5.195000 2.060000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.072800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.840000 0.835000 1.010000 ;
        RECT 0.085000 1.010000 0.255000 2.320000 ;
        RECT 0.085000 2.320000 2.435000 2.400000 ;
        RECT 0.085000 2.400000 4.135000 2.490000 ;
        RECT 0.665000 0.255000 2.575000 0.425000 ;
        RECT 0.665000 0.425000 0.835000 0.840000 ;
        RECT 2.045000 2.060000 2.435000 2.320000 ;
        RECT 2.045000 2.490000 4.135000 2.570000 ;
        RECT 2.045000 2.570000 2.435000 2.980000 ;
        RECT 2.190000 0.425000 2.575000 0.500000 ;
        RECT 3.805000 2.570000 4.135000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.280000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.245000 5.280000 3.415000 ;
      RECT 0.115000  0.085000 0.495000 0.670000 ;
      RECT 0.115000  2.660000 0.445000 3.245000 ;
      RECT 0.425000  1.180000 0.835000 1.550000 ;
      RECT 0.650000  1.820000 1.175000 2.150000 ;
      RECT 1.005000  0.635000 1.450000 1.010000 ;
      RECT 1.005000  1.010000 2.585000 1.180000 ;
      RECT 1.005000  1.180000 1.175000 1.820000 ;
      RECT 1.230000  2.660000 1.875000 3.245000 ;
      RECT 1.680000  0.595000 2.010000 0.670000 ;
      RECT 1.680000  0.670000 5.165000 0.840000 ;
      RECT 1.915000  1.180000 2.585000 1.550000 ;
      RECT 2.640000  2.740000 2.970000 3.245000 ;
      RECT 2.755000  0.350000 3.085000 0.670000 ;
      RECT 2.755000  0.840000 3.085000 1.010000 ;
      RECT 3.260000  2.740000 3.600000 2.905000 ;
      RECT 3.260000  2.905000 4.635000 3.075000 ;
      RECT 3.265000  0.085000 3.600000 0.500000 ;
      RECT 3.780000  0.490000 4.110000 0.670000 ;
      RECT 4.305000  2.400000 4.635000 2.905000 ;
      RECT 4.310000  0.085000 4.655000 0.500000 ;
      RECT 4.805000  2.400000 5.135000 3.245000 ;
      RECT 4.835000  0.490000 5.165000 0.670000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  1.210000 0.805000 1.380000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  1.210000 3.205000 1.380000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
    LAYER met1 ;
      RECT 0.575000 1.180000 0.865000 1.225000 ;
      RECT 0.575000 1.225000 3.265000 1.365000 ;
      RECT 0.575000 1.365000 0.865000 1.410000 ;
      RECT 2.975000 1.180000 3.265000 1.225000 ;
      RECT 2.975000 1.365000 3.265000 1.410000 ;
  END
END sky130_fd_sc_hs__xnor2_2
MACRO sky130_fd_sc_hs__xnor2_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAPARTIALMETALSIDEAREA  2.779000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.350000 5.835000 1.775000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.560000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 1.350000 2.155000 1.680000 ;
        RECT 1.985000 1.680000 2.155000 1.945000 ;
        RECT 1.985000 1.945000 6.535000 2.115000 ;
        RECT 6.365000 1.350000 8.155000 1.765000 ;
        RECT 6.365000 1.765000 6.535000 1.945000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.474200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.545000 2.285000 7.655000 2.455000 ;
        RECT 3.035000 0.595000 3.365000 1.010000 ;
        RECT 3.035000 1.010000 8.495000 1.180000 ;
        RECT 4.060000 0.595000 4.390000 1.010000 ;
        RECT 7.325000 1.935000 8.555000 2.105000 ;
        RECT 7.325000 2.105000 7.655000 2.285000 ;
        RECT 7.325000 2.455000 7.655000 2.735000 ;
        RECT 8.225000 2.105000 8.555000 2.735000 ;
        RECT 8.325000 1.180000 8.495000 1.935000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.120000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.120000 0.085000 ;
      RECT 0.000000  3.245000 9.120000 3.415000 ;
      RECT 0.115000  0.350000 0.365000 0.980000 ;
      RECT 0.115000  0.980000 1.375000 1.150000 ;
      RECT 0.115000  1.820000 0.365000 3.245000 ;
      RECT 0.545000  0.085000 0.875000 0.810000 ;
      RECT 0.545000  1.320000 1.315000 1.650000 ;
      RECT 0.565000  1.820000 0.895000 1.950000 ;
      RECT 0.565000  1.950000 1.795000 2.120000 ;
      RECT 0.565000  2.120000 0.895000 2.700000 ;
      RECT 1.045000  0.350000 2.305000 0.600000 ;
      RECT 1.045000  0.600000 1.375000 0.980000 ;
      RECT 1.085000  1.650000 1.315000 1.780000 ;
      RECT 1.095000  2.290000 1.265000 3.245000 ;
      RECT 1.465000  2.120000 1.795000 2.625000 ;
      RECT 1.465000  2.625000 4.590000 2.795000 ;
      RECT 1.545000  0.770000 1.875000 1.010000 ;
      RECT 1.545000  1.010000 2.565000 1.180000 ;
      RECT 2.000000  2.965000 2.340000 3.245000 ;
      RECT 2.395000  1.180000 2.565000 1.350000 ;
      RECT 2.395000  1.350000 4.085000 1.680000 ;
      RECT 2.535000  0.255000 4.890000 0.425000 ;
      RECT 2.535000  0.425000 2.865000 0.840000 ;
      RECT 3.080000  2.965000 3.410000 3.245000 ;
      RECT 3.535000  0.425000 3.865000 0.840000 ;
      RECT 3.580000  2.795000 4.590000 2.955000 ;
      RECT 4.560000  0.425000 4.890000 0.670000 ;
      RECT 4.560000  0.670000 9.005000 0.840000 ;
      RECT 4.810000  2.625000 7.125000 2.795000 ;
      RECT 4.810000  2.795000 5.060000 2.980000 ;
      RECT 5.070000  0.085000 5.400000 0.500000 ;
      RECT 5.265000  2.965000 5.600000 3.245000 ;
      RECT 5.580000  0.350000 5.910000 0.670000 ;
      RECT 5.805000  2.795000 6.135000 2.980000 ;
      RECT 6.090000  0.085000 6.420000 0.500000 ;
      RECT 6.340000  2.965000 6.670000 3.245000 ;
      RECT 6.600000  0.350000 6.930000 0.670000 ;
      RECT 6.875000  2.795000 7.125000 2.905000 ;
      RECT 6.875000  2.905000 9.005000 3.075000 ;
      RECT 7.110000  0.085000 7.475000 0.500000 ;
      RECT 7.655000  0.350000 7.985000 0.670000 ;
      RECT 7.855000  2.275000 8.025000 2.905000 ;
      RECT 8.165000  0.085000 8.495000 0.500000 ;
      RECT 8.675000  0.350000 9.005000 0.670000 ;
      RECT 8.675000  0.840000 9.005000 1.130000 ;
      RECT 8.755000  1.935000 9.005000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  1.580000 1.285000 1.750000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  1.580000 4.645000 1.750000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
    LAYER met1 ;
      RECT 1.055000 1.550000 1.345000 1.595000 ;
      RECT 1.055000 1.595000 4.705000 1.735000 ;
      RECT 1.055000 1.735000 1.345000 1.780000 ;
      RECT 4.415000 1.550000 4.705000 1.595000 ;
      RECT 4.415000 1.735000 4.705000 1.780000 ;
  END
END sky130_fd_sc_hs__xnor2_4
MACRO sky130_fd_sc_hs__xnor3_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.845000 1.425000 7.205000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.693000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.705000 1.350000 4.375000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.995000 1.350000 1.325000 1.780000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.530100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.440000 0.445000 1.170000 ;
        RECT 0.085000 1.170000 0.255000 1.840000 ;
        RECT 0.085000 1.840000 0.355000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.425000  1.340000 0.785000 1.670000 ;
      RECT 0.555000  2.290000 0.805000 3.245000 ;
      RECT 0.615000  0.660000 1.665000 0.830000 ;
      RECT 0.615000  0.830000 0.785000 1.340000 ;
      RECT 0.615000  1.670000 0.785000 1.950000 ;
      RECT 0.615000  1.950000 1.145000 2.120000 ;
      RECT 0.625000  0.085000 0.955000 0.490000 ;
      RECT 0.975000  2.120000 1.145000 2.905000 ;
      RECT 0.975000  2.905000 2.655000 3.075000 ;
      RECT 1.135000  1.000000 1.665000 1.170000 ;
      RECT 1.315000  1.950000 1.665000 2.500000 ;
      RECT 1.495000  0.255000 2.665000 0.425000 ;
      RECT 1.495000  0.425000 1.665000 0.660000 ;
      RECT 1.495000  1.170000 1.665000 1.580000 ;
      RECT 1.495000  1.580000 2.845000 1.750000 ;
      RECT 1.495000  1.750000 1.665000 1.950000 ;
      RECT 1.835000  0.595000 2.165000 1.140000 ;
      RECT 1.835000  1.140000 3.185000 1.310000 ;
      RECT 1.835000  1.310000 2.275000 1.410000 ;
      RECT 1.875000  1.950000 2.125000 2.370000 ;
      RECT 1.875000  2.370000 5.265000 2.540000 ;
      RECT 1.875000  2.540000 2.125000 2.735000 ;
      RECT 2.325000  2.710000 2.655000 2.905000 ;
      RECT 2.335000  0.425000 2.665000 0.970000 ;
      RECT 2.515000  1.480000 2.845000 1.580000 ;
      RECT 2.515000  1.750000 2.845000 1.810000 ;
      RECT 2.835000  0.350000 3.165000 0.670000 ;
      RECT 2.835000  0.670000 6.535000 0.765000 ;
      RECT 2.835000  0.765000 5.180000 0.840000 ;
      RECT 2.835000  0.840000 3.525000 0.970000 ;
      RECT 2.850000  2.030000 3.185000 2.200000 ;
      RECT 3.015000  1.310000 3.185000 2.030000 ;
      RECT 3.355000  0.970000 3.525000 2.370000 ;
      RECT 3.395000  0.085000 3.725000 0.500000 ;
      RECT 3.395000  2.710000 3.725000 3.245000 ;
      RECT 3.905000  1.010000 4.715000 1.180000 ;
      RECT 3.920000  1.950000 4.715000 2.200000 ;
      RECT 4.465000  0.255000 7.035000 0.425000 ;
      RECT 4.465000  0.425000 4.840000 0.500000 ;
      RECT 4.490000  2.710000 4.820000 2.905000 ;
      RECT 4.490000  2.905000 7.090000 3.075000 ;
      RECT 4.545000  1.180000 4.715000 1.355000 ;
      RECT 4.545000  1.355000 5.045000 1.685000 ;
      RECT 4.545000  1.685000 4.715000 1.950000 ;
      RECT 5.010000  0.595000 6.535000 0.670000 ;
      RECT 5.015000  1.855000 5.265000 2.370000 ;
      RECT 5.015000  2.540000 5.265000 2.575000 ;
      RECT 5.020000  1.015000 5.485000 1.180000 ;
      RECT 5.020000  1.180000 5.605000 1.185000 ;
      RECT 5.315000  1.185000 5.605000 1.410000 ;
      RECT 5.435000  1.410000 5.605000 1.765000 ;
      RECT 5.435000  1.765000 6.250000 1.935000 ;
      RECT 5.550000  2.105000 5.880000 2.565000 ;
      RECT 5.550000  2.565000 6.590000 2.735000 ;
      RECT 5.775000  0.935000 6.085000 1.425000 ;
      RECT 5.775000  1.425000 6.590000 1.595000 ;
      RECT 6.080000  1.935000 6.250000 2.395000 ;
      RECT 6.255000  0.765000 6.535000 1.210000 ;
      RECT 6.420000  1.595000 6.590000 2.565000 ;
      RECT 6.705000  0.425000 7.035000 1.085000 ;
      RECT 6.705000  1.085000 7.620000 1.255000 ;
      RECT 6.760000  1.950000 7.620000 2.120000 ;
      RECT 6.760000  2.120000 7.090000 2.905000 ;
      RECT 7.205000  0.085000 7.615000 0.915000 ;
      RECT 7.260000  2.290000 7.590000 3.245000 ;
      RECT 7.415000  1.255000 7.620000 1.425000 ;
      RECT 7.415000  1.425000 7.665000 1.755000 ;
      RECT 7.415000  1.755000 7.620000 1.950000 ;
      RECT 7.790000  2.190000 8.075000 2.930000 ;
      RECT 7.795000  0.585000 8.075000 1.255000 ;
      RECT 7.835000  1.255000 8.075000 2.190000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  1.210000 2.245000 1.380000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  1.210000 5.605000 1.380000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  1.210000 6.085000 1.380000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  1.210000 8.005000 1.380000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
    LAYER met1 ;
      RECT 2.015000 1.180000 2.305000 1.225000 ;
      RECT 2.015000 1.225000 5.665000 1.365000 ;
      RECT 2.015000 1.365000 2.305000 1.410000 ;
      RECT 5.375000 1.180000 5.665000 1.225000 ;
      RECT 5.375000 1.365000 5.665000 1.410000 ;
      RECT 5.855000 1.180000 6.145000 1.225000 ;
      RECT 5.855000 1.225000 8.065000 1.365000 ;
      RECT 5.855000 1.365000 6.145000 1.410000 ;
      RECT 7.775000 1.180000 8.065000 1.225000 ;
      RECT 7.775000 1.365000 8.065000 1.410000 ;
  END
END sky130_fd_sc_hs__xnor3_1
MACRO sky130_fd_sc_hs__xnor3_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955000 1.375000 1.315000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.693000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.735000 1.350000 4.405000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.845000 1.350000 7.175000 1.780000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.750000 1.840000 8.095000 2.980000 ;
        RECT 7.765000 0.440000 8.095000 1.170000 ;
        RECT 7.925000 1.170000 8.095000 1.840000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
      RECT 0.000000  3.245000 8.640000 3.415000 ;
      RECT 0.085000  0.385000 0.405000 1.065000 ;
      RECT 0.085000  1.065000 0.325000 2.290000 ;
      RECT 0.085000  2.290000 0.445000 2.885000 ;
      RECT 0.495000  1.235000 0.745000 1.950000 ;
      RECT 0.495000  1.950000 1.375000 2.120000 ;
      RECT 0.575000  1.035000 1.345000 1.205000 ;
      RECT 0.575000  1.205000 0.745000 1.235000 ;
      RECT 0.585000  0.085000 0.915000 0.865000 ;
      RECT 0.645000  2.305000 0.925000 3.245000 ;
      RECT 1.095000  0.255000 3.530000 0.425000 ;
      RECT 1.095000  0.425000 1.345000 1.035000 ;
      RECT 1.095000  2.120000 1.375000 2.905000 ;
      RECT 1.095000  2.905000 3.675000 3.075000 ;
      RECT 1.545000  1.165000 2.385000 1.380000 ;
      RECT 1.545000  1.380000 1.715000 2.565000 ;
      RECT 1.545000  2.565000 2.605000 2.735000 ;
      RECT 1.625000  0.595000 2.725000 0.615000 ;
      RECT 1.625000  0.615000 5.160000 0.765000 ;
      RECT 1.625000  0.765000 1.955000 0.995000 ;
      RECT 1.885000  1.550000 2.755000 1.720000 ;
      RECT 1.885000  1.720000 2.105000 2.395000 ;
      RECT 2.135000  0.935000 2.385000 1.165000 ;
      RECT 2.275000  1.890000 2.605000 2.565000 ;
      RECT 2.555000  0.765000 5.160000 0.785000 ;
      RECT 2.555000  0.955000 2.985000 1.285000 ;
      RECT 2.555000  1.285000 2.755000 1.550000 ;
      RECT 2.835000  1.875000 3.145000 2.370000 ;
      RECT 2.835000  2.370000 4.755000 2.395000 ;
      RECT 2.835000  2.395000 6.320000 2.540000 ;
      RECT 2.835000  2.540000 3.065000 2.620000 ;
      RECT 3.155000  1.375000 3.565000 1.705000 ;
      RECT 3.200000  0.425000 3.530000 0.445000 ;
      RECT 3.345000  2.710000 3.675000 2.905000 ;
      RECT 3.395000  0.955000 4.090000 1.125000 ;
      RECT 3.395000  1.125000 3.565000 1.375000 ;
      RECT 3.395000  1.705000 3.565000 1.950000 ;
      RECT 3.395000  1.950000 4.255000 2.200000 ;
      RECT 4.270000  0.085000 4.600000 0.445000 ;
      RECT 4.455000  2.735000 4.785000 3.245000 ;
      RECT 4.585000  0.785000 5.160000 0.965000 ;
      RECT 4.585000  0.965000 4.755000 2.370000 ;
      RECT 4.585000  2.540000 6.320000 2.565000 ;
      RECT 4.830000  0.350000 5.160000 0.615000 ;
      RECT 4.925000  1.135000 6.160000 1.305000 ;
      RECT 4.925000  1.305000 5.155000 1.975000 ;
      RECT 4.925000  1.975000 5.335000 2.225000 ;
      RECT 5.325000  1.475000 6.675000 1.805000 ;
      RECT 5.330000  0.255000 6.500000 0.425000 ;
      RECT 5.330000  0.425000 5.660000 0.965000 ;
      RECT 5.535000  2.735000 5.865000 2.905000 ;
      RECT 5.535000  2.905000 7.210000 3.075000 ;
      RECT 5.830000  0.595000 6.160000 1.135000 ;
      RECT 6.070000  1.975000 6.320000 2.395000 ;
      RECT 6.070000  2.565000 6.320000 2.735000 ;
      RECT 6.330000  0.425000 6.500000 0.660000 ;
      RECT 6.330000  0.660000 7.060000 0.830000 ;
      RECT 6.390000  1.000000 6.720000 1.170000 ;
      RECT 6.390000  1.170000 6.675000 1.475000 ;
      RECT 6.505000  1.805000 6.675000 1.950000 ;
      RECT 6.505000  1.950000 6.870000 2.500000 ;
      RECT 6.890000  0.830000 7.060000 1.010000 ;
      RECT 6.890000  1.010000 7.580000 1.180000 ;
      RECT 6.900000  0.085000 7.585000 0.490000 ;
      RECT 7.040000  1.950000 7.580000 2.120000 ;
      RECT 7.040000  2.120000 7.210000 2.905000 ;
      RECT 7.230000  0.490000 7.585000 0.840000 ;
      RECT 7.380000  2.290000 7.550000 3.245000 ;
      RECT 7.410000  1.180000 7.580000 1.340000 ;
      RECT 7.410000  1.340000 7.755000 1.670000 ;
      RECT 7.410000  1.670000 7.580000 1.950000 ;
      RECT 8.275000  0.085000 8.525000 1.250000 ;
      RECT 8.280000  1.820000 8.530000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  1.210000 0.325000 1.380000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  1.210000 1.765000 1.380000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  1.210000 2.725000 1.380000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  1.210000 5.125000 1.380000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
    LAYER met1 ;
      RECT 0.095000 1.180000 0.385000 1.225000 ;
      RECT 0.095000 1.225000 1.825000 1.365000 ;
      RECT 0.095000 1.365000 0.385000 1.410000 ;
      RECT 1.535000 1.180000 1.825000 1.225000 ;
      RECT 1.535000 1.365000 1.825000 1.410000 ;
      RECT 2.495000 1.180000 2.785000 1.225000 ;
      RECT 2.495000 1.225000 5.185000 1.365000 ;
      RECT 2.495000 1.365000 2.785000 1.410000 ;
      RECT 4.895000 1.180000 5.185000 1.225000 ;
      RECT 4.895000 1.365000 5.185000 1.410000 ;
  END
END sky130_fd_sc_hs__xnor3_2
MACRO sky130_fd_sc_hs__xnor3_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.915000 1.375000 1.315000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.693000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.940000 1.350000 4.270000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.780000 1.350000 7.110000 1.780000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.280000 1.840000 8.640000 2.980000 ;
        RECT 8.345000 0.470000 8.675000 1.170000 ;
        RECT 8.470000 1.170000 8.675000 1.420000 ;
        RECT 8.470000 1.420000 9.535000 1.625000 ;
        RECT 8.470000 1.625000 8.640000 1.840000 ;
        RECT 9.180000 1.625000 9.535000 2.980000 ;
        RECT 9.205000 0.440000 9.535000 1.420000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.085000  0.365000  0.495000 0.865000 ;
      RECT 0.085000  0.865000  0.285000 1.845000 ;
      RECT 0.085000  1.845000  0.365000 2.885000 ;
      RECT 0.455000  1.035000  1.425000 1.205000 ;
      RECT 0.455000  1.205000  0.705000 1.465000 ;
      RECT 0.535000  1.465000  0.705000 1.950000 ;
      RECT 0.535000  1.950000  1.395000 2.120000 ;
      RECT 0.565000  2.290000  0.895000 3.245000 ;
      RECT 0.665000  0.085000  0.995000 0.865000 ;
      RECT 1.065000  2.120000  1.395000 2.905000 ;
      RECT 1.065000  2.905000  3.680000 3.075000 ;
      RECT 1.175000  0.255000  3.530000 0.425000 ;
      RECT 1.175000  0.425000  1.425000 1.035000 ;
      RECT 1.565000  1.375000  1.765000 2.565000 ;
      RECT 1.565000  2.565000  2.725000 2.735000 ;
      RECT 1.595000  1.165000  2.385000 1.335000 ;
      RECT 1.595000  1.335000  1.765000 1.375000 ;
      RECT 1.625000  0.595000  2.725000 0.615000 ;
      RECT 1.625000  0.615000  5.160000 0.765000 ;
      RECT 1.625000  0.765000  1.955000 0.995000 ;
      RECT 1.935000  1.505000  2.755000 1.675000 ;
      RECT 1.935000  1.675000  2.245000 2.120000 ;
      RECT 1.935000  2.120000  2.135000 2.155000 ;
      RECT 2.135000  0.935000  2.385000 1.165000 ;
      RECT 2.305000  2.290000  2.725000 2.565000 ;
      RECT 2.555000  0.765000  5.160000 0.785000 ;
      RECT 2.555000  0.955000  3.020000 1.205000 ;
      RECT 2.555000  1.205000  2.755000 1.505000 ;
      RECT 2.895000  1.875000  3.145000 2.370000 ;
      RECT 2.895000  2.370000  4.610000 2.390000 ;
      RECT 2.895000  2.390000  6.270000 2.540000 ;
      RECT 2.895000  2.540000  3.145000 2.545000 ;
      RECT 2.995000  1.375000  3.770000 1.705000 ;
      RECT 3.200000  0.425000  3.530000 0.445000 ;
      RECT 3.350000  2.710000  3.680000 2.905000 ;
      RECT 3.600000  0.955000  4.090000 1.125000 ;
      RECT 3.600000  1.125000  3.770000 1.375000 ;
      RECT 3.600000  1.705000  3.770000 1.950000 ;
      RECT 3.600000  1.950000  4.270000 2.200000 ;
      RECT 4.270000  0.085000  4.600000 0.445000 ;
      RECT 4.390000  2.730000  4.720000 3.245000 ;
      RECT 4.440000  0.785000  5.160000 1.030000 ;
      RECT 4.440000  1.030000  4.610000 2.370000 ;
      RECT 4.440000  2.540000  6.270000 2.560000 ;
      RECT 4.780000  1.210000  6.160000 1.380000 ;
      RECT 4.780000  1.380000  4.950000 1.950000 ;
      RECT 4.780000  1.950000  5.280000 2.220000 ;
      RECT 4.830000  0.350000  5.160000 0.615000 ;
      RECT 5.120000  1.550000  6.610000 1.720000 ;
      RECT 5.120000  1.720000  5.450000 1.780000 ;
      RECT 5.330000  0.255000  6.500000 0.425000 ;
      RECT 5.330000  0.425000  5.660000 1.010000 ;
      RECT 5.405000  1.180000  6.160000 1.210000 ;
      RECT 5.485000  2.730000  5.815000 2.905000 ;
      RECT 5.485000  2.905000  7.315000 3.075000 ;
      RECT 5.830000  0.595000  6.160000 1.180000 ;
      RECT 6.020000  1.970000  6.270000 2.390000 ;
      RECT 6.020000  2.560000  6.270000 2.735000 ;
      RECT 6.330000  0.425000  6.500000 0.660000 ;
      RECT 6.330000  0.660000  7.060000 0.830000 ;
      RECT 6.390000  1.000000  6.720000 1.170000 ;
      RECT 6.390000  1.170000  6.610000 1.550000 ;
      RECT 6.440000  1.720000  6.610000 1.990000 ;
      RECT 6.440000  1.990000  6.960000 2.500000 ;
      RECT 6.890000  0.830000  7.060000 1.010000 ;
      RECT 6.890000  1.010000  7.490000 1.180000 ;
      RECT 6.900000  0.085000  8.165000 0.490000 ;
      RECT 7.130000  1.950000  7.490000 2.120000 ;
      RECT 7.130000  2.120000  7.315000 2.905000 ;
      RECT 7.230000  0.490000  8.165000 0.840000 ;
      RECT 7.320000  1.180000  7.490000 1.340000 ;
      RECT 7.320000  1.340000  8.300000 1.670000 ;
      RECT 7.320000  1.670000  7.490000 1.950000 ;
      RECT 7.485000  2.290000  8.110000 3.245000 ;
      RECT 7.685000  1.840000  8.110000 2.290000 ;
      RECT 7.915000  0.840000  8.165000 1.170000 ;
      RECT 8.810000  1.820000  8.980000 3.245000 ;
      RECT 8.855000  0.085000  9.025000 1.250000 ;
      RECT 9.710000  1.820000  9.960000 3.245000 ;
      RECT 9.715000  0.085000  9.965000 1.250000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  1.950000 0.325000 2.120000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  1.950000 1.765000 2.120000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  1.950000 2.245000 2.120000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  1.950000 5.125000 2.120000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
    LAYER met1 ;
      RECT 0.095000 1.920000 0.385000 1.965000 ;
      RECT 0.095000 1.965000 1.825000 2.105000 ;
      RECT 0.095000 2.105000 0.385000 2.150000 ;
      RECT 1.535000 1.920000 1.825000 1.965000 ;
      RECT 1.535000 2.105000 1.825000 2.150000 ;
      RECT 2.015000 1.920000 2.305000 1.965000 ;
      RECT 2.015000 1.965000 5.185000 2.105000 ;
      RECT 2.015000 2.105000 2.305000 2.150000 ;
      RECT 4.895000 1.920000 5.185000 1.965000 ;
      RECT 4.895000 2.105000 5.185000 2.150000 ;
  END
END sky130_fd_sc_hs__xnor3_4
MACRO sky130_fd_sc_hs__xor2_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.512000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.775000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.512000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.285000 1.365000 2.845000 1.695000 ;
        RECT 2.515000 1.350000 2.845000 1.365000 ;
        RECT 2.515000 1.695000 2.845000 1.780000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.697200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 0.415000 2.970000 0.980000 ;
        RECT 2.525000 0.980000 3.755000 1.150000 ;
        RECT 3.365000 1.820000 3.755000 2.980000 ;
        RECT 3.585000 1.150000 3.755000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.175000  0.085000 0.775000 0.990000 ;
      RECT 0.325000  1.940000 0.655000 3.245000 ;
      RECT 0.945000  0.710000 1.640000 1.040000 ;
      RECT 0.945000  1.040000 1.115000 1.950000 ;
      RECT 0.945000  1.950000 3.195000 2.120000 ;
      RECT 0.945000  2.120000 1.525000 2.980000 ;
      RECT 1.755000  2.290000 3.195000 2.460000 ;
      RECT 1.755000  2.460000 2.085000 2.980000 ;
      RECT 1.820000  0.085000 2.150000 1.195000 ;
      RECT 2.255000  2.650000 2.695000 3.245000 ;
      RECT 2.865000  2.460000 3.195000 2.980000 ;
      RECT 3.025000  1.320000 3.415000 1.650000 ;
      RECT 3.025000  1.650000 3.195000 1.950000 ;
      RECT 3.210000  0.085000 3.540000 0.745000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__xor2_1
MACRO sky130_fd_sc_hs__xor2_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.804000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.585000 1.165000 0.915000 1.620000 ;
        RECT 0.585000 1.620000 2.515000 1.790000 ;
        RECT 1.845000 1.350000 2.515000 1.620000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.804000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.155000 1.010000 4.145000 1.180000 ;
        RECT 1.155000 1.180000 1.485000 1.450000 ;
        RECT 3.485000 1.180000 4.145000 1.550000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.754100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.025000 1.850000 4.685000 2.020000 ;
        RECT 3.025000 2.020000 3.195000 2.735000 ;
        RECT 3.330000 0.595000 3.660000 0.670000 ;
        RECT 3.330000 0.670000 4.685000 0.840000 ;
        RECT 4.355000 0.350000 4.685000 0.670000 ;
        RECT 4.355000 0.840000 4.685000 1.850000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.115000  0.085000 0.710000 0.500000 ;
      RECT 0.115000  2.300000 0.445000 3.245000 ;
      RECT 0.245000  0.670000 1.220000 0.840000 ;
      RECT 0.245000  0.840000 0.415000 1.960000 ;
      RECT 0.245000  1.960000 2.855000 2.130000 ;
      RECT 0.890000  0.350000 1.220000 0.670000 ;
      RECT 1.065000  2.130000 1.315000 2.980000 ;
      RECT 1.390000  0.085000 1.720000 0.840000 ;
      RECT 1.545000  2.300000 2.825000 2.470000 ;
      RECT 1.545000  2.470000 1.795000 2.980000 ;
      RECT 1.970000  0.350000 2.300000 0.670000 ;
      RECT 1.970000  0.670000 3.160000 0.840000 ;
      RECT 1.995000  2.640000 2.325000 3.245000 ;
      RECT 2.480000  0.085000 2.820000 0.500000 ;
      RECT 2.495000  2.470000 2.825000 2.905000 ;
      RECT 2.495000  2.905000 3.675000 3.075000 ;
      RECT 2.685000  1.350000 3.125000 1.680000 ;
      RECT 2.685000  1.680000 2.855000 1.960000 ;
      RECT 2.990000  0.255000 4.175000 0.425000 ;
      RECT 2.990000  0.425000 3.160000 0.670000 ;
      RECT 3.395000  2.190000 4.685000 2.360000 ;
      RECT 3.395000  2.360000 3.675000 2.905000 ;
      RECT 3.840000  0.425000 4.175000 0.500000 ;
      RECT 3.845000  2.530000 4.175000 3.245000 ;
      RECT 4.345000  2.360000 4.685000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_hs__xor2_2
MACRO sky130_fd_sc_hs__xor2_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.638000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.440000 1.420000 1.110000 1.750000 ;
        RECT 0.515000 0.580000 1.445000 0.600000 ;
        RECT 0.515000 0.600000 3.040000 0.750000 ;
        RECT 0.515000 0.750000 0.685000 1.420000 ;
        RECT 1.275000 0.750000 3.040000 0.770000 ;
        RECT 2.870000 0.770000 3.040000 1.020000 ;
        RECT 2.870000 1.020000 3.935000 1.190000 ;
        RECT 3.765000 1.190000 3.935000 1.350000 ;
        RECT 3.765000 1.350000 5.635000 1.520000 ;
        RECT 3.965000 1.520000 5.635000 1.775000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.638000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.030000 1.470000 2.360000 1.850000 ;
        RECT 2.030000 1.850000 3.655000 1.945000 ;
        RECT 2.030000 1.945000 5.975000 2.020000 ;
        RECT 3.485000 2.020000 5.975000 2.115000 ;
        RECT 5.805000 1.550000 8.165000 1.780000 ;
        RECT 5.805000 1.780000 5.975000 1.945000 ;
        RECT 5.885000 1.350000 8.165000 1.550000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  1.504500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.985000 2.190000 3.315000 2.285000 ;
        RECT 2.985000 2.285000 6.315000 2.455000 ;
        RECT 2.985000 2.455000 3.315000 2.735000 ;
        RECT 3.210000 0.470000 3.540000 0.680000 ;
        RECT 3.210000 0.680000 4.275000 0.850000 ;
        RECT 3.885000 2.455000 4.215000 2.735000 ;
        RECT 4.105000 0.850000 4.275000 1.010000 ;
        RECT 4.105000 1.010000 8.505000 1.180000 ;
        RECT 6.145000 1.950000 8.505000 2.120000 ;
        RECT 6.145000 2.120000 6.315000 2.285000 ;
        RECT 6.835000 0.595000 7.165000 1.010000 ;
        RECT 7.845000 0.595000 8.015000 1.010000 ;
        RECT 8.335000 1.180000 8.505000 1.950000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
      RECT 0.000000  3.245000 8.640000 3.415000 ;
      RECT 0.095000  0.085000 0.345000 1.250000 ;
      RECT 0.160000  1.920000 1.360000 2.090000 ;
      RECT 0.160000  2.090000 0.490000 2.980000 ;
      RECT 0.690000  2.260000 0.940000 3.245000 ;
      RECT 0.855000  0.920000 1.105000 0.940000 ;
      RECT 0.855000  0.940000 2.700000 1.190000 ;
      RECT 0.855000  1.190000 1.105000 1.250000 ;
      RECT 1.110000  2.090000 1.360000 2.905000 ;
      RECT 1.110000  2.905000 2.340000 3.075000 ;
      RECT 1.285000  0.085000 1.615000 0.410000 ;
      RECT 1.560000  1.190000 1.810000 2.735000 ;
      RECT 2.010000  2.190000 2.340000 2.905000 ;
      RECT 2.415000  0.085000 2.745000 0.430000 ;
      RECT 2.530000  1.190000 2.700000 1.360000 ;
      RECT 2.530000  1.360000 3.595000 1.680000 ;
      RECT 2.535000  2.190000 2.785000 2.905000 ;
      RECT 2.535000  2.905000 4.665000 3.075000 ;
      RECT 3.515000  2.625000 3.685000 2.905000 ;
      RECT 3.720000  0.085000 4.135000 0.510000 ;
      RECT 4.415000  2.625000 6.655000 2.795000 ;
      RECT 4.415000  2.795000 4.665000 2.905000 ;
      RECT 4.445000  0.350000 4.695000 0.670000 ;
      RECT 4.445000  0.670000 6.655000 0.840000 ;
      RECT 4.855000  2.965000 5.185000 3.245000 ;
      RECT 4.875000  0.085000 5.205000 0.500000 ;
      RECT 5.375000  2.795000 5.705000 2.980000 ;
      RECT 5.385000  0.350000 5.715000 0.670000 ;
      RECT 5.890000  2.965000 6.220000 3.245000 ;
      RECT 5.895000  0.085000 6.225000 0.500000 ;
      RECT 6.405000  0.255000 8.525000 0.425000 ;
      RECT 6.405000  0.425000 6.655000 0.670000 ;
      RECT 6.485000  2.290000 8.535000 2.460000 ;
      RECT 6.485000  2.460000 6.655000 2.625000 ;
      RECT 6.485000  2.795000 6.655000 2.980000 ;
      RECT 6.855000  2.630000 7.105000 3.245000 ;
      RECT 7.305000  2.460000 7.635000 2.980000 ;
      RECT 7.335000  0.425000 7.665000 0.840000 ;
      RECT 7.835000  2.630000 8.005000 3.245000 ;
      RECT 8.195000  0.425000 8.525000 0.840000 ;
      RECT 8.205000  2.460000 8.535000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
  END
END sky130_fd_sc_hs__xor2_4
MACRO sky130_fd_sc_hs__xor3_1
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.960000 1.180000 1.285000 1.750000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.693000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.920000 1.350000 5.250000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.875000 1.180000 7.205000 1.685000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.755000 0.400000 9.005000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.120000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.120000 0.085000 ;
      RECT 0.000000  3.245000 9.120000 3.415000 ;
      RECT 0.085000  0.650000 0.445000 0.660000 ;
      RECT 0.085000  0.660000 1.965000 0.830000 ;
      RECT 0.085000  0.830000 0.445000 1.300000 ;
      RECT 0.085000  1.300000 0.255000 2.260000 ;
      RECT 0.085000  2.260000 0.600000 2.980000 ;
      RECT 0.425000  1.470000 0.750000 1.920000 ;
      RECT 0.425000  1.920000 1.625000 1.940000 ;
      RECT 0.425000  1.940000 1.700000 2.090000 ;
      RECT 0.625000  0.085000 1.195000 0.490000 ;
      RECT 0.770000  2.260000 1.100000 3.245000 ;
      RECT 1.370000  2.090000 1.700000 2.905000 ;
      RECT 1.370000  2.905000 3.895000 3.075000 ;
      RECT 1.455000  1.000000 1.625000 1.920000 ;
      RECT 1.795000  0.830000 1.965000 1.260000 ;
      RECT 1.795000  1.260000 2.760000 1.430000 ;
      RECT 1.930000  1.940000 2.260000 2.565000 ;
      RECT 1.930000  2.565000 3.555000 2.735000 ;
      RECT 2.135000  0.290000 3.215000 0.460000 ;
      RECT 2.135000  0.460000 2.385000 1.090000 ;
      RECT 2.430000  1.430000 2.760000 2.395000 ;
      RECT 2.590000  0.630000 2.850000 1.090000 ;
      RECT 2.590000  1.090000 2.760000 1.260000 ;
      RECT 2.965000  1.875000 3.215000 2.395000 ;
      RECT 3.020000  0.460000 3.215000 1.875000 ;
      RECT 3.385000  0.255000 5.145000 0.425000 ;
      RECT 3.385000  0.425000 3.555000 2.565000 ;
      RECT 3.725000  0.595000 4.805000 0.765000 ;
      RECT 3.725000  0.765000 3.895000 1.435000 ;
      RECT 3.725000  1.435000 4.055000 1.735000 ;
      RECT 3.725000  1.905000 4.395000 2.755000 ;
      RECT 3.725000  2.755000 3.895000 2.905000 ;
      RECT 4.065000  0.935000 4.395000 1.265000 ;
      RECT 4.225000  1.265000 4.395000 1.905000 ;
      RECT 4.580000  0.765000 4.805000 1.130000 ;
      RECT 4.580000  1.130000 4.750000 2.980000 ;
      RECT 4.950000  1.950000 5.200000 3.245000 ;
      RECT 4.975000  0.425000 5.145000 0.850000 ;
      RECT 4.975000  0.850000 6.025000 1.020000 ;
      RECT 5.315000  0.085000 5.565000 0.680000 ;
      RECT 5.405000  1.950000 5.625000 1.990000 ;
      RECT 5.405000  1.990000 5.855000 2.840000 ;
      RECT 5.420000  1.190000 6.365000 1.360000 ;
      RECT 5.420000  1.360000 5.625000 1.950000 ;
      RECT 5.775000  0.255000 7.645000 0.425000 ;
      RECT 5.775000  0.425000 6.025000 0.850000 ;
      RECT 5.805000  1.530000 6.195000 1.820000 ;
      RECT 6.025000  1.820000 6.195000 2.905000 ;
      RECT 6.025000  2.905000 7.605000 3.075000 ;
      RECT 6.195000  0.595000 7.305000 0.765000 ;
      RECT 6.195000  0.765000 6.365000 1.190000 ;
      RECT 6.365000  1.550000 6.705000 2.735000 ;
      RECT 6.535000  0.935000 6.705000 1.550000 ;
      RECT 6.875000  1.855000 7.645000 2.025000 ;
      RECT 6.875000  2.025000 7.205000 2.735000 ;
      RECT 6.885000  0.765000 7.305000 0.925000 ;
      RECT 7.435000  2.195000 7.985000 2.525000 ;
      RECT 7.435000  2.525000 7.605000 2.905000 ;
      RECT 7.475000  0.425000 7.645000 1.855000 ;
      RECT 7.815000  0.400000 8.065000 0.860000 ;
      RECT 7.815000  0.860000 7.985000 2.195000 ;
      RECT 8.225000  1.950000 8.555000 3.245000 ;
      RECT 8.245000  0.085000 8.575000 1.180000 ;
      RECT 8.255000  1.350000 8.585000 1.780000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  1.580000 3.205000 1.750000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  1.580000 5.605000 1.750000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  1.580000 6.565000 1.750000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  1.580000 8.485000 1.750000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
    LAYER met1 ;
      RECT 2.975000 1.550000 3.265000 1.595000 ;
      RECT 2.975000 1.595000 5.665000 1.735000 ;
      RECT 2.975000 1.735000 3.265000 1.780000 ;
      RECT 5.375000 1.550000 5.665000 1.595000 ;
      RECT 5.375000 1.735000 5.665000 1.780000 ;
      RECT 6.335000 1.550000 6.625000 1.595000 ;
      RECT 6.335000 1.595000 8.545000 1.735000 ;
      RECT 6.335000 1.735000 6.625000 1.780000 ;
      RECT 8.255000 1.550000 8.545000 1.595000 ;
      RECT 8.255000 1.735000 8.545000 1.780000 ;
  END
END sky130_fd_sc_hs__xor3_1
MACRO sky130_fd_sc_hs__xor3_2
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.600000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955000 1.180000 1.285000 1.750000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.693000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.920000 1.180000 5.250000 1.550000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.875000 1.180000 7.125000 1.685000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.705000 0.370000 9.035000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.600000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.600000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.600000 0.085000 ;
      RECT 0.000000  3.245000 9.600000 3.415000 ;
      RECT 0.085000  0.650000 0.445000 0.660000 ;
      RECT 0.085000  0.660000 1.965000 0.830000 ;
      RECT 0.085000  0.830000 0.445000 1.275000 ;
      RECT 0.085000  1.275000 0.255000 2.260000 ;
      RECT 0.085000  2.260000 0.595000 2.955000 ;
      RECT 0.425000  1.445000 0.745000 1.920000 ;
      RECT 0.425000  1.920000 1.625000 2.075000 ;
      RECT 0.425000  2.075000 1.640000 2.090000 ;
      RECT 0.625000  0.085000 1.195000 0.490000 ;
      RECT 0.765000  2.260000 1.095000 3.245000 ;
      RECT 1.310000  2.090000 1.640000 2.905000 ;
      RECT 1.310000  2.905000 3.895000 3.075000 ;
      RECT 1.455000  1.000000 1.625000 1.920000 ;
      RECT 1.795000  0.830000 1.965000 1.395000 ;
      RECT 1.795000  1.395000 2.680000 1.565000 ;
      RECT 1.850000  2.075000 2.180000 2.565000 ;
      RECT 1.850000  2.565000 3.555000 2.735000 ;
      RECT 2.135000  0.425000 3.215000 0.595000 ;
      RECT 2.135000  0.595000 2.305000 1.225000 ;
      RECT 2.350000  1.565000 2.680000 2.395000 ;
      RECT 2.510000  0.765000 2.875000 1.225000 ;
      RECT 2.510000  1.225000 2.680000 1.395000 ;
      RECT 2.885000  1.875000 3.215000 2.395000 ;
      RECT 3.045000  0.595000 3.215000 1.875000 ;
      RECT 3.385000  0.255000 5.145000 0.425000 ;
      RECT 3.385000  0.425000 3.555000 2.565000 ;
      RECT 3.725000  0.595000 4.805000 0.765000 ;
      RECT 3.725000  0.765000 3.895000 1.435000 ;
      RECT 3.725000  1.435000 4.055000 1.735000 ;
      RECT 3.725000  1.905000 4.395000 2.755000 ;
      RECT 3.725000  2.755000 3.895000 2.905000 ;
      RECT 4.065000  0.935000 4.395000 1.265000 ;
      RECT 4.225000  1.265000 4.395000 1.905000 ;
      RECT 4.580000  0.765000 4.805000 1.010000 ;
      RECT 4.580000  1.010000 4.750000 2.980000 ;
      RECT 4.950000  1.820000 5.200000 3.245000 ;
      RECT 4.975000  0.425000 5.145000 0.675000 ;
      RECT 4.975000  0.675000 6.025000 0.845000 ;
      RECT 5.315000  0.085000 5.565000 0.505000 ;
      RECT 5.405000  1.920000 5.840000 2.980000 ;
      RECT 5.510000  1.015000 6.365000 1.185000 ;
      RECT 5.510000  1.185000 5.680000 1.920000 ;
      RECT 5.775000  0.255000 7.605000 0.425000 ;
      RECT 5.775000  0.425000 6.025000 0.675000 ;
      RECT 5.850000  1.355000 6.180000 1.685000 ;
      RECT 6.010000  1.685000 6.180000 2.905000 ;
      RECT 6.010000  2.905000 7.450000 3.075000 ;
      RECT 6.195000  0.595000 7.265000 0.765000 ;
      RECT 6.195000  0.765000 6.365000 1.015000 ;
      RECT 6.350000  1.355000 6.705000 1.525000 ;
      RECT 6.350000  1.525000 6.600000 2.700000 ;
      RECT 6.535000  0.935000 6.705000 1.355000 ;
      RECT 6.785000  1.855000 7.465000 2.025000 ;
      RECT 6.785000  2.025000 7.050000 2.690000 ;
      RECT 6.885000  0.765000 7.265000 0.925000 ;
      RECT 7.280000  2.195000 7.805000 2.500000 ;
      RECT 7.280000  2.500000 7.450000 2.905000 ;
      RECT 7.295000  1.095000 7.605000 1.265000 ;
      RECT 7.295000  1.265000 7.465000 1.855000 ;
      RECT 7.435000  0.425000 7.605000 1.095000 ;
      RECT 7.635000  1.435000 8.025000 1.605000 ;
      RECT 7.635000  1.605000 7.805000 2.195000 ;
      RECT 7.775000  0.370000 8.025000 1.435000 ;
      RECT 7.975000  1.820000 8.145000 2.320000 ;
      RECT 7.975000  2.320000 8.530000 3.245000 ;
      RECT 8.195000  1.320000 8.525000 1.650000 ;
      RECT 8.205000  0.085000 8.535000 1.150000 ;
      RECT 8.315000  1.650000 8.525000 2.150000 ;
      RECT 9.215000  0.085000 9.465000 1.150000 ;
      RECT 9.235000  1.820000 9.485000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  1.950000 3.205000 2.120000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  1.950000 5.605000 2.120000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  1.950000 6.565000 2.120000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  1.950000 8.485000 2.120000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
    LAYER met1 ;
      RECT 2.975000 1.920000 3.265000 1.965000 ;
      RECT 2.975000 1.965000 5.665000 2.105000 ;
      RECT 2.975000 2.105000 3.265000 2.150000 ;
      RECT 5.375000 1.920000 5.665000 1.965000 ;
      RECT 5.375000 2.105000 5.665000 2.150000 ;
      RECT 6.335000 1.920000 6.625000 1.965000 ;
      RECT 6.335000 1.965000 8.545000 2.105000 ;
      RECT 6.335000 2.105000 6.625000 2.150000 ;
      RECT 8.255000 1.920000 8.545000 1.965000 ;
      RECT 8.255000 2.105000 8.545000 2.150000 ;
  END
END sky130_fd_sc_hs__xor3_2
MACRO sky130_fd_sc_hs__xor3_4
  CLASS CORE ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.56000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.910000 1.180000 1.285000 1.670000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.693000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.910000 1.180000 5.240000 1.550000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.810000 1.450000 7.070000 1.780000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.685000 1.820000 9.125000 2.980000 ;
        RECT 8.830000 0.350000 9.160000 1.085000 ;
        RECT 8.955000 1.085000 9.160000 1.300000 ;
        RECT 8.955000 1.300000 9.940000 1.470000 ;
        RECT 8.955000 1.470000 9.125000 1.820000 ;
        RECT 9.665000 1.470000 9.940000 1.550000 ;
        RECT 9.665000 1.550000 9.995000 2.980000 ;
        RECT 9.690000 0.350000 9.940000 1.300000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.560000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.560000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 10.560000 0.085000 ;
      RECT  0.000000  3.245000 10.560000 3.415000 ;
      RECT  0.085000  0.570000  0.445000 0.580000 ;
      RECT  0.085000  0.580000  1.965000 0.750000 ;
      RECT  0.085000  0.750000  0.445000 1.250000 ;
      RECT  0.085000  1.250000  0.255000 2.180000 ;
      RECT  0.085000  2.180000  0.365000 2.980000 ;
      RECT  0.425000  1.470000  0.700000 1.840000 ;
      RECT  0.425000  1.840000  1.625000 2.010000 ;
      RECT  0.565000  2.180000  0.895000 3.245000 ;
      RECT  0.625000  0.085000  1.035000 0.410000 ;
      RECT  1.065000  2.010000  1.395000 2.905000 ;
      RECT  1.065000  2.905000  3.825000 3.075000 ;
      RECT  1.455000  0.920000  1.625000 1.840000 ;
      RECT  1.600000  2.180000  1.930000 2.565000 ;
      RECT  1.600000  2.565000  3.485000 2.735000 ;
      RECT  1.795000  0.750000  1.965000 1.420000 ;
      RECT  1.795000  1.420000  2.805000 1.590000 ;
      RECT  2.135000  0.450000  3.145000 0.620000 ;
      RECT  2.135000  0.620000  2.385000 1.250000 ;
      RECT  2.135000  1.590000  2.385000 2.395000 ;
      RECT  2.555000  0.790000  2.805000 1.420000 ;
      RECT  2.555000  1.875000  3.145000 2.395000 ;
      RECT  2.975000  0.620000  3.145000 1.875000 ;
      RECT  3.315000  0.255000  5.080000 0.425000 ;
      RECT  3.315000  0.425000  3.485000 2.565000 ;
      RECT  3.655000  0.595000  4.740000 0.765000 ;
      RECT  3.655000  0.765000  3.825000 1.435000 ;
      RECT  3.655000  1.435000  3.985000 1.735000 ;
      RECT  3.655000  1.905000  4.325000 2.755000 ;
      RECT  3.655000  2.755000  3.825000 2.905000 ;
      RECT  3.995000  0.935000  4.325000 1.265000 ;
      RECT  4.155000  1.265000  4.325000 1.905000 ;
      RECT  4.535000  0.765000  4.740000 1.130000 ;
      RECT  4.535000  1.130000  4.705000 2.980000 ;
      RECT  4.905000  1.820000  5.235000 3.245000 ;
      RECT  4.910000  0.425000  5.080000 0.780000 ;
      RECT  4.910000  0.780000  5.960000 0.950000 ;
      RECT  5.250000  0.085000  5.500000 0.610000 ;
      RECT  5.405000  1.920000  5.795000 2.800000 ;
      RECT  5.435000  1.120000  6.300000 1.290000 ;
      RECT  5.435000  1.290000  5.605000 1.920000 ;
      RECT  5.710000  0.255000  7.410000 0.425000 ;
      RECT  5.710000  0.425000  5.960000 0.780000 ;
      RECT  5.775000  1.460000  6.135000 1.750000 ;
      RECT  5.965000  1.750000  6.135000 2.905000 ;
      RECT  5.965000  2.905000  7.500000 3.075000 ;
      RECT  6.130000  0.595000  7.070000 0.765000 ;
      RECT  6.130000  0.765000  6.300000 1.120000 ;
      RECT  6.305000  1.920000  6.640000 2.735000 ;
      RECT  6.470000  0.935000  6.640000 1.920000 ;
      RECT  6.820000  0.765000  7.070000 1.275000 ;
      RECT  6.835000  1.950000  7.410000 2.120000 ;
      RECT  6.835000  2.120000  7.085000 2.735000 ;
      RECT  7.240000  0.425000  7.410000 1.950000 ;
      RECT  7.330000  2.290000  7.750000 2.710000 ;
      RECT  7.330000  2.710000  7.500000 2.905000 ;
      RECT  7.580000  0.415000  8.150000 0.745000 ;
      RECT  7.580000  0.745000  7.750000 2.290000 ;
      RECT  7.920000  1.255000  8.785000 1.585000 ;
      RECT  7.945000  1.820000  8.115000 2.330000 ;
      RECT  7.945000  2.330000  8.500000 3.245000 ;
      RECT  8.285000  1.585000  8.515000 2.150000 ;
      RECT  8.330000  0.085000  8.660000 1.085000 ;
      RECT  9.295000  1.820000  9.465000 3.245000 ;
      RECT  9.340000  0.085000  9.510000 1.130000 ;
      RECT 10.120000  0.085000 10.450000 1.130000 ;
      RECT 10.195000  1.820000 10.445000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  1.950000  2.725000 2.120000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  1.950000  5.605000 2.120000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  1.950000  6.565000 2.120000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  1.950000  8.485000 2.120000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
    LAYER met1 ;
      RECT 2.495000 1.920000 2.785000 1.965000 ;
      RECT 2.495000 1.965000 5.665000 2.105000 ;
      RECT 2.495000 2.105000 2.785000 2.150000 ;
      RECT 5.375000 1.920000 5.665000 1.965000 ;
      RECT 5.375000 2.105000 5.665000 2.150000 ;
      RECT 6.335000 1.920000 6.625000 1.965000 ;
      RECT 6.335000 1.965000 8.545000 2.105000 ;
      RECT 6.335000 2.105000 6.625000 2.150000 ;
      RECT 8.255000 1.920000 8.545000 1.965000 ;
      RECT 8.255000 2.105000 8.545000 2.150000 ;
  END
END sky130_fd_sc_hs__xor3_4
END LIBRARY
