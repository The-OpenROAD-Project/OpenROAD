../sky130_temp_sensor/HEADER.lef