VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
	DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

USEMINSPACING OBS OFF ;

PROPERTYDEFINITIONS
LAYER LEF58_TYPE STRING ;
LAYER LEF58_SPACING STRING ;
LAYER LEF58_WIDTH STRING ;
LAYER LEF58_AREA STRING ;
LAYER LEF58_MINENCLOSEDAREA STRING ;
END PROPERTYDEFINITIONS

LAYER metal1
	TYPE ROUTING ;
	DIRECTION HORIZONTAL ;
	PITCH 1 ;
	WIDTH 1 ;
END metal1

MACRO MACRO_CELL
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 10 BY 10 ;
  SYMMETRY X Y R90 ;
  PIN VDD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0 5 0 5 ;
    END
  END VDD
  PIN GND
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0 5 0 5 ;
    END
  END GND
  PIN IN_REG[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0 5 0 5 ;
    END
  END IN_REG[0]
  PIN IN_REG[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0 5 0 5 ;
    END
  END IN_REG[1]
  PIN OUT_REG[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0 5 0 5 ;
    END
  END OUT_REG[0]
  PIN OUT_REG[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0 5 0 5 ;
    END
  END OUT_REG[1]
END MACRO_CELL

END LIBRARY
