VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.1 ;

LAYER M1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 ;
  WIDTH 0.1 ;
  OFFSET 0.1 ;
  AREA 0.042 ;
END M1

LAYER M2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 ;
  WIDTH 0.1 ;
  OFFSET 0.1 ;
  AREA 0.052 ;
END M2

LAYER nwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE NWELL ;" ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE PWELL ;" ;
END pwell

SITE site1
  CLASS CORE ;
  SIZE 50 BY 20 ;
END site1

MACRO snl_bufx1
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
END snl_bufx1

MACRO snl_bufx2
 SIZE 50 BY 20 ;
 PIN Z DIRECTION OUTPUT ; END Z
 PIN A DIRECTION INPUT ; END A
 PIN VDD DIRECTION INOUT ; USE POWER ; END VDD
 PIN VSS DIRECTION INOUT ; USE GROUND ; END VSS
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.090 0.085 0.345 0.885 ;
        RECT 1.015 0.085 1.345 0.465 ;
        RECT 3.220 0.085 3.550 0.485 ;
        RECT 0.000 -0.085 4.140 0.085 ;
    END
  END VGND
  # power/ground PINs
  PIN VNB
    DIRECTION INPUT ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.135 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INPUT ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.090 1.495 0.345 2.635 ;
        RECT 1.160 1.835 1.380 2.635 ;
        RECT 2.125 2.255 2.455 2.635 ;
    END
  END VPWR
END snl_bufx2

END LIBRARY
