# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_io__top_ground_hvc_wpad
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 200 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    ANTENNAPARTIALMETALSIDEAREA  111.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 1.270000 56.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 53.125000 75.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    ANTENNAPARTIALMETALSIDEAREA  111.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 1.270000 51.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 48.365000 75.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN G_PAD
    ANTENNAPARTIALMETALSIDEAREA  284.1730 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 36.645000 139.325000 37.970000 145.935000 ;
    END
  END G_PAD
  PIN DRN_HVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 15.620000 185.295000 74.290000 190.015000 ;
        RECT 16.805000  47.455000 74.290000  54.765000 ;
        RECT 16.805000 139.455000 74.290000 146.710000 ;
        RECT 16.805000 162.455000 74.290000 171.155000 ;
        RECT 16.875000 146.710000 74.290000 146.780000 ;
        RECT 16.945000 146.780000 74.290000 146.850000 ;
        RECT 17.015000 146.850000 74.290000 146.920000 ;
        RECT 17.085000 146.920000 74.290000 146.990000 ;
        RECT 17.155000 146.990000 74.290000 147.060000 ;
        RECT 17.225000 147.060000 74.290000 147.130000 ;
        RECT 17.295000 147.130000 74.290000 147.200000 ;
        RECT 17.365000 147.200000 74.290000 147.270000 ;
        RECT 17.435000 147.270000 74.290000 147.340000 ;
        RECT 17.505000 147.340000 74.290000 147.410000 ;
        RECT 17.530000  54.765000 74.290000  54.835000 ;
        RECT 17.575000 147.410000 74.290000 147.480000 ;
        RECT 17.600000  54.835000 74.290000  54.905000 ;
        RECT 17.645000 147.480000 74.290000 147.550000 ;
        RECT 17.670000  54.905000 74.290000  54.975000 ;
        RECT 17.715000 147.550000 74.290000 147.620000 ;
        RECT 17.740000  54.975000 74.290000  55.045000 ;
        RECT 17.785000 147.620000 74.290000 147.690000 ;
        RECT 17.810000  55.045000 74.290000  55.115000 ;
        RECT 17.855000 147.690000 74.290000 147.760000 ;
        RECT 17.880000  55.115000 74.290000  55.185000 ;
        RECT 17.925000 147.760000 74.290000 147.830000 ;
        RECT 17.950000  55.185000 74.290000  55.255000 ;
        RECT 17.995000 147.830000 74.290000 147.900000 ;
        RECT 18.020000  55.255000 74.290000  55.325000 ;
        RECT 18.065000 147.900000 74.290000 147.970000 ;
        RECT 18.090000  55.325000 74.290000  55.395000 ;
        RECT 18.135000 147.970000 74.290000 148.040000 ;
        RECT 18.160000  55.395000 74.290000  55.465000 ;
        RECT 18.205000 148.040000 74.290000 148.110000 ;
        RECT 18.230000  55.465000 74.290000  55.535000 ;
        RECT 18.250000 148.110000 74.290000 148.155000 ;
        RECT 18.300000  55.535000 74.290000  55.605000 ;
        RECT 18.370000  55.605000 74.290000  55.675000 ;
        RECT 18.410000  74.155000 74.290000  74.415000 ;
        RECT 18.440000  55.675000 74.290000  55.745000 ;
        RECT 18.510000  55.745000 74.290000  55.815000 ;
        RECT 18.580000  55.815000 74.290000  55.885000 ;
        RECT 18.650000  55.885000 74.290000  55.955000 ;
        RECT 18.720000  55.955000 74.290000  56.025000 ;
        RECT 18.790000  56.025000 74.290000  56.095000 ;
        RECT 18.850000  56.095000 74.290000  56.155000 ;
        RECT 23.690000  74.415000 74.290000  74.485000 ;
        RECT 23.700000  74.105000 74.290000  74.155000 ;
        RECT 23.760000  74.485000 74.290000  74.555000 ;
        RECT 23.770000  74.035000 74.290000  74.105000 ;
        RECT 23.830000  74.555000 74.290000  74.625000 ;
        RECT 23.840000  73.965000 74.290000  74.035000 ;
        RECT 23.900000  74.625000 74.290000  74.695000 ;
        RECT 23.910000  73.895000 74.290000  73.965000 ;
        RECT 23.970000  74.695000 74.290000  74.765000 ;
        RECT 23.980000  73.825000 74.290000  73.895000 ;
        RECT 24.040000  74.765000 74.290000  74.835000 ;
        RECT 24.050000  73.755000 74.290000  73.825000 ;
        RECT 24.110000  74.835000 74.290000  74.905000 ;
        RECT 24.120000  73.685000 74.290000  73.755000 ;
        RECT 24.180000  74.905000 74.290000  74.975000 ;
        RECT 24.190000  73.615000 74.290000  73.685000 ;
        RECT 24.250000  74.975000 74.290000  75.045000 ;
        RECT 24.260000  73.545000 74.290000  73.615000 ;
        RECT 24.320000  75.045000 74.290000  75.115000 ;
        RECT 24.330000  73.475000 74.290000  73.545000 ;
        RECT 24.390000  75.115000 74.290000  75.185000 ;
        RECT 24.400000  73.405000 74.290000  73.475000 ;
        RECT 24.460000  75.185000 74.290000  75.255000 ;
        RECT 24.470000  73.335000 74.290000  73.405000 ;
        RECT 24.530000  75.255000 74.290000  75.325000 ;
        RECT 24.540000  73.265000 74.290000  73.335000 ;
        RECT 24.600000  75.325000 74.290000  75.395000 ;
        RECT 24.610000  73.195000 74.290000  73.265000 ;
        RECT 24.670000  75.395000 74.290000  75.465000 ;
        RECT 24.680000  73.125000 74.290000  73.195000 ;
        RECT 24.740000  75.465000 74.290000  75.535000 ;
        RECT 24.750000  73.055000 74.290000  73.125000 ;
        RECT 24.810000  75.535000 74.290000  75.605000 ;
        RECT 24.820000  70.455000 74.290000  72.985000 ;
        RECT 24.820000  72.985000 74.290000  73.055000 ;
        RECT 24.820000  75.605000 74.290000  75.615000 ;
        RECT 24.820000  75.615000 74.290000  79.155000 ;
        RECT 24.820000  93.455000 74.290000 102.155000 ;
        RECT 24.820000 116.455000 74.290000 125.155000 ;
        RECT 37.890000  12.295000 74.290000  25.660000 ;
        RECT 46.750000  12.265000 74.290000  12.295000 ;
        RECT 46.820000  12.195000 74.290000  12.265000 ;
        RECT 46.890000  12.125000 74.290000  12.195000 ;
        RECT 46.960000  12.055000 74.290000  12.125000 ;
        RECT 47.030000  11.985000 74.290000  12.055000 ;
        RECT 47.100000  11.915000 74.290000  11.985000 ;
        RECT 47.170000  11.845000 74.290000  11.915000 ;
        RECT 47.240000  11.775000 74.290000  11.845000 ;
        RECT 47.310000  11.705000 74.290000  11.775000 ;
        RECT 47.380000  11.635000 74.290000  11.705000 ;
        RECT 47.450000  11.565000 74.290000  11.635000 ;
        RECT 47.520000  11.495000 74.290000  11.565000 ;
        RECT 47.590000  11.425000 74.290000  11.495000 ;
        RECT 47.660000  11.355000 74.290000  11.425000 ;
        RECT 47.730000  11.285000 74.290000  11.355000 ;
        RECT 47.800000  11.215000 74.290000  11.285000 ;
        RECT 47.870000  11.145000 74.290000  11.215000 ;
        RECT 47.940000  11.075000 74.290000  11.145000 ;
        RECT 48.010000  11.005000 74.290000  11.075000 ;
        RECT 48.080000  10.935000 74.290000  11.005000 ;
        RECT 48.150000  10.865000 74.290000  10.935000 ;
        RECT 48.220000  10.795000 74.290000  10.865000 ;
        RECT 48.290000  10.725000 74.290000  10.795000 ;
        RECT 48.360000  10.655000 74.290000  10.725000 ;
        RECT 48.430000  10.585000 74.290000  10.655000 ;
        RECT 48.500000  10.515000 74.290000  10.585000 ;
        RECT 48.570000  10.445000 74.290000  10.515000 ;
        RECT 48.640000  10.375000 74.290000  10.445000 ;
        RECT 48.710000  10.305000 74.290000  10.375000 ;
        RECT 48.780000  10.235000 74.290000  10.305000 ;
        RECT 48.850000  10.165000 74.290000  10.235000 ;
        RECT 48.920000  10.095000 74.290000  10.165000 ;
        RECT 48.990000  10.025000 74.290000  10.095000 ;
        RECT 49.060000   9.955000 74.290000  10.025000 ;
        RECT 49.130000   9.885000 74.290000   9.955000 ;
        RECT 49.200000   9.815000 74.290000   9.885000 ;
        RECT 49.270000   9.745000 74.290000   9.815000 ;
        RECT 49.340000   9.675000 74.290000   9.745000 ;
        RECT 49.410000   9.605000 74.290000   9.675000 ;
        RECT 49.480000   9.535000 74.290000   9.605000 ;
        RECT 49.550000   9.465000 74.290000   9.535000 ;
        RECT 49.620000   9.395000 74.290000   9.465000 ;
        RECT 49.690000   9.325000 74.290000   9.395000 ;
        RECT 49.760000   9.255000 74.290000   9.325000 ;
        RECT 49.830000   9.185000 74.290000   9.255000 ;
        RECT 49.900000   9.115000 74.290000   9.185000 ;
        RECT 49.970000   9.045000 74.290000   9.115000 ;
        RECT 50.040000   8.975000 74.290000   9.045000 ;
        RECT 50.110000   8.905000 74.290000   8.975000 ;
        RECT 50.180000   8.835000 74.290000   8.905000 ;
        RECT 50.250000   8.765000 74.290000   8.835000 ;
        RECT 50.320000   8.695000 74.290000   8.765000 ;
        RECT 50.390000   0.000000 74.290000   8.625000 ;
        RECT 50.390000   8.625000 74.290000   8.695000 ;
        RECT 55.885000  25.660000 74.290000  25.730000 ;
        RECT 55.955000  25.730000 74.290000  25.800000 ;
        RECT 56.025000  25.800000 74.290000  25.870000 ;
        RECT 56.095000  25.870000 74.290000  25.940000 ;
        RECT 56.165000  25.940000 74.290000  26.010000 ;
        RECT 56.235000  26.010000 74.290000  26.080000 ;
        RECT 56.305000  26.080000 74.290000  26.150000 ;
        RECT 56.375000  26.150000 74.290000  26.220000 ;
        RECT 56.445000  26.220000 74.290000  26.290000 ;
        RECT 56.515000  26.290000 74.290000  26.360000 ;
        RECT 56.585000  26.360000 74.290000  26.430000 ;
        RECT 56.655000  26.430000 74.290000  26.500000 ;
        RECT 56.725000  26.500000 74.290000  26.570000 ;
        RECT 56.795000  26.570000 74.290000  26.640000 ;
        RECT 56.865000  26.640000 74.290000  26.710000 ;
        RECT 56.935000  26.710000 74.290000  26.780000 ;
        RECT 57.005000  26.780000 74.290000  26.850000 ;
        RECT 57.075000  26.850000 74.290000  26.920000 ;
        RECT 57.145000  26.920000 74.290000  26.990000 ;
        RECT 57.215000  26.990000 74.290000  27.060000 ;
        RECT 57.285000  27.060000 74.290000  27.130000 ;
        RECT 57.355000  27.130000 74.290000  27.200000 ;
        RECT 57.425000  27.200000 74.290000  27.270000 ;
        RECT 57.495000  27.270000 74.290000  27.340000 ;
        RECT 57.540000  47.390000 74.290000  47.455000 ;
        RECT 57.540000  70.420000 74.290000  70.455000 ;
        RECT 57.540000 116.390000 74.290000 116.455000 ;
        RECT 57.540000 139.425000 74.290000 139.455000 ;
        RECT 57.540000 162.440000 74.290000 162.455000 ;
        RECT 57.555000 148.155000 74.290000 148.225000 ;
        RECT 57.565000  27.340000 74.290000  27.410000 ;
        RECT 57.595000  56.155000 74.290000  56.225000 ;
        RECT 57.610000  47.320000 74.290000  47.390000 ;
        RECT 57.610000  70.350000 74.290000  70.420000 ;
        RECT 57.610000  93.410000 74.290000  93.455000 ;
        RECT 57.610000 116.320000 74.290000 116.390000 ;
        RECT 57.610000 139.355000 74.290000 139.425000 ;
        RECT 57.610000 162.370000 74.290000 162.440000 ;
        RECT 57.625000  79.155000 74.290000  79.225000 ;
        RECT 57.625000 102.155000 74.290000 102.225000 ;
        RECT 57.625000 125.155000 74.290000 125.225000 ;
        RECT 57.625000 148.225000 74.290000 148.295000 ;
        RECT 57.635000  27.410000 74.290000  27.480000 ;
        RECT 57.635000 171.155000 74.290000 171.225000 ;
        RECT 57.665000  56.225000 74.290000  56.295000 ;
        RECT 57.680000  47.250000 74.290000  47.320000 ;
        RECT 57.680000  70.280000 74.290000  70.350000 ;
        RECT 57.680000  93.340000 74.290000  93.410000 ;
        RECT 57.680000 116.250000 74.290000 116.320000 ;
        RECT 57.680000 139.285000 74.290000 139.355000 ;
        RECT 57.680000 162.300000 74.290000 162.370000 ;
        RECT 57.695000  79.225000 74.290000  79.295000 ;
        RECT 57.695000 102.225000 74.290000 102.295000 ;
        RECT 57.695000 125.225000 74.290000 125.295000 ;
        RECT 57.695000 148.295000 74.290000 148.365000 ;
        RECT 57.705000  27.480000 74.290000  27.550000 ;
        RECT 57.705000 171.225000 74.290000 171.295000 ;
        RECT 57.735000  56.295000 74.290000  56.365000 ;
        RECT 57.750000  47.180000 74.290000  47.250000 ;
        RECT 57.750000  70.210000 74.290000  70.280000 ;
        RECT 57.750000  93.270000 74.290000  93.340000 ;
        RECT 57.750000 116.180000 74.290000 116.250000 ;
        RECT 57.750000 139.215000 74.290000 139.285000 ;
        RECT 57.750000 162.230000 74.290000 162.300000 ;
        RECT 57.765000  79.295000 74.290000  79.365000 ;
        RECT 57.765000 102.295000 74.290000 102.365000 ;
        RECT 57.765000 125.295000 74.290000 125.365000 ;
        RECT 57.765000 148.365000 74.290000 148.435000 ;
        RECT 57.775000  27.550000 74.290000  27.620000 ;
        RECT 57.775000 171.295000 74.290000 171.365000 ;
        RECT 57.805000  56.365000 74.290000  56.435000 ;
        RECT 57.820000  47.110000 74.290000  47.180000 ;
        RECT 57.820000  70.140000 74.290000  70.210000 ;
        RECT 57.820000  93.200000 74.290000  93.270000 ;
        RECT 57.820000 116.110000 74.290000 116.180000 ;
        RECT 57.820000 139.145000 74.290000 139.215000 ;
        RECT 57.820000 162.160000 74.290000 162.230000 ;
        RECT 57.835000  79.365000 74.290000  79.435000 ;
        RECT 57.835000 102.365000 74.290000 102.435000 ;
        RECT 57.835000 125.365000 74.290000 125.435000 ;
        RECT 57.835000 148.435000 74.290000 148.505000 ;
        RECT 57.845000  27.620000 74.290000  27.690000 ;
        RECT 57.845000 171.365000 74.290000 171.435000 ;
        RECT 57.875000  56.435000 74.290000  56.505000 ;
        RECT 57.890000  47.040000 74.290000  47.110000 ;
        RECT 57.890000  70.070000 74.290000  70.140000 ;
        RECT 57.890000  93.130000 74.290000  93.200000 ;
        RECT 57.890000 116.040000 74.290000 116.110000 ;
        RECT 57.890000 139.075000 74.290000 139.145000 ;
        RECT 57.890000 162.090000 74.290000 162.160000 ;
        RECT 57.905000  79.435000 74.290000  79.505000 ;
        RECT 57.905000 102.435000 74.290000 102.505000 ;
        RECT 57.905000 125.435000 74.290000 125.505000 ;
        RECT 57.905000 148.505000 74.290000 148.575000 ;
        RECT 57.915000  27.690000 74.290000  27.760000 ;
        RECT 57.915000 171.435000 74.290000 171.505000 ;
        RECT 57.945000  56.505000 74.290000  56.575000 ;
        RECT 57.960000  46.970000 74.290000  47.040000 ;
        RECT 57.960000  70.000000 74.290000  70.070000 ;
        RECT 57.960000  93.060000 74.290000  93.130000 ;
        RECT 57.960000 115.970000 74.290000 116.040000 ;
        RECT 57.960000 139.005000 74.290000 139.075000 ;
        RECT 57.960000 162.020000 74.290000 162.090000 ;
        RECT 57.975000  79.505000 74.290000  79.575000 ;
        RECT 57.975000 102.505000 74.290000 102.575000 ;
        RECT 57.975000 125.505000 74.290000 125.575000 ;
        RECT 57.975000 148.575000 74.290000 148.645000 ;
        RECT 57.985000  27.760000 74.290000  27.830000 ;
        RECT 57.985000 171.505000 74.290000 171.575000 ;
        RECT 58.015000  56.575000 74.290000  56.645000 ;
        RECT 58.030000  46.900000 74.290000  46.970000 ;
        RECT 58.030000  69.930000 74.290000  70.000000 ;
        RECT 58.030000  92.990000 74.290000  93.060000 ;
        RECT 58.030000 115.900000 74.290000 115.970000 ;
        RECT 58.030000 138.935000 74.290000 139.005000 ;
        RECT 58.030000 161.950000 74.290000 162.020000 ;
        RECT 58.045000  79.575000 74.290000  79.645000 ;
        RECT 58.045000 102.575000 74.290000 102.645000 ;
        RECT 58.045000 125.575000 74.290000 125.645000 ;
        RECT 58.045000 148.645000 74.290000 148.715000 ;
        RECT 58.055000  27.830000 74.290000  27.900000 ;
        RECT 58.055000 171.575000 74.290000 171.645000 ;
        RECT 58.085000  56.645000 74.290000  56.715000 ;
        RECT 58.100000  46.830000 74.290000  46.900000 ;
        RECT 58.100000  69.860000 74.290000  69.930000 ;
        RECT 58.100000  92.920000 74.290000  92.990000 ;
        RECT 58.100000 115.830000 74.290000 115.900000 ;
        RECT 58.100000 138.865000 74.290000 138.935000 ;
        RECT 58.100000 161.880000 74.290000 161.950000 ;
        RECT 58.115000  79.645000 74.290000  79.715000 ;
        RECT 58.115000 102.645000 74.290000 102.715000 ;
        RECT 58.115000 125.645000 74.290000 125.715000 ;
        RECT 58.115000 148.715000 74.290000 148.785000 ;
        RECT 58.125000  27.900000 74.290000  27.970000 ;
        RECT 58.125000 171.645000 74.290000 171.715000 ;
        RECT 58.155000  56.715000 74.290000  56.785000 ;
        RECT 58.170000  46.760000 74.290000  46.830000 ;
        RECT 58.170000  69.790000 74.290000  69.860000 ;
        RECT 58.170000  92.850000 74.290000  92.920000 ;
        RECT 58.170000 115.760000 74.290000 115.830000 ;
        RECT 58.170000 138.795000 74.290000 138.865000 ;
        RECT 58.170000 161.810000 74.290000 161.880000 ;
        RECT 58.185000  79.715000 74.290000  79.785000 ;
        RECT 58.185000 102.715000 74.290000 102.785000 ;
        RECT 58.185000 125.715000 74.290000 125.785000 ;
        RECT 58.185000 148.785000 74.290000 148.855000 ;
        RECT 58.195000  27.970000 74.290000  28.040000 ;
        RECT 58.195000 171.715000 74.290000 171.785000 ;
        RECT 58.225000  56.785000 74.290000  56.855000 ;
        RECT 58.240000  46.690000 74.290000  46.760000 ;
        RECT 58.240000  69.720000 74.290000  69.790000 ;
        RECT 58.240000  92.780000 74.290000  92.850000 ;
        RECT 58.240000 115.690000 74.290000 115.760000 ;
        RECT 58.240000 138.725000 74.290000 138.795000 ;
        RECT 58.240000 161.740000 74.290000 161.810000 ;
        RECT 58.255000  79.785000 74.290000  79.855000 ;
        RECT 58.255000 102.785000 74.290000 102.855000 ;
        RECT 58.255000 125.785000 74.290000 125.855000 ;
        RECT 58.255000 148.855000 74.290000 148.925000 ;
        RECT 58.265000  28.040000 74.290000  28.110000 ;
        RECT 58.265000 171.785000 74.290000 171.855000 ;
        RECT 58.295000  56.855000 74.290000  56.925000 ;
        RECT 58.310000  46.620000 74.290000  46.690000 ;
        RECT 58.310000  69.650000 74.290000  69.720000 ;
        RECT 58.310000  92.710000 74.290000  92.780000 ;
        RECT 58.310000 115.620000 74.290000 115.690000 ;
        RECT 58.310000 138.655000 74.290000 138.725000 ;
        RECT 58.310000 161.670000 74.290000 161.740000 ;
        RECT 58.325000  79.855000 74.290000  79.925000 ;
        RECT 58.325000 102.855000 74.290000 102.925000 ;
        RECT 58.325000 125.855000 74.290000 125.925000 ;
        RECT 58.325000 148.925000 74.290000 148.995000 ;
        RECT 58.335000  28.110000 74.290000  28.180000 ;
        RECT 58.335000 171.855000 74.290000 171.925000 ;
        RECT 58.365000  56.925000 74.290000  56.995000 ;
        RECT 58.380000  46.550000 74.290000  46.620000 ;
        RECT 58.380000  69.580000 74.290000  69.650000 ;
        RECT 58.380000  92.640000 74.290000  92.710000 ;
        RECT 58.380000 115.550000 74.290000 115.620000 ;
        RECT 58.380000 138.585000 74.290000 138.655000 ;
        RECT 58.380000 161.600000 74.290000 161.670000 ;
        RECT 58.395000  79.925000 74.290000  79.995000 ;
        RECT 58.395000 102.925000 74.290000 102.995000 ;
        RECT 58.395000 125.925000 74.290000 125.995000 ;
        RECT 58.395000 148.995000 74.290000 149.065000 ;
        RECT 58.405000  28.180000 74.290000  28.250000 ;
        RECT 58.405000 171.925000 74.290000 171.995000 ;
        RECT 58.435000  56.995000 74.290000  57.065000 ;
        RECT 58.450000  46.480000 74.290000  46.550000 ;
        RECT 58.450000  69.510000 74.290000  69.580000 ;
        RECT 58.450000  92.570000 74.290000  92.640000 ;
        RECT 58.450000 115.480000 74.290000 115.550000 ;
        RECT 58.450000 138.515000 74.290000 138.585000 ;
        RECT 58.450000 161.530000 74.290000 161.600000 ;
        RECT 58.465000  79.995000 74.290000  80.065000 ;
        RECT 58.465000 102.995000 74.290000 103.065000 ;
        RECT 58.465000 125.995000 74.290000 126.065000 ;
        RECT 58.465000 149.065000 74.290000 149.135000 ;
        RECT 58.475000  28.250000 74.290000  28.320000 ;
        RECT 58.475000 171.995000 74.290000 172.065000 ;
        RECT 58.505000  57.065000 74.290000  57.135000 ;
        RECT 58.520000  46.410000 74.290000  46.480000 ;
        RECT 58.520000  69.440000 74.290000  69.510000 ;
        RECT 58.520000  92.500000 74.290000  92.570000 ;
        RECT 58.520000 115.410000 74.290000 115.480000 ;
        RECT 58.520000 138.445000 74.290000 138.515000 ;
        RECT 58.520000 161.460000 74.290000 161.530000 ;
        RECT 58.535000  80.065000 74.290000  80.135000 ;
        RECT 58.535000 103.065000 74.290000 103.135000 ;
        RECT 58.535000 126.065000 74.290000 126.135000 ;
        RECT 58.535000 149.135000 74.290000 149.205000 ;
        RECT 58.545000  28.320000 74.290000  28.390000 ;
        RECT 58.545000 172.065000 74.290000 172.135000 ;
        RECT 58.575000  57.135000 74.290000  57.205000 ;
        RECT 58.590000  46.340000 74.290000  46.410000 ;
        RECT 58.590000  69.370000 74.290000  69.440000 ;
        RECT 58.590000  92.430000 74.290000  92.500000 ;
        RECT 58.590000 115.340000 74.290000 115.410000 ;
        RECT 58.590000 138.375000 74.290000 138.445000 ;
        RECT 58.590000 161.390000 74.290000 161.460000 ;
        RECT 58.605000  80.135000 74.290000  80.205000 ;
        RECT 58.605000 103.135000 74.290000 103.205000 ;
        RECT 58.605000 126.135000 74.290000 126.205000 ;
        RECT 58.605000 149.205000 74.290000 149.275000 ;
        RECT 58.615000  28.390000 74.290000  28.460000 ;
        RECT 58.615000 172.135000 74.290000 172.205000 ;
        RECT 58.645000  57.205000 74.290000  57.275000 ;
        RECT 58.660000  46.270000 74.290000  46.340000 ;
        RECT 58.660000  69.300000 74.290000  69.370000 ;
        RECT 58.660000  92.360000 74.290000  92.430000 ;
        RECT 58.660000 115.270000 74.290000 115.340000 ;
        RECT 58.660000 138.305000 74.290000 138.375000 ;
        RECT 58.660000 161.320000 74.290000 161.390000 ;
        RECT 58.675000  80.205000 74.290000  80.275000 ;
        RECT 58.675000 103.205000 74.290000 103.275000 ;
        RECT 58.675000 126.205000 74.290000 126.275000 ;
        RECT 58.675000 149.275000 74.290000 149.345000 ;
        RECT 58.685000  28.460000 74.290000  28.530000 ;
        RECT 58.685000 172.205000 74.290000 172.275000 ;
        RECT 58.715000  57.275000 74.290000  57.345000 ;
        RECT 58.730000  46.200000 74.290000  46.270000 ;
        RECT 58.730000  69.230000 74.290000  69.300000 ;
        RECT 58.730000  92.290000 74.290000  92.360000 ;
        RECT 58.730000 115.200000 74.290000 115.270000 ;
        RECT 58.730000 138.235000 74.290000 138.305000 ;
        RECT 58.730000 161.250000 74.290000 161.320000 ;
        RECT 58.730000 185.260000 74.290000 185.295000 ;
        RECT 58.745000  80.275000 74.290000  80.345000 ;
        RECT 58.745000 103.275000 74.290000 103.345000 ;
        RECT 58.745000 126.275000 74.290000 126.345000 ;
        RECT 58.745000 149.345000 74.290000 149.415000 ;
        RECT 58.755000  28.530000 74.290000  28.600000 ;
        RECT 58.755000 172.275000 74.290000 172.345000 ;
        RECT 58.785000  57.345000 74.290000  57.415000 ;
        RECT 58.800000  46.130000 74.290000  46.200000 ;
        RECT 58.800000  69.160000 74.290000  69.230000 ;
        RECT 58.800000  92.220000 74.290000  92.290000 ;
        RECT 58.800000 115.130000 74.290000 115.200000 ;
        RECT 58.800000 138.165000 74.290000 138.235000 ;
        RECT 58.800000 161.180000 74.290000 161.250000 ;
        RECT 58.800000 185.190000 74.290000 185.260000 ;
        RECT 58.815000  80.345000 74.290000  80.415000 ;
        RECT 58.815000 103.345000 74.290000 103.415000 ;
        RECT 58.815000 126.345000 74.290000 126.415000 ;
        RECT 58.815000 149.415000 74.290000 149.485000 ;
        RECT 58.825000  28.600000 74.290000  28.670000 ;
        RECT 58.825000 172.345000 74.290000 172.415000 ;
        RECT 58.855000  57.415000 74.290000  57.485000 ;
        RECT 58.870000  46.060000 74.290000  46.130000 ;
        RECT 58.870000  69.090000 74.290000  69.160000 ;
        RECT 58.870000  92.150000 74.290000  92.220000 ;
        RECT 58.870000 115.060000 74.290000 115.130000 ;
        RECT 58.870000 138.095000 74.290000 138.165000 ;
        RECT 58.870000 161.110000 74.290000 161.180000 ;
        RECT 58.870000 185.120000 74.290000 185.190000 ;
        RECT 58.885000  80.415000 74.290000  80.485000 ;
        RECT 58.885000 103.415000 74.290000 103.485000 ;
        RECT 58.885000 126.415000 74.290000 126.485000 ;
        RECT 58.885000 149.485000 74.290000 149.555000 ;
        RECT 58.895000  28.670000 74.290000  28.740000 ;
        RECT 58.895000 172.415000 74.290000 172.485000 ;
        RECT 58.925000  57.485000 74.290000  57.555000 ;
        RECT 58.940000  45.990000 74.290000  46.060000 ;
        RECT 58.940000  69.020000 74.290000  69.090000 ;
        RECT 58.940000  92.080000 74.290000  92.150000 ;
        RECT 58.940000 114.990000 74.290000 115.060000 ;
        RECT 58.940000 138.025000 74.290000 138.095000 ;
        RECT 58.940000 161.040000 74.290000 161.110000 ;
        RECT 58.940000 185.050000 74.290000 185.120000 ;
        RECT 58.955000  80.485000 74.290000  80.555000 ;
        RECT 58.955000 103.485000 74.290000 103.555000 ;
        RECT 58.955000 126.485000 74.290000 126.555000 ;
        RECT 58.955000 149.555000 74.290000 149.625000 ;
        RECT 58.965000  28.740000 74.290000  28.810000 ;
        RECT 58.965000 172.485000 74.290000 172.555000 ;
        RECT 58.995000  57.555000 74.290000  57.625000 ;
        RECT 59.010000  45.920000 74.290000  45.990000 ;
        RECT 59.010000  68.950000 74.290000  69.020000 ;
        RECT 59.010000  92.010000 74.290000  92.080000 ;
        RECT 59.010000 114.920000 74.290000 114.990000 ;
        RECT 59.010000 137.955000 74.290000 138.025000 ;
        RECT 59.010000 160.970000 74.290000 161.040000 ;
        RECT 59.010000 184.980000 74.290000 185.050000 ;
        RECT 59.025000  80.555000 74.290000  80.625000 ;
        RECT 59.025000 103.555000 74.290000 103.625000 ;
        RECT 59.025000 126.555000 74.290000 126.625000 ;
        RECT 59.025000 149.625000 74.290000 149.695000 ;
        RECT 59.035000  28.810000 74.290000  28.880000 ;
        RECT 59.035000 172.555000 74.290000 172.625000 ;
        RECT 59.065000  57.625000 74.290000  57.695000 ;
        RECT 59.080000  45.850000 74.290000  45.920000 ;
        RECT 59.080000  68.880000 74.290000  68.950000 ;
        RECT 59.080000  91.940000 74.290000  92.010000 ;
        RECT 59.080000 114.850000 74.290000 114.920000 ;
        RECT 59.080000 137.885000 74.290000 137.955000 ;
        RECT 59.080000 160.900000 74.290000 160.970000 ;
        RECT 59.080000 184.910000 74.290000 184.980000 ;
        RECT 59.095000  80.625000 74.290000  80.695000 ;
        RECT 59.095000 103.625000 74.290000 103.695000 ;
        RECT 59.095000 126.625000 74.290000 126.695000 ;
        RECT 59.095000 149.695000 74.290000 149.765000 ;
        RECT 59.105000  28.880000 74.290000  28.950000 ;
        RECT 59.105000 172.625000 74.290000 172.695000 ;
        RECT 59.135000  57.695000 74.290000  57.765000 ;
        RECT 59.150000  45.780000 74.290000  45.850000 ;
        RECT 59.150000  68.810000 74.290000  68.880000 ;
        RECT 59.150000  91.870000 74.290000  91.940000 ;
        RECT 59.150000 114.780000 74.290000 114.850000 ;
        RECT 59.150000 137.815000 74.290000 137.885000 ;
        RECT 59.150000 160.830000 74.290000 160.900000 ;
        RECT 59.150000 184.840000 74.290000 184.910000 ;
        RECT 59.165000  80.695000 74.290000  80.765000 ;
        RECT 59.165000 103.695000 74.290000 103.765000 ;
        RECT 59.165000 126.695000 74.290000 126.765000 ;
        RECT 59.165000 149.765000 74.290000 149.835000 ;
        RECT 59.175000  28.950000 74.290000  29.020000 ;
        RECT 59.175000 172.695000 74.290000 172.765000 ;
        RECT 59.205000  57.765000 74.290000  57.835000 ;
        RECT 59.220000  45.710000 74.290000  45.780000 ;
        RECT 59.220000  68.740000 74.290000  68.810000 ;
        RECT 59.220000  91.800000 74.290000  91.870000 ;
        RECT 59.220000 114.710000 74.290000 114.780000 ;
        RECT 59.220000 137.745000 74.290000 137.815000 ;
        RECT 59.220000 160.760000 74.290000 160.830000 ;
        RECT 59.220000 184.770000 74.290000 184.840000 ;
        RECT 59.235000  80.765000 74.290000  80.835000 ;
        RECT 59.235000 103.765000 74.290000 103.835000 ;
        RECT 59.235000 126.765000 74.290000 126.835000 ;
        RECT 59.235000 149.835000 74.290000 149.905000 ;
        RECT 59.245000  29.020000 74.290000  29.090000 ;
        RECT 59.245000 172.765000 74.290000 172.835000 ;
        RECT 59.275000  57.835000 74.290000  57.905000 ;
        RECT 59.290000  45.640000 74.290000  45.710000 ;
        RECT 59.290000  68.670000 74.290000  68.740000 ;
        RECT 59.290000  91.730000 74.290000  91.800000 ;
        RECT 59.290000 114.640000 74.290000 114.710000 ;
        RECT 59.290000 137.675000 74.290000 137.745000 ;
        RECT 59.290000 160.690000 74.290000 160.760000 ;
        RECT 59.290000 184.700000 74.290000 184.770000 ;
        RECT 59.305000  80.835000 74.290000  80.905000 ;
        RECT 59.305000 103.835000 74.290000 103.905000 ;
        RECT 59.305000 126.835000 74.290000 126.905000 ;
        RECT 59.305000 149.905000 74.290000 149.975000 ;
        RECT 59.315000  29.090000 74.290000  29.160000 ;
        RECT 59.315000 172.835000 74.290000 172.905000 ;
        RECT 59.345000  57.905000 74.290000  57.975000 ;
        RECT 59.360000  45.570000 74.290000  45.640000 ;
        RECT 59.360000  68.600000 74.290000  68.670000 ;
        RECT 59.360000  91.660000 74.290000  91.730000 ;
        RECT 59.360000 114.570000 74.290000 114.640000 ;
        RECT 59.360000 137.605000 74.290000 137.675000 ;
        RECT 59.360000 160.620000 74.290000 160.690000 ;
        RECT 59.360000 184.630000 74.290000 184.700000 ;
        RECT 59.375000  80.905000 74.290000  80.975000 ;
        RECT 59.375000 103.905000 74.290000 103.975000 ;
        RECT 59.375000 126.905000 74.290000 126.975000 ;
        RECT 59.375000 149.975000 74.290000 150.045000 ;
        RECT 59.385000  29.160000 74.290000  29.230000 ;
        RECT 59.385000 172.905000 74.290000 172.975000 ;
        RECT 59.415000  57.975000 74.290000  58.045000 ;
        RECT 59.430000  45.500000 74.290000  45.570000 ;
        RECT 59.430000  68.530000 74.290000  68.600000 ;
        RECT 59.430000  91.590000 74.290000  91.660000 ;
        RECT 59.430000 114.500000 74.290000 114.570000 ;
        RECT 59.430000 137.535000 74.290000 137.605000 ;
        RECT 59.430000 160.550000 74.290000 160.620000 ;
        RECT 59.430000 184.560000 74.290000 184.630000 ;
        RECT 59.445000  80.975000 74.290000  81.045000 ;
        RECT 59.445000 103.975000 74.290000 104.045000 ;
        RECT 59.445000 126.975000 74.290000 127.045000 ;
        RECT 59.445000 150.045000 74.290000 150.115000 ;
        RECT 59.455000  29.230000 74.290000  29.300000 ;
        RECT 59.455000 172.975000 74.290000 173.045000 ;
        RECT 59.485000  58.045000 74.290000  58.115000 ;
        RECT 59.500000  45.430000 74.290000  45.500000 ;
        RECT 59.500000  68.460000 74.290000  68.530000 ;
        RECT 59.500000  91.520000 74.290000  91.590000 ;
        RECT 59.500000 114.430000 74.290000 114.500000 ;
        RECT 59.500000 137.465000 74.290000 137.535000 ;
        RECT 59.500000 160.480000 74.290000 160.550000 ;
        RECT 59.500000 184.490000 74.290000 184.560000 ;
        RECT 59.515000  81.045000 74.290000  81.115000 ;
        RECT 59.515000 104.045000 74.290000 104.115000 ;
        RECT 59.515000 127.045000 74.290000 127.115000 ;
        RECT 59.515000 150.115000 74.290000 150.185000 ;
        RECT 59.525000  29.300000 74.290000  29.370000 ;
        RECT 59.525000 173.045000 74.290000 173.115000 ;
        RECT 59.555000  58.115000 74.290000  58.185000 ;
        RECT 59.570000  45.360000 74.290000  45.430000 ;
        RECT 59.570000  68.390000 74.290000  68.460000 ;
        RECT 59.570000  91.450000 74.290000  91.520000 ;
        RECT 59.570000 114.360000 74.290000 114.430000 ;
        RECT 59.570000 137.395000 74.290000 137.465000 ;
        RECT 59.570000 160.410000 74.290000 160.480000 ;
        RECT 59.570000 184.420000 74.290000 184.490000 ;
        RECT 59.585000  81.115000 74.290000  81.185000 ;
        RECT 59.585000 104.115000 74.290000 104.185000 ;
        RECT 59.585000 127.115000 74.290000 127.185000 ;
        RECT 59.585000 150.185000 74.290000 150.255000 ;
        RECT 59.595000  29.370000 74.290000  29.440000 ;
        RECT 59.595000 173.115000 74.290000 173.185000 ;
        RECT 59.625000  58.185000 74.290000  58.255000 ;
        RECT 59.640000  45.290000 74.290000  45.360000 ;
        RECT 59.640000  68.320000 74.290000  68.390000 ;
        RECT 59.640000  91.380000 74.290000  91.450000 ;
        RECT 59.640000 114.290000 74.290000 114.360000 ;
        RECT 59.640000 137.325000 74.290000 137.395000 ;
        RECT 59.640000 160.340000 74.290000 160.410000 ;
        RECT 59.640000 184.350000 74.290000 184.420000 ;
        RECT 59.655000  81.185000 74.290000  81.255000 ;
        RECT 59.655000 104.185000 74.290000 104.255000 ;
        RECT 59.655000 127.185000 74.290000 127.255000 ;
        RECT 59.655000 150.255000 74.290000 150.325000 ;
        RECT 59.665000  29.440000 74.290000  29.510000 ;
        RECT 59.665000 173.185000 74.290000 173.255000 ;
        RECT 59.695000  58.255000 74.290000  58.325000 ;
        RECT 59.710000  45.220000 74.290000  45.290000 ;
        RECT 59.710000  68.250000 74.290000  68.320000 ;
        RECT 59.710000  91.310000 74.290000  91.380000 ;
        RECT 59.710000 114.220000 74.290000 114.290000 ;
        RECT 59.710000 137.255000 74.290000 137.325000 ;
        RECT 59.710000 160.270000 74.290000 160.340000 ;
        RECT 59.710000 184.280000 74.290000 184.350000 ;
        RECT 59.725000  81.255000 74.290000  81.325000 ;
        RECT 59.725000 104.255000 74.290000 104.325000 ;
        RECT 59.725000 127.255000 74.290000 127.325000 ;
        RECT 59.725000 150.325000 74.290000 150.395000 ;
        RECT 59.735000  29.510000 74.290000  29.580000 ;
        RECT 59.735000 173.255000 74.290000 173.325000 ;
        RECT 59.765000  58.325000 74.290000  58.395000 ;
        RECT 59.780000  45.150000 74.290000  45.220000 ;
        RECT 59.780000  68.180000 74.290000  68.250000 ;
        RECT 59.780000  91.240000 74.290000  91.310000 ;
        RECT 59.780000 114.150000 74.290000 114.220000 ;
        RECT 59.780000 137.185000 74.290000 137.255000 ;
        RECT 59.780000 160.200000 74.290000 160.270000 ;
        RECT 59.780000 184.210000 74.290000 184.280000 ;
        RECT 59.795000  81.325000 74.290000  81.395000 ;
        RECT 59.795000 104.325000 74.290000 104.395000 ;
        RECT 59.795000 127.325000 74.290000 127.395000 ;
        RECT 59.795000 150.395000 74.290000 150.465000 ;
        RECT 59.805000  29.580000 74.290000  29.650000 ;
        RECT 59.805000 173.325000 74.290000 173.395000 ;
        RECT 59.835000  58.395000 74.290000  58.465000 ;
        RECT 59.850000  45.080000 74.290000  45.150000 ;
        RECT 59.850000  68.110000 74.290000  68.180000 ;
        RECT 59.850000  91.170000 74.290000  91.240000 ;
        RECT 59.850000 114.080000 74.290000 114.150000 ;
        RECT 59.850000 137.115000 74.290000 137.185000 ;
        RECT 59.850000 160.130000 74.290000 160.200000 ;
        RECT 59.850000 184.140000 74.290000 184.210000 ;
        RECT 59.865000  81.395000 74.290000  81.465000 ;
        RECT 59.865000 104.395000 74.290000 104.465000 ;
        RECT 59.865000 127.395000 74.290000 127.465000 ;
        RECT 59.865000 150.465000 74.290000 150.535000 ;
        RECT 59.875000  29.650000 74.290000  29.720000 ;
        RECT 59.875000 173.395000 74.290000 173.465000 ;
        RECT 59.905000  58.465000 74.290000  58.535000 ;
        RECT 59.920000  45.010000 74.290000  45.080000 ;
        RECT 59.920000  68.040000 74.290000  68.110000 ;
        RECT 59.920000  91.100000 74.290000  91.170000 ;
        RECT 59.920000 114.010000 74.290000 114.080000 ;
        RECT 59.920000 137.045000 74.290000 137.115000 ;
        RECT 59.920000 160.060000 74.290000 160.130000 ;
        RECT 59.920000 184.070000 74.290000 184.140000 ;
        RECT 59.935000  81.465000 74.290000  81.535000 ;
        RECT 59.935000 104.465000 74.290000 104.535000 ;
        RECT 59.935000 127.465000 74.290000 127.535000 ;
        RECT 59.935000 150.535000 74.290000 150.605000 ;
        RECT 59.945000  29.720000 74.290000  29.790000 ;
        RECT 59.945000 173.465000 74.290000 173.535000 ;
        RECT 59.975000  58.535000 74.290000  58.605000 ;
        RECT 59.990000  44.940000 74.290000  45.010000 ;
        RECT 59.990000  67.970000 74.290000  68.040000 ;
        RECT 59.990000  91.030000 74.290000  91.100000 ;
        RECT 59.990000 113.940000 74.290000 114.010000 ;
        RECT 59.990000 136.975000 74.290000 137.045000 ;
        RECT 59.990000 159.990000 74.290000 160.060000 ;
        RECT 59.990000 184.000000 74.290000 184.070000 ;
        RECT 60.005000  81.535000 74.290000  81.605000 ;
        RECT 60.005000 104.535000 74.290000 104.605000 ;
        RECT 60.005000 127.535000 74.290000 127.605000 ;
        RECT 60.005000 150.605000 74.290000 150.675000 ;
        RECT 60.015000  29.790000 74.290000  29.860000 ;
        RECT 60.015000 173.535000 74.290000 173.605000 ;
        RECT 60.045000  58.605000 74.290000  58.675000 ;
        RECT 60.060000  44.870000 74.290000  44.940000 ;
        RECT 60.060000  67.900000 74.290000  67.970000 ;
        RECT 60.060000  90.960000 74.290000  91.030000 ;
        RECT 60.060000 113.870000 74.290000 113.940000 ;
        RECT 60.060000 136.905000 74.290000 136.975000 ;
        RECT 60.060000 159.920000 74.290000 159.990000 ;
        RECT 60.060000 183.930000 74.290000 184.000000 ;
        RECT 60.075000  81.605000 74.290000  81.675000 ;
        RECT 60.075000 104.605000 74.290000 104.675000 ;
        RECT 60.075000 127.605000 74.290000 127.675000 ;
        RECT 60.075000 150.675000 74.290000 150.745000 ;
        RECT 60.085000  29.860000 74.290000  29.930000 ;
        RECT 60.085000 173.605000 74.290000 173.675000 ;
        RECT 60.115000  58.675000 74.290000  58.745000 ;
        RECT 60.130000  44.800000 74.290000  44.870000 ;
        RECT 60.130000  67.830000 74.290000  67.900000 ;
        RECT 60.130000  90.890000 74.290000  90.960000 ;
        RECT 60.130000 113.800000 74.290000 113.870000 ;
        RECT 60.130000 136.835000 74.290000 136.905000 ;
        RECT 60.130000 159.850000 74.290000 159.920000 ;
        RECT 60.130000 183.860000 74.290000 183.930000 ;
        RECT 60.145000  81.675000 74.290000  81.745000 ;
        RECT 60.145000 104.675000 74.290000 104.745000 ;
        RECT 60.145000 127.675000 74.290000 127.745000 ;
        RECT 60.145000 150.745000 74.290000 150.815000 ;
        RECT 60.155000  29.930000 74.290000  30.000000 ;
        RECT 60.155000 173.675000 74.290000 173.745000 ;
        RECT 60.185000  58.745000 74.290000  58.815000 ;
        RECT 60.200000  44.730000 74.290000  44.800000 ;
        RECT 60.200000  67.760000 74.290000  67.830000 ;
        RECT 60.200000  90.820000 74.290000  90.890000 ;
        RECT 60.200000 113.730000 74.290000 113.800000 ;
        RECT 60.200000 136.765000 74.290000 136.835000 ;
        RECT 60.200000 159.780000 74.290000 159.850000 ;
        RECT 60.200000 183.790000 74.290000 183.860000 ;
        RECT 60.215000  81.745000 74.290000  81.815000 ;
        RECT 60.215000 104.745000 74.290000 104.815000 ;
        RECT 60.215000 127.745000 74.290000 127.815000 ;
        RECT 60.215000 150.815000 74.290000 150.885000 ;
        RECT 60.225000  30.000000 74.290000  30.070000 ;
        RECT 60.225000 173.745000 74.290000 173.815000 ;
        RECT 60.255000  58.815000 74.290000  58.885000 ;
        RECT 60.270000  44.660000 74.290000  44.730000 ;
        RECT 60.270000  67.690000 74.290000  67.760000 ;
        RECT 60.270000  90.750000 74.290000  90.820000 ;
        RECT 60.270000 113.660000 74.290000 113.730000 ;
        RECT 60.270000 136.695000 74.290000 136.765000 ;
        RECT 60.270000 159.710000 74.290000 159.780000 ;
        RECT 60.270000 183.720000 74.290000 183.790000 ;
        RECT 60.285000  81.815000 74.290000  81.885000 ;
        RECT 60.285000 104.815000 74.290000 104.885000 ;
        RECT 60.285000 127.815000 74.290000 127.885000 ;
        RECT 60.285000 150.885000 74.290000 150.955000 ;
        RECT 60.295000  30.070000 74.290000  30.140000 ;
        RECT 60.295000 173.815000 74.290000 173.885000 ;
        RECT 60.325000  58.885000 74.290000  58.955000 ;
        RECT 60.340000  44.590000 74.290000  44.660000 ;
        RECT 60.340000  67.620000 74.290000  67.690000 ;
        RECT 60.340000  90.680000 74.290000  90.750000 ;
        RECT 60.340000 113.590000 74.290000 113.660000 ;
        RECT 60.340000 136.625000 74.290000 136.695000 ;
        RECT 60.340000 159.640000 74.290000 159.710000 ;
        RECT 60.340000 183.650000 74.290000 183.720000 ;
        RECT 60.355000  81.885000 74.290000  81.955000 ;
        RECT 60.355000 104.885000 74.290000 104.955000 ;
        RECT 60.355000 127.885000 74.290000 127.955000 ;
        RECT 60.355000 150.955000 74.290000 151.025000 ;
        RECT 60.365000  30.140000 74.290000  30.210000 ;
        RECT 60.365000 173.885000 74.290000 173.955000 ;
        RECT 60.395000  58.955000 74.290000  59.025000 ;
        RECT 60.410000  44.520000 74.290000  44.590000 ;
        RECT 60.410000  67.550000 74.290000  67.620000 ;
        RECT 60.410000  90.610000 74.290000  90.680000 ;
        RECT 60.410000 113.520000 74.290000 113.590000 ;
        RECT 60.410000 136.555000 74.290000 136.625000 ;
        RECT 60.410000 159.570000 74.290000 159.640000 ;
        RECT 60.410000 183.580000 74.290000 183.650000 ;
        RECT 60.425000  81.955000 74.290000  82.025000 ;
        RECT 60.425000 104.955000 74.290000 105.025000 ;
        RECT 60.425000 127.955000 74.290000 128.025000 ;
        RECT 60.425000 151.025000 74.290000 151.095000 ;
        RECT 60.435000  30.210000 74.290000  30.280000 ;
        RECT 60.435000 173.955000 74.290000 174.025000 ;
        RECT 60.465000  59.025000 74.290000  59.095000 ;
        RECT 60.480000  44.450000 74.290000  44.520000 ;
        RECT 60.480000  67.480000 74.290000  67.550000 ;
        RECT 60.480000  90.540000 74.290000  90.610000 ;
        RECT 60.480000 113.450000 74.290000 113.520000 ;
        RECT 60.480000 136.485000 74.290000 136.555000 ;
        RECT 60.480000 159.500000 74.290000 159.570000 ;
        RECT 60.480000 183.510000 74.290000 183.580000 ;
        RECT 60.495000  82.025000 74.290000  82.095000 ;
        RECT 60.495000 105.025000 74.290000 105.095000 ;
        RECT 60.495000 128.025000 74.290000 128.095000 ;
        RECT 60.495000 151.095000 74.290000 151.165000 ;
        RECT 60.505000  30.280000 74.290000  30.350000 ;
        RECT 60.505000 174.025000 74.290000 174.095000 ;
        RECT 60.535000  59.095000 74.290000  59.165000 ;
        RECT 60.550000  44.380000 74.290000  44.450000 ;
        RECT 60.550000  67.410000 74.290000  67.480000 ;
        RECT 60.550000  90.470000 74.290000  90.540000 ;
        RECT 60.550000 113.380000 74.290000 113.450000 ;
        RECT 60.550000 136.415000 74.290000 136.485000 ;
        RECT 60.550000 159.430000 74.290000 159.500000 ;
        RECT 60.550000 183.440000 74.290000 183.510000 ;
        RECT 60.565000  82.095000 74.290000  82.165000 ;
        RECT 60.565000 105.095000 74.290000 105.165000 ;
        RECT 60.565000 128.095000 74.290000 128.165000 ;
        RECT 60.565000 151.165000 74.290000 151.235000 ;
        RECT 60.575000  30.350000 74.290000  30.420000 ;
        RECT 60.575000 174.095000 74.290000 174.165000 ;
        RECT 60.605000  59.165000 74.290000  59.235000 ;
        RECT 60.620000  44.310000 74.290000  44.380000 ;
        RECT 60.620000  67.340000 74.290000  67.410000 ;
        RECT 60.620000  90.400000 74.290000  90.470000 ;
        RECT 60.620000 113.310000 74.290000 113.380000 ;
        RECT 60.620000 136.345000 74.290000 136.415000 ;
        RECT 60.620000 159.360000 74.290000 159.430000 ;
        RECT 60.620000 183.370000 74.290000 183.440000 ;
        RECT 60.635000  82.165000 74.290000  82.235000 ;
        RECT 60.635000 105.165000 74.290000 105.235000 ;
        RECT 60.635000 128.165000 74.290000 128.235000 ;
        RECT 60.635000 151.235000 74.290000 151.305000 ;
        RECT 60.645000  30.420000 74.290000  30.490000 ;
        RECT 60.645000 174.165000 74.290000 174.235000 ;
        RECT 60.675000  59.235000 74.290000  59.305000 ;
        RECT 60.690000  44.240000 74.290000  44.310000 ;
        RECT 60.690000  67.270000 74.290000  67.340000 ;
        RECT 60.690000  90.330000 74.290000  90.400000 ;
        RECT 60.690000 113.240000 74.290000 113.310000 ;
        RECT 60.690000 136.275000 74.290000 136.345000 ;
        RECT 60.690000 159.290000 74.290000 159.360000 ;
        RECT 60.690000 183.300000 74.290000 183.370000 ;
        RECT 60.705000  82.235000 74.290000  82.305000 ;
        RECT 60.705000 105.235000 74.290000 105.305000 ;
        RECT 60.705000 128.235000 74.290000 128.305000 ;
        RECT 60.705000 151.305000 74.290000 151.375000 ;
        RECT 60.715000  30.490000 74.290000  30.560000 ;
        RECT 60.715000 174.235000 74.290000 174.305000 ;
        RECT 60.745000  59.305000 74.290000  59.375000 ;
        RECT 60.760000  44.170000 74.290000  44.240000 ;
        RECT 60.760000  67.200000 74.290000  67.270000 ;
        RECT 60.760000  90.260000 74.290000  90.330000 ;
        RECT 60.760000 113.170000 74.290000 113.240000 ;
        RECT 60.760000 136.205000 74.290000 136.275000 ;
        RECT 60.760000 159.220000 74.290000 159.290000 ;
        RECT 60.760000 183.230000 74.290000 183.300000 ;
        RECT 60.775000  82.305000 74.290000  82.375000 ;
        RECT 60.775000 105.305000 74.290000 105.375000 ;
        RECT 60.775000 128.305000 74.290000 128.375000 ;
        RECT 60.775000 151.375000 74.290000 151.445000 ;
        RECT 60.785000  30.560000 74.290000  30.630000 ;
        RECT 60.785000 174.305000 74.290000 174.375000 ;
        RECT 60.815000  59.375000 74.290000  59.445000 ;
        RECT 60.830000  44.100000 74.290000  44.170000 ;
        RECT 60.830000  67.130000 74.290000  67.200000 ;
        RECT 60.830000  90.190000 74.290000  90.260000 ;
        RECT 60.830000 113.100000 74.290000 113.170000 ;
        RECT 60.830000 136.135000 74.290000 136.205000 ;
        RECT 60.830000 159.150000 74.290000 159.220000 ;
        RECT 60.830000 183.160000 74.290000 183.230000 ;
        RECT 60.845000  82.375000 74.290000  82.445000 ;
        RECT 60.845000 105.375000 74.290000 105.445000 ;
        RECT 60.845000 128.375000 74.290000 128.445000 ;
        RECT 60.845000 151.445000 74.290000 151.515000 ;
        RECT 60.855000  30.630000 74.290000  30.700000 ;
        RECT 60.855000 174.375000 74.290000 174.445000 ;
        RECT 60.885000  59.445000 74.290000  59.515000 ;
        RECT 60.900000  44.030000 74.290000  44.100000 ;
        RECT 60.900000  67.060000 74.290000  67.130000 ;
        RECT 60.900000  90.120000 74.290000  90.190000 ;
        RECT 60.900000 113.030000 74.290000 113.100000 ;
        RECT 60.900000 136.065000 74.290000 136.135000 ;
        RECT 60.900000 159.080000 74.290000 159.150000 ;
        RECT 60.900000 183.090000 74.290000 183.160000 ;
        RECT 60.915000  82.445000 74.290000  82.515000 ;
        RECT 60.915000 105.445000 74.290000 105.515000 ;
        RECT 60.915000 128.445000 74.290000 128.515000 ;
        RECT 60.915000 151.515000 74.290000 151.585000 ;
        RECT 60.925000  30.700000 74.290000  30.770000 ;
        RECT 60.925000 174.445000 74.290000 174.515000 ;
        RECT 60.955000  59.515000 74.290000  59.585000 ;
        RECT 60.970000  43.960000 74.290000  44.030000 ;
        RECT 60.970000  66.990000 74.290000  67.060000 ;
        RECT 60.970000  90.050000 74.290000  90.120000 ;
        RECT 60.970000 112.960000 74.290000 113.030000 ;
        RECT 60.970000 135.995000 74.290000 136.065000 ;
        RECT 60.970000 159.010000 74.290000 159.080000 ;
        RECT 60.970000 183.020000 74.290000 183.090000 ;
        RECT 60.985000  82.515000 74.290000  82.585000 ;
        RECT 60.985000 105.515000 74.290000 105.585000 ;
        RECT 60.985000 128.515000 74.290000 128.585000 ;
        RECT 60.985000 151.585000 74.290000 151.655000 ;
        RECT 60.995000  30.770000 74.290000  30.840000 ;
        RECT 60.995000 174.515000 74.290000 174.585000 ;
        RECT 61.025000  59.585000 74.290000  59.655000 ;
        RECT 61.040000  43.890000 74.290000  43.960000 ;
        RECT 61.040000  66.920000 74.290000  66.990000 ;
        RECT 61.040000  89.980000 74.290000  90.050000 ;
        RECT 61.040000 112.890000 74.290000 112.960000 ;
        RECT 61.040000 135.925000 74.290000 135.995000 ;
        RECT 61.040000 158.940000 74.290000 159.010000 ;
        RECT 61.040000 182.950000 74.290000 183.020000 ;
        RECT 61.055000  82.585000 74.290000  82.655000 ;
        RECT 61.055000 105.585000 74.290000 105.655000 ;
        RECT 61.055000 128.585000 74.290000 128.655000 ;
        RECT 61.055000 151.655000 74.290000 151.725000 ;
        RECT 61.065000  30.840000 74.290000  30.910000 ;
        RECT 61.065000 174.585000 74.290000 174.655000 ;
        RECT 61.095000  59.655000 74.290000  59.725000 ;
        RECT 61.110000  30.910000 74.290000  30.955000 ;
        RECT 61.110000  30.955000 74.290000  43.820000 ;
        RECT 61.110000  43.820000 74.290000  43.890000 ;
        RECT 61.110000  59.725000 74.290000  59.740000 ;
        RECT 61.110000  59.740000 74.290000  66.850000 ;
        RECT 61.110000  66.850000 74.290000  66.920000 ;
        RECT 61.110000  82.655000 74.290000  82.710000 ;
        RECT 61.110000  82.710000 74.290000  89.910000 ;
        RECT 61.110000  89.910000 74.290000  89.980000 ;
        RECT 61.110000 105.655000 74.290000 105.710000 ;
        RECT 61.110000 105.710000 74.290000 112.820000 ;
        RECT 61.110000 112.820000 74.290000 112.890000 ;
        RECT 61.110000 128.655000 74.290000 128.710000 ;
        RECT 61.110000 128.710000 74.290000 135.855000 ;
        RECT 61.110000 135.855000 74.290000 135.925000 ;
        RECT 61.110000 151.725000 74.290000 151.780000 ;
        RECT 61.110000 151.780000 74.290000 158.870000 ;
        RECT 61.110000 158.870000 74.290000 158.940000 ;
        RECT 61.110000 174.655000 74.290000 174.700000 ;
        RECT 61.110000 174.700000 74.290000 182.880000 ;
        RECT 61.110000 182.880000 74.290000 182.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000   0.000000 48.890000  96.150000 ;
        RECT 37.890000  96.150000 48.890000  96.300000 ;
        RECT 37.890000  96.300000 49.040000  96.450000 ;
        RECT 37.890000  96.450000 49.190000  96.600000 ;
        RECT 37.890000  96.600000 49.340000  96.750000 ;
        RECT 37.890000  96.750000 49.490000  96.900000 ;
        RECT 37.890000  96.900000 49.640000  97.050000 ;
        RECT 37.890000  97.050000 49.790000  97.200000 ;
        RECT 37.890000  97.200000 49.940000  97.350000 ;
        RECT 37.890000  97.350000 50.090000  97.500000 ;
        RECT 37.890000  97.500000 50.240000  97.650000 ;
        RECT 37.890000  97.650000 50.390000  97.800000 ;
        RECT 37.890000  97.800000 50.540000  97.950000 ;
        RECT 37.890000  97.950000 50.690000  98.100000 ;
        RECT 37.890000  98.100000 50.840000  98.250000 ;
        RECT 37.890000  98.250000 50.990000  98.300000 ;
        RECT 37.890000  98.300000 51.040000  99.505000 ;
        RECT 37.890000  99.505000 43.400000  99.655000 ;
        RECT 37.890000  99.655000 43.250000  99.805000 ;
        RECT 37.890000  99.805000 43.100000  99.955000 ;
        RECT 37.890000  99.955000 42.950000 100.105000 ;
        RECT 37.890000 100.105000 42.840000 100.215000 ;
        RECT 37.890000 100.215000 42.840000 102.135000 ;
        RECT 37.890000 102.135000 42.840000 102.285000 ;
        RECT 37.890000 102.285000 42.990000 102.435000 ;
        RECT 37.890000 102.435000 43.140000 102.585000 ;
        RECT 37.890000 102.585000 43.290000 102.735000 ;
        RECT 37.890000 102.735000 43.440000 102.885000 ;
        RECT 37.890000 102.885000 43.590000 103.035000 ;
        RECT 37.890000 103.035000 43.740000 103.185000 ;
        RECT 37.890000 103.185000 43.890000 103.335000 ;
        RECT 37.890000 103.335000 44.040000 103.485000 ;
        RECT 37.890000 103.485000 44.190000 103.635000 ;
        RECT 37.890000 103.635000 44.340000 103.785000 ;
        RECT 37.890000 103.785000 44.490000 103.935000 ;
        RECT 37.890000 103.935000 44.640000 104.085000 ;
        RECT 37.890000 104.085000 44.790000 104.235000 ;
        RECT 37.890000 104.235000 44.940000 104.385000 ;
        RECT 37.890000 104.385000 45.090000 104.535000 ;
        RECT 37.890000 104.535000 45.240000 104.685000 ;
        RECT 37.890000 104.685000 45.390000 104.835000 ;
        RECT 37.890000 104.835000 45.540000 104.985000 ;
        RECT 37.890000 104.985000 45.690000 105.135000 ;
        RECT 37.890000 105.135000 45.840000 105.285000 ;
        RECT 37.890000 105.285000 45.990000 105.435000 ;
        RECT 37.890000 105.435000 46.140000 105.585000 ;
        RECT 37.890000 105.585000 46.290000 105.655000 ;
        RECT 37.965000 175.350000 48.855000 190.020000 ;
        RECT 38.040000 105.655000 46.360000 105.805000 ;
        RECT 38.055000 175.260000 48.855000 175.350000 ;
        RECT 38.190000 105.805000 46.510000 105.955000 ;
        RECT 38.205000 175.110000 48.855000 175.260000 ;
        RECT 38.340000 105.955000 46.660000 106.105000 ;
        RECT 38.355000 174.960000 48.855000 175.110000 ;
        RECT 38.490000 106.105000 46.810000 106.255000 ;
        RECT 38.505000 174.810000 48.855000 174.960000 ;
        RECT 38.640000 106.255000 46.960000 106.405000 ;
        RECT 38.655000 174.660000 48.855000 174.810000 ;
        RECT 38.790000 106.405000 47.110000 106.555000 ;
        RECT 38.805000 174.510000 48.855000 174.660000 ;
        RECT 38.940000 106.555000 47.260000 106.705000 ;
        RECT 38.955000 174.360000 48.855000 174.510000 ;
        RECT 39.090000 106.705000 47.410000 106.855000 ;
        RECT 39.105000 174.210000 48.855000 174.360000 ;
        RECT 39.240000 106.855000 47.560000 107.005000 ;
        RECT 39.255000 174.060000 48.855000 174.210000 ;
        RECT 39.390000 107.005000 47.710000 107.155000 ;
        RECT 39.405000 173.910000 48.855000 174.060000 ;
        RECT 39.540000 107.155000 47.860000 107.305000 ;
        RECT 39.555000 173.760000 48.855000 173.910000 ;
        RECT 39.690000 107.305000 48.010000 107.455000 ;
        RECT 39.705000 173.610000 48.855000 173.760000 ;
        RECT 39.840000 107.455000 48.160000 107.605000 ;
        RECT 39.855000 173.460000 48.855000 173.610000 ;
        RECT 39.990000 107.605000 48.310000 107.755000 ;
        RECT 40.005000 173.310000 48.855000 173.460000 ;
        RECT 40.140000 107.755000 48.460000 107.905000 ;
        RECT 40.155000 173.160000 48.855000 173.310000 ;
        RECT 40.290000 107.905000 48.610000 108.055000 ;
        RECT 40.305000 173.010000 48.855000 173.160000 ;
        RECT 40.385000 108.055000 48.760000 108.150000 ;
        RECT 40.455000 172.860000 48.855000 173.010000 ;
        RECT 40.535000 108.150000 48.855000 108.300000 ;
        RECT 40.605000 172.710000 48.855000 172.860000 ;
        RECT 40.685000 108.300000 48.855000 108.450000 ;
        RECT 40.755000 172.560000 48.855000 172.710000 ;
        RECT 40.835000 108.450000 48.855000 108.600000 ;
        RECT 40.905000 172.410000 48.855000 172.560000 ;
        RECT 40.985000 108.600000 48.855000 108.750000 ;
        RECT 41.055000 172.260000 48.855000 172.410000 ;
        RECT 41.135000 108.750000 48.855000 108.900000 ;
        RECT 41.205000 172.110000 48.855000 172.260000 ;
        RECT 41.285000 108.900000 48.855000 109.050000 ;
        RECT 41.355000 171.960000 48.855000 172.110000 ;
        RECT 41.435000 109.050000 48.855000 109.200000 ;
        RECT 41.505000 171.810000 48.855000 171.960000 ;
        RECT 41.585000 109.200000 48.855000 109.350000 ;
        RECT 41.655000 171.660000 48.855000 171.810000 ;
        RECT 41.735000 109.350000 48.855000 109.500000 ;
        RECT 41.805000 171.510000 48.855000 171.660000 ;
        RECT 41.885000 109.500000 48.855000 109.650000 ;
        RECT 41.955000 171.360000 48.855000 171.510000 ;
        RECT 42.035000 109.650000 48.855000 109.800000 ;
        RECT 42.105000 171.210000 48.855000 171.360000 ;
        RECT 42.185000 109.800000 48.855000 109.950000 ;
        RECT 42.255000 171.060000 48.855000 171.210000 ;
        RECT 42.335000 109.950000 48.855000 110.100000 ;
        RECT 42.405000 170.910000 48.855000 171.060000 ;
        RECT 42.485000 110.100000 48.855000 110.250000 ;
        RECT 42.555000 170.760000 48.855000 170.910000 ;
        RECT 42.635000 110.250000 48.855000 110.400000 ;
        RECT 42.705000 170.610000 48.855000 170.760000 ;
        RECT 42.785000 110.400000 48.855000 110.550000 ;
        RECT 42.855000 110.550000 48.855000 110.620000 ;
        RECT 42.855000 110.620000 48.855000 170.460000 ;
        RECT 42.855000 170.460000 48.855000 170.610000 ;
        RECT 44.655000  99.505000 51.040000  99.610000 ;
        RECT 44.760000  99.610000 51.040000  99.715000 ;
        RECT 44.910000  99.715000 51.040000  99.865000 ;
        RECT 45.060000  99.865000 51.190000 100.015000 ;
        RECT 45.210000 100.015000 51.340000 100.165000 ;
        RECT 45.260000 100.165000 51.490000 100.215000 ;
        RECT 45.260000 100.215000 51.540000 100.365000 ;
        RECT 45.260000 100.365000 51.690000 100.515000 ;
        RECT 45.260000 100.515000 51.840000 100.665000 ;
        RECT 45.260000 100.665000 51.990000 100.815000 ;
        RECT 45.260000 100.815000 52.140000 100.965000 ;
        RECT 45.260000 100.965000 52.290000 101.115000 ;
        RECT 45.260000 101.115000 52.440000 101.265000 ;
        RECT 45.260000 101.265000 52.590000 101.415000 ;
        RECT 45.260000 101.415000 52.740000 101.565000 ;
        RECT 45.260000 101.565000 52.890000 101.715000 ;
        RECT 45.260000 101.715000 53.040000 101.865000 ;
        RECT 45.260000 101.865000 53.190000 102.015000 ;
        RECT 45.260000 102.015000 53.340000 102.165000 ;
        RECT 45.260000 102.165000 53.490000 102.315000 ;
        RECT 45.260000 102.315000 53.640000 102.415000 ;
        RECT 45.410000 102.415000 53.740000 102.565000 ;
        RECT 45.560000 102.565000 53.890000 102.715000 ;
        RECT 45.710000 102.715000 54.040000 102.865000 ;
        RECT 45.860000 102.865000 54.190000 103.015000 ;
        RECT 46.010000 103.015000 54.340000 103.165000 ;
        RECT 46.160000 103.165000 54.490000 103.315000 ;
        RECT 46.310000 103.315000 54.640000 103.465000 ;
        RECT 46.460000 103.465000 54.790000 103.615000 ;
        RECT 46.610000 103.615000 54.940000 103.765000 ;
        RECT 46.760000 103.765000 55.090000 103.915000 ;
        RECT 46.910000 103.915000 55.240000 104.065000 ;
        RECT 47.060000 104.065000 55.390000 104.215000 ;
        RECT 47.210000 104.215000 55.540000 104.365000 ;
        RECT 47.360000 104.365000 55.690000 104.515000 ;
        RECT 47.510000 104.515000 55.840000 104.665000 ;
        RECT 47.660000 104.665000 55.990000 104.815000 ;
        RECT 47.810000 104.815000 56.140000 104.965000 ;
        RECT 47.960000 104.965000 56.290000 105.115000 ;
        RECT 48.110000 105.115000 56.440000 105.265000 ;
        RECT 48.260000 105.265000 56.590000 105.415000 ;
        RECT 48.410000 105.415000 56.740000 105.565000 ;
        RECT 48.560000 105.565000 56.890000 105.715000 ;
        RECT 48.710000 105.715000 57.040000 105.865000 ;
        RECT 48.860000 105.865000 57.190000 106.015000 ;
        RECT 49.010000 106.015000 57.340000 106.165000 ;
        RECT 49.160000 106.165000 57.490000 106.315000 ;
        RECT 49.310000 106.315000 57.640000 106.465000 ;
        RECT 49.460000 106.465000 57.790000 106.615000 ;
        RECT 49.610000 106.615000 57.940000 106.765000 ;
        RECT 49.760000 106.765000 58.090000 106.915000 ;
        RECT 49.775000 172.645000 59.285000 173.020000 ;
        RECT 49.775000 173.020000 59.285000 173.170000 ;
        RECT 49.775000 173.170000 59.435000 173.320000 ;
        RECT 49.775000 173.320000 59.585000 173.470000 ;
        RECT 49.775000 173.470000 59.735000 173.620000 ;
        RECT 49.775000 173.620000 59.885000 173.770000 ;
        RECT 49.775000 173.770000 60.035000 173.920000 ;
        RECT 49.775000 173.920000 60.185000 174.070000 ;
        RECT 49.775000 174.070000 60.335000 174.220000 ;
        RECT 49.775000 174.220000 60.485000 174.370000 ;
        RECT 49.775000 174.370000 60.635000 174.520000 ;
        RECT 49.775000 174.520000 60.785000 174.670000 ;
        RECT 49.775000 174.670000 60.935000 174.680000 ;
        RECT 49.775000 174.680000 60.945000 190.040000 ;
        RECT 49.835000 172.585000 59.285000 172.645000 ;
        RECT 49.910000 106.915000 58.240000 107.065000 ;
        RECT 49.985000 172.435000 59.285000 172.585000 ;
        RECT 50.060000 107.065000 58.390000 107.215000 ;
        RECT 50.135000 172.285000 59.285000 172.435000 ;
        RECT 50.210000 107.215000 58.540000 107.365000 ;
        RECT 50.285000 172.135000 59.285000 172.285000 ;
        RECT 50.360000 107.365000 58.690000 107.515000 ;
        RECT 50.435000 171.985000 59.285000 172.135000 ;
        RECT 50.510000 107.515000 58.840000 107.665000 ;
        RECT 50.585000 171.835000 59.285000 171.985000 ;
        RECT 50.660000 107.665000 58.990000 107.815000 ;
        RECT 50.735000 171.685000 59.285000 171.835000 ;
        RECT 50.805000 107.815000 59.140000 107.960000 ;
        RECT 50.885000 171.535000 59.285000 171.685000 ;
        RECT 50.955000 107.960000 59.285000 108.110000 ;
        RECT 51.035000 171.385000 59.285000 171.535000 ;
        RECT 51.105000 108.110000 59.285000 108.260000 ;
        RECT 51.185000 171.235000 59.285000 171.385000 ;
        RECT 51.255000 108.260000 59.285000 108.410000 ;
        RECT 51.335000 171.085000 59.285000 171.235000 ;
        RECT 51.405000 108.410000 59.285000 108.560000 ;
        RECT 51.485000 170.935000 59.285000 171.085000 ;
        RECT 51.555000 108.560000 59.285000 108.710000 ;
        RECT 51.635000 170.785000 59.285000 170.935000 ;
        RECT 51.705000 108.710000 59.285000 108.860000 ;
        RECT 51.785000 170.635000 59.285000 170.785000 ;
        RECT 51.855000 108.860000 59.285000 109.010000 ;
        RECT 51.935000 170.485000 59.285000 170.635000 ;
        RECT 52.005000 109.010000 59.285000 109.160000 ;
        RECT 52.085000 170.335000 59.285000 170.485000 ;
        RECT 52.155000 109.160000 59.285000 109.310000 ;
        RECT 52.235000 170.185000 59.285000 170.335000 ;
        RECT 52.305000 109.310000 59.285000 109.460000 ;
        RECT 52.385000 170.035000 59.285000 170.185000 ;
        RECT 52.455000 109.460000 59.285000 109.610000 ;
        RECT 52.535000 169.885000 59.285000 170.035000 ;
        RECT 52.605000 109.610000 59.285000 109.760000 ;
        RECT 52.685000 169.735000 59.285000 169.885000 ;
        RECT 52.755000 109.760000 59.285000 109.910000 ;
        RECT 52.835000 169.585000 59.285000 169.735000 ;
        RECT 52.905000 109.910000 59.285000 110.060000 ;
        RECT 52.985000 169.435000 59.285000 169.585000 ;
        RECT 53.055000 110.060000 59.285000 110.210000 ;
        RECT 53.135000 169.285000 59.285000 169.435000 ;
        RECT 53.205000 110.210000 59.285000 110.360000 ;
        RECT 53.285000 110.360000 59.285000 110.440000 ;
        RECT 53.285000 110.440000 59.285000 169.135000 ;
        RECT 53.285000 169.135000 59.285000 169.285000 ;
    END
  END DRN_HVC
  PIN G_CORE
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.495000   0.000000 24.395000  36.510000 ;
        RECT 0.495000  46.960000 24.395000  90.500000 ;
        RECT 0.495000  90.500000 24.245000  90.650000 ;
        RECT 0.495000  90.650000 24.095000  90.800000 ;
        RECT 0.495000  90.800000 23.945000  90.950000 ;
        RECT 0.495000  90.950000 23.795000  91.100000 ;
        RECT 0.495000  91.100000 23.645000  91.250000 ;
        RECT 0.495000  91.250000 23.495000  91.400000 ;
        RECT 0.495000  91.400000 23.345000  91.550000 ;
        RECT 0.495000  91.550000 23.195000  91.700000 ;
        RECT 0.495000  91.700000 23.045000  91.850000 ;
        RECT 0.495000  91.850000 22.895000  92.000000 ;
        RECT 0.495000  92.000000 22.745000  92.150000 ;
        RECT 0.495000  92.150000 22.595000  92.300000 ;
        RECT 0.495000  92.300000 22.445000  92.450000 ;
        RECT 0.495000  92.450000 22.295000  92.600000 ;
        RECT 0.495000  92.600000 22.145000  92.750000 ;
        RECT 0.495000  92.750000 21.995000  92.900000 ;
        RECT 0.495000  92.900000 21.845000  93.050000 ;
        RECT 0.495000  93.050000 21.695000  93.200000 ;
        RECT 0.495000  93.200000 21.545000  93.350000 ;
        RECT 0.495000  93.350000 21.395000  93.500000 ;
        RECT 0.495000  93.500000 21.245000  93.650000 ;
        RECT 0.495000  93.650000 21.095000  93.800000 ;
        RECT 0.495000  93.800000 20.945000  93.950000 ;
        RECT 0.495000  93.950000 20.795000  94.100000 ;
        RECT 0.495000  94.100000 20.645000  94.250000 ;
        RECT 0.495000  94.250000 20.495000  94.400000 ;
        RECT 0.495000  94.400000 20.345000  94.550000 ;
        RECT 0.495000  94.550000 20.195000  94.700000 ;
        RECT 0.495000  94.700000 20.045000  94.850000 ;
        RECT 0.495000  94.850000 19.895000  95.000000 ;
        RECT 0.495000  95.000000 19.745000  95.150000 ;
        RECT 0.495000  95.150000 19.595000  95.300000 ;
        RECT 0.495000  95.300000 19.445000  95.450000 ;
        RECT 0.495000  95.450000 19.295000  95.600000 ;
        RECT 0.495000  95.600000 19.145000  95.750000 ;
        RECT 0.495000  95.750000 18.995000  95.900000 ;
        RECT 0.495000  95.900000 18.845000  96.050000 ;
        RECT 0.495000  96.050000 18.695000  96.200000 ;
        RECT 0.495000  96.200000 18.545000  96.350000 ;
        RECT 0.495000  96.350000 18.395000  96.500000 ;
        RECT 0.495000  96.500000 18.245000  96.650000 ;
        RECT 0.495000  96.650000 18.095000  96.800000 ;
        RECT 0.495000  96.800000 17.945000  96.950000 ;
        RECT 0.495000  96.950000 17.795000  97.100000 ;
        RECT 0.495000  97.100000 17.645000  97.250000 ;
        RECT 0.495000  97.250000 17.495000  97.400000 ;
        RECT 0.495000  97.400000 17.345000  97.550000 ;
        RECT 0.495000  97.550000 17.195000  97.700000 ;
        RECT 0.495000  97.700000 17.045000  97.850000 ;
        RECT 0.495000  97.850000 16.895000  98.000000 ;
        RECT 0.495000  98.000000 16.745000  98.150000 ;
        RECT 0.495000  98.150000 16.595000  98.300000 ;
        RECT 0.495000  98.300000 16.445000  98.450000 ;
        RECT 0.495000  98.450000 16.295000  98.600000 ;
        RECT 0.495000  98.600000 16.145000  98.750000 ;
        RECT 0.495000  98.750000 15.995000  98.900000 ;
        RECT 0.495000  98.900000 15.845000  99.050000 ;
        RECT 0.495000  99.050000 15.695000  99.200000 ;
        RECT 0.495000  99.200000 15.545000  99.350000 ;
        RECT 0.495000  99.350000 15.395000  99.500000 ;
        RECT 0.495000  99.500000 15.245000  99.650000 ;
        RECT 0.495000  99.650000 15.095000  99.800000 ;
        RECT 0.495000  99.800000 14.945000  99.950000 ;
        RECT 0.495000  99.950000 14.795000 100.100000 ;
        RECT 0.495000 100.100000 14.645000 100.250000 ;
        RECT 0.495000 100.250000 14.495000 100.400000 ;
        RECT 0.495000 100.400000 14.345000 100.550000 ;
        RECT 0.495000 100.550000 14.195000 100.700000 ;
        RECT 0.495000 100.700000 14.045000 100.850000 ;
        RECT 0.495000 100.850000 13.895000 101.000000 ;
        RECT 0.495000 101.000000 13.745000 101.150000 ;
        RECT 0.495000 101.150000 13.595000 101.300000 ;
        RECT 0.495000 101.300000 13.500000 101.395000 ;
        RECT 0.495000 101.395000 13.500000 173.155000 ;
        RECT 0.520000  46.935000 24.395000  46.960000 ;
        RECT 0.645000  36.510000 24.395000  36.660000 ;
        RECT 0.670000  46.785000 24.395000  46.935000 ;
        RECT 0.795000  36.660000 24.395000  36.810000 ;
        RECT 0.820000  46.635000 24.395000  46.785000 ;
        RECT 0.945000  36.810000 24.395000  36.960000 ;
        RECT 0.970000  36.960000 24.395000  36.985000 ;
        RECT 0.970000  36.985000 24.395000  46.485000 ;
        RECT 0.970000  46.485000 24.395000  46.635000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390000   0.000000 74.290000  90.185000 ;
        RECT 50.540000  90.185000 74.290000  90.335000 ;
        RECT 50.690000  90.335000 74.290000  90.485000 ;
        RECT 50.840000  90.485000 74.290000  90.635000 ;
        RECT 50.990000  90.635000 74.290000  90.785000 ;
        RECT 51.140000  90.785000 74.290000  90.935000 ;
        RECT 51.290000  90.935000 74.290000  91.085000 ;
        RECT 51.440000  91.085000 74.290000  91.235000 ;
        RECT 51.590000  91.235000 74.290000  91.385000 ;
        RECT 51.740000  91.385000 74.290000  91.535000 ;
        RECT 51.890000  91.535000 74.290000  91.685000 ;
        RECT 52.040000  91.685000 74.290000  91.835000 ;
        RECT 52.190000  91.835000 74.290000  91.985000 ;
        RECT 52.340000  91.985000 74.290000  92.135000 ;
        RECT 52.490000  92.135000 74.290000  92.285000 ;
        RECT 52.640000  92.285000 74.290000  92.435000 ;
        RECT 52.790000  92.435000 74.290000  92.585000 ;
        RECT 52.940000  92.585000 74.290000  92.735000 ;
        RECT 53.090000  92.735000 74.290000  92.885000 ;
        RECT 53.240000  92.885000 74.290000  93.035000 ;
        RECT 53.390000  93.035000 74.290000  93.185000 ;
        RECT 53.540000  93.185000 74.290000  93.335000 ;
        RECT 53.690000  93.335000 74.290000  93.485000 ;
        RECT 53.840000  93.485000 74.290000  93.635000 ;
        RECT 53.990000  93.635000 74.290000  93.785000 ;
        RECT 54.140000  93.785000 74.290000  93.935000 ;
        RECT 54.290000  93.935000 74.290000  94.085000 ;
        RECT 54.440000  94.085000 74.290000  94.235000 ;
        RECT 54.590000  94.235000 74.290000  94.385000 ;
        RECT 54.740000  94.385000 74.290000  94.535000 ;
        RECT 54.890000  94.535000 74.290000  94.685000 ;
        RECT 55.040000  94.685000 74.290000  94.835000 ;
        RECT 55.190000  94.835000 74.290000  94.985000 ;
        RECT 55.340000  94.985000 74.290000  95.135000 ;
        RECT 55.490000  95.135000 74.290000  95.285000 ;
        RECT 55.640000  95.285000 74.290000  95.435000 ;
        RECT 55.790000  95.435000 74.290000  95.585000 ;
        RECT 55.940000  95.585000 74.290000  95.735000 ;
        RECT 56.090000  95.735000 74.290000  95.885000 ;
        RECT 56.240000  95.885000 74.290000  96.035000 ;
        RECT 56.390000  96.035000 74.290000  96.185000 ;
        RECT 56.540000  96.185000 74.290000  96.335000 ;
        RECT 56.690000  96.335000 74.290000  96.485000 ;
        RECT 56.840000  96.485000 74.290000  96.635000 ;
        RECT 56.990000  96.635000 74.290000  96.785000 ;
        RECT 57.140000  96.785000 74.290000  96.935000 ;
        RECT 57.290000  96.935000 74.290000  97.085000 ;
        RECT 57.440000  97.085000 74.290000  97.235000 ;
        RECT 57.590000  97.235000 74.290000  97.385000 ;
        RECT 57.740000  97.385000 74.290000  97.535000 ;
        RECT 57.890000  97.535000 74.290000  97.685000 ;
        RECT 58.040000  97.685000 74.290000  97.835000 ;
        RECT 58.190000  97.835000 74.290000  97.985000 ;
        RECT 58.340000  97.985000 74.290000  98.135000 ;
        RECT 58.490000  98.135000 74.290000  98.285000 ;
        RECT 58.640000  98.285000 74.290000  98.435000 ;
        RECT 58.790000  98.435000 74.290000  98.585000 ;
        RECT 58.940000  98.585000 74.290000  98.735000 ;
        RECT 59.090000  98.735000 74.290000  98.885000 ;
        RECT 59.240000  98.885000 74.290000  99.035000 ;
        RECT 59.390000  99.035000 74.290000  99.185000 ;
        RECT 59.540000  99.185000 74.290000  99.335000 ;
        RECT 59.690000  99.335000 74.290000  99.485000 ;
        RECT 59.840000  99.485000 74.290000  99.635000 ;
        RECT 59.990000  99.635000 74.290000  99.785000 ;
        RECT 60.140000  99.785000 74.290000  99.935000 ;
        RECT 60.290000  99.935000 74.290000 100.085000 ;
        RECT 60.440000 100.085000 74.290000 100.235000 ;
        RECT 60.590000 100.235000 74.290000 100.385000 ;
        RECT 60.740000 100.385000 74.290000 100.535000 ;
        RECT 60.890000 100.535000 74.290000 100.685000 ;
        RECT 61.040000 100.685000 74.290000 100.835000 ;
        RECT 61.190000 100.835000 74.290000 100.985000 ;
        RECT 61.340000 100.985000 74.290000 101.135000 ;
        RECT 61.490000 101.135000 74.290000 101.285000 ;
        RECT 61.500000 101.285000 74.290000 101.295000 ;
        RECT 61.500000 101.295000 74.290000 173.320000 ;
    END
  END G_CORE
  PIN OGC_HVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 25.895000 0.000000 27.895000 0.535000 ;
    END
  END OGC_HVC
  PIN SRC_BDY_HVC
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT  0.495000   0.000000 24.395000   2.055000 ;
        RECT  0.565000   2.055000 24.395000   2.125000 ;
        RECT  0.635000   2.125000 24.395000   2.195000 ;
        RECT  0.705000   2.195000 24.395000   2.265000 ;
        RECT  0.775000   2.265000 24.395000   2.335000 ;
        RECT  0.845000   2.335000 24.395000   2.405000 ;
        RECT  0.915000   2.405000 24.395000   2.475000 ;
        RECT  0.985000   2.475000 24.395000   2.545000 ;
        RECT  1.005000   2.545000 24.395000   2.565000 ;
        RECT  1.005000   2.565000 24.395000   8.595000 ;
        RECT  1.005000   8.595000 24.395000   8.665000 ;
        RECT  1.005000   8.665000 24.465000   8.735000 ;
        RECT  1.005000   8.735000 24.535000   8.805000 ;
        RECT  1.005000   8.805000 24.605000   8.875000 ;
        RECT  1.005000   8.875000 24.675000   8.945000 ;
        RECT  1.005000   8.945000 24.745000   9.015000 ;
        RECT  1.005000   9.015000 24.815000   9.085000 ;
        RECT  1.005000   9.085000 24.885000   9.155000 ;
        RECT  1.005000   9.155000 24.955000   9.225000 ;
        RECT  1.005000   9.225000 25.025000   9.295000 ;
        RECT  1.005000   9.295000 25.095000   9.365000 ;
        RECT  1.005000   9.365000 25.165000   9.435000 ;
        RECT  1.005000   9.435000 25.235000   9.505000 ;
        RECT  1.005000   9.505000 25.305000   9.575000 ;
        RECT  1.005000   9.575000 25.375000   9.645000 ;
        RECT  1.005000   9.645000 25.445000   9.715000 ;
        RECT  1.005000   9.715000 25.515000   9.785000 ;
        RECT  1.005000   9.785000 25.585000   9.855000 ;
        RECT  1.005000   9.855000 25.655000   9.925000 ;
        RECT  1.005000   9.925000 25.725000   9.995000 ;
        RECT  1.005000   9.995000 25.795000  10.065000 ;
        RECT  1.005000  10.065000 25.865000  10.135000 ;
        RECT  1.005000  10.135000 25.935000  10.205000 ;
        RECT  1.005000  10.205000 26.005000  10.275000 ;
        RECT  1.005000  10.275000 26.075000  10.345000 ;
        RECT  1.005000  10.345000 26.145000  10.415000 ;
        RECT  1.005000  10.415000 26.215000  10.485000 ;
        RECT  1.005000  10.485000 26.285000  10.555000 ;
        RECT  1.005000  10.555000 26.355000  10.625000 ;
        RECT  1.005000  10.625000 26.425000  10.695000 ;
        RECT  1.005000  10.695000 26.495000  10.765000 ;
        RECT  1.005000  10.765000 26.565000  10.835000 ;
        RECT  1.005000  10.835000 26.635000  10.905000 ;
        RECT  1.005000  10.905000 26.705000  10.975000 ;
        RECT  1.005000  10.975000 26.775000  11.045000 ;
        RECT  1.005000  11.045000 26.845000  11.115000 ;
        RECT  1.005000  11.115000 26.915000  11.185000 ;
        RECT  1.005000  11.185000 26.985000  11.255000 ;
        RECT  1.005000  11.255000 27.055000  11.325000 ;
        RECT  1.005000  11.325000 27.125000  11.395000 ;
        RECT  1.005000  11.395000 27.195000  11.465000 ;
        RECT  1.005000  11.465000 27.265000  11.535000 ;
        RECT  1.005000  11.535000 27.335000  11.605000 ;
        RECT  1.005000  11.605000 27.405000  11.675000 ;
        RECT  1.005000  11.675000 27.475000  11.745000 ;
        RECT  1.005000  11.745000 27.545000  11.815000 ;
        RECT  1.005000  11.815000 27.615000  11.885000 ;
        RECT  1.005000  11.885000 27.685000  11.955000 ;
        RECT  1.005000  11.955000 27.755000  12.025000 ;
        RECT  1.005000  12.025000 27.825000  12.095000 ;
        RECT  1.005000  12.095000 27.895000  12.165000 ;
        RECT  1.005000  12.165000 27.965000  12.235000 ;
        RECT  1.005000  12.235000 28.035000  12.305000 ;
        RECT  1.005000  12.305000 28.105000  12.375000 ;
        RECT  1.005000  12.375000 28.175000  12.400000 ;
        RECT  1.005000  12.400000 36.895000  25.700000 ;
        RECT  1.005000  25.700000 18.750000  25.770000 ;
        RECT  1.005000  25.770000 18.680000  25.840000 ;
        RECT  1.005000  25.840000 18.610000  25.910000 ;
        RECT  1.005000  25.910000 18.540000  25.980000 ;
        RECT  1.005000  25.980000 18.470000  26.050000 ;
        RECT  1.005000  26.050000 18.400000  26.120000 ;
        RECT  1.005000  26.120000 18.330000  26.190000 ;
        RECT  1.005000  26.190000 18.260000  26.260000 ;
        RECT  1.005000  26.260000 18.190000  26.330000 ;
        RECT  1.005000  26.330000 18.120000  26.400000 ;
        RECT  1.005000  26.400000 18.050000  26.470000 ;
        RECT  1.005000  26.470000 17.980000  26.540000 ;
        RECT  1.005000  26.540000 17.910000  26.610000 ;
        RECT  1.005000  26.610000 17.840000  26.680000 ;
        RECT  1.005000  26.680000 17.770000  26.750000 ;
        RECT  1.005000  26.750000 17.700000  26.820000 ;
        RECT  1.005000  26.820000 17.630000  26.890000 ;
        RECT  1.005000  26.890000 17.560000  26.960000 ;
        RECT  1.005000  26.960000 17.490000  27.030000 ;
        RECT  1.005000  27.030000 17.420000  27.100000 ;
        RECT  1.005000  27.100000 17.350000  27.170000 ;
        RECT  1.005000  27.170000 17.280000  27.240000 ;
        RECT  1.005000  27.240000 17.210000  27.310000 ;
        RECT  1.005000  27.310000 17.140000  27.380000 ;
        RECT  1.005000  27.380000 17.070000  27.450000 ;
        RECT  1.005000  27.450000 17.000000  27.520000 ;
        RECT  1.005000  27.520000 16.930000  27.590000 ;
        RECT  1.005000  27.590000 16.860000  27.660000 ;
        RECT  1.005000  27.660000 16.790000  27.730000 ;
        RECT  1.005000  27.730000 16.720000  27.800000 ;
        RECT  1.005000  27.800000 16.650000  27.870000 ;
        RECT  1.005000  27.870000 16.580000  27.940000 ;
        RECT  1.005000  27.940000 16.510000  28.010000 ;
        RECT  1.005000  28.010000 16.440000  28.080000 ;
        RECT  1.005000  28.080000 16.370000  28.150000 ;
        RECT  1.005000  28.150000 16.300000  28.220000 ;
        RECT  1.005000  28.220000 16.230000  28.290000 ;
        RECT  1.005000  28.290000 16.160000  28.360000 ;
        RECT  1.005000  28.360000 16.090000  28.430000 ;
        RECT  1.005000  28.430000 16.020000  28.500000 ;
        RECT  1.005000  28.500000 15.950000  28.570000 ;
        RECT  1.005000  28.570000 15.880000  28.640000 ;
        RECT  1.005000  28.640000 15.810000  28.710000 ;
        RECT  1.005000  28.710000 15.740000  28.780000 ;
        RECT  1.005000  28.780000 15.670000  28.850000 ;
        RECT  1.005000  28.850000 15.600000  28.920000 ;
        RECT  1.005000  28.920000 15.530000  28.990000 ;
        RECT  1.005000  28.990000 15.460000  29.060000 ;
        RECT  1.005000  29.060000 15.390000  29.130000 ;
        RECT  1.005000  29.130000 15.320000  29.200000 ;
        RECT  1.005000  29.200000 15.250000  29.270000 ;
        RECT  1.005000  29.270000 15.205000  29.315000 ;
        RECT  1.005000  29.315000 15.205000  35.665000 ;
        RECT  1.005000  35.665000 15.205000  35.735000 ;
        RECT  1.005000  35.735000 15.275000  35.805000 ;
        RECT  1.005000  35.805000 15.345000  35.875000 ;
        RECT  1.005000  35.875000 15.415000  35.945000 ;
        RECT  1.005000  35.945000 15.485000  36.015000 ;
        RECT  1.005000  36.015000 15.555000  36.085000 ;
        RECT  1.005000  36.085000 15.625000  36.155000 ;
        RECT  1.005000  36.155000 15.695000  36.225000 ;
        RECT  1.005000  36.225000 15.765000  36.295000 ;
        RECT  1.005000  36.295000 15.835000  36.365000 ;
        RECT  1.005000  36.365000 15.905000  36.435000 ;
        RECT  1.005000  36.435000 15.975000  36.505000 ;
        RECT  1.005000  36.505000 16.045000  36.575000 ;
        RECT  1.005000  36.575000 16.115000  36.640000 ;
        RECT  1.005000  47.130000 14.120000  54.215000 ;
        RECT  1.005000  54.215000 14.120000  54.285000 ;
        RECT  1.005000  54.285000 14.190000  54.355000 ;
        RECT  1.005000  54.355000 14.260000  54.425000 ;
        RECT  1.005000  54.425000 14.330000  54.495000 ;
        RECT  1.005000  54.495000 14.400000  54.565000 ;
        RECT  1.005000  54.565000 14.470000  54.635000 ;
        RECT  1.005000  54.635000 14.540000  54.705000 ;
        RECT  1.005000  54.705000 14.610000  54.775000 ;
        RECT  1.005000  54.775000 14.680000  54.845000 ;
        RECT  1.005000  54.845000 14.750000  54.915000 ;
        RECT  1.005000  54.915000 14.820000  54.985000 ;
        RECT  1.005000  54.985000 14.890000  55.055000 ;
        RECT  1.005000  55.055000 14.960000  55.125000 ;
        RECT  1.005000  55.125000 15.030000  55.195000 ;
        RECT  1.005000  55.195000 15.100000  55.265000 ;
        RECT  1.005000  55.265000 15.170000  55.335000 ;
        RECT  1.005000  55.335000 15.240000  55.405000 ;
        RECT  1.005000  55.405000 15.310000  55.475000 ;
        RECT  1.005000  55.475000 15.380000  55.545000 ;
        RECT  1.005000  55.545000 15.450000  55.615000 ;
        RECT  1.005000  55.615000 15.520000  55.685000 ;
        RECT  1.005000  55.685000 15.590000  55.755000 ;
        RECT  1.005000  55.755000 15.660000  55.825000 ;
        RECT  1.005000  55.825000 15.730000  55.895000 ;
        RECT  1.005000  55.895000 15.800000  55.965000 ;
        RECT  1.005000  55.965000 15.870000  56.035000 ;
        RECT  1.005000  56.035000 15.940000  56.105000 ;
        RECT  1.005000  56.105000 16.010000  56.175000 ;
        RECT  1.005000  56.175000 16.080000  56.245000 ;
        RECT  1.005000  56.245000 16.150000  56.315000 ;
        RECT  1.005000  56.315000 16.220000  56.385000 ;
        RECT  1.005000  56.385000 16.290000  56.455000 ;
        RECT  1.005000  56.455000 16.360000  56.525000 ;
        RECT  1.005000  56.525000 16.430000  56.595000 ;
        RECT  1.005000  56.595000 16.500000  56.665000 ;
        RECT  1.005000  56.665000 16.570000  56.735000 ;
        RECT  1.005000  56.735000 16.640000  56.805000 ;
        RECT  1.005000  56.805000 16.710000  56.875000 ;
        RECT  1.005000  56.875000 16.780000  56.945000 ;
        RECT  1.005000  56.945000 16.850000  57.015000 ;
        RECT  1.005000  57.015000 16.920000  57.085000 ;
        RECT  1.005000  57.085000 16.990000  57.155000 ;
        RECT  1.005000  57.155000 17.060000  57.225000 ;
        RECT  1.005000  57.225000 17.130000  57.295000 ;
        RECT  1.005000  57.295000 17.200000  57.365000 ;
        RECT  1.005000  57.365000 17.270000  57.435000 ;
        RECT  1.005000  57.435000 17.340000  57.505000 ;
        RECT  1.005000  57.505000 17.410000  57.575000 ;
        RECT  1.005000  57.575000 17.480000  57.645000 ;
        RECT  1.005000  57.645000 17.550000  57.715000 ;
        RECT  1.005000  57.715000 17.620000  57.780000 ;
        RECT  1.005000  57.780000 56.710000  66.480000 ;
        RECT  1.005000  66.480000 17.595000  66.550000 ;
        RECT  1.005000  66.550000 17.525000  66.620000 ;
        RECT  1.005000  66.620000 17.455000  66.690000 ;
        RECT  1.005000  66.690000 17.385000  66.760000 ;
        RECT  1.005000  66.760000 17.315000  66.830000 ;
        RECT  1.005000  66.830000 17.245000  66.900000 ;
        RECT  1.005000  66.900000 17.175000  66.970000 ;
        RECT  1.005000  66.970000 17.105000  67.040000 ;
        RECT  1.005000  67.040000 17.035000  67.110000 ;
        RECT  1.005000  67.110000 16.965000  67.180000 ;
        RECT  1.005000  67.180000 16.895000  67.250000 ;
        RECT  1.005000  67.250000 16.825000  67.320000 ;
        RECT  1.005000  67.320000 16.755000  67.390000 ;
        RECT  1.005000  67.390000 16.685000  67.460000 ;
        RECT  1.005000  67.460000 16.615000  67.530000 ;
        RECT  1.005000  67.530000 16.545000  67.600000 ;
        RECT  1.005000  67.600000 16.475000  67.670000 ;
        RECT  1.005000  67.670000 16.405000  67.740000 ;
        RECT  1.005000  67.740000 16.335000  67.810000 ;
        RECT  1.005000  67.810000 16.265000  67.880000 ;
        RECT  1.005000  67.880000 16.195000  67.950000 ;
        RECT  1.005000  67.950000 16.125000  68.020000 ;
        RECT  1.005000  68.020000 16.055000  68.090000 ;
        RECT  1.005000  68.090000 15.985000  68.160000 ;
        RECT  1.005000  68.160000 15.915000  68.230000 ;
        RECT  1.005000  68.230000 15.845000  68.300000 ;
        RECT  1.005000  68.300000 15.775000  68.370000 ;
        RECT  1.005000  68.370000 15.705000  68.440000 ;
        RECT  1.005000  68.440000 15.635000  68.510000 ;
        RECT  1.005000  68.510000 15.565000  68.580000 ;
        RECT  1.005000  68.580000 15.495000  68.650000 ;
        RECT  1.005000  68.650000 15.425000  68.720000 ;
        RECT  1.005000  68.720000 15.355000  68.790000 ;
        RECT  1.005000  68.790000 15.285000  68.860000 ;
        RECT  1.005000  68.860000 15.215000  68.930000 ;
        RECT  1.005000  68.930000 15.145000  69.000000 ;
        RECT  1.005000  69.000000 15.075000  69.070000 ;
        RECT  1.005000  69.070000 15.005000  69.140000 ;
        RECT  1.005000  69.140000 14.935000  69.210000 ;
        RECT  1.005000  69.210000 14.865000  69.280000 ;
        RECT  1.005000  69.280000 14.795000  69.350000 ;
        RECT  1.005000  69.350000 14.725000  69.420000 ;
        RECT  1.005000  69.420000 14.655000  69.490000 ;
        RECT  1.005000  69.490000 14.585000  69.560000 ;
        RECT  1.005000  69.560000 14.515000  69.630000 ;
        RECT  1.005000  69.630000 14.445000  69.700000 ;
        RECT  1.005000  69.700000 14.375000  69.770000 ;
        RECT  1.005000  69.770000 14.305000  69.840000 ;
        RECT  1.005000  69.840000 14.235000  69.910000 ;
        RECT  1.005000  69.910000 14.165000  69.980000 ;
        RECT  1.005000  69.980000 14.120000  70.025000 ;
        RECT  1.005000  70.025000 14.120000  77.240000 ;
        RECT  1.005000  77.240000 14.120000  77.310000 ;
        RECT  1.005000  77.310000 14.190000  77.380000 ;
        RECT  1.005000  77.380000 14.260000  77.450000 ;
        RECT  1.005000  77.450000 14.330000  77.520000 ;
        RECT  1.005000  77.520000 14.400000  77.590000 ;
        RECT  1.005000  77.590000 14.470000  77.660000 ;
        RECT  1.005000  77.660000 14.540000  77.730000 ;
        RECT  1.005000  77.730000 14.610000  77.800000 ;
        RECT  1.005000  77.800000 14.680000  77.870000 ;
        RECT  1.005000  77.870000 14.750000  77.940000 ;
        RECT  1.005000  77.940000 14.820000  78.010000 ;
        RECT  1.005000  78.010000 14.890000  78.080000 ;
        RECT  1.005000  78.080000 14.960000  78.150000 ;
        RECT  1.005000  78.150000 15.030000  78.220000 ;
        RECT  1.005000  78.220000 15.100000  78.290000 ;
        RECT  1.005000  78.290000 15.170000  78.360000 ;
        RECT  1.005000  78.360000 15.240000  78.430000 ;
        RECT  1.005000  78.430000 15.310000  78.500000 ;
        RECT  1.005000  78.500000 15.380000  78.570000 ;
        RECT  1.005000  78.570000 15.450000  78.640000 ;
        RECT  1.005000  78.640000 15.520000  78.710000 ;
        RECT  1.005000  78.710000 15.590000  78.780000 ;
        RECT  1.005000  78.780000 15.660000  78.850000 ;
        RECT  1.005000  78.850000 15.730000  78.920000 ;
        RECT  1.005000  78.920000 15.800000  78.990000 ;
        RECT  1.005000  78.990000 15.870000  79.060000 ;
        RECT  1.005000  79.060000 15.940000  79.130000 ;
        RECT  1.005000  79.130000 16.010000  79.200000 ;
        RECT  1.005000  79.200000 16.080000  79.270000 ;
        RECT  1.005000  79.270000 16.150000  79.340000 ;
        RECT  1.005000  79.340000 16.220000  79.410000 ;
        RECT  1.005000  79.410000 16.290000  79.480000 ;
        RECT  1.005000  79.480000 16.360000  79.550000 ;
        RECT  1.005000  79.550000 16.430000  79.620000 ;
        RECT  1.005000  79.620000 16.500000  79.690000 ;
        RECT  1.005000  79.690000 16.570000  79.760000 ;
        RECT  1.005000  79.760000 16.640000  79.830000 ;
        RECT  1.005000  79.830000 16.710000  79.900000 ;
        RECT  1.005000  79.900000 16.780000  79.970000 ;
        RECT  1.005000  79.970000 16.850000  80.040000 ;
        RECT  1.005000  80.040000 16.920000  80.110000 ;
        RECT  1.005000  80.110000 16.990000  80.180000 ;
        RECT  1.005000  80.180000 17.060000  80.250000 ;
        RECT  1.005000  80.250000 17.130000  80.320000 ;
        RECT  1.005000  80.320000 17.200000  80.390000 ;
        RECT  1.005000  80.390000 17.270000  80.460000 ;
        RECT  1.005000  80.460000 17.340000  80.530000 ;
        RECT  1.005000  80.530000 17.410000  80.600000 ;
        RECT  1.005000  80.600000 17.480000  80.670000 ;
        RECT  1.005000  80.670000 17.550000  80.740000 ;
        RECT  1.005000  80.740000 17.620000  80.780000 ;
        RECT  1.005000  80.780000 56.705000  89.480000 ;
        RECT  1.005000  89.480000 17.595000  89.550000 ;
        RECT  1.005000  89.550000 17.525000  89.620000 ;
        RECT  1.005000  89.620000 17.455000  89.690000 ;
        RECT  1.005000  89.690000 17.385000  89.760000 ;
        RECT  1.005000  89.760000 17.315000  89.830000 ;
        RECT  1.005000  89.830000 17.245000  89.900000 ;
        RECT  1.005000  89.900000 17.175000  89.970000 ;
        RECT  1.005000  89.970000 17.105000  90.040000 ;
        RECT  1.005000  90.040000 17.035000  90.110000 ;
        RECT  1.005000  90.110000 16.965000  90.180000 ;
        RECT  1.005000  90.180000 16.895000  90.250000 ;
        RECT  1.005000  90.250000 16.825000  90.320000 ;
        RECT  1.005000  90.320000 16.755000  90.390000 ;
        RECT  1.005000  90.390000 16.685000  90.460000 ;
        RECT  1.005000  90.460000 16.615000  90.530000 ;
        RECT  1.005000  90.530000 16.545000  90.600000 ;
        RECT  1.005000  90.600000 16.475000  90.670000 ;
        RECT  1.005000  90.670000 16.405000  90.740000 ;
        RECT  1.005000  90.740000 16.335000  90.810000 ;
        RECT  1.005000  90.810000 16.265000  90.880000 ;
        RECT  1.005000  90.880000 16.195000  90.950000 ;
        RECT  1.005000  90.950000 16.125000  91.020000 ;
        RECT  1.005000  91.020000 16.055000  91.090000 ;
        RECT  1.005000  91.090000 15.985000  91.160000 ;
        RECT  1.005000  91.160000 15.915000  91.230000 ;
        RECT  1.005000  91.230000 15.845000  91.300000 ;
        RECT  1.005000  91.300000 15.775000  91.370000 ;
        RECT  1.005000  91.370000 15.705000  91.440000 ;
        RECT  1.005000  91.440000 15.635000  91.510000 ;
        RECT  1.005000  91.510000 15.565000  91.580000 ;
        RECT  1.005000  91.580000 15.495000  91.650000 ;
        RECT  1.005000  91.650000 15.425000  91.720000 ;
        RECT  1.005000  91.720000 15.355000  91.790000 ;
        RECT  1.005000  91.790000 15.285000  91.860000 ;
        RECT  1.005000  91.860000 15.215000  91.930000 ;
        RECT  1.005000  91.930000 15.145000  92.000000 ;
        RECT  1.005000  92.000000 15.075000  92.070000 ;
        RECT  1.005000  92.070000 15.005000  92.140000 ;
        RECT  1.005000  92.140000 14.935000  92.210000 ;
        RECT  1.005000  92.210000 14.865000  92.280000 ;
        RECT  1.005000  92.280000 14.795000  92.350000 ;
        RECT  1.005000  92.350000 14.725000  92.420000 ;
        RECT  1.005000  92.420000 14.655000  92.490000 ;
        RECT  1.005000  92.490000 14.585000  92.560000 ;
        RECT  1.005000  92.560000 14.515000  92.630000 ;
        RECT  1.005000  92.630000 14.445000  92.700000 ;
        RECT  1.005000  92.700000 14.375000  92.770000 ;
        RECT  1.005000  92.770000 14.305000  92.840000 ;
        RECT  1.005000  92.840000 14.235000  92.910000 ;
        RECT  1.005000  92.910000 14.165000  92.980000 ;
        RECT  1.005000  92.980000 14.120000  93.025000 ;
        RECT  1.005000  93.025000 14.120000 100.240000 ;
        RECT  1.005000 100.240000 14.120000 100.310000 ;
        RECT  1.005000 100.310000 14.190000 100.380000 ;
        RECT  1.005000 100.380000 14.260000 100.450000 ;
        RECT  1.005000 100.450000 14.330000 100.520000 ;
        RECT  1.005000 100.520000 14.400000 100.590000 ;
        RECT  1.005000 100.590000 14.470000 100.660000 ;
        RECT  1.005000 100.660000 14.540000 100.730000 ;
        RECT  1.005000 100.730000 14.610000 100.800000 ;
        RECT  1.005000 100.800000 14.680000 100.870000 ;
        RECT  1.005000 100.870000 14.750000 100.940000 ;
        RECT  1.005000 100.940000 14.820000 101.010000 ;
        RECT  1.005000 101.010000 14.890000 101.080000 ;
        RECT  1.005000 101.080000 14.960000 101.150000 ;
        RECT  1.005000 101.150000 15.030000 101.220000 ;
        RECT  1.005000 101.220000 15.100000 101.290000 ;
        RECT  1.005000 101.290000 15.170000 101.360000 ;
        RECT  1.005000 101.360000 15.240000 101.430000 ;
        RECT  1.005000 101.430000 15.310000 101.500000 ;
        RECT  1.005000 101.500000 15.380000 101.570000 ;
        RECT  1.005000 101.570000 15.450000 101.640000 ;
        RECT  1.005000 101.640000 15.520000 101.710000 ;
        RECT  1.005000 101.710000 15.590000 101.780000 ;
        RECT  1.005000 101.780000 15.660000 101.850000 ;
        RECT  1.005000 101.850000 15.730000 101.920000 ;
        RECT  1.005000 101.920000 15.800000 101.990000 ;
        RECT  1.005000 101.990000 15.870000 102.060000 ;
        RECT  1.005000 102.060000 15.940000 102.130000 ;
        RECT  1.005000 102.130000 16.010000 102.200000 ;
        RECT  1.005000 102.200000 16.080000 102.270000 ;
        RECT  1.005000 102.270000 16.150000 102.340000 ;
        RECT  1.005000 102.340000 16.220000 102.410000 ;
        RECT  1.005000 102.410000 16.290000 102.480000 ;
        RECT  1.005000 102.480000 16.360000 102.550000 ;
        RECT  1.005000 102.550000 16.430000 102.620000 ;
        RECT  1.005000 102.620000 16.500000 102.690000 ;
        RECT  1.005000 102.690000 16.570000 102.760000 ;
        RECT  1.005000 102.760000 16.640000 102.830000 ;
        RECT  1.005000 102.830000 16.710000 102.900000 ;
        RECT  1.005000 102.900000 16.780000 102.970000 ;
        RECT  1.005000 102.970000 16.850000 103.040000 ;
        RECT  1.005000 103.040000 16.920000 103.110000 ;
        RECT  1.005000 103.110000 16.990000 103.180000 ;
        RECT  1.005000 103.180000 17.060000 103.250000 ;
        RECT  1.005000 103.250000 17.130000 103.320000 ;
        RECT  1.005000 103.320000 17.200000 103.390000 ;
        RECT  1.005000 103.390000 17.270000 103.460000 ;
        RECT  1.005000 103.460000 17.340000 103.530000 ;
        RECT  1.005000 103.530000 17.410000 103.600000 ;
        RECT  1.005000 103.600000 17.480000 103.670000 ;
        RECT  1.005000 103.670000 17.550000 103.740000 ;
        RECT  1.005000 103.740000 17.620000 103.780000 ;
        RECT  1.005000 103.780000 56.705000 112.480000 ;
        RECT  1.005000 112.480000 17.635000 112.550000 ;
        RECT  1.005000 112.550000 17.565000 112.620000 ;
        RECT  1.005000 112.620000 17.495000 112.690000 ;
        RECT  1.005000 112.690000 17.425000 112.760000 ;
        RECT  1.005000 112.760000 17.355000 112.830000 ;
        RECT  1.005000 112.830000 17.285000 112.900000 ;
        RECT  1.005000 112.900000 17.215000 112.970000 ;
        RECT  1.005000 112.970000 17.145000 113.040000 ;
        RECT  1.005000 113.040000 17.075000 113.110000 ;
        RECT  1.005000 113.110000 17.005000 113.180000 ;
        RECT  1.005000 113.180000 16.935000 113.250000 ;
        RECT  1.005000 113.250000 16.865000 113.320000 ;
        RECT  1.005000 113.320000 16.795000 113.390000 ;
        RECT  1.005000 113.390000 16.725000 113.460000 ;
        RECT  1.005000 113.460000 16.655000 113.530000 ;
        RECT  1.005000 113.530000 16.585000 113.600000 ;
        RECT  1.005000 113.600000 16.515000 113.670000 ;
        RECT  1.005000 113.670000 16.445000 113.740000 ;
        RECT  1.005000 113.740000 16.375000 113.810000 ;
        RECT  1.005000 113.810000 16.305000 113.880000 ;
        RECT  1.005000 113.880000 16.235000 113.950000 ;
        RECT  1.005000 113.950000 16.165000 114.020000 ;
        RECT  1.005000 114.020000 16.095000 114.090000 ;
        RECT  1.005000 114.090000 16.025000 114.160000 ;
        RECT  1.005000 114.160000 15.955000 114.230000 ;
        RECT  1.005000 114.230000 15.885000 114.300000 ;
        RECT  1.005000 114.300000 15.815000 114.370000 ;
        RECT  1.005000 114.370000 15.745000 114.440000 ;
        RECT  1.005000 114.440000 15.675000 114.510000 ;
        RECT  1.005000 114.510000 15.605000 114.580000 ;
        RECT  1.005000 114.580000 15.535000 114.650000 ;
        RECT  1.005000 114.650000 15.465000 114.720000 ;
        RECT  1.005000 114.720000 15.395000 114.790000 ;
        RECT  1.005000 114.790000 15.325000 114.860000 ;
        RECT  1.005000 114.860000 15.255000 114.930000 ;
        RECT  1.005000 114.930000 15.185000 115.000000 ;
        RECT  1.005000 115.000000 15.115000 115.070000 ;
        RECT  1.005000 115.070000 15.045000 115.140000 ;
        RECT  1.005000 115.140000 14.975000 115.210000 ;
        RECT  1.005000 115.210000 14.905000 115.280000 ;
        RECT  1.005000 115.280000 14.835000 115.350000 ;
        RECT  1.005000 115.350000 14.765000 115.420000 ;
        RECT  1.005000 115.420000 14.695000 115.490000 ;
        RECT  1.005000 115.490000 14.625000 115.560000 ;
        RECT  1.005000 115.560000 14.555000 115.630000 ;
        RECT  1.005000 115.630000 14.485000 115.700000 ;
        RECT  1.005000 115.700000 14.415000 115.770000 ;
        RECT  1.005000 115.770000 14.345000 115.840000 ;
        RECT  1.005000 115.840000 14.275000 115.910000 ;
        RECT  1.005000 115.910000 14.205000 115.980000 ;
        RECT  1.005000 115.980000 14.135000 116.050000 ;
        RECT  1.005000 116.050000 14.120000 116.065000 ;
        RECT  1.005000 116.065000 14.120000 123.145000 ;
        RECT  1.005000 123.145000 14.120000 123.215000 ;
        RECT  1.005000 123.215000 14.190000 123.285000 ;
        RECT  1.005000 123.285000 14.260000 123.355000 ;
        RECT  1.005000 123.355000 14.330000 123.425000 ;
        RECT  1.005000 123.425000 14.400000 123.495000 ;
        RECT  1.005000 123.495000 14.470000 123.565000 ;
        RECT  1.005000 123.565000 14.540000 123.635000 ;
        RECT  1.005000 123.635000 14.610000 123.705000 ;
        RECT  1.005000 123.705000 14.680000 123.775000 ;
        RECT  1.005000 123.775000 14.750000 123.845000 ;
        RECT  1.005000 123.845000 14.820000 123.915000 ;
        RECT  1.005000 123.915000 14.890000 123.985000 ;
        RECT  1.005000 123.985000 14.960000 124.055000 ;
        RECT  1.005000 124.055000 15.030000 124.125000 ;
        RECT  1.005000 124.125000 15.100000 124.195000 ;
        RECT  1.005000 124.195000 15.170000 124.265000 ;
        RECT  1.005000 124.265000 15.240000 124.335000 ;
        RECT  1.005000 124.335000 15.310000 124.405000 ;
        RECT  1.005000 124.405000 15.380000 124.475000 ;
        RECT  1.005000 124.475000 15.450000 124.545000 ;
        RECT  1.005000 124.545000 15.520000 124.615000 ;
        RECT  1.005000 124.615000 15.590000 124.685000 ;
        RECT  1.005000 124.685000 15.660000 124.755000 ;
        RECT  1.005000 124.755000 15.730000 124.825000 ;
        RECT  1.005000 124.825000 15.800000 124.895000 ;
        RECT  1.005000 124.895000 15.870000 124.965000 ;
        RECT  1.005000 124.965000 15.940000 125.035000 ;
        RECT  1.005000 125.035000 16.010000 125.105000 ;
        RECT  1.005000 125.105000 16.080000 125.175000 ;
        RECT  1.005000 125.175000 16.150000 125.245000 ;
        RECT  1.005000 125.245000 16.220000 125.315000 ;
        RECT  1.005000 125.315000 16.290000 125.385000 ;
        RECT  1.005000 125.385000 16.360000 125.455000 ;
        RECT  1.005000 125.455000 16.430000 125.525000 ;
        RECT  1.005000 125.525000 16.500000 125.595000 ;
        RECT  1.005000 125.595000 16.570000 125.665000 ;
        RECT  1.005000 125.665000 16.640000 125.735000 ;
        RECT  1.005000 125.735000 16.710000 125.805000 ;
        RECT  1.005000 125.805000 16.780000 125.875000 ;
        RECT  1.005000 125.875000 16.850000 125.945000 ;
        RECT  1.005000 125.945000 16.920000 126.015000 ;
        RECT  1.005000 126.015000 16.990000 126.085000 ;
        RECT  1.005000 126.085000 17.060000 126.155000 ;
        RECT  1.005000 126.155000 17.130000 126.225000 ;
        RECT  1.005000 126.225000 17.200000 126.295000 ;
        RECT  1.005000 126.295000 17.270000 126.365000 ;
        RECT  1.005000 126.365000 17.340000 126.435000 ;
        RECT  1.005000 126.435000 17.410000 126.505000 ;
        RECT  1.005000 126.505000 17.480000 126.575000 ;
        RECT  1.005000 126.575000 17.550000 126.645000 ;
        RECT  1.005000 126.645000 17.620000 126.715000 ;
        RECT  1.005000 126.715000 17.690000 126.780000 ;
        RECT  1.005000 126.780000 56.705000 135.480000 ;
        RECT  1.005000 135.480000 17.740000 135.550000 ;
        RECT  1.005000 135.550000 17.670000 135.620000 ;
        RECT  1.005000 135.620000 17.600000 135.690000 ;
        RECT  1.005000 135.690000 17.530000 135.760000 ;
        RECT  1.005000 135.760000 17.460000 135.830000 ;
        RECT  1.005000 135.830000 17.390000 135.900000 ;
        RECT  1.005000 135.900000 17.320000 135.970000 ;
        RECT  1.005000 135.970000 17.250000 136.040000 ;
        RECT  1.005000 136.040000 17.180000 136.110000 ;
        RECT  1.005000 136.110000 17.110000 136.180000 ;
        RECT  1.005000 136.180000 17.040000 136.250000 ;
        RECT  1.005000 136.250000 16.970000 136.320000 ;
        RECT  1.005000 136.320000 16.900000 136.390000 ;
        RECT  1.005000 136.390000 16.830000 136.460000 ;
        RECT  1.005000 136.460000 16.760000 136.530000 ;
        RECT  1.005000 136.530000 16.690000 136.600000 ;
        RECT  1.005000 136.600000 16.620000 136.670000 ;
        RECT  1.005000 136.670000 16.550000 136.740000 ;
        RECT  1.005000 136.740000 16.480000 136.810000 ;
        RECT  1.005000 136.810000 16.410000 136.880000 ;
        RECT  1.005000 136.880000 16.340000 136.950000 ;
        RECT  1.005000 136.950000 16.270000 137.020000 ;
        RECT  1.005000 137.020000 16.200000 137.090000 ;
        RECT  1.005000 137.090000 16.130000 137.160000 ;
        RECT  1.005000 137.160000 16.060000 137.230000 ;
        RECT  1.005000 137.230000 15.990000 137.300000 ;
        RECT  1.005000 137.300000 15.920000 137.370000 ;
        RECT  1.005000 137.370000 15.850000 137.440000 ;
        RECT  1.005000 137.440000 15.780000 137.510000 ;
        RECT  1.005000 137.510000 15.710000 137.580000 ;
        RECT  1.005000 137.580000 15.640000 137.650000 ;
        RECT  1.005000 137.650000 15.570000 137.720000 ;
        RECT  1.005000 137.720000 15.500000 137.790000 ;
        RECT  1.005000 137.790000 15.430000 137.860000 ;
        RECT  1.005000 137.860000 15.360000 137.930000 ;
        RECT  1.005000 137.930000 15.290000 138.000000 ;
        RECT  1.005000 138.000000 15.220000 138.070000 ;
        RECT  1.005000 138.070000 15.150000 138.140000 ;
        RECT  1.005000 138.140000 15.080000 138.210000 ;
        RECT  1.005000 138.210000 15.010000 138.280000 ;
        RECT  1.005000 138.280000 14.940000 138.350000 ;
        RECT  1.005000 138.350000 14.870000 138.420000 ;
        RECT  1.005000 138.420000 14.800000 138.490000 ;
        RECT  1.005000 138.490000 14.730000 138.560000 ;
        RECT  1.005000 138.560000 14.660000 138.630000 ;
        RECT  1.005000 138.630000 14.590000 138.700000 ;
        RECT  1.005000 138.700000 14.520000 138.770000 ;
        RECT  1.005000 138.770000 14.450000 138.840000 ;
        RECT  1.005000 138.840000 14.380000 138.910000 ;
        RECT  1.005000 138.910000 14.310000 138.980000 ;
        RECT  1.005000 138.980000 14.240000 139.050000 ;
        RECT  1.005000 139.050000 14.170000 139.120000 ;
        RECT  1.005000 139.120000 14.120000 139.170000 ;
        RECT  1.005000 139.170000 14.120000 146.215000 ;
        RECT  1.005000 146.215000 14.120000 146.285000 ;
        RECT  1.005000 146.285000 14.190000 146.355000 ;
        RECT  1.005000 146.355000 14.260000 146.425000 ;
        RECT  1.005000 146.425000 14.330000 146.495000 ;
        RECT  1.005000 146.495000 14.400000 146.565000 ;
        RECT  1.005000 146.565000 14.470000 146.635000 ;
        RECT  1.005000 146.635000 14.540000 146.705000 ;
        RECT  1.005000 146.705000 14.610000 146.775000 ;
        RECT  1.005000 146.775000 14.680000 146.845000 ;
        RECT  1.005000 146.845000 14.750000 146.915000 ;
        RECT  1.005000 146.915000 14.820000 146.985000 ;
        RECT  1.005000 146.985000 14.890000 147.055000 ;
        RECT  1.005000 147.055000 14.960000 147.125000 ;
        RECT  1.005000 147.125000 15.030000 147.195000 ;
        RECT  1.005000 147.195000 15.100000 147.265000 ;
        RECT  1.005000 147.265000 15.170000 147.335000 ;
        RECT  1.005000 147.335000 15.240000 147.405000 ;
        RECT  1.005000 147.405000 15.310000 147.475000 ;
        RECT  1.005000 147.475000 15.380000 147.545000 ;
        RECT  1.005000 147.545000 15.450000 147.615000 ;
        RECT  1.005000 147.615000 15.520000 147.685000 ;
        RECT  1.005000 147.685000 15.590000 147.755000 ;
        RECT  1.005000 147.755000 15.660000 147.825000 ;
        RECT  1.005000 147.825000 15.730000 147.895000 ;
        RECT  1.005000 147.895000 15.800000 147.965000 ;
        RECT  1.005000 147.965000 15.870000 148.035000 ;
        RECT  1.005000 148.035000 15.940000 148.105000 ;
        RECT  1.005000 148.105000 16.010000 148.175000 ;
        RECT  1.005000 148.175000 16.080000 148.245000 ;
        RECT  1.005000 148.245000 16.150000 148.315000 ;
        RECT  1.005000 148.315000 16.220000 148.385000 ;
        RECT  1.005000 148.385000 16.290000 148.455000 ;
        RECT  1.005000 148.455000 16.360000 148.525000 ;
        RECT  1.005000 148.525000 16.430000 148.595000 ;
        RECT  1.005000 148.595000 16.500000 148.665000 ;
        RECT  1.005000 148.665000 16.570000 148.735000 ;
        RECT  1.005000 148.735000 16.640000 148.805000 ;
        RECT  1.005000 148.805000 16.710000 148.875000 ;
        RECT  1.005000 148.875000 16.780000 148.945000 ;
        RECT  1.005000 148.945000 16.850000 149.015000 ;
        RECT  1.005000 149.015000 16.920000 149.085000 ;
        RECT  1.005000 149.085000 16.990000 149.155000 ;
        RECT  1.005000 149.155000 17.060000 149.225000 ;
        RECT  1.005000 149.225000 17.130000 149.295000 ;
        RECT  1.005000 149.295000 17.200000 149.365000 ;
        RECT  1.005000 149.365000 17.270000 149.435000 ;
        RECT  1.005000 149.435000 17.340000 149.505000 ;
        RECT  1.005000 149.505000 17.410000 149.575000 ;
        RECT  1.005000 149.575000 17.480000 149.645000 ;
        RECT  1.005000 149.645000 17.550000 149.715000 ;
        RECT  1.005000 149.715000 17.620000 149.780000 ;
        RECT  1.005000 149.780000 56.705000 158.480000 ;
        RECT  1.005000 158.480000 17.650000 158.550000 ;
        RECT  1.005000 158.550000 17.580000 158.620000 ;
        RECT  1.005000 158.620000 17.510000 158.690000 ;
        RECT  1.005000 158.690000 17.440000 158.760000 ;
        RECT  1.005000 158.760000 17.370000 158.830000 ;
        RECT  1.005000 158.830000 17.300000 158.900000 ;
        RECT  1.005000 158.900000 17.230000 158.970000 ;
        RECT  1.005000 158.970000 17.160000 159.040000 ;
        RECT  1.005000 159.040000 17.090000 159.110000 ;
        RECT  1.005000 159.110000 17.020000 159.180000 ;
        RECT  1.005000 159.180000 16.950000 159.250000 ;
        RECT  1.005000 159.250000 16.880000 159.320000 ;
        RECT  1.005000 159.320000 16.810000 159.390000 ;
        RECT  1.005000 159.390000 16.740000 159.460000 ;
        RECT  1.005000 159.460000 16.670000 159.530000 ;
        RECT  1.005000 159.530000 16.600000 159.600000 ;
        RECT  1.005000 159.600000 16.530000 159.670000 ;
        RECT  1.005000 159.670000 16.460000 159.740000 ;
        RECT  1.005000 159.740000 16.390000 159.810000 ;
        RECT  1.005000 159.810000 16.320000 159.880000 ;
        RECT  1.005000 159.880000 16.250000 159.950000 ;
        RECT  1.005000 159.950000 16.180000 160.020000 ;
        RECT  1.005000 160.020000 16.110000 160.090000 ;
        RECT  1.005000 160.090000 16.040000 160.160000 ;
        RECT  1.005000 160.160000 15.970000 160.230000 ;
        RECT  1.005000 160.230000 15.900000 160.300000 ;
        RECT  1.005000 160.300000 15.830000 160.370000 ;
        RECT  1.005000 160.370000 15.760000 160.440000 ;
        RECT  1.005000 160.440000 15.690000 160.510000 ;
        RECT  1.005000 160.510000 15.620000 160.580000 ;
        RECT  1.005000 160.580000 15.550000 160.650000 ;
        RECT  1.005000 160.650000 15.480000 160.720000 ;
        RECT  1.005000 160.720000 15.410000 160.790000 ;
        RECT  1.005000 160.790000 15.340000 160.860000 ;
        RECT  1.005000 160.860000 15.270000 160.930000 ;
        RECT  1.005000 160.930000 15.200000 161.000000 ;
        RECT  1.005000 161.000000 15.130000 161.070000 ;
        RECT  1.005000 161.070000 15.060000 161.140000 ;
        RECT  1.005000 161.140000 14.990000 161.210000 ;
        RECT  1.005000 161.210000 14.920000 161.280000 ;
        RECT  1.005000 161.280000 14.850000 161.350000 ;
        RECT  1.005000 161.350000 14.780000 161.420000 ;
        RECT  1.005000 161.420000 14.710000 161.490000 ;
        RECT  1.005000 161.490000 14.640000 161.560000 ;
        RECT  1.005000 161.560000 14.570000 161.630000 ;
        RECT  1.005000 161.630000 14.500000 161.700000 ;
        RECT  1.005000 161.700000 14.430000 161.770000 ;
        RECT  1.005000 161.770000 14.360000 161.840000 ;
        RECT  1.005000 161.840000 14.290000 161.910000 ;
        RECT  1.005000 161.910000 14.220000 161.980000 ;
        RECT  1.005000 161.980000 14.150000 162.050000 ;
        RECT  1.005000 162.050000 14.120000 162.080000 ;
        RECT  1.005000 162.080000 14.120000 169.220000 ;
        RECT  1.005000 169.220000 14.120000 169.290000 ;
        RECT  1.005000 169.290000 14.190000 169.360000 ;
        RECT  1.005000 169.360000 14.260000 169.430000 ;
        RECT  1.005000 169.430000 14.330000 169.500000 ;
        RECT  1.005000 169.500000 14.400000 169.570000 ;
        RECT  1.005000 169.570000 14.470000 169.640000 ;
        RECT  1.005000 169.640000 14.540000 169.710000 ;
        RECT  1.005000 169.710000 14.610000 169.780000 ;
        RECT  1.005000 169.780000 14.680000 169.850000 ;
        RECT  1.005000 169.850000 14.750000 169.920000 ;
        RECT  1.005000 169.920000 14.820000 169.990000 ;
        RECT  1.005000 169.990000 14.890000 170.060000 ;
        RECT  1.005000 170.060000 14.960000 170.130000 ;
        RECT  1.005000 170.130000 15.030000 170.200000 ;
        RECT  1.005000 170.200000 15.100000 170.270000 ;
        RECT  1.005000 170.270000 15.170000 170.340000 ;
        RECT  1.005000 170.340000 15.240000 170.410000 ;
        RECT  1.005000 170.410000 15.310000 170.480000 ;
        RECT  1.005000 170.480000 15.380000 170.550000 ;
        RECT  1.005000 170.550000 15.450000 170.620000 ;
        RECT  1.005000 170.620000 15.520000 170.690000 ;
        RECT  1.005000 170.690000 15.590000 170.760000 ;
        RECT  1.005000 170.760000 15.660000 170.830000 ;
        RECT  1.005000 170.830000 15.730000 170.900000 ;
        RECT  1.005000 170.900000 15.800000 170.970000 ;
        RECT  1.005000 170.970000 15.870000 171.040000 ;
        RECT  1.005000 171.040000 15.940000 171.110000 ;
        RECT  1.005000 171.110000 16.010000 171.180000 ;
        RECT  1.005000 171.180000 16.080000 171.250000 ;
        RECT  1.005000 171.250000 16.150000 171.320000 ;
        RECT  1.005000 171.320000 16.220000 171.390000 ;
        RECT  1.005000 171.390000 16.290000 171.460000 ;
        RECT  1.005000 171.460000 16.360000 171.530000 ;
        RECT  1.005000 171.530000 16.430000 171.600000 ;
        RECT  1.005000 171.600000 16.500000 171.670000 ;
        RECT  1.005000 171.670000 16.570000 171.740000 ;
        RECT  1.005000 171.740000 16.640000 171.810000 ;
        RECT  1.005000 171.810000 16.710000 171.880000 ;
        RECT  1.005000 171.880000 16.780000 171.950000 ;
        RECT  1.005000 171.950000 16.850000 172.020000 ;
        RECT  1.005000 172.020000 16.920000 172.090000 ;
        RECT  1.005000 172.090000 16.990000 172.160000 ;
        RECT  1.005000 172.160000 17.060000 172.230000 ;
        RECT  1.005000 172.230000 17.130000 172.300000 ;
        RECT  1.005000 172.300000 17.200000 172.370000 ;
        RECT  1.005000 172.370000 17.270000 172.440000 ;
        RECT  1.005000 172.440000 17.340000 172.510000 ;
        RECT  1.005000 172.510000 17.410000 172.580000 ;
        RECT  1.005000 172.580000 17.480000 172.650000 ;
        RECT  1.005000 172.650000 17.550000 172.720000 ;
        RECT  1.005000 172.720000 17.620000 172.780000 ;
        RECT  1.005000 172.780000 57.960000 181.480000 ;
        RECT  1.005000 181.480000 17.625000 181.550000 ;
        RECT  1.005000 181.550000 17.555000 181.620000 ;
        RECT  1.005000 181.620000 17.485000 181.690000 ;
        RECT  1.005000 181.690000 17.415000 181.760000 ;
        RECT  1.005000 181.760000 17.345000 181.830000 ;
        RECT  1.005000 181.830000 17.275000 181.900000 ;
        RECT  1.005000 181.900000 17.205000 181.970000 ;
        RECT  1.005000 181.970000 17.135000 182.040000 ;
        RECT  1.005000 182.040000 17.065000 182.110000 ;
        RECT  1.005000 182.110000 16.995000 182.180000 ;
        RECT  1.005000 182.180000 16.925000 182.250000 ;
        RECT  1.005000 182.250000 16.855000 182.320000 ;
        RECT  1.005000 182.320000 16.785000 182.390000 ;
        RECT  1.005000 182.390000 16.715000 182.460000 ;
        RECT  1.005000 182.460000 16.645000 182.530000 ;
        RECT  1.005000 182.530000 16.575000 182.600000 ;
        RECT  1.005000 182.600000 16.505000 182.670000 ;
        RECT  1.005000 182.670000 16.435000 182.740000 ;
        RECT  1.005000 182.740000 16.365000 182.810000 ;
        RECT  1.005000 182.810000 16.295000 182.880000 ;
        RECT  1.005000 182.880000 16.225000 182.950000 ;
        RECT  1.005000 182.950000 16.155000 183.020000 ;
        RECT  1.005000 183.020000 16.085000 183.090000 ;
        RECT  1.005000 183.090000 16.015000 183.160000 ;
        RECT  1.005000 183.160000 15.945000 183.230000 ;
        RECT  1.005000 183.230000 15.875000 183.300000 ;
        RECT  1.005000 183.300000 15.805000 183.370000 ;
        RECT  1.005000 183.370000 15.735000 183.440000 ;
        RECT  1.005000 183.440000 15.665000 183.510000 ;
        RECT  1.005000 183.510000 15.595000 183.580000 ;
        RECT  1.005000 183.580000 15.525000 183.650000 ;
        RECT  1.005000 183.650000 15.455000 183.720000 ;
        RECT  1.005000 183.720000 15.385000 183.790000 ;
        RECT  1.005000 183.790000 15.315000 183.860000 ;
        RECT  1.005000 183.860000 15.245000 183.930000 ;
        RECT  1.005000 183.930000 15.175000 184.000000 ;
        RECT  1.005000 184.000000 15.105000 184.070000 ;
        RECT  1.005000 184.070000 15.035000 184.140000 ;
        RECT  1.005000 184.140000 14.965000 184.210000 ;
        RECT  1.005000 184.210000 14.895000 184.280000 ;
        RECT  1.005000 184.280000 14.825000 184.350000 ;
        RECT  1.005000 184.350000 14.755000 184.420000 ;
        RECT  1.005000 184.420000 14.685000 184.490000 ;
        RECT  1.005000 184.490000 14.615000 184.560000 ;
        RECT  1.005000 184.560000 14.545000 184.630000 ;
        RECT  1.005000 184.630000 14.475000 184.700000 ;
        RECT  1.005000 184.700000 14.405000 184.770000 ;
        RECT  1.005000 184.770000 14.335000 184.840000 ;
        RECT  1.005000 184.840000 14.265000 184.910000 ;
        RECT  1.005000 184.910000 14.195000 184.980000 ;
        RECT  1.005000 184.980000 14.125000 185.050000 ;
        RECT  1.005000 185.050000 14.120000 185.055000 ;
        RECT  1.005000 185.055000 14.120000 189.585000 ;
        RECT  1.005000 189.585000 14.120000 189.655000 ;
        RECT  1.005000 189.655000 14.190000 189.725000 ;
        RECT  1.005000 189.725000 14.260000 189.795000 ;
        RECT  1.005000 189.795000 14.330000 189.865000 ;
        RECT  1.005000 189.865000 14.400000 189.935000 ;
        RECT  1.005000 189.935000 14.470000 190.005000 ;
        RECT  1.005000 190.005000 14.540000 190.075000 ;
        RECT  1.005000 190.075000 14.610000 190.145000 ;
        RECT  1.005000 190.145000 14.680000 190.215000 ;
        RECT  1.005000 190.215000 14.750000 190.285000 ;
        RECT  1.005000 190.285000 14.820000 190.355000 ;
        RECT  1.005000 190.355000 14.890000 190.425000 ;
        RECT  1.005000 190.425000 14.960000 190.495000 ;
        RECT  1.005000 190.495000 15.030000 190.560000 ;
        RECT  1.005000 190.560000 67.200000 195.075000 ;
        RECT  1.010000  47.125000 14.120000  47.130000 ;
        RECT  1.045000  36.640000 16.180000  36.680000 ;
        RECT  1.050000  47.085000 14.120000  47.125000 ;
        RECT  1.085000  36.680000 16.220000  36.720000 ;
        RECT  1.090000  36.720000 16.260000  36.725000 ;
        RECT  1.090000  36.725000 16.265000  36.795000 ;
        RECT  1.090000  36.795000 16.335000  36.865000 ;
        RECT  1.090000  36.865000 16.405000  36.935000 ;
        RECT  1.090000  36.935000 16.475000  37.005000 ;
        RECT  1.090000  37.005000 16.545000  37.075000 ;
        RECT  1.090000  37.075000 16.615000  37.145000 ;
        RECT  1.090000  37.145000 16.685000  37.215000 ;
        RECT  1.090000  37.215000 16.755000  37.285000 ;
        RECT  1.090000  37.285000 16.825000  37.355000 ;
        RECT  1.090000  37.355000 16.895000  37.425000 ;
        RECT  1.090000  37.425000 16.965000  37.495000 ;
        RECT  1.090000  37.495000 17.035000  37.565000 ;
        RECT  1.090000  37.565000 17.105000  37.635000 ;
        RECT  1.090000  37.635000 17.175000  37.705000 ;
        RECT  1.090000  37.705000 17.245000  37.775000 ;
        RECT  1.090000  37.775000 17.315000  37.845000 ;
        RECT  1.090000  37.845000 17.385000  37.915000 ;
        RECT  1.090000  37.915000 17.455000  37.985000 ;
        RECT  1.090000  37.985000 17.525000  38.055000 ;
        RECT  1.090000  38.055000 17.595000  38.125000 ;
        RECT  1.090000  38.125000 17.665000  38.195000 ;
        RECT  1.090000  38.195000 17.735000  38.265000 ;
        RECT  1.090000  38.265000 17.805000  38.335000 ;
        RECT  1.090000  38.335000 17.875000  38.405000 ;
        RECT  1.090000  38.405000 17.945000  38.475000 ;
        RECT  1.090000  38.475000 18.015000  38.545000 ;
        RECT  1.090000  38.545000 18.085000  38.615000 ;
        RECT  1.090000  38.615000 18.155000  38.685000 ;
        RECT  1.090000  38.685000 18.225000  38.755000 ;
        RECT  1.090000  38.755000 18.295000  38.825000 ;
        RECT  1.090000  38.825000 18.365000  38.895000 ;
        RECT  1.090000  38.895000 18.435000  38.965000 ;
        RECT  1.090000  38.965000 18.505000  39.035000 ;
        RECT  1.090000  39.035000 18.575000  39.105000 ;
        RECT  1.090000  39.105000 18.645000  39.175000 ;
        RECT  1.090000  39.175000 18.715000  39.245000 ;
        RECT  1.090000  39.245000 18.785000  39.315000 ;
        RECT  1.090000  39.315000 18.855000  39.385000 ;
        RECT  1.090000  39.385000 18.925000  39.455000 ;
        RECT  1.090000  39.455000 18.995000  39.525000 ;
        RECT  1.090000  39.525000 19.065000  39.595000 ;
        RECT  1.090000  39.595000 19.135000  39.665000 ;
        RECT  1.090000  39.665000 19.205000  39.735000 ;
        RECT  1.090000  39.735000 19.275000  39.805000 ;
        RECT  1.090000  39.805000 19.345000  39.875000 ;
        RECT  1.090000  39.875000 19.415000  39.945000 ;
        RECT  1.090000  39.945000 19.485000  40.015000 ;
        RECT  1.090000  40.015000 19.555000  40.085000 ;
        RECT  1.090000  40.085000 19.625000  40.155000 ;
        RECT  1.090000  40.155000 19.695000  40.225000 ;
        RECT  1.090000  40.225000 19.765000  40.295000 ;
        RECT  1.090000  40.295000 19.835000  40.350000 ;
        RECT  1.090000  40.350000 56.160000  40.420000 ;
        RECT  1.090000  40.420000 56.090000  40.490000 ;
        RECT  1.090000  40.490000 56.020000  40.560000 ;
        RECT  1.090000  40.560000 55.950000  40.630000 ;
        RECT  1.090000  40.630000 55.880000  40.700000 ;
        RECT  1.090000  40.700000 55.810000  40.770000 ;
        RECT  1.090000  40.770000 55.740000  40.840000 ;
        RECT  1.090000  40.840000 55.670000  40.910000 ;
        RECT  1.090000  40.910000 55.600000  40.980000 ;
        RECT  1.090000  40.980000 55.530000  41.050000 ;
        RECT  1.090000  41.050000 55.460000  41.120000 ;
        RECT  1.090000  41.120000 55.390000  41.190000 ;
        RECT  1.090000  41.190000 55.320000  41.260000 ;
        RECT  1.090000  41.260000 55.250000  41.330000 ;
        RECT  1.090000  41.330000 55.180000  41.400000 ;
        RECT  1.090000  41.400000 55.110000  41.470000 ;
        RECT  1.090000  41.470000 55.040000  41.540000 ;
        RECT  1.090000  41.540000 54.970000  41.610000 ;
        RECT  1.090000  41.610000 54.900000  41.680000 ;
        RECT  1.090000  41.680000 54.830000  41.750000 ;
        RECT  1.090000  41.750000 54.760000  41.820000 ;
        RECT  1.090000  41.820000 54.690000  41.890000 ;
        RECT  1.090000  41.890000 54.620000  41.960000 ;
        RECT  1.090000  41.960000 54.550000  42.030000 ;
        RECT  1.090000  42.030000 54.480000  42.100000 ;
        RECT  1.090000  42.100000 54.410000  42.170000 ;
        RECT  1.090000  42.170000 54.340000  42.240000 ;
        RECT  1.090000  42.240000 54.270000  42.310000 ;
        RECT  1.090000  42.310000 54.200000  42.380000 ;
        RECT  1.090000  42.380000 16.985000  42.450000 ;
        RECT  1.090000  42.450000 16.915000  42.520000 ;
        RECT  1.090000  42.520000 16.845000  42.590000 ;
        RECT  1.090000  42.590000 16.775000  42.660000 ;
        RECT  1.090000  42.660000 16.705000  42.730000 ;
        RECT  1.090000  42.730000 16.635000  42.800000 ;
        RECT  1.090000  42.800000 16.565000  42.870000 ;
        RECT  1.090000  42.870000 16.495000  42.940000 ;
        RECT  1.090000  42.940000 16.425000  43.010000 ;
        RECT  1.090000  43.010000 16.355000  43.080000 ;
        RECT  1.090000  43.080000 16.285000  43.150000 ;
        RECT  1.090000  43.150000 16.215000  43.220000 ;
        RECT  1.090000  43.220000 16.145000  43.290000 ;
        RECT  1.090000  43.290000 16.075000  43.360000 ;
        RECT  1.090000  43.360000 16.005000  43.430000 ;
        RECT  1.090000  43.430000 15.935000  43.500000 ;
        RECT  1.090000  43.500000 15.865000  43.570000 ;
        RECT  1.090000  43.570000 15.795000  43.640000 ;
        RECT  1.090000  43.640000 15.725000  43.710000 ;
        RECT  1.090000  43.710000 15.655000  43.780000 ;
        RECT  1.090000  43.780000 15.585000  43.850000 ;
        RECT  1.090000  43.850000 15.515000  43.920000 ;
        RECT  1.090000  43.920000 15.445000  43.990000 ;
        RECT  1.090000  43.990000 15.375000  44.060000 ;
        RECT  1.090000  44.060000 15.305000  44.130000 ;
        RECT  1.090000  44.130000 15.235000  44.200000 ;
        RECT  1.090000  44.200000 15.165000  44.270000 ;
        RECT  1.090000  44.270000 15.095000  44.340000 ;
        RECT  1.090000  44.340000 15.025000  44.410000 ;
        RECT  1.090000  44.410000 14.955000  44.480000 ;
        RECT  1.090000  44.480000 14.885000  44.550000 ;
        RECT  1.090000  44.550000 14.815000  44.620000 ;
        RECT  1.090000  44.620000 14.745000  44.690000 ;
        RECT  1.090000  44.690000 14.675000  44.760000 ;
        RECT  1.090000  44.760000 14.605000  44.830000 ;
        RECT  1.090000  44.830000 14.535000  44.900000 ;
        RECT  1.090000  44.900000 14.465000  44.970000 ;
        RECT  1.090000  44.970000 14.395000  45.040000 ;
        RECT  1.090000  45.040000 14.325000  45.110000 ;
        RECT  1.090000  45.110000 14.255000  45.180000 ;
        RECT  1.090000  45.180000 14.185000  45.250000 ;
        RECT  1.090000  45.250000 14.120000  45.315000 ;
        RECT  1.090000  45.315000 14.120000  47.045000 ;
        RECT  1.090000  47.045000 14.120000  47.085000 ;
        RECT 52.630000  40.295000 56.230000  40.350000 ;
        RECT 52.700000  40.225000 56.285000  40.295000 ;
        RECT 52.770000  40.155000 56.355000  40.225000 ;
        RECT 52.840000  40.085000 56.425000  40.155000 ;
        RECT 52.910000  40.015000 56.495000  40.085000 ;
        RECT 52.980000  39.945000 56.565000  40.015000 ;
        RECT 53.050000  39.875000 56.635000  39.945000 ;
        RECT 53.120000  39.805000 56.705000  39.875000 ;
        RECT 53.190000  39.735000 56.775000  39.805000 ;
        RECT 53.260000  39.665000 56.845000  39.735000 ;
        RECT 53.270000  39.655000 56.915000  39.665000 ;
        RECT 53.340000  39.585000 56.915000  39.655000 ;
        RECT 53.410000  39.515000 56.915000  39.585000 ;
        RECT 53.480000  39.445000 56.915000  39.515000 ;
        RECT 53.550000  39.375000 56.915000  39.445000 ;
        RECT 53.620000  39.305000 56.915000  39.375000 ;
        RECT 53.690000  39.235000 56.915000  39.305000 ;
        RECT 53.760000  39.165000 56.915000  39.235000 ;
        RECT 53.830000  39.095000 56.915000  39.165000 ;
        RECT 53.900000  39.025000 56.915000  39.095000 ;
        RECT 53.970000  38.955000 56.915000  39.025000 ;
        RECT 54.040000  38.885000 56.915000  38.955000 ;
        RECT 54.110000  38.815000 56.915000  38.885000 ;
        RECT 54.180000  38.745000 56.915000  38.815000 ;
        RECT 54.250000  38.675000 56.915000  38.745000 ;
        RECT 54.320000  38.605000 56.915000  38.675000 ;
        RECT 54.390000  38.535000 56.915000  38.605000 ;
        RECT 54.460000  38.465000 56.915000  38.535000 ;
        RECT 54.530000  38.395000 56.915000  38.465000 ;
        RECT 54.600000  38.325000 56.915000  38.395000 ;
        RECT 54.670000  36.115000 56.915000  38.255000 ;
        RECT 54.670000  38.255000 56.915000  38.325000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.050000 172.755000 25.010000 195.100000 ;
        RECT 14.055000 172.750000 25.010000 172.755000 ;
        RECT 14.110000 172.695000 25.010000 172.750000 ;
        RECT 14.165000 172.640000 25.010000 172.695000 ;
        RECT 14.300000 172.505000 24.875000 172.640000 ;
        RECT 14.450000 172.355000 24.725000 172.505000 ;
        RECT 14.600000 172.205000 24.575000 172.355000 ;
        RECT 14.750000 172.055000 24.425000 172.205000 ;
        RECT 14.900000 171.905000 24.275000 172.055000 ;
        RECT 15.050000 171.755000 24.125000 171.905000 ;
        RECT 15.200000 171.605000 23.975000 171.755000 ;
        RECT 15.350000 171.455000 23.825000 171.605000 ;
        RECT 15.500000 102.200000 23.830000 102.350000 ;
        RECT 15.500000 102.350000 23.680000 102.500000 ;
        RECT 15.500000 102.500000 23.530000 102.650000 ;
        RECT 15.500000 102.650000 23.380000 102.800000 ;
        RECT 15.500000 102.800000 23.230000 102.950000 ;
        RECT 15.500000 102.950000 23.080000 103.100000 ;
        RECT 15.500000 103.100000 22.930000 103.250000 ;
        RECT 15.500000 103.250000 22.780000 103.400000 ;
        RECT 15.500000 103.400000 22.630000 103.550000 ;
        RECT 15.500000 103.550000 22.480000 103.700000 ;
        RECT 15.500000 103.700000 22.330000 103.850000 ;
        RECT 15.500000 103.850000 22.180000 104.000000 ;
        RECT 15.500000 104.000000 22.030000 104.150000 ;
        RECT 15.500000 104.150000 21.880000 104.300000 ;
        RECT 15.500000 104.300000 21.730000 104.450000 ;
        RECT 15.500000 104.450000 21.580000 104.600000 ;
        RECT 15.500000 104.600000 21.500000 104.680000 ;
        RECT 15.500000 104.680000 21.500000 169.130000 ;
        RECT 15.500000 169.130000 21.500000 169.280000 ;
        RECT 15.500000 169.280000 21.650000 169.430000 ;
        RECT 15.500000 169.430000 21.800000 169.580000 ;
        RECT 15.500000 169.580000 21.950000 169.730000 ;
        RECT 15.500000 169.730000 22.100000 169.880000 ;
        RECT 15.500000 169.880000 22.250000 170.030000 ;
        RECT 15.500000 170.030000 22.400000 170.180000 ;
        RECT 15.500000 170.180000 22.550000 170.330000 ;
        RECT 15.500000 170.330000 22.700000 170.480000 ;
        RECT 15.500000 170.480000 22.850000 170.630000 ;
        RECT 15.500000 170.630000 23.000000 170.780000 ;
        RECT 15.500000 170.780000 23.150000 170.930000 ;
        RECT 15.500000 170.930000 23.300000 171.080000 ;
        RECT 15.500000 171.080000 23.450000 171.230000 ;
        RECT 15.500000 171.230000 23.600000 171.305000 ;
        RECT 15.500000 171.305000 23.675000 171.455000 ;
        RECT 15.645000 102.055000 23.980000 102.200000 ;
        RECT 15.795000 101.905000 24.125000 102.055000 ;
        RECT 15.945000 101.755000 24.275000 101.905000 ;
        RECT 16.095000 101.605000 24.425000 101.755000 ;
        RECT 16.245000 101.455000 24.575000 101.605000 ;
        RECT 16.395000 101.305000 24.725000 101.455000 ;
        RECT 16.545000 101.155000 24.875000 101.305000 ;
        RECT 16.695000 101.005000 25.025000 101.155000 ;
        RECT 16.845000 100.855000 25.175000 101.005000 ;
        RECT 16.995000 100.705000 25.325000 100.855000 ;
        RECT 17.145000 100.555000 25.475000 100.705000 ;
        RECT 17.295000 100.405000 25.625000 100.555000 ;
        RECT 17.445000 100.255000 25.775000 100.405000 ;
        RECT 17.595000 100.105000 25.925000 100.255000 ;
        RECT 17.745000  99.955000 26.075000 100.105000 ;
        RECT 17.895000  99.805000 26.225000  99.955000 ;
        RECT 18.045000  99.655000 26.375000  99.805000 ;
        RECT 18.195000  99.505000 26.525000  99.655000 ;
        RECT 18.345000  99.355000 26.675000  99.505000 ;
        RECT 18.495000  99.205000 26.825000  99.355000 ;
        RECT 18.645000  99.055000 26.975000  99.205000 ;
        RECT 18.795000  98.905000 27.125000  99.055000 ;
        RECT 18.945000  98.755000 27.275000  98.905000 ;
        RECT 19.095000  98.605000 27.425000  98.755000 ;
        RECT 19.245000  98.455000 27.575000  98.605000 ;
        RECT 19.395000  98.305000 27.725000  98.455000 ;
        RECT 19.545000  98.155000 27.875000  98.305000 ;
        RECT 19.695000  98.005000 28.025000  98.155000 ;
        RECT 19.845000  97.855000 28.175000  98.005000 ;
        RECT 19.995000  97.705000 28.325000  97.855000 ;
        RECT 20.145000  97.555000 28.475000  97.705000 ;
        RECT 20.295000  97.405000 28.625000  97.555000 ;
        RECT 20.445000  97.255000 28.775000  97.405000 ;
        RECT 20.595000  97.105000 28.925000  97.255000 ;
        RECT 20.745000  96.955000 29.075000  97.105000 ;
        RECT 20.895000  96.805000 29.225000  96.955000 ;
        RECT 21.045000  96.655000 29.375000  96.805000 ;
        RECT 21.195000  96.505000 29.525000  96.655000 ;
        RECT 21.345000  96.355000 29.525000  96.505000 ;
        RECT 21.495000  96.205000 29.525000  96.355000 ;
        RECT 21.645000  96.055000 29.525000  96.205000 ;
        RECT 21.795000  95.905000 29.525000  96.055000 ;
        RECT 21.945000  95.755000 29.525000  95.905000 ;
        RECT 22.095000  95.605000 29.525000  95.755000 ;
        RECT 22.245000  95.455000 29.525000  95.605000 ;
        RECT 22.395000  95.305000 29.525000  95.455000 ;
        RECT 22.545000  95.155000 29.525000  95.305000 ;
        RECT 22.695000  95.005000 29.525000  95.155000 ;
        RECT 22.845000  94.855000 29.525000  95.005000 ;
        RECT 22.995000  94.705000 29.525000  94.855000 ;
        RECT 23.145000  94.555000 29.525000  94.705000 ;
        RECT 23.295000  94.405000 29.525000  94.555000 ;
        RECT 23.445000  94.255000 29.525000  94.405000 ;
        RECT 23.595000  94.105000 29.525000  94.255000 ;
        RECT 23.745000  92.540000 29.935000  92.690000 ;
        RECT 23.745000  92.690000 29.785000  92.840000 ;
        RECT 23.745000  92.840000 29.635000  92.990000 ;
        RECT 23.745000  92.990000 29.525000  93.100000 ;
        RECT 23.745000  93.100000 29.525000  93.955000 ;
        RECT 23.745000  93.955000 29.525000  94.105000 ;
        RECT 23.820000  92.465000 30.085000  92.540000 ;
        RECT 23.895000  92.390000 30.160000  92.465000 ;
        RECT 23.945000  92.340000 36.895000  92.390000 ;
        RECT 24.095000  92.190000 36.895000  92.340000 ;
        RECT 24.245000  92.040000 36.895000  92.190000 ;
        RECT 24.395000  91.890000 36.895000  92.040000 ;
        RECT 24.545000  91.740000 36.895000  91.890000 ;
        RECT 24.695000  91.590000 36.895000  91.740000 ;
        RECT 24.845000  91.440000 36.895000  91.590000 ;
        RECT 24.995000  91.290000 36.895000  91.440000 ;
        RECT 25.145000  91.140000 36.895000  91.290000 ;
        RECT 25.295000  90.990000 36.895000  91.140000 ;
        RECT 25.445000  90.840000 36.895000  90.990000 ;
        RECT 25.595000  90.690000 36.895000  90.840000 ;
        RECT 25.745000  90.540000 36.895000  90.690000 ;
        RECT 25.895000   0.000000 36.895000  90.390000 ;
        RECT 25.895000  90.390000 36.895000  90.540000 ;
        RECT 25.930000 102.390000 34.250000 102.540000 ;
        RECT 25.930000 102.540000 34.100000 102.690000 ;
        RECT 25.930000 102.690000 33.950000 102.840000 ;
        RECT 25.930000 102.840000 33.800000 102.990000 ;
        RECT 25.930000 102.990000 33.650000 103.140000 ;
        RECT 25.930000 103.140000 33.500000 103.290000 ;
        RECT 25.930000 103.290000 33.350000 103.440000 ;
        RECT 25.930000 103.440000 33.200000 103.590000 ;
        RECT 25.930000 103.590000 33.050000 103.740000 ;
        RECT 25.930000 103.740000 32.900000 103.890000 ;
        RECT 25.930000 103.890000 32.750000 104.040000 ;
        RECT 25.930000 104.040000 32.600000 104.190000 ;
        RECT 25.930000 104.190000 32.450000 104.340000 ;
        RECT 25.930000 104.340000 32.300000 104.490000 ;
        RECT 25.930000 104.490000 32.150000 104.640000 ;
        RECT 25.930000 104.640000 32.000000 104.790000 ;
        RECT 25.930000 104.790000 31.930000 104.860000 ;
        RECT 25.930000 104.860000 31.930000 170.460000 ;
        RECT 25.930000 170.460000 31.930000 170.610000 ;
        RECT 25.930000 170.610000 32.080000 170.760000 ;
        RECT 25.930000 170.760000 32.230000 170.910000 ;
        RECT 25.930000 170.910000 32.380000 171.060000 ;
        RECT 25.930000 171.060000 32.530000 171.210000 ;
        RECT 25.930000 171.210000 32.680000 171.360000 ;
        RECT 25.930000 171.360000 32.830000 171.510000 ;
        RECT 25.930000 171.510000 32.980000 171.660000 ;
        RECT 25.930000 171.660000 33.130000 171.810000 ;
        RECT 25.930000 171.810000 33.280000 171.960000 ;
        RECT 25.930000 171.960000 33.430000 172.110000 ;
        RECT 25.930000 172.110000 33.580000 172.260000 ;
        RECT 25.930000 172.260000 33.730000 172.410000 ;
        RECT 25.930000 172.410000 33.880000 172.560000 ;
        RECT 25.930000 172.560000 34.030000 172.710000 ;
        RECT 25.930000 172.710000 34.180000 172.860000 ;
        RECT 25.930000 172.860000 34.330000 173.010000 ;
        RECT 25.930000 173.010000 34.480000 173.160000 ;
        RECT 25.930000 173.160000 34.630000 173.310000 ;
        RECT 25.930000 173.310000 34.780000 173.460000 ;
        RECT 25.930000 173.460000 34.930000 173.610000 ;
        RECT 25.930000 173.610000 35.080000 173.760000 ;
        RECT 25.930000 173.760000 35.230000 173.910000 ;
        RECT 25.930000 173.910000 35.380000 174.060000 ;
        RECT 25.930000 174.060000 35.530000 174.210000 ;
        RECT 25.930000 174.210000 35.680000 174.360000 ;
        RECT 25.930000 174.360000 35.830000 174.510000 ;
        RECT 25.930000 174.510000 35.980000 174.660000 ;
        RECT 25.930000 174.660000 36.130000 174.810000 ;
        RECT 25.930000 174.810000 36.280000 174.960000 ;
        RECT 25.930000 174.960000 36.430000 175.110000 ;
        RECT 25.930000 175.110000 36.580000 175.260000 ;
        RECT 25.930000 175.260000 36.730000 175.350000 ;
        RECT 25.930000 175.350000 36.820000 195.100000 ;
        RECT 26.025000 102.295000 34.400000 102.390000 ;
        RECT 26.175000 102.145000 34.495000 102.295000 ;
        RECT 26.325000 101.995000 34.645000 102.145000 ;
        RECT 26.475000 101.845000 34.795000 101.995000 ;
        RECT 26.625000 101.695000 34.945000 101.845000 ;
        RECT 26.775000 101.545000 35.095000 101.695000 ;
        RECT 26.925000 101.395000 35.245000 101.545000 ;
        RECT 27.075000 101.245000 35.395000 101.395000 ;
        RECT 27.225000 101.095000 35.545000 101.245000 ;
        RECT 27.375000 100.945000 35.695000 101.095000 ;
        RECT 27.525000 100.795000 35.845000 100.945000 ;
        RECT 27.675000 100.645000 35.995000 100.795000 ;
        RECT 27.825000 100.495000 36.145000 100.645000 ;
        RECT 27.975000 100.345000 36.295000 100.495000 ;
        RECT 28.125000 100.195000 36.445000 100.345000 ;
        RECT 28.275000 100.045000 36.595000 100.195000 ;
        RECT 28.425000  99.895000 36.745000 100.045000 ;
        RECT 28.495000  99.825000 36.895000  99.895000 ;
        RECT 28.645000  99.675000 36.895000  99.825000 ;
        RECT 28.795000  99.525000 36.895000  99.675000 ;
        RECT 28.945000  99.375000 36.895000  99.525000 ;
        RECT 29.095000  99.225000 36.895000  99.375000 ;
        RECT 29.245000  99.075000 36.895000  99.225000 ;
        RECT 29.395000  98.925000 36.895000  99.075000 ;
        RECT 29.545000  98.775000 36.895000  98.925000 ;
        RECT 29.695000  98.625000 36.895000  98.775000 ;
        RECT 29.845000  98.475000 36.895000  98.625000 ;
        RECT 29.995000  98.325000 36.895000  98.475000 ;
        RECT 30.145000  98.175000 36.895000  98.325000 ;
        RECT 30.295000  98.025000 36.895000  98.175000 ;
        RECT 30.445000  97.875000 36.895000  98.025000 ;
        RECT 30.595000  97.725000 36.895000  97.875000 ;
        RECT 30.745000  97.575000 36.895000  97.725000 ;
        RECT 30.895000  97.425000 36.895000  97.575000 ;
        RECT 31.045000  97.275000 36.895000  97.425000 ;
        RECT 31.195000  97.125000 36.895000  97.275000 ;
        RECT 31.345000  96.975000 36.895000  97.125000 ;
        RECT 31.385000  92.390000 36.895000  92.540000 ;
        RECT 31.495000  96.825000 36.895000  96.975000 ;
        RECT 31.535000  92.540000 36.895000  92.690000 ;
        RECT 31.645000  96.675000 36.895000  96.825000 ;
        RECT 31.685000  92.690000 36.895000  92.840000 ;
        RECT 31.795000  96.525000 36.895000  96.675000 ;
        RECT 31.835000  92.840000 36.895000  92.990000 ;
        RECT 31.945000  92.990000 36.895000  93.100000 ;
        RECT 31.945000  93.100000 36.895000  96.375000 ;
        RECT 31.945000  96.375000 36.895000  96.525000 ;
    END
  END SRC_BDY_HVC
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 8.885000 1.270000 13.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 8.885000 75.000000 13.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 8.985000 1.270000 13.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 8.985000 75.000000 13.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2.035000 1.270000 7.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 2.035000 75.000000 7.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 2.135000 1.270000 7.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 2.135000 75.000000 7.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 14.935000 0.965000 18.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035000 14.935000 75.000000 18.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 15.035000 0.965000 18.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 15.035000 75.000000 18.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 19.785000 1.270000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 70.035000 1.270000 95.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 19.785000 75.000000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 70.035000 75.000000 95.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 19.885000 1.270000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 70.035000 1.270000 94.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 19.885000 75.000000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 70.035000 75.000000 94.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 64.085000 1.270000 68.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 64.085000 75.000000 68.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 64.185000 1.270000 68.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 64.185000 75.000000 68.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 36.735000 1.270000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 47.735000 1.270000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 51.645000 1.270000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 56.405000 1.270000 56.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 36.735000 75.000000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 47.735000 75.000000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.645000 75.000000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 56.405000 75.000000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 36.840000 1.270000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 47.735000 1.270000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 36.840000 75.000000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 47.735000 75.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 41.585000 1.270000 46.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 41.585000 75.000000 46.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 41.685000 1.270000 46.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 41.685000 75.000000 46.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 25.835000 1.270000 30.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 25.835000 75.000000 30.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 25.935000 1.270000 30.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 25.935000 75.000000 30.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 58.235000 1.270000 62.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 58.235000 75.000000 62.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 58.335000 1.270000 62.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 58.335000 75.000000 62.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 31.885000 1.270000 35.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 31.885000 75.000000 35.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 31.985000 1.270000 35.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 31.985000 75.000000 35.235000 ;
    END
  END VSWITCH
  OBS
    LAYER li1 ;
      RECT  1.145000  43.280000  1.315000  43.810000 ;
      RECT  3.100000  27.160000 48.200000  28.030000 ;
      RECT  3.100000  28.030000  4.020000  38.695000 ;
      RECT  3.100000  38.695000 48.200000  39.565000 ;
      RECT  3.130000  27.140000 48.200000  27.160000 ;
      RECT  3.130000  39.565000 48.200000  39.585000 ;
      RECT  4.735000  29.230000 45.955000  29.430000 ;
      RECT  4.735000  29.430000  4.905000  37.425000 ;
      RECT  4.735000  37.425000 45.955000  37.595000 ;
      RECT  6.115000  33.340000  6.285000  36.490000 ;
      RECT  6.340000  36.970000 45.060000  37.230000 ;
      RECT  6.895000  29.775000  7.065000  32.860000 ;
      RECT  7.675000  33.335000  7.845000  36.490000 ;
      RECT  8.050000  43.270000  8.580000  43.440000 ;
      RECT  8.455000  29.770000  8.625000  32.860000 ;
      RECT  8.510000 162.655000 10.360000 169.150000 ;
      RECT  9.135000  43.505000 70.125000  44.755000 ;
      RECT  9.135000  44.755000 10.385000  71.570000 ;
      RECT  9.135000  71.570000 21.085000  72.820000 ;
      RECT  9.150000 169.400000 10.400000 198.445000 ;
      RECT  9.150000 198.445000 70.125000 199.695000 ;
      RECT  9.170000 133.350000 20.990000 134.540000 ;
      RECT  9.170000 134.540000 10.360000 162.655000 ;
      RECT  9.170000 169.150000 10.360000 169.400000 ;
      RECT  9.200000 133.205000 14.190000 133.350000 ;
      RECT  9.235000  33.340000  9.405000  36.490000 ;
      RECT  9.405000  74.180000  9.935000  74.350000 ;
      RECT 10.015000  29.775000 10.185000  32.860000 ;
      RECT 10.770000 162.655000 11.975000 169.905000 ;
      RECT 10.795000  33.335000 10.965000  36.490000 ;
      RECT 11.100000 170.415000 11.990000 196.835000 ;
      RECT 11.100000 196.835000 68.155000 197.725000 ;
      RECT 11.105000  45.460000 68.155000  46.350000 ;
      RECT 11.105000  46.350000 11.995000  69.975000 ;
      RECT 11.105000  69.975000 22.680000  70.865000 ;
      RECT 11.125000 135.315000 22.660000 136.165000 ;
      RECT 11.125000 136.165000 12.100000 158.915000 ;
      RECT 11.125000 158.915000 11.975000 162.655000 ;
      RECT 11.125000 169.905000 11.975000 170.415000 ;
      RECT 11.575000  29.770000 11.745000  32.860000 ;
      RECT 12.065000   1.000000 70.650000   1.890000 ;
      RECT 12.065000   1.890000 13.045000  22.230000 ;
      RECT 12.065000  22.230000 56.085000  22.350000 ;
      RECT 12.065000  22.350000 56.105000  23.240000 ;
      RECT 12.355000  33.340000 12.525000  36.490000 ;
      RECT 12.400000 159.555000 64.500000 161.990000 ;
      RECT 12.830000 182.570000 66.685000 184.990000 ;
      RECT 13.085000  46.815000 64.500000  46.990000 ;
      RECT 13.085000  46.990000 13.255000  67.965000 ;
      RECT 13.090000  46.740000 64.500000  46.815000 ;
      RECT 13.135000  29.775000 13.305000  32.860000 ;
      RECT 13.915000  33.335000 14.085000  36.490000 ;
      RECT 14.385000  47.160000 15.415000  66.930000 ;
      RECT 14.385000 139.160000 15.415000 158.930000 ;
      RECT 14.385000 162.160000 15.415000 181.930000 ;
      RECT 14.385000 185.160000 15.435000 195.185000 ;
      RECT 14.695000  29.770000 14.865000  32.860000 ;
      RECT 15.475000  33.340000 15.645000  36.490000 ;
      RECT 15.705000  67.340000 64.500000  68.995000 ;
      RECT 15.780000 136.540000 64.500000 138.990000 ;
      RECT 15.780000 159.340000 64.500000 159.555000 ;
      RECT 15.780000 182.340000 66.685000 182.570000 ;
      RECT 15.780000 195.370000 16.490000 195.540000 ;
      RECT 16.255000  29.770000 16.425000  32.860000 ;
      RECT 17.035000  33.335000 17.205000  36.490000 ;
      RECT 17.790000 195.370000 18.500000 195.540000 ;
      RECT 17.815000  29.770000 17.985000  32.860000 ;
      RECT 17.835000 133.145000 20.990000 133.350000 ;
      RECT 18.470000  74.200000 19.000000  74.370000 ;
      RECT 18.595000  33.340000 18.765000  36.490000 ;
      RECT 18.985000  47.515000 19.875000  66.855000 ;
      RECT 18.985000 139.515000 19.875000 158.810000 ;
      RECT 18.985000 162.515000 19.875000 181.810000 ;
      RECT 18.985000 185.515000 19.875000 195.075000 ;
      RECT 19.375000  29.775000 19.545000  32.860000 ;
      RECT 19.565000  97.500000 20.990000 133.145000 ;
      RECT 19.800000  72.820000 21.085000  96.895000 ;
      RECT 19.800000  96.895000 20.990000  97.500000 ;
      RECT 20.155000  33.335000 20.325000  36.490000 ;
      RECT 20.380000 195.370000 21.090000 195.540000 ;
      RECT 20.935000  29.770000 21.105000  32.860000 ;
      RECT 21.715000  33.340000 21.885000  36.490000 ;
      RECT 21.790000  70.865000 22.680000  97.450000 ;
      RECT 21.810000  97.450000 22.660000 135.315000 ;
      RECT 22.390000 195.370000 23.100000 195.540000 ;
      RECT 22.495000  29.775000 22.665000  32.860000 ;
      RECT 23.025000  90.495000 64.500000  92.990000 ;
      RECT 23.055000 113.340000 64.500000 115.990000 ;
      RECT 23.275000  33.335000 23.445000  36.490000 ;
      RECT 23.510000  68.995000 64.500000  69.990000 ;
      RECT 23.585000  47.515000 24.475000  66.810000 ;
      RECT 23.585000  70.160000 24.615000  89.930000 ;
      RECT 23.585000  93.160000 24.615000 112.930000 ;
      RECT 23.585000 116.160000 24.615000 135.930000 ;
      RECT 23.585000 139.515000 24.475000 158.765000 ;
      RECT 23.585000 162.515000 24.475000 181.765000 ;
      RECT 23.585000 185.515000 24.475000 195.030000 ;
      RECT 24.055000  29.770000 24.225000  32.860000 ;
      RECT 24.835000  33.340000 25.005000  36.490000 ;
      RECT 24.980000  90.370000 64.500000  90.495000 ;
      RECT 24.980000 136.370000 64.500000 136.540000 ;
      RECT 24.980000 195.370000 25.690000 195.540000 ;
      RECT 25.615000  29.775000 25.785000  32.860000 ;
      RECT 25.670000  90.340000 64.500000  90.370000 ;
      RECT 25.670000 136.340000 64.500000 136.370000 ;
      RECT 26.395000  33.335000 26.565000  36.490000 ;
      RECT 26.990000 195.370000 27.700000 195.540000 ;
      RECT 27.175000  29.770000 27.345000  32.860000 ;
      RECT 27.955000  33.340000 28.125000  36.490000 ;
      RECT 28.185000  47.515000 29.075000  66.810000 ;
      RECT 28.185000  70.515000 29.075000  89.810000 ;
      RECT 28.185000  93.515000 29.075000 112.855000 ;
      RECT 28.185000 116.515000 29.075000 135.810000 ;
      RECT 28.185000 139.515000 29.075000 158.765000 ;
      RECT 28.185000 162.515000 29.075000 181.765000 ;
      RECT 28.185000 185.515000 29.075000 195.030000 ;
      RECT 28.735000  29.775000 28.905000  32.860000 ;
      RECT 29.515000  33.335000 29.685000  36.490000 ;
      RECT 29.580000 195.370000 30.290000 195.540000 ;
      RECT 30.295000  29.770000 30.465000  32.860000 ;
      RECT 31.075000  33.340000 31.245000  36.490000 ;
      RECT 31.590000 195.370000 32.300000 195.540000 ;
      RECT 31.855000  29.775000 32.025000  32.860000 ;
      RECT 32.635000  33.335000 32.805000  36.490000 ;
      RECT 32.785000  47.515000 33.675000  66.810000 ;
      RECT 32.785000  70.515000 33.675000  89.765000 ;
      RECT 32.785000  93.515000 33.675000 112.810000 ;
      RECT 32.785000 116.515000 33.675000 135.765000 ;
      RECT 32.785000 139.515000 33.675000 158.765000 ;
      RECT 32.785000 162.515000 33.675000 181.765000 ;
      RECT 32.785000 185.515000 33.675000 195.030000 ;
      RECT 33.415000  29.770000 33.585000  32.860000 ;
      RECT 34.180000 195.370000 34.890000 195.540000 ;
      RECT 34.195000  33.340000 34.365000  36.490000 ;
      RECT 34.975000  29.775000 35.145000  32.860000 ;
      RECT 35.755000  33.335000 35.925000  36.490000 ;
      RECT 36.190000 195.370000 36.900000 195.540000 ;
      RECT 36.535000  29.770000 36.705000  32.860000 ;
      RECT 37.315000  33.340000 37.485000  36.490000 ;
      RECT 37.385000  47.515000 38.275000  66.810000 ;
      RECT 37.385000  70.515000 38.275000  89.765000 ;
      RECT 37.385000  93.515000 38.275000 112.810000 ;
      RECT 37.385000 116.515000 38.275000 135.765000 ;
      RECT 37.385000 139.515000 38.275000 158.765000 ;
      RECT 37.385000 162.515000 38.275000 181.765000 ;
      RECT 37.385000 185.515000 38.275000 195.030000 ;
      RECT 38.095000  29.775000 38.265000  32.860000 ;
      RECT 38.780000 195.370000 39.490000 195.540000 ;
      RECT 38.875000  33.335000 39.045000  36.490000 ;
      RECT 39.655000  29.770000 39.825000  32.860000 ;
      RECT 40.435000  33.335000 40.605000  36.490000 ;
      RECT 40.790000 195.370000 41.500000 195.540000 ;
      RECT 41.215000  29.770000 41.385000  32.860000 ;
      RECT 41.985000  47.515000 42.875000  66.810000 ;
      RECT 41.985000  70.515000 42.875000  89.765000 ;
      RECT 41.985000  93.515000 42.875000 112.810000 ;
      RECT 41.985000 116.515000 42.875000 135.765000 ;
      RECT 41.985000 139.515000 42.875000 158.765000 ;
      RECT 41.985000 162.515000 42.875000 181.765000 ;
      RECT 41.985000 185.515000 42.875000 195.030000 ;
      RECT 41.995000  33.340000 42.165000  36.490000 ;
      RECT 42.775000  29.775000 42.945000  32.860000 ;
      RECT 43.380000 195.370000 44.090000 195.540000 ;
      RECT 43.555000  33.335000 43.725000  36.490000 ;
      RECT 44.335000  29.770000 44.505000  32.860000 ;
      RECT 45.115000  33.340000 45.285000  36.490000 ;
      RECT 45.390000 195.370000 46.100000 195.540000 ;
      RECT 45.755000  29.430000 45.955000  37.425000 ;
      RECT 46.585000  47.515000 47.475000  66.810000 ;
      RECT 46.585000  70.515000 47.475000  89.765000 ;
      RECT 46.585000  93.515000 47.475000 112.810000 ;
      RECT 46.585000 116.515000 47.475000 135.765000 ;
      RECT 46.585000 139.515000 47.475000 158.765000 ;
      RECT 46.585000 162.515000 47.475000 181.765000 ;
      RECT 46.585000 185.515000 47.475000 195.030000 ;
      RECT 47.310000  28.030000 48.200000  29.215000 ;
      RECT 47.310000  29.525000 48.200000  38.695000 ;
      RECT 47.330000  29.215000 48.180000  29.525000 ;
      RECT 47.980000 195.370000 48.690000 195.540000 ;
      RECT 49.990000 195.370000 50.700000 195.540000 ;
      RECT 51.185000  47.515000 52.075000  66.810000 ;
      RECT 51.185000  70.515000 52.075000  89.765000 ;
      RECT 51.185000  93.515000 52.075000 112.810000 ;
      RECT 51.185000 116.515000 52.075000 135.765000 ;
      RECT 51.185000 139.515000 52.075000 158.765000 ;
      RECT 51.185000 162.515000 52.075000 181.765000 ;
      RECT 51.185000 185.515000 52.075000 195.030000 ;
      RECT 52.320000  29.300000 68.865000  31.060000 ;
      RECT 52.320000  31.060000 53.210000  41.455000 ;
      RECT 52.320000  41.455000 68.865000  42.495000 ;
      RECT 52.580000 195.370000 53.290000 195.540000 ;
      RECT 53.960000  31.835000 67.140000  32.005000 ;
      RECT 53.960000  32.005000 54.130000  40.410000 ;
      RECT 53.960000  40.410000 67.140000  40.580000 ;
      RECT 54.590000 195.370000 55.300000 195.540000 ;
      RECT 54.695000  36.190000 54.865000  39.290000 ;
      RECT 54.940000  39.770000 66.335000  39.940000 ;
      RECT 55.215000  23.240000 56.105000  28.345000 ;
      RECT 55.215000  28.345000 70.630000  29.300000 ;
      RECT 55.465000  32.620000 55.635000  35.770000 ;
      RECT 55.785000  47.515000 56.675000  66.810000 ;
      RECT 55.785000  70.515000 56.675000  89.765000 ;
      RECT 55.785000  93.515000 56.675000 112.810000 ;
      RECT 55.785000 116.515000 56.675000 135.765000 ;
      RECT 55.785000 139.515000 56.675000 158.765000 ;
      RECT 55.785000 162.515000 56.675000 181.765000 ;
      RECT 55.785000 185.515000 56.675000 195.140000 ;
      RECT 56.255000  36.190000 56.425000  39.290000 ;
      RECT 56.820000  23.480000 57.050000  27.485000 ;
      RECT 56.820000  27.485000 62.810000  27.715000 ;
      RECT 56.850000  21.465000 57.020000  23.480000 ;
      RECT 57.025000  32.620000 57.195000  35.770000 ;
      RECT 57.180000 195.370000 57.890000 195.540000 ;
      RECT 57.555000  23.480000 57.785000  26.430000 ;
      RECT 57.815000  21.735000 61.815000  21.965000 ;
      RECT 57.815000  36.190000 57.985000  39.290000 ;
      RECT 58.585000  32.620000 58.755000  35.770000 ;
      RECT 59.190000 195.370000 59.900000 195.540000 ;
      RECT 59.375000  36.190000 59.545000  39.290000 ;
      RECT 60.145000  32.620000 60.315000  35.770000 ;
      RECT 60.385000  47.515000 61.275000  66.810000 ;
      RECT 60.385000  70.515000 61.275000  89.765000 ;
      RECT 60.385000  93.515000 61.275000 112.810000 ;
      RECT 60.385000 116.515000 61.275000 135.765000 ;
      RECT 60.385000 139.515000 61.275000 158.765000 ;
      RECT 60.385000 162.515000 61.275000 181.765000 ;
      RECT 60.385000 185.515000 61.275000 195.140000 ;
      RECT 60.935000  36.190000 61.105000  39.290000 ;
      RECT 61.705000  32.620000 61.875000  35.770000 ;
      RECT 61.780000 195.370000 62.490000 195.540000 ;
      RECT 61.850000  23.480000 62.080000  26.430000 ;
      RECT 62.495000  36.190000 62.665000  39.290000 ;
      RECT 62.580000  23.480000 62.810000  27.485000 ;
      RECT 62.610000  21.465000 62.780000  23.480000 ;
      RECT 63.265000  32.620000 63.435000  35.770000 ;
      RECT 63.790000 195.370000 64.500000 195.540000 ;
      RECT 64.055000  36.190000 64.225000  39.290000 ;
      RECT 64.825000  32.620000 64.995000  35.770000 ;
      RECT 64.845000  47.160000 65.875000  66.930000 ;
      RECT 64.845000  70.160000 65.875000  72.950000 ;
      RECT 64.845000  87.140000 65.875000  89.930000 ;
      RECT 64.845000  93.160000 65.875000  95.950000 ;
      RECT 64.845000 110.145000 65.875000 112.935000 ;
      RECT 64.845000 116.160000 65.875000 118.950000 ;
      RECT 64.845000 133.140000 65.875000 135.930000 ;
      RECT 64.845000 139.160000 65.875000 158.930000 ;
      RECT 64.845000 162.160000 65.875000 181.930000 ;
      RECT 64.845000 185.160000 65.875000 195.180000 ;
      RECT 64.985000  72.950000 65.875000  87.140000 ;
      RECT 64.985000  95.950000 65.875000 110.145000 ;
      RECT 64.985000 118.950000 65.875000 133.140000 ;
      RECT 65.615000  36.190000 65.785000  39.290000 ;
      RECT 66.385000  32.620000 66.555000  35.770000 ;
      RECT 66.935000  32.005000 67.140000  36.065000 ;
      RECT 66.935000  36.275000 67.140000  40.410000 ;
      RECT 66.970000  36.065000 67.140000  36.275000 ;
      RECT 67.265000  46.350000 68.155000 101.315000 ;
      RECT 67.265000 166.045000 68.155000 196.835000 ;
      RECT 67.290000 101.315000 68.140000 101.710000 ;
      RECT 67.290000 101.710000 68.155000 165.645000 ;
      RECT 67.290000 165.645000 68.140000 166.045000 ;
      RECT 67.975000  31.060000 68.865000  40.480000 ;
      RECT 67.975000  41.315000 68.865000  41.455000 ;
      RECT 68.000000  40.480000 68.830000  41.315000 ;
      RECT 68.875000  44.755000 70.125000  45.995000 ;
      RECT 68.875000  46.185000 70.125000 198.445000 ;
      RECT 68.905000  45.995000 70.095000  46.185000 ;
      RECT 69.740000  22.520000 70.630000  28.345000 ;
      RECT 69.760000   1.890000 70.650000   2.770000 ;
      RECT 69.765000   3.845000 70.630000   8.915000 ;
      RECT 69.765000   9.845000 70.630000  14.915000 ;
      RECT 69.765000  16.165000 70.630000  21.235000 ;
      RECT 69.780000   2.770000 70.630000   3.845000 ;
      RECT 69.780000   8.915000 70.630000   9.845000 ;
      RECT 69.780000  14.915000 70.630000  16.165000 ;
      RECT 69.780000  21.235000 70.630000  22.520000 ;
      RECT 70.470000  42.820000 71.055000  42.990000 ;
      RECT 70.725000  42.735000 71.055000  42.820000 ;
      RECT 72.245000 199.210000 72.775000 199.380000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 75.000000 200.000000 ;
    LAYER met2 ;
      RECT  0.000000   0.000000  0.215000   2.170000 ;
      RECT  0.000000   0.000000  0.215000   2.170000 ;
      RECT  0.000000   2.170000  0.215000   2.240000 ;
      RECT  0.000000   2.170000  0.725000   2.680000 ;
      RECT  0.000000   2.240000  0.285000   2.310000 ;
      RECT  0.000000   2.310000  0.355000   2.380000 ;
      RECT  0.000000   2.380000  0.425000   2.450000 ;
      RECT  0.000000   2.450000  0.495000   2.520000 ;
      RECT  0.000000   2.520000  0.565000   2.590000 ;
      RECT  0.000000   2.590000  0.635000   2.660000 ;
      RECT  0.000000   2.660000  0.705000   2.680000 ;
      RECT  0.000000   2.680000  0.725000  36.755000 ;
      RECT  0.000000   2.680000  0.725000  36.755000 ;
      RECT  0.000000  36.755000  0.725000  36.800000 ;
      RECT  0.000000  36.755000  0.810000  36.840000 ;
      RECT  0.000000  36.800000  0.770000  36.840000 ;
      RECT  0.000000  36.840000  0.810000  46.930000 ;
      RECT  0.000000  36.840000  0.810000  46.930000 ;
      RECT  0.000000  46.930000  0.725000  47.015000 ;
      RECT  0.000000  46.930000  0.770000  46.970000 ;
      RECT  0.000000  46.970000  0.730000  47.010000 ;
      RECT  0.000000  47.010000  0.725000  47.015000 ;
      RECT  0.000000  47.015000  0.725000 195.355000 ;
      RECT  0.000000  47.015000  0.725000 195.355000 ;
      RECT  0.000000 195.355000 67.480000 200.000000 ;
      RECT  0.000000 195.355000 75.000000 200.000000 ;
      RECT 14.400000  45.430000 57.415000  47.315000 ;
      RECT 14.400000  45.430000 59.035000  45.500000 ;
      RECT 14.400000  45.430000 59.035000  45.500000 ;
      RECT 14.400000  45.500000 58.965000  45.570000 ;
      RECT 14.400000  45.500000 58.965000  45.570000 ;
      RECT 14.400000  45.570000 58.895000  45.640000 ;
      RECT 14.400000  45.570000 58.895000  45.640000 ;
      RECT 14.400000  45.640000 58.825000  45.710000 ;
      RECT 14.400000  45.640000 58.825000  45.710000 ;
      RECT 14.400000  45.710000 58.755000  45.780000 ;
      RECT 14.400000  45.710000 58.755000  45.780000 ;
      RECT 14.400000  45.780000 58.685000  45.850000 ;
      RECT 14.400000  45.780000 58.685000  45.850000 ;
      RECT 14.400000  45.850000 58.615000  45.920000 ;
      RECT 14.400000  45.850000 58.615000  45.920000 ;
      RECT 14.400000  45.920000 58.545000  45.990000 ;
      RECT 14.400000  45.920000 58.545000  45.990000 ;
      RECT 14.400000  45.990000 58.475000  46.060000 ;
      RECT 14.400000  45.990000 58.475000  46.060000 ;
      RECT 14.400000  46.060000 58.405000  46.130000 ;
      RECT 14.400000  46.060000 58.405000  46.130000 ;
      RECT 14.400000  46.130000 58.335000  46.200000 ;
      RECT 14.400000  46.130000 58.335000  46.200000 ;
      RECT 14.400000  46.200000 58.265000  46.270000 ;
      RECT 14.400000  46.200000 58.265000  46.270000 ;
      RECT 14.400000  46.270000 58.195000  46.340000 ;
      RECT 14.400000  46.270000 58.195000  46.340000 ;
      RECT 14.400000  46.340000 58.125000  46.410000 ;
      RECT 14.400000  46.340000 58.125000  46.410000 ;
      RECT 14.400000  46.410000 58.055000  46.480000 ;
      RECT 14.400000  46.410000 58.055000  46.480000 ;
      RECT 14.400000  46.480000 57.985000  46.550000 ;
      RECT 14.400000  46.480000 57.985000  46.550000 ;
      RECT 14.400000  46.550000 57.915000  46.620000 ;
      RECT 14.400000  46.550000 57.915000  46.620000 ;
      RECT 14.400000  46.620000 57.845000  46.690000 ;
      RECT 14.400000  46.620000 57.845000  46.690000 ;
      RECT 14.400000  46.690000 57.775000  46.760000 ;
      RECT 14.400000  46.690000 57.775000  46.760000 ;
      RECT 14.400000  46.760000 57.705000  46.830000 ;
      RECT 14.400000  46.760000 57.705000  46.830000 ;
      RECT 14.400000  46.830000 57.635000  46.900000 ;
      RECT 14.400000  46.830000 57.635000  46.900000 ;
      RECT 14.400000  46.900000 57.565000  46.970000 ;
      RECT 14.400000  46.900000 57.565000  46.970000 ;
      RECT 14.400000  46.970000 57.495000  47.040000 ;
      RECT 14.400000  46.970000 57.495000  47.040000 ;
      RECT 14.400000  47.040000 57.425000  47.110000 ;
      RECT 14.400000  47.040000 57.425000  47.110000 ;
      RECT 14.400000  47.110000 57.360000  47.175000 ;
      RECT 14.400000  47.110000 57.360000  47.175000 ;
      RECT 14.400000  47.175000 16.525000  54.100000 ;
      RECT 14.400000  47.315000 16.665000  54.100000 ;
      RECT 14.400000  54.100000 16.665000  54.905000 ;
      RECT 14.400000  70.140000 57.405000  70.160000 ;
      RECT 14.400000  70.140000 57.405000  70.160000 ;
      RECT 14.400000  70.140000 57.445000  70.315000 ;
      RECT 14.400000  70.160000 57.390000  70.175000 ;
      RECT 14.400000  70.160000 57.390000  70.175000 ;
      RECT 14.400000  70.175000 24.540000  72.870000 ;
      RECT 14.400000  70.315000 24.680000  72.925000 ;
      RECT 14.400000  72.870000 24.470000  72.940000 ;
      RECT 14.400000  72.870000 24.470000  72.940000 ;
      RECT 14.400000  72.925000 23.590000  74.015000 ;
      RECT 14.400000  72.940000 24.400000  73.010000 ;
      RECT 14.400000  72.940000 24.400000  73.010000 ;
      RECT 14.400000  73.010000 24.330000  73.080000 ;
      RECT 14.400000  73.010000 24.330000  73.080000 ;
      RECT 14.400000  73.080000 24.260000  73.150000 ;
      RECT 14.400000  73.080000 24.260000  73.150000 ;
      RECT 14.400000  73.150000 24.190000  73.220000 ;
      RECT 14.400000  73.150000 24.190000  73.220000 ;
      RECT 14.400000  73.220000 24.120000  73.290000 ;
      RECT 14.400000  73.220000 24.120000  73.290000 ;
      RECT 14.400000  73.290000 24.050000  73.360000 ;
      RECT 14.400000  73.290000 24.050000  73.360000 ;
      RECT 14.400000  73.360000 23.980000  73.430000 ;
      RECT 14.400000  73.360000 23.980000  73.430000 ;
      RECT 14.400000  73.430000 23.910000  73.500000 ;
      RECT 14.400000  73.430000 23.910000  73.500000 ;
      RECT 14.400000  73.500000 23.840000  73.570000 ;
      RECT 14.400000  73.500000 23.840000  73.570000 ;
      RECT 14.400000  73.570000 23.770000  73.640000 ;
      RECT 14.400000  73.570000 23.770000  73.640000 ;
      RECT 14.400000  73.640000 23.700000  73.710000 ;
      RECT 14.400000  73.640000 23.700000  73.710000 ;
      RECT 14.400000  73.710000 23.630000  73.780000 ;
      RECT 14.400000  73.710000 23.630000  73.780000 ;
      RECT 14.400000  73.780000 23.560000  73.850000 ;
      RECT 14.400000  73.780000 23.560000  73.850000 ;
      RECT 14.400000  73.850000 23.535000  73.875000 ;
      RECT 14.400000  73.850000 23.535000  73.875000 ;
      RECT 14.400000  73.875000 18.130000  74.695000 ;
      RECT 14.400000  74.015000 18.270000  74.555000 ;
      RECT 14.400000  74.555000 24.680000  75.675000 ;
      RECT 14.400000  74.695000 23.505000  74.765000 ;
      RECT 14.400000  74.695000 23.505000  74.765000 ;
      RECT 14.400000  74.765000 23.575000  74.835000 ;
      RECT 14.400000  74.765000 23.575000  74.835000 ;
      RECT 14.400000  74.835000 23.645000  74.905000 ;
      RECT 14.400000  74.835000 23.645000  74.905000 ;
      RECT 14.400000  74.905000 23.715000  74.975000 ;
      RECT 14.400000  74.905000 23.715000  74.975000 ;
      RECT 14.400000  74.975000 23.785000  75.045000 ;
      RECT 14.400000  74.975000 23.785000  75.045000 ;
      RECT 14.400000  75.045000 23.855000  75.115000 ;
      RECT 14.400000  75.045000 23.855000  75.115000 ;
      RECT 14.400000  75.115000 23.925000  75.185000 ;
      RECT 14.400000  75.115000 23.925000  75.185000 ;
      RECT 14.400000  75.185000 23.995000  75.255000 ;
      RECT 14.400000  75.185000 23.995000  75.255000 ;
      RECT 14.400000  75.255000 24.065000  75.325000 ;
      RECT 14.400000  75.255000 24.065000  75.325000 ;
      RECT 14.400000  75.325000 24.135000  75.395000 ;
      RECT 14.400000  75.325000 24.135000  75.395000 ;
      RECT 14.400000  75.395000 24.205000  75.465000 ;
      RECT 14.400000  75.395000 24.205000  75.465000 ;
      RECT 14.400000  75.465000 24.275000  75.535000 ;
      RECT 14.400000  75.465000 24.275000  75.535000 ;
      RECT 14.400000  75.535000 24.345000  75.605000 ;
      RECT 14.400000  75.535000 24.345000  75.605000 ;
      RECT 14.400000  75.605000 24.415000  75.675000 ;
      RECT 14.400000  75.605000 24.415000  75.675000 ;
      RECT 14.400000  75.675000 24.485000  75.730000 ;
      RECT 14.400000  75.675000 24.485000  75.730000 ;
      RECT 14.400000  75.675000 24.680000  77.125000 ;
      RECT 14.400000  75.730000 24.540000  77.125000 ;
      RECT 14.400000  77.125000 24.680000  79.295000 ;
      RECT 14.400000  93.140000 57.465000  93.160000 ;
      RECT 14.400000  93.140000 57.465000  93.160000 ;
      RECT 14.400000  93.140000 57.505000  93.315000 ;
      RECT 14.400000  93.160000 57.450000  93.175000 ;
      RECT 14.400000  93.160000 57.450000  93.175000 ;
      RECT 14.400000  93.175000 24.540000 100.125000 ;
      RECT 14.400000  93.315000 24.680000 100.125000 ;
      RECT 14.400000 100.125000 24.680000 102.295000 ;
      RECT 14.400000 116.180000 24.540000 123.030000 ;
      RECT 14.400000 116.180000 57.415000 116.315000 ;
      RECT 14.400000 116.315000 24.680000 123.030000 ;
      RECT 14.400000 123.030000 24.680000 125.295000 ;
      RECT 14.400000 139.285000 16.525000 146.100000 ;
      RECT 14.400000 139.285000 57.450000 139.315000 ;
      RECT 14.400000 139.315000 16.665000 146.100000 ;
      RECT 14.400000 146.100000 16.665000 146.770000 ;
      RECT 14.400000 162.195000 16.525000 169.105000 ;
      RECT 14.400000 162.195000 57.465000 162.315000 ;
      RECT 14.400000 162.315000 16.665000 169.105000 ;
      RECT 14.400000 169.105000 16.665000 171.295000 ;
      RECT 14.400000 185.170000 15.340000 189.470000 ;
      RECT 14.400000 185.170000 15.480000 189.470000 ;
      RECT 14.400000 189.470000 15.480000 190.155000 ;
      RECT 14.405000 116.175000 24.540000 116.180000 ;
      RECT 14.405000 116.175000 24.540000 116.180000 ;
      RECT 14.410000 162.185000 16.525000 162.195000 ;
      RECT 14.415000 185.155000 15.340000 185.170000 ;
      RECT 14.415000 185.155000 15.480000 185.170000 ;
      RECT 14.420000  70.120000 57.425000  70.140000 ;
      RECT 14.420000  70.120000 57.425000  70.140000 ;
      RECT 14.420000 162.175000 16.525000 162.185000 ;
      RECT 14.445000  45.385000 59.105000  45.430000 ;
      RECT 14.445000  45.385000 59.105000  45.430000 ;
      RECT 14.455000  93.085000 57.485000  93.140000 ;
      RECT 14.455000  93.085000 57.485000  93.140000 ;
      RECT 14.455000 139.230000 16.525000 139.285000 ;
      RECT 14.460000 116.120000 57.360000 116.175000 ;
      RECT 14.460000 116.120000 57.360000 116.175000 ;
      RECT 14.470000  54.100000 16.525000  54.170000 ;
      RECT 14.470000  77.125000 24.540000  77.195000 ;
      RECT 14.470000  77.125000 24.540000  77.195000 ;
      RECT 14.470000 100.125000 24.540000 100.195000 ;
      RECT 14.470000 100.125000 24.540000 100.195000 ;
      RECT 14.470000 123.030000 24.540000 123.100000 ;
      RECT 14.470000 123.030000 24.540000 123.100000 ;
      RECT 14.470000 146.100000 16.525000 146.170000 ;
      RECT 14.470000 169.105000 16.525000 169.175000 ;
      RECT 14.470000 189.470000 15.340000 189.540000 ;
      RECT 14.475000 162.120000 57.410000 162.175000 ;
      RECT 14.475000 162.120000 57.410000 162.175000 ;
      RECT 14.485000 185.085000 15.340000 185.155000 ;
      RECT 14.490000  70.050000 57.445000  70.120000 ;
      RECT 14.490000  70.050000 57.445000  70.120000 ;
      RECT 14.510000 139.175000 16.525000 139.230000 ;
      RECT 14.515000  45.315000 59.150000  45.385000 ;
      RECT 14.515000  45.315000 59.150000  45.385000 ;
      RECT 14.525000  93.015000 57.540000  93.085000 ;
      RECT 14.525000  93.015000 57.540000  93.085000 ;
      RECT 14.530000 116.050000 57.415000 116.120000 ;
      RECT 14.530000 116.050000 57.415000 116.120000 ;
      RECT 14.540000  54.170000 16.525000  54.240000 ;
      RECT 14.540000  77.195000 24.540000  77.265000 ;
      RECT 14.540000  77.195000 24.540000  77.265000 ;
      RECT 14.540000 100.195000 24.540000 100.265000 ;
      RECT 14.540000 100.195000 24.540000 100.265000 ;
      RECT 14.540000 123.100000 24.540000 123.170000 ;
      RECT 14.540000 123.100000 24.540000 123.170000 ;
      RECT 14.540000 146.170000 16.525000 146.240000 ;
      RECT 14.540000 169.175000 16.525000 169.245000 ;
      RECT 14.540000 189.540000 15.340000 189.610000 ;
      RECT 14.545000 162.050000 57.465000 162.120000 ;
      RECT 14.545000 162.050000 57.465000 162.120000 ;
      RECT 14.555000 185.015000 15.340000 185.085000 ;
      RECT 14.560000  69.980000 57.515000  70.050000 ;
      RECT 14.560000  69.980000 57.515000  70.050000 ;
      RECT 14.565000 139.120000 57.395000 139.175000 ;
      RECT 14.565000 139.120000 57.395000 139.175000 ;
      RECT 14.565000 185.005000 58.580000 185.015000 ;
      RECT 14.585000  45.245000 59.220000  45.315000 ;
      RECT 14.585000  45.245000 59.220000  45.315000 ;
      RECT 14.595000  92.945000 57.610000  93.015000 ;
      RECT 14.595000  92.945000 57.610000  93.015000 ;
      RECT 14.600000 115.980000 57.485000 116.050000 ;
      RECT 14.600000 115.980000 57.485000 116.050000 ;
      RECT 14.610000  54.240000 16.525000  54.310000 ;
      RECT 14.610000  77.265000 24.540000  77.335000 ;
      RECT 14.610000  77.265000 24.540000  77.335000 ;
      RECT 14.610000 100.265000 24.540000 100.335000 ;
      RECT 14.610000 100.265000 24.540000 100.335000 ;
      RECT 14.610000 123.170000 24.540000 123.240000 ;
      RECT 14.610000 123.170000 24.540000 123.240000 ;
      RECT 14.610000 146.240000 16.525000 146.310000 ;
      RECT 14.610000 169.245000 16.525000 169.315000 ;
      RECT 14.610000 189.610000 15.340000 189.680000 ;
      RECT 14.615000 161.980000 57.535000 162.050000 ;
      RECT 14.615000 161.980000 57.535000 162.050000 ;
      RECT 14.630000  69.910000 57.585000  69.980000 ;
      RECT 14.630000  69.910000 57.585000  69.980000 ;
      RECT 14.635000 139.050000 57.450000 139.120000 ;
      RECT 14.635000 139.050000 57.450000 139.120000 ;
      RECT 14.635000 184.935000 58.590000 185.005000 ;
      RECT 14.655000  45.175000 59.290000  45.245000 ;
      RECT 14.655000  45.175000 59.290000  45.245000 ;
      RECT 14.665000  92.875000 57.680000  92.945000 ;
      RECT 14.665000  92.875000 57.680000  92.945000 ;
      RECT 14.670000 115.910000 57.555000 115.980000 ;
      RECT 14.670000 115.910000 57.555000 115.980000 ;
      RECT 14.680000  54.310000 16.525000  54.380000 ;
      RECT 14.680000  77.335000 24.540000  77.405000 ;
      RECT 14.680000  77.335000 24.540000  77.405000 ;
      RECT 14.680000 100.335000 24.540000 100.405000 ;
      RECT 14.680000 100.335000 24.540000 100.405000 ;
      RECT 14.680000 123.240000 24.540000 123.310000 ;
      RECT 14.680000 123.240000 24.540000 123.310000 ;
      RECT 14.680000 146.310000 16.525000 146.380000 ;
      RECT 14.680000 169.315000 16.525000 169.385000 ;
      RECT 14.680000 189.680000 15.340000 189.750000 ;
      RECT 14.685000 161.910000 57.605000 161.980000 ;
      RECT 14.685000 161.910000 57.605000 161.980000 ;
      RECT 14.700000  69.840000 57.655000  69.910000 ;
      RECT 14.700000  69.840000 57.655000  69.910000 ;
      RECT 14.705000 138.980000 57.520000 139.050000 ;
      RECT 14.705000 138.980000 57.520000 139.050000 ;
      RECT 14.705000 184.865000 58.660000 184.935000 ;
      RECT 14.725000  45.105000 59.360000  45.175000 ;
      RECT 14.725000  45.105000 59.360000  45.175000 ;
      RECT 14.735000  92.805000 57.750000  92.875000 ;
      RECT 14.735000  92.805000 57.750000  92.875000 ;
      RECT 14.740000 115.840000 57.625000 115.910000 ;
      RECT 14.740000 115.840000 57.625000 115.910000 ;
      RECT 14.750000  54.380000 16.525000  54.450000 ;
      RECT 14.750000  77.405000 24.540000  77.475000 ;
      RECT 14.750000  77.405000 24.540000  77.475000 ;
      RECT 14.750000 100.405000 24.540000 100.475000 ;
      RECT 14.750000 100.405000 24.540000 100.475000 ;
      RECT 14.750000 123.310000 24.540000 123.380000 ;
      RECT 14.750000 123.310000 24.540000 123.380000 ;
      RECT 14.750000 146.380000 16.525000 146.450000 ;
      RECT 14.750000 169.385000 16.525000 169.455000 ;
      RECT 14.750000 189.750000 15.340000 189.820000 ;
      RECT 14.755000 161.840000 57.675000 161.910000 ;
      RECT 14.755000 161.840000 57.675000 161.910000 ;
      RECT 14.770000  69.770000 57.725000  69.840000 ;
      RECT 14.770000  69.770000 57.725000  69.840000 ;
      RECT 14.775000 138.910000 57.590000 138.980000 ;
      RECT 14.775000 138.910000 57.590000 138.980000 ;
      RECT 14.775000 184.795000 58.730000 184.865000 ;
      RECT 14.795000  45.035000 59.430000  45.105000 ;
      RECT 14.795000  45.035000 59.430000  45.105000 ;
      RECT 14.805000  92.735000 57.820000  92.805000 ;
      RECT 14.805000  92.735000 57.820000  92.805000 ;
      RECT 14.810000 115.770000 57.695000 115.840000 ;
      RECT 14.810000 115.770000 57.695000 115.840000 ;
      RECT 14.820000  54.450000 16.525000  54.520000 ;
      RECT 14.820000  77.475000 24.540000  77.545000 ;
      RECT 14.820000  77.475000 24.540000  77.545000 ;
      RECT 14.820000 100.475000 24.540000 100.545000 ;
      RECT 14.820000 100.475000 24.540000 100.545000 ;
      RECT 14.820000 123.380000 24.540000 123.450000 ;
      RECT 14.820000 123.380000 24.540000 123.450000 ;
      RECT 14.820000 146.450000 16.525000 146.520000 ;
      RECT 14.820000 169.455000 16.525000 169.525000 ;
      RECT 14.820000 189.820000 15.340000 189.890000 ;
      RECT 14.825000 161.770000 57.745000 161.840000 ;
      RECT 14.825000 161.770000 57.745000 161.840000 ;
      RECT 14.840000  69.700000 57.795000  69.770000 ;
      RECT 14.840000  69.700000 57.795000  69.770000 ;
      RECT 14.845000 138.840000 57.660000 138.910000 ;
      RECT 14.845000 138.840000 57.660000 138.910000 ;
      RECT 14.845000 184.725000 58.800000 184.795000 ;
      RECT 14.865000  44.965000 59.500000  45.035000 ;
      RECT 14.865000  44.965000 59.500000  45.035000 ;
      RECT 14.875000  92.665000 57.890000  92.735000 ;
      RECT 14.875000  92.665000 57.890000  92.735000 ;
      RECT 14.880000 115.700000 57.765000 115.770000 ;
      RECT 14.880000 115.700000 57.765000 115.770000 ;
      RECT 14.890000  54.520000 16.525000  54.590000 ;
      RECT 14.890000  77.545000 24.540000  77.615000 ;
      RECT 14.890000  77.545000 24.540000  77.615000 ;
      RECT 14.890000 100.545000 24.540000 100.615000 ;
      RECT 14.890000 100.545000 24.540000 100.615000 ;
      RECT 14.890000 123.450000 24.540000 123.520000 ;
      RECT 14.890000 123.450000 24.540000 123.520000 ;
      RECT 14.890000 146.520000 16.525000 146.590000 ;
      RECT 14.890000 169.525000 16.525000 169.595000 ;
      RECT 14.890000 189.890000 15.340000 189.960000 ;
      RECT 14.895000 161.700000 57.815000 161.770000 ;
      RECT 14.895000 161.700000 57.815000 161.770000 ;
      RECT 14.910000  69.630000 57.865000  69.700000 ;
      RECT 14.910000  69.630000 57.865000  69.700000 ;
      RECT 14.915000 138.770000 57.730000 138.840000 ;
      RECT 14.915000 138.770000 57.730000 138.840000 ;
      RECT 14.915000 184.655000 58.870000 184.725000 ;
      RECT 14.935000  44.895000 59.570000  44.965000 ;
      RECT 14.935000  44.895000 59.570000  44.965000 ;
      RECT 14.945000  92.595000 57.960000  92.665000 ;
      RECT 14.945000  92.595000 57.960000  92.665000 ;
      RECT 14.950000 115.630000 57.835000 115.700000 ;
      RECT 14.950000 115.630000 57.835000 115.700000 ;
      RECT 14.960000  54.590000 16.525000  54.660000 ;
      RECT 14.960000  77.615000 24.540000  77.685000 ;
      RECT 14.960000  77.615000 24.540000  77.685000 ;
      RECT 14.960000 100.615000 24.540000 100.685000 ;
      RECT 14.960000 100.615000 24.540000 100.685000 ;
      RECT 14.960000 123.520000 24.540000 123.590000 ;
      RECT 14.960000 123.520000 24.540000 123.590000 ;
      RECT 14.960000 146.590000 16.525000 146.660000 ;
      RECT 14.960000 169.595000 16.525000 169.665000 ;
      RECT 14.960000 189.960000 15.340000 190.030000 ;
      RECT 14.965000 161.630000 57.885000 161.700000 ;
      RECT 14.965000 161.630000 57.885000 161.700000 ;
      RECT 14.980000  69.560000 57.935000  69.630000 ;
      RECT 14.980000  69.560000 57.935000  69.630000 ;
      RECT 14.985000 138.700000 57.800000 138.770000 ;
      RECT 14.985000 138.700000 57.800000 138.770000 ;
      RECT 14.985000 184.585000 58.940000 184.655000 ;
      RECT 15.005000  44.825000 59.640000  44.895000 ;
      RECT 15.005000  44.825000 59.640000  44.895000 ;
      RECT 15.015000  92.525000 58.030000  92.595000 ;
      RECT 15.015000  92.525000 58.030000  92.595000 ;
      RECT 15.020000 115.560000 57.905000 115.630000 ;
      RECT 15.020000 115.560000 57.905000 115.630000 ;
      RECT 15.030000  54.660000 16.525000  54.730000 ;
      RECT 15.030000  77.685000 24.540000  77.755000 ;
      RECT 15.030000  77.685000 24.540000  77.755000 ;
      RECT 15.030000 100.685000 24.540000 100.755000 ;
      RECT 15.030000 100.685000 24.540000 100.755000 ;
      RECT 15.030000 123.590000 24.540000 123.660000 ;
      RECT 15.030000 123.590000 24.540000 123.660000 ;
      RECT 15.030000 146.660000 16.525000 146.730000 ;
      RECT 15.030000 169.665000 16.525000 169.735000 ;
      RECT 15.030000 190.030000 15.340000 190.100000 ;
      RECT 15.035000 161.560000 57.955000 161.630000 ;
      RECT 15.035000 161.560000 57.955000 161.630000 ;
      RECT 15.050000  69.490000 58.005000  69.560000 ;
      RECT 15.050000  69.490000 58.005000  69.560000 ;
      RECT 15.055000 138.630000 57.870000 138.700000 ;
      RECT 15.055000 138.630000 57.870000 138.700000 ;
      RECT 15.055000 184.515000 59.010000 184.585000 ;
      RECT 15.070000 146.770000 18.190000 148.295000 ;
      RECT 15.075000  44.755000 59.710000  44.825000 ;
      RECT 15.075000  44.755000 59.710000  44.825000 ;
      RECT 15.085000  92.455000 58.100000  92.525000 ;
      RECT 15.085000  92.455000 58.100000  92.525000 ;
      RECT 15.085000 190.155000 75.000000 190.280000 ;
      RECT 15.090000 115.490000 57.975000 115.560000 ;
      RECT 15.090000 115.490000 57.975000 115.560000 ;
      RECT 15.100000  54.730000 16.525000  54.800000 ;
      RECT 15.100000  77.755000 24.540000  77.825000 ;
      RECT 15.100000  77.755000 24.540000  77.825000 ;
      RECT 15.100000 100.755000 24.540000 100.825000 ;
      RECT 15.100000 100.755000 24.540000 100.825000 ;
      RECT 15.100000 123.660000 24.540000 123.730000 ;
      RECT 15.100000 123.660000 24.540000 123.730000 ;
      RECT 15.100000 146.730000 16.525000 146.800000 ;
      RECT 15.100000 169.735000 16.525000 169.805000 ;
      RECT 15.100000 190.100000 15.340000 190.170000 ;
      RECT 15.105000 161.490000 58.025000 161.560000 ;
      RECT 15.105000 161.490000 58.025000 161.560000 ;
      RECT 15.120000  69.420000 58.075000  69.490000 ;
      RECT 15.120000  69.420000 58.075000  69.490000 ;
      RECT 15.125000 138.560000 57.940000 138.630000 ;
      RECT 15.125000 138.560000 57.940000 138.630000 ;
      RECT 15.125000 146.800000 16.525000 146.825000 ;
      RECT 15.125000 184.445000 59.080000 184.515000 ;
      RECT 15.145000  44.685000 59.780000  44.755000 ;
      RECT 15.145000  44.685000 59.780000  44.755000 ;
      RECT 15.155000  92.385000 58.170000  92.455000 ;
      RECT 15.155000  92.385000 58.170000  92.455000 ;
      RECT 15.160000 115.420000 58.045000 115.490000 ;
      RECT 15.160000 115.420000 58.045000 115.490000 ;
      RECT 15.170000  54.800000 16.525000  54.870000 ;
      RECT 15.170000  77.825000 24.540000  77.895000 ;
      RECT 15.170000  77.825000 24.540000  77.895000 ;
      RECT 15.170000 100.825000 24.540000 100.895000 ;
      RECT 15.170000 100.825000 24.540000 100.895000 ;
      RECT 15.170000 123.730000 24.540000 123.800000 ;
      RECT 15.170000 123.730000 24.540000 123.800000 ;
      RECT 15.170000 169.805000 16.525000 169.875000 ;
      RECT 15.170000 190.170000 15.340000 190.240000 ;
      RECT 15.175000 161.420000 58.095000 161.490000 ;
      RECT 15.175000 161.420000 58.095000 161.490000 ;
      RECT 15.190000  69.350000 58.145000  69.420000 ;
      RECT 15.190000  69.350000 58.145000  69.420000 ;
      RECT 15.195000 138.490000 58.010000 138.560000 ;
      RECT 15.195000 138.490000 58.010000 138.560000 ;
      RECT 15.195000 146.825000 16.525000 146.895000 ;
      RECT 15.195000 184.375000 59.150000 184.445000 ;
      RECT 15.205000  54.905000 18.790000  56.295000 ;
      RECT 15.210000 190.240000 15.340000 190.280000 ;
      RECT 15.215000  44.615000 59.850000  44.685000 ;
      RECT 15.215000  44.615000 59.850000  44.685000 ;
      RECT 15.225000  92.315000 58.240000  92.385000 ;
      RECT 15.225000  92.315000 58.240000  92.385000 ;
      RECT 15.230000 115.350000 58.115000 115.420000 ;
      RECT 15.230000 115.350000 58.115000 115.420000 ;
      RECT 15.240000  54.870000 16.525000  54.940000 ;
      RECT 15.240000  77.895000 24.540000  77.965000 ;
      RECT 15.240000  77.895000 24.540000  77.965000 ;
      RECT 15.240000 100.895000 24.540000 100.965000 ;
      RECT 15.240000 100.895000 24.540000 100.965000 ;
      RECT 15.240000 123.800000 24.540000 123.870000 ;
      RECT 15.240000 123.800000 24.540000 123.870000 ;
      RECT 15.240000 169.875000 16.525000 169.945000 ;
      RECT 15.245000 161.350000 58.165000 161.420000 ;
      RECT 15.245000 161.350000 58.165000 161.420000 ;
      RECT 15.260000  69.280000 58.215000  69.350000 ;
      RECT 15.260000  69.280000 58.215000  69.350000 ;
      RECT 15.265000 138.420000 58.080000 138.490000 ;
      RECT 15.265000 138.420000 58.080000 138.490000 ;
      RECT 15.265000 146.895000 16.595000 146.965000 ;
      RECT 15.265000 184.305000 59.220000 184.375000 ;
      RECT 15.285000  44.545000 59.920000  44.615000 ;
      RECT 15.285000  44.545000 59.920000  44.615000 ;
      RECT 15.295000  92.245000 58.310000  92.315000 ;
      RECT 15.295000  92.245000 58.310000  92.315000 ;
      RECT 15.300000 115.280000 58.185000 115.350000 ;
      RECT 15.300000 115.280000 58.185000 115.350000 ;
      RECT 15.310000  54.940000 16.525000  55.010000 ;
      RECT 15.310000  77.965000 24.540000  78.035000 ;
      RECT 15.310000  77.965000 24.540000  78.035000 ;
      RECT 15.310000 100.965000 24.540000 101.035000 ;
      RECT 15.310000 100.965000 24.540000 101.035000 ;
      RECT 15.310000 123.870000 24.540000 123.940000 ;
      RECT 15.310000 123.870000 24.540000 123.940000 ;
      RECT 15.310000 169.945000 16.525000 170.015000 ;
      RECT 15.315000 161.280000 58.235000 161.350000 ;
      RECT 15.315000 161.280000 58.235000 161.350000 ;
      RECT 15.330000  69.210000 58.285000  69.280000 ;
      RECT 15.330000  69.210000 58.285000  69.280000 ;
      RECT 15.335000 138.350000 58.150000 138.420000 ;
      RECT 15.335000 138.350000 58.150000 138.420000 ;
      RECT 15.335000 146.965000 16.665000 147.035000 ;
      RECT 15.335000 184.235000 59.290000 184.305000 ;
      RECT 15.345000  55.010000 16.525000  55.045000 ;
      RECT 15.355000  44.475000 59.990000  44.545000 ;
      RECT 15.355000  44.475000 59.990000  44.545000 ;
      RECT 15.365000  92.175000 58.380000  92.245000 ;
      RECT 15.365000  92.175000 58.380000  92.245000 ;
      RECT 15.370000 115.210000 58.255000 115.280000 ;
      RECT 15.370000 115.210000 58.255000 115.280000 ;
      RECT 15.380000  78.035000 24.540000  78.105000 ;
      RECT 15.380000  78.035000 24.540000  78.105000 ;
      RECT 15.380000 101.035000 24.540000 101.105000 ;
      RECT 15.380000 101.035000 24.540000 101.105000 ;
      RECT 15.380000 123.940000 24.540000 124.010000 ;
      RECT 15.380000 123.940000 24.540000 124.010000 ;
      RECT 15.380000 170.015000 16.525000 170.085000 ;
      RECT 15.385000 161.210000 58.305000 161.280000 ;
      RECT 15.385000 161.210000 58.305000 161.280000 ;
      RECT 15.400000  69.140000 58.355000  69.210000 ;
      RECT 15.400000  69.140000 58.355000  69.210000 ;
      RECT 15.405000 138.280000 58.220000 138.350000 ;
      RECT 15.405000 138.280000 58.220000 138.350000 ;
      RECT 15.405000 147.035000 16.735000 147.105000 ;
      RECT 15.405000 184.165000 59.360000 184.235000 ;
      RECT 15.415000  55.045000 17.345000  55.115000 ;
      RECT 15.425000  44.405000 60.060000  44.475000 ;
      RECT 15.425000  44.405000 60.060000  44.475000 ;
      RECT 15.435000  92.105000 58.450000  92.175000 ;
      RECT 15.435000  92.105000 58.450000  92.175000 ;
      RECT 15.440000 115.140000 58.325000 115.210000 ;
      RECT 15.440000 115.140000 58.325000 115.210000 ;
      RECT 15.450000  78.105000 24.540000  78.175000 ;
      RECT 15.450000  78.105000 24.540000  78.175000 ;
      RECT 15.450000 101.105000 24.540000 101.175000 ;
      RECT 15.450000 101.105000 24.540000 101.175000 ;
      RECT 15.450000 124.010000 24.540000 124.080000 ;
      RECT 15.450000 124.010000 24.540000 124.080000 ;
      RECT 15.450000 170.085000 16.525000 170.155000 ;
      RECT 15.455000 161.140000 58.375000 161.210000 ;
      RECT 15.455000 161.140000 58.375000 161.210000 ;
      RECT 15.470000  69.070000 58.425000  69.140000 ;
      RECT 15.470000  69.070000 58.425000  69.140000 ;
      RECT 15.475000 138.210000 58.290000 138.280000 ;
      RECT 15.475000 138.210000 58.290000 138.280000 ;
      RECT 15.475000 147.105000 16.805000 147.175000 ;
      RECT 15.475000 184.095000 59.430000 184.165000 ;
      RECT 15.485000  29.430000 59.190000  29.500000 ;
      RECT 15.485000  29.430000 59.190000  29.500000 ;
      RECT 15.485000  29.430000 60.970000  31.015000 ;
      RECT 15.485000  29.500000 59.260000  29.570000 ;
      RECT 15.485000  29.500000 59.260000  29.570000 ;
      RECT 15.485000  29.570000 59.330000  29.640000 ;
      RECT 15.485000  29.570000 59.330000  29.640000 ;
      RECT 15.485000  29.640000 59.400000  29.710000 ;
      RECT 15.485000  29.640000 59.400000  29.710000 ;
      RECT 15.485000  29.710000 59.470000  29.780000 ;
      RECT 15.485000  29.710000 59.470000  29.780000 ;
      RECT 15.485000  29.780000 59.540000  29.850000 ;
      RECT 15.485000  29.780000 59.540000  29.850000 ;
      RECT 15.485000  29.850000 59.610000  29.920000 ;
      RECT 15.485000  29.850000 59.610000  29.920000 ;
      RECT 15.485000  29.920000 59.680000  29.990000 ;
      RECT 15.485000  29.920000 59.680000  29.990000 ;
      RECT 15.485000  29.990000 59.750000  30.060000 ;
      RECT 15.485000  29.990000 59.750000  30.060000 ;
      RECT 15.485000  30.060000 59.820000  30.130000 ;
      RECT 15.485000  30.060000 59.820000  30.130000 ;
      RECT 15.485000  30.130000 59.890000  30.200000 ;
      RECT 15.485000  30.130000 59.890000  30.200000 ;
      RECT 15.485000  30.200000 59.960000  30.270000 ;
      RECT 15.485000  30.200000 59.960000  30.270000 ;
      RECT 15.485000  30.270000 60.030000  30.340000 ;
      RECT 15.485000  30.270000 60.030000  30.340000 ;
      RECT 15.485000  30.340000 60.100000  30.410000 ;
      RECT 15.485000  30.340000 60.100000  30.410000 ;
      RECT 15.485000  30.410000 60.170000  30.480000 ;
      RECT 15.485000  30.410000 60.170000  30.480000 ;
      RECT 15.485000  30.480000 60.240000  30.550000 ;
      RECT 15.485000  30.480000 60.240000  30.550000 ;
      RECT 15.485000  30.550000 60.310000  30.620000 ;
      RECT 15.485000  30.550000 60.310000  30.620000 ;
      RECT 15.485000  30.620000 60.380000  30.690000 ;
      RECT 15.485000  30.620000 60.380000  30.690000 ;
      RECT 15.485000  30.690000 60.450000  30.760000 ;
      RECT 15.485000  30.690000 60.450000  30.760000 ;
      RECT 15.485000  30.760000 60.520000  30.830000 ;
      RECT 15.485000  30.760000 60.520000  30.830000 ;
      RECT 15.485000  30.830000 60.590000  30.900000 ;
      RECT 15.485000  30.830000 60.590000  30.900000 ;
      RECT 15.485000  30.900000 60.660000  30.970000 ;
      RECT 15.485000  30.900000 60.660000  30.970000 ;
      RECT 15.485000  30.970000 60.730000  31.040000 ;
      RECT 15.485000  30.970000 60.730000  31.040000 ;
      RECT 15.485000  31.015000 60.970000  35.550000 ;
      RECT 15.485000  31.040000 60.800000  31.070000 ;
      RECT 15.485000  31.040000 60.800000  31.070000 ;
      RECT 15.485000  31.070000 60.830000  35.550000 ;
      RECT 15.485000  35.550000 60.970000  35.975000 ;
      RECT 15.485000  55.115000 17.415000  55.185000 ;
      RECT 15.495000  44.335000 60.130000  44.405000 ;
      RECT 15.495000  44.335000 60.130000  44.405000 ;
      RECT 15.505000  29.410000 59.170000  29.430000 ;
      RECT 15.505000  29.410000 59.170000  29.430000 ;
      RECT 15.505000  92.035000 58.520000  92.105000 ;
      RECT 15.505000  92.035000 58.520000  92.105000 ;
      RECT 15.510000 115.070000 58.395000 115.140000 ;
      RECT 15.510000 115.070000 58.395000 115.140000 ;
      RECT 15.520000  78.175000 24.540000  78.245000 ;
      RECT 15.520000  78.175000 24.540000  78.245000 ;
      RECT 15.520000 101.175000 24.540000 101.245000 ;
      RECT 15.520000 101.175000 24.540000 101.245000 ;
      RECT 15.520000 124.080000 24.540000 124.150000 ;
      RECT 15.520000 124.080000 24.540000 124.150000 ;
      RECT 15.520000 170.155000 16.525000 170.225000 ;
      RECT 15.525000 161.070000 58.445000 161.140000 ;
      RECT 15.525000 161.070000 58.445000 161.140000 ;
      RECT 15.540000  69.000000 58.495000  69.070000 ;
      RECT 15.540000  69.000000 58.495000  69.070000 ;
      RECT 15.545000 138.140000 58.360000 138.210000 ;
      RECT 15.545000 138.140000 58.360000 138.210000 ;
      RECT 15.545000 147.175000 16.875000 147.245000 ;
      RECT 15.545000 184.025000 59.500000 184.095000 ;
      RECT 15.555000  35.550000 60.830000  35.620000 ;
      RECT 15.555000  35.550000 60.830000  35.620000 ;
      RECT 15.555000  55.185000 17.485000  55.255000 ;
      RECT 15.565000  44.265000 60.200000  44.335000 ;
      RECT 15.565000  44.265000 60.200000  44.335000 ;
      RECT 15.575000  29.340000 59.100000  29.410000 ;
      RECT 15.575000  29.340000 59.100000  29.410000 ;
      RECT 15.575000  91.965000 58.590000  92.035000 ;
      RECT 15.575000  91.965000 58.590000  92.035000 ;
      RECT 15.580000 115.000000 58.465000 115.070000 ;
      RECT 15.580000 115.000000 58.465000 115.070000 ;
      RECT 15.590000  78.245000 24.540000  78.315000 ;
      RECT 15.590000  78.245000 24.540000  78.315000 ;
      RECT 15.590000 101.245000 24.540000 101.315000 ;
      RECT 15.590000 101.245000 24.540000 101.315000 ;
      RECT 15.590000 124.150000 24.540000 124.220000 ;
      RECT 15.590000 124.150000 24.540000 124.220000 ;
      RECT 15.590000 170.225000 16.525000 170.295000 ;
      RECT 15.595000 161.000000 58.515000 161.070000 ;
      RECT 15.595000 161.000000 58.515000 161.070000 ;
      RECT 15.610000  68.930000 58.565000  69.000000 ;
      RECT 15.610000  68.930000 58.565000  69.000000 ;
      RECT 15.615000 138.070000 58.430000 138.140000 ;
      RECT 15.615000 138.070000 58.430000 138.140000 ;
      RECT 15.615000 147.245000 16.945000 147.315000 ;
      RECT 15.615000 183.955000 59.570000 184.025000 ;
      RECT 15.625000  35.620000 60.830000  35.690000 ;
      RECT 15.625000  35.620000 60.830000  35.690000 ;
      RECT 15.625000  55.255000 17.555000  55.325000 ;
      RECT 15.635000  44.195000 60.270000  44.265000 ;
      RECT 15.635000  44.195000 60.270000  44.265000 ;
      RECT 15.645000  29.270000 59.030000  29.340000 ;
      RECT 15.645000  29.270000 59.030000  29.340000 ;
      RECT 15.645000  91.895000 58.660000  91.965000 ;
      RECT 15.645000  91.895000 58.660000  91.965000 ;
      RECT 15.650000 114.930000 58.535000 115.000000 ;
      RECT 15.650000 114.930000 58.535000 115.000000 ;
      RECT 15.660000  78.315000 24.540000  78.385000 ;
      RECT 15.660000  78.315000 24.540000  78.385000 ;
      RECT 15.660000 101.315000 24.540000 101.385000 ;
      RECT 15.660000 101.315000 24.540000 101.385000 ;
      RECT 15.660000 124.220000 24.540000 124.290000 ;
      RECT 15.660000 124.220000 24.540000 124.290000 ;
      RECT 15.660000 170.295000 16.525000 170.365000 ;
      RECT 15.665000 160.930000 58.585000 161.000000 ;
      RECT 15.665000 160.930000 58.585000 161.000000 ;
      RECT 15.680000  68.860000 58.635000  68.930000 ;
      RECT 15.680000  68.860000 58.635000  68.930000 ;
      RECT 15.685000 138.000000 58.500000 138.070000 ;
      RECT 15.685000 138.000000 58.500000 138.070000 ;
      RECT 15.685000 147.315000 17.015000 147.385000 ;
      RECT 15.685000 183.885000 59.640000 183.955000 ;
      RECT 15.695000  35.690000 60.830000  35.760000 ;
      RECT 15.695000  35.690000 60.830000  35.760000 ;
      RECT 15.695000  55.325000 17.625000  55.395000 ;
      RECT 15.705000  44.125000 60.340000  44.195000 ;
      RECT 15.705000  44.125000 60.340000  44.195000 ;
      RECT 15.715000  29.200000 58.960000  29.270000 ;
      RECT 15.715000  29.200000 58.960000  29.270000 ;
      RECT 15.715000  91.825000 58.730000  91.895000 ;
      RECT 15.715000  91.825000 58.730000  91.895000 ;
      RECT 15.720000 114.860000 58.605000 114.930000 ;
      RECT 15.720000 114.860000 58.605000 114.930000 ;
      RECT 15.730000  78.385000 24.540000  78.455000 ;
      RECT 15.730000  78.385000 24.540000  78.455000 ;
      RECT 15.730000 101.385000 24.540000 101.455000 ;
      RECT 15.730000 101.385000 24.540000 101.455000 ;
      RECT 15.730000 124.290000 24.540000 124.360000 ;
      RECT 15.730000 124.290000 24.540000 124.360000 ;
      RECT 15.730000 170.365000 16.525000 170.435000 ;
      RECT 15.735000 160.860000 58.655000 160.930000 ;
      RECT 15.735000 160.860000 58.655000 160.930000 ;
      RECT 15.750000  68.790000 58.705000  68.860000 ;
      RECT 15.750000  68.790000 58.705000  68.860000 ;
      RECT 15.755000 137.930000 58.570000 138.000000 ;
      RECT 15.755000 137.930000 58.570000 138.000000 ;
      RECT 15.755000 147.385000 17.085000 147.455000 ;
      RECT 15.755000 183.815000 59.710000 183.885000 ;
      RECT 15.765000  35.760000 60.830000  35.830000 ;
      RECT 15.765000  35.760000 60.830000  35.830000 ;
      RECT 15.765000  55.395000 17.695000  55.465000 ;
      RECT 15.770000  35.830000 60.830000  35.835000 ;
      RECT 15.770000  35.830000 60.830000  35.835000 ;
      RECT 15.775000  44.055000 60.410000  44.125000 ;
      RECT 15.775000  44.055000 60.410000  44.125000 ;
      RECT 15.785000  29.130000 58.890000  29.200000 ;
      RECT 15.785000  29.130000 58.890000  29.200000 ;
      RECT 15.785000  91.755000 58.800000  91.825000 ;
      RECT 15.785000  91.755000 58.800000  91.825000 ;
      RECT 15.790000 114.790000 58.675000 114.860000 ;
      RECT 15.790000 114.790000 58.675000 114.860000 ;
      RECT 15.800000  78.455000 24.540000  78.525000 ;
      RECT 15.800000  78.455000 24.540000  78.525000 ;
      RECT 15.800000 101.455000 24.540000 101.525000 ;
      RECT 15.800000 101.455000 24.540000 101.525000 ;
      RECT 15.800000 124.360000 24.540000 124.430000 ;
      RECT 15.800000 124.360000 24.540000 124.430000 ;
      RECT 15.800000 170.435000 16.525000 170.505000 ;
      RECT 15.805000 160.790000 58.725000 160.860000 ;
      RECT 15.805000 160.790000 58.725000 160.860000 ;
      RECT 15.820000  68.720000 58.775000  68.790000 ;
      RECT 15.820000  68.720000 58.775000  68.790000 ;
      RECT 15.825000 137.860000 58.640000 137.930000 ;
      RECT 15.825000 137.860000 58.640000 137.930000 ;
      RECT 15.825000 147.455000 17.155000 147.525000 ;
      RECT 15.825000 183.745000 59.780000 183.815000 ;
      RECT 15.835000  55.465000 17.765000  55.535000 ;
      RECT 15.840000  35.835000 54.390000  35.905000 ;
      RECT 15.840000  35.835000 54.390000  35.905000 ;
      RECT 15.845000  43.985000 60.480000  44.055000 ;
      RECT 15.845000  43.985000 60.480000  44.055000 ;
      RECT 15.855000  29.060000 58.820000  29.130000 ;
      RECT 15.855000  29.060000 58.820000  29.130000 ;
      RECT 15.855000  91.685000 58.870000  91.755000 ;
      RECT 15.855000  91.685000 58.870000  91.755000 ;
      RECT 15.860000 114.720000 58.745000 114.790000 ;
      RECT 15.860000 114.720000 58.745000 114.790000 ;
      RECT 15.870000  78.525000 24.540000  78.595000 ;
      RECT 15.870000  78.525000 24.540000  78.595000 ;
      RECT 15.870000 101.525000 24.540000 101.595000 ;
      RECT 15.870000 101.525000 24.540000 101.595000 ;
      RECT 15.870000 124.430000 24.540000 124.500000 ;
      RECT 15.870000 124.430000 24.540000 124.500000 ;
      RECT 15.870000 170.505000 16.525000 170.575000 ;
      RECT 15.875000 160.720000 58.795000 160.790000 ;
      RECT 15.875000 160.720000 58.795000 160.790000 ;
      RECT 15.890000  68.650000 58.845000  68.720000 ;
      RECT 15.890000  68.650000 58.845000  68.720000 ;
      RECT 15.895000 137.790000 58.710000 137.860000 ;
      RECT 15.895000 137.790000 58.710000 137.860000 ;
      RECT 15.895000 147.525000 17.225000 147.595000 ;
      RECT 15.895000 183.675000 59.850000 183.745000 ;
      RECT 15.905000  55.535000 17.835000  55.605000 ;
      RECT 15.910000  35.905000 54.390000  35.975000 ;
      RECT 15.910000  35.905000 54.390000  35.975000 ;
      RECT 15.910000  35.975000 54.530000  38.195000 ;
      RECT 15.915000  43.915000 60.550000  43.985000 ;
      RECT 15.915000  43.915000 60.550000  43.985000 ;
      RECT 15.925000  28.990000 58.750000  29.060000 ;
      RECT 15.925000  28.990000 58.750000  29.060000 ;
      RECT 15.925000  91.615000 58.940000  91.685000 ;
      RECT 15.925000  91.615000 58.940000  91.685000 ;
      RECT 15.930000 114.650000 58.815000 114.720000 ;
      RECT 15.930000 114.650000 58.815000 114.720000 ;
      RECT 15.940000  78.595000 24.540000  78.665000 ;
      RECT 15.940000  78.595000 24.540000  78.665000 ;
      RECT 15.940000 101.595000 24.540000 101.665000 ;
      RECT 15.940000 101.595000 24.540000 101.665000 ;
      RECT 15.940000 124.500000 24.540000 124.570000 ;
      RECT 15.940000 124.500000 24.540000 124.570000 ;
      RECT 15.940000 170.575000 16.525000 170.645000 ;
      RECT 15.945000 160.650000 58.865000 160.720000 ;
      RECT 15.945000 160.650000 58.865000 160.720000 ;
      RECT 15.960000  68.580000 58.915000  68.650000 ;
      RECT 15.960000  68.580000 58.915000  68.650000 ;
      RECT 15.965000 137.720000 58.780000 137.790000 ;
      RECT 15.965000 137.720000 58.780000 137.790000 ;
      RECT 15.965000 147.595000 17.295000 147.665000 ;
      RECT 15.965000 183.605000 59.920000 183.675000 ;
      RECT 15.975000  55.605000 17.905000  55.675000 ;
      RECT 15.980000  35.975000 54.390000  36.045000 ;
      RECT 15.980000  35.975000 54.390000  36.045000 ;
      RECT 15.985000  43.845000 60.620000  43.915000 ;
      RECT 15.985000  43.845000 60.620000  43.915000 ;
      RECT 15.995000  28.920000 58.680000  28.990000 ;
      RECT 15.995000  28.920000 58.680000  28.990000 ;
      RECT 15.995000  91.545000 59.010000  91.615000 ;
      RECT 15.995000  91.545000 59.010000  91.615000 ;
      RECT 16.000000 114.580000 58.885000 114.650000 ;
      RECT 16.000000 114.580000 58.885000 114.650000 ;
      RECT 16.010000  78.665000 24.540000  78.735000 ;
      RECT 16.010000  78.665000 24.540000  78.735000 ;
      RECT 16.010000 101.665000 24.540000 101.735000 ;
      RECT 16.010000 101.665000 24.540000 101.735000 ;
      RECT 16.010000 124.570000 24.540000 124.640000 ;
      RECT 16.010000 124.570000 24.540000 124.640000 ;
      RECT 16.010000 170.645000 16.525000 170.715000 ;
      RECT 16.015000 160.580000 58.935000 160.650000 ;
      RECT 16.015000 160.580000 58.935000 160.650000 ;
      RECT 16.030000  68.510000 58.985000  68.580000 ;
      RECT 16.030000  68.510000 58.985000  68.580000 ;
      RECT 16.035000 137.650000 58.850000 137.720000 ;
      RECT 16.035000 137.650000 58.850000 137.720000 ;
      RECT 16.035000 147.665000 17.365000 147.735000 ;
      RECT 16.035000 183.535000 59.990000 183.605000 ;
      RECT 16.045000  55.675000 17.975000  55.745000 ;
      RECT 16.050000  36.045000 54.390000  36.115000 ;
      RECT 16.050000  36.045000 54.390000  36.115000 ;
      RECT 16.055000  43.775000 60.690000  43.845000 ;
      RECT 16.055000  43.775000 60.690000  43.845000 ;
      RECT 16.065000  28.850000 58.610000  28.920000 ;
      RECT 16.065000  28.850000 58.610000  28.920000 ;
      RECT 16.065000  91.475000 59.080000  91.545000 ;
      RECT 16.065000  91.475000 59.080000  91.545000 ;
      RECT 16.070000  43.760000 59.300000  45.430000 ;
      RECT 16.070000 114.510000 58.955000 114.580000 ;
      RECT 16.070000 114.510000 58.955000 114.580000 ;
      RECT 16.080000  78.735000 24.540000  78.805000 ;
      RECT 16.080000  78.735000 24.540000  78.805000 ;
      RECT 16.080000 101.735000 24.540000 101.805000 ;
      RECT 16.080000 101.735000 24.540000 101.805000 ;
      RECT 16.080000 124.640000 24.540000 124.710000 ;
      RECT 16.080000 124.640000 24.540000 124.710000 ;
      RECT 16.080000 170.715000 16.525000 170.785000 ;
      RECT 16.085000 160.510000 59.005000 160.580000 ;
      RECT 16.085000 160.510000 59.005000 160.580000 ;
      RECT 16.100000  68.440000 59.055000  68.510000 ;
      RECT 16.100000  68.440000 59.055000  68.510000 ;
      RECT 16.105000 137.580000 58.920000 137.650000 ;
      RECT 16.105000 137.580000 58.920000 137.650000 ;
      RECT 16.105000 147.735000 17.435000 147.805000 ;
      RECT 16.105000 183.465000 60.060000 183.535000 ;
      RECT 16.115000  55.745000 18.045000  55.815000 ;
      RECT 16.120000  36.115000 54.390000  36.185000 ;
      RECT 16.120000  36.115000 54.390000  36.185000 ;
      RECT 16.125000  43.705000 60.760000  43.775000 ;
      RECT 16.125000  43.705000 60.760000  43.775000 ;
      RECT 16.135000  28.780000 58.540000  28.850000 ;
      RECT 16.135000  28.780000 58.540000  28.850000 ;
      RECT 16.135000  91.405000 59.150000  91.475000 ;
      RECT 16.135000  91.405000 59.150000  91.475000 ;
      RECT 16.140000 114.440000 59.025000 114.510000 ;
      RECT 16.140000 114.440000 59.025000 114.510000 ;
      RECT 16.150000  78.805000 24.540000  78.875000 ;
      RECT 16.150000  78.805000 24.540000  78.875000 ;
      RECT 16.150000 101.805000 24.540000 101.875000 ;
      RECT 16.150000 101.805000 24.540000 101.875000 ;
      RECT 16.150000 124.710000 24.540000 124.780000 ;
      RECT 16.150000 124.710000 24.540000 124.780000 ;
      RECT 16.150000 170.785000 16.525000 170.855000 ;
      RECT 16.155000 160.440000 59.075000 160.510000 ;
      RECT 16.155000 160.440000 59.075000 160.510000 ;
      RECT 16.170000  68.370000 59.125000  68.440000 ;
      RECT 16.170000  68.370000 59.125000  68.440000 ;
      RECT 16.175000 137.510000 58.990000 137.580000 ;
      RECT 16.175000 137.510000 58.990000 137.580000 ;
      RECT 16.175000 147.805000 17.505000 147.875000 ;
      RECT 16.175000 183.395000 60.130000 183.465000 ;
      RECT 16.185000  55.815000 18.115000  55.885000 ;
      RECT 16.190000  36.185000 54.390000  36.255000 ;
      RECT 16.190000  36.185000 54.390000  36.255000 ;
      RECT 16.190000  43.640000 60.830000  43.705000 ;
      RECT 16.190000  43.640000 60.830000  43.705000 ;
      RECT 16.205000  28.710000 58.470000  28.780000 ;
      RECT 16.205000  28.710000 58.470000  28.780000 ;
      RECT 16.205000  91.335000 59.220000  91.405000 ;
      RECT 16.205000  91.335000 59.220000  91.405000 ;
      RECT 16.210000 114.370000 59.095000 114.440000 ;
      RECT 16.210000 114.370000 59.095000 114.440000 ;
      RECT 16.220000  78.875000 24.540000  78.945000 ;
      RECT 16.220000  78.875000 24.540000  78.945000 ;
      RECT 16.220000 101.875000 24.540000 101.945000 ;
      RECT 16.220000 101.875000 24.540000 101.945000 ;
      RECT 16.220000 124.780000 24.540000 124.850000 ;
      RECT 16.220000 124.780000 24.540000 124.850000 ;
      RECT 16.220000 170.855000 16.525000 170.925000 ;
      RECT 16.225000 160.370000 59.145000 160.440000 ;
      RECT 16.225000 160.370000 59.145000 160.440000 ;
      RECT 16.240000  68.300000 59.195000  68.370000 ;
      RECT 16.240000  68.300000 59.195000  68.370000 ;
      RECT 16.245000 137.440000 59.060000 137.510000 ;
      RECT 16.245000 137.440000 59.060000 137.510000 ;
      RECT 16.245000 147.875000 17.575000 147.945000 ;
      RECT 16.245000 183.325000 60.200000 183.395000 ;
      RECT 16.255000  55.885000 18.185000  55.955000 ;
      RECT 16.260000  36.255000 54.390000  36.325000 ;
      RECT 16.260000  36.255000 54.390000  36.325000 ;
      RECT 16.260000  43.570000 60.830000  43.640000 ;
      RECT 16.260000  43.570000 60.830000  43.640000 ;
      RECT 16.275000  28.640000 58.400000  28.710000 ;
      RECT 16.275000  28.640000 58.400000  28.710000 ;
      RECT 16.275000  91.265000 59.290000  91.335000 ;
      RECT 16.275000  91.265000 59.290000  91.335000 ;
      RECT 16.280000 114.300000 59.165000 114.370000 ;
      RECT 16.280000 114.300000 59.165000 114.370000 ;
      RECT 16.290000  78.945000 24.540000  79.015000 ;
      RECT 16.290000  78.945000 24.540000  79.015000 ;
      RECT 16.290000 101.945000 24.540000 102.015000 ;
      RECT 16.290000 101.945000 24.540000 102.015000 ;
      RECT 16.290000 124.850000 24.540000 124.920000 ;
      RECT 16.290000 124.850000 24.540000 124.920000 ;
      RECT 16.290000 170.925000 16.525000 170.995000 ;
      RECT 16.295000 160.300000 59.215000 160.370000 ;
      RECT 16.295000 160.300000 59.215000 160.370000 ;
      RECT 16.310000  68.230000 59.265000  68.300000 ;
      RECT 16.310000  68.230000 59.265000  68.300000 ;
      RECT 16.315000 137.370000 59.130000 137.440000 ;
      RECT 16.315000 137.370000 59.130000 137.440000 ;
      RECT 16.315000 147.945000 17.645000 148.015000 ;
      RECT 16.315000 183.255000 60.270000 183.325000 ;
      RECT 16.325000  55.955000 18.255000  56.025000 ;
      RECT 16.330000  36.325000 54.390000  36.395000 ;
      RECT 16.330000  36.325000 54.390000  36.395000 ;
      RECT 16.330000  43.500000 60.830000  43.570000 ;
      RECT 16.330000  43.500000 60.830000  43.570000 ;
      RECT 16.345000  28.570000 58.330000  28.640000 ;
      RECT 16.345000  28.570000 58.330000  28.640000 ;
      RECT 16.345000  91.195000 59.360000  91.265000 ;
      RECT 16.345000  91.195000 59.360000  91.265000 ;
      RECT 16.350000 114.230000 59.235000 114.300000 ;
      RECT 16.350000 114.230000 59.235000 114.300000 ;
      RECT 16.360000  79.015000 24.540000  79.085000 ;
      RECT 16.360000  79.015000 24.540000  79.085000 ;
      RECT 16.360000 102.015000 24.540000 102.085000 ;
      RECT 16.360000 102.015000 24.540000 102.085000 ;
      RECT 16.360000 124.920000 24.540000 124.990000 ;
      RECT 16.360000 124.920000 24.540000 124.990000 ;
      RECT 16.360000 170.995000 16.525000 171.065000 ;
      RECT 16.365000 160.230000 59.285000 160.300000 ;
      RECT 16.365000 160.230000 59.285000 160.300000 ;
      RECT 16.380000  68.160000 59.335000  68.230000 ;
      RECT 16.380000  68.160000 59.335000  68.230000 ;
      RECT 16.385000 137.300000 59.200000 137.370000 ;
      RECT 16.385000 137.300000 59.200000 137.370000 ;
      RECT 16.385000 148.015000 17.715000 148.085000 ;
      RECT 16.385000 183.185000 60.340000 183.255000 ;
      RECT 16.395000  56.025000 18.325000  56.095000 ;
      RECT 16.400000  36.395000 54.390000  36.465000 ;
      RECT 16.400000  36.395000 54.390000  36.465000 ;
      RECT 16.400000  43.430000 60.830000  43.500000 ;
      RECT 16.400000  43.430000 60.830000  43.500000 ;
      RECT 16.415000  28.500000 58.260000  28.570000 ;
      RECT 16.415000  28.500000 58.260000  28.570000 ;
      RECT 16.415000  91.125000 59.430000  91.195000 ;
      RECT 16.415000  91.125000 59.430000  91.195000 ;
      RECT 16.420000 114.160000 59.305000 114.230000 ;
      RECT 16.420000 114.160000 59.305000 114.230000 ;
      RECT 16.430000  79.085000 24.540000  79.155000 ;
      RECT 16.430000  79.085000 24.540000  79.155000 ;
      RECT 16.430000 102.085000 24.540000 102.155000 ;
      RECT 16.430000 102.085000 24.540000 102.155000 ;
      RECT 16.430000 124.990000 24.540000 125.060000 ;
      RECT 16.430000 124.990000 24.540000 125.060000 ;
      RECT 16.430000 171.065000 16.525000 171.135000 ;
      RECT 16.435000 160.160000 59.355000 160.230000 ;
      RECT 16.435000 160.160000 59.355000 160.230000 ;
      RECT 16.450000  68.090000 59.405000  68.160000 ;
      RECT 16.450000  68.090000 59.405000  68.160000 ;
      RECT 16.455000 137.230000 59.270000 137.300000 ;
      RECT 16.455000 137.230000 59.270000 137.300000 ;
      RECT 16.455000 148.085000 17.785000 148.155000 ;
      RECT 16.455000 183.115000 60.410000 183.185000 ;
      RECT 16.465000  56.095000 18.395000  56.165000 ;
      RECT 16.470000  36.465000 54.390000  36.535000 ;
      RECT 16.470000  36.465000 54.390000  36.535000 ;
      RECT 16.470000  43.360000 60.830000  43.430000 ;
      RECT 16.470000  43.360000 60.830000  43.430000 ;
      RECT 16.485000  28.430000 58.190000  28.500000 ;
      RECT 16.485000  28.430000 58.190000  28.500000 ;
      RECT 16.485000  91.055000 59.500000  91.125000 ;
      RECT 16.485000  91.055000 59.500000  91.125000 ;
      RECT 16.490000 114.090000 59.375000 114.160000 ;
      RECT 16.490000 114.090000 59.375000 114.160000 ;
      RECT 16.500000  79.155000 24.540000  79.225000 ;
      RECT 16.500000  79.155000 24.540000  79.225000 ;
      RECT 16.500000 102.155000 24.540000 102.225000 ;
      RECT 16.500000 102.155000 24.540000 102.225000 ;
      RECT 16.500000 125.060000 24.540000 125.130000 ;
      RECT 16.500000 125.060000 24.540000 125.130000 ;
      RECT 16.500000 171.135000 16.525000 171.205000 ;
      RECT 16.505000 160.090000 59.425000 160.160000 ;
      RECT 16.505000 160.090000 59.425000 160.160000 ;
      RECT 16.520000  68.020000 59.475000  68.090000 ;
      RECT 16.520000  68.020000 59.475000  68.090000 ;
      RECT 16.525000 137.160000 59.340000 137.230000 ;
      RECT 16.525000 137.160000 59.340000 137.230000 ;
      RECT 16.525000 148.155000 17.855000 148.225000 ;
      RECT 16.525000 183.045000 60.480000 183.115000 ;
      RECT 16.535000  56.165000 18.465000  56.235000 ;
      RECT 16.540000  36.535000 54.390000  36.605000 ;
      RECT 16.540000  36.535000 54.390000  36.605000 ;
      RECT 16.540000  43.290000 60.830000  43.360000 ;
      RECT 16.540000  43.290000 60.830000  43.360000 ;
      RECT 16.555000  28.360000 58.120000  28.430000 ;
      RECT 16.555000  28.360000 58.120000  28.430000 ;
      RECT 16.555000  90.985000 59.570000  91.055000 ;
      RECT 16.555000  90.985000 59.570000  91.055000 ;
      RECT 16.560000 114.020000 59.445000 114.090000 ;
      RECT 16.560000 114.020000 59.445000 114.090000 ;
      RECT 16.570000  79.225000 24.540000  79.295000 ;
      RECT 16.570000  79.225000 24.540000  79.295000 ;
      RECT 16.570000  79.295000 58.700000  80.500000 ;
      RECT 16.570000 102.225000 24.540000 102.295000 ;
      RECT 16.570000 102.225000 24.540000 102.295000 ;
      RECT 16.570000 102.295000 58.700000 103.500000 ;
      RECT 16.570000 125.130000 24.540000 125.200000 ;
      RECT 16.570000 125.130000 24.540000 125.200000 ;
      RECT 16.575000 160.020000 59.495000 160.090000 ;
      RECT 16.575000 160.020000 59.495000 160.090000 ;
      RECT 16.590000  67.950000 59.545000  68.020000 ;
      RECT 16.590000  67.950000 59.545000  68.020000 ;
      RECT 16.590000 171.295000 58.710000 172.500000 ;
      RECT 16.595000  56.295000 58.670000  57.500000 ;
      RECT 16.595000 137.090000 59.410000 137.160000 ;
      RECT 16.595000 137.090000 59.410000 137.160000 ;
      RECT 16.595000 148.225000 17.925000 148.295000 ;
      RECT 16.595000 148.295000 58.630000 149.500000 ;
      RECT 16.595000 182.975000 60.550000 183.045000 ;
      RECT 16.605000  56.235000 18.535000  56.305000 ;
      RECT 16.610000  36.605000 54.390000  36.675000 ;
      RECT 16.610000  36.605000 54.390000  36.675000 ;
      RECT 16.610000  43.220000 60.830000  43.290000 ;
      RECT 16.610000  43.220000 60.830000  43.290000 ;
      RECT 16.625000  28.290000 58.050000  28.360000 ;
      RECT 16.625000  28.290000 58.050000  28.360000 ;
      RECT 16.625000  90.915000 59.640000  90.985000 ;
      RECT 16.625000  90.915000 59.640000  90.985000 ;
      RECT 16.630000 113.950000 59.515000 114.020000 ;
      RECT 16.630000 113.950000 59.515000 114.020000 ;
      RECT 16.640000  79.295000 24.540000  79.365000 ;
      RECT 16.640000  79.295000 24.540000  79.365000 ;
      RECT 16.640000 102.295000 24.540000 102.365000 ;
      RECT 16.640000 102.295000 24.540000 102.365000 ;
      RECT 16.640000 125.200000 24.540000 125.270000 ;
      RECT 16.640000 125.200000 24.540000 125.270000 ;
      RECT 16.645000 159.950000 59.565000 160.020000 ;
      RECT 16.645000 159.950000 59.565000 160.020000 ;
      RECT 16.660000  67.880000 59.615000  67.950000 ;
      RECT 16.660000  67.880000 59.615000  67.950000 ;
      RECT 16.665000 125.295000 58.700000 126.500000 ;
      RECT 16.665000 137.020000 59.480000 137.090000 ;
      RECT 16.665000 137.020000 59.480000 137.090000 ;
      RECT 16.665000 148.295000 17.995000 148.365000 ;
      RECT 16.665000 182.905000 60.620000 182.975000 ;
      RECT 16.675000  56.305000 18.605000  56.375000 ;
      RECT 16.680000  36.675000 54.390000  36.745000 ;
      RECT 16.680000  36.675000 54.390000  36.745000 ;
      RECT 16.680000  43.150000 60.830000  43.220000 ;
      RECT 16.680000  43.150000 60.830000  43.220000 ;
      RECT 16.695000  28.220000 57.980000  28.290000 ;
      RECT 16.695000  28.220000 57.980000  28.290000 ;
      RECT 16.695000  90.845000 59.710000  90.915000 ;
      RECT 16.695000  90.845000 59.710000  90.915000 ;
      RECT 16.700000 113.880000 59.585000 113.950000 ;
      RECT 16.700000 113.880000 59.585000 113.950000 ;
      RECT 16.710000  79.365000 24.540000  79.435000 ;
      RECT 16.710000  79.365000 24.540000  79.435000 ;
      RECT 16.710000 102.365000 24.540000 102.435000 ;
      RECT 16.710000 102.365000 24.540000 102.435000 ;
      RECT 16.710000 125.270000 24.540000 125.340000 ;
      RECT 16.710000 125.270000 24.540000 125.340000 ;
      RECT 16.715000 159.880000 59.635000 159.950000 ;
      RECT 16.715000 159.880000 59.635000 159.950000 ;
      RECT 16.730000  67.810000 59.685000  67.880000 ;
      RECT 16.730000  67.810000 59.685000  67.880000 ;
      RECT 16.735000  56.375000 18.675000  56.435000 ;
      RECT 16.735000 136.950000 59.550000 137.020000 ;
      RECT 16.735000 136.950000 59.550000 137.020000 ;
      RECT 16.735000 148.365000 18.065000 148.435000 ;
      RECT 16.735000 182.835000 60.690000 182.905000 ;
      RECT 16.750000  36.745000 54.390000  36.815000 ;
      RECT 16.750000  36.745000 54.390000  36.815000 ;
      RECT 16.750000  43.080000 60.830000  43.150000 ;
      RECT 16.750000  43.080000 60.830000  43.150000 ;
      RECT 16.750000 182.820000 58.635000 185.155000 ;
      RECT 16.765000  28.150000 57.910000  28.220000 ;
      RECT 16.765000  28.150000 57.910000  28.220000 ;
      RECT 16.765000  90.775000 59.780000  90.845000 ;
      RECT 16.765000  90.775000 59.780000  90.845000 ;
      RECT 16.770000 113.810000 59.655000 113.880000 ;
      RECT 16.770000 113.810000 59.655000 113.880000 ;
      RECT 16.780000  79.435000 24.540000  79.505000 ;
      RECT 16.780000  79.435000 24.540000  79.505000 ;
      RECT 16.780000  79.435000 57.440000  79.505000 ;
      RECT 16.780000 102.435000 24.540000 102.505000 ;
      RECT 16.780000 102.435000 24.540000 102.505000 ;
      RECT 16.780000 102.435000 57.440000 102.505000 ;
      RECT 16.780000 125.340000 24.540000 125.410000 ;
      RECT 16.780000 125.340000 24.540000 125.410000 ;
      RECT 16.785000 159.810000 59.705000 159.880000 ;
      RECT 16.785000 159.810000 59.705000 159.880000 ;
      RECT 16.800000  67.740000 59.755000  67.810000 ;
      RECT 16.800000  67.740000 59.755000  67.810000 ;
      RECT 16.800000 171.435000 57.450000 171.505000 ;
      RECT 16.805000  56.435000 57.410000  56.505000 ;
      RECT 16.805000 125.410000 24.540000 125.435000 ;
      RECT 16.805000 125.410000 24.540000 125.435000 ;
      RECT 16.805000 136.880000 59.620000 136.950000 ;
      RECT 16.805000 136.880000 59.620000 136.950000 ;
      RECT 16.805000 148.435000 57.370000 148.505000 ;
      RECT 16.805000 182.765000 60.760000 182.835000 ;
      RECT 16.820000  36.815000 54.390000  36.885000 ;
      RECT 16.820000  36.815000 54.390000  36.885000 ;
      RECT 16.820000  43.010000 60.830000  43.080000 ;
      RECT 16.820000  43.010000 60.830000  43.080000 ;
      RECT 16.830000 182.740000 60.830000 182.765000 ;
      RECT 16.835000  28.080000 57.840000  28.150000 ;
      RECT 16.835000  28.080000 57.840000  28.150000 ;
      RECT 16.835000  90.705000 59.850000  90.775000 ;
      RECT 16.835000  90.705000 59.850000  90.775000 ;
      RECT 16.840000 113.740000 59.725000 113.810000 ;
      RECT 16.840000 113.740000 59.725000 113.810000 ;
      RECT 16.850000  79.505000 24.540000  79.575000 ;
      RECT 16.850000  79.505000 24.540000  79.575000 ;
      RECT 16.850000  79.505000 57.510000  79.575000 ;
      RECT 16.850000 102.505000 24.540000 102.575000 ;
      RECT 16.850000 102.505000 24.540000 102.575000 ;
      RECT 16.850000 102.505000 57.510000 102.575000 ;
      RECT 16.855000 159.740000 59.775000 159.810000 ;
      RECT 16.855000 159.740000 59.775000 159.810000 ;
      RECT 16.870000  67.670000 59.825000  67.740000 ;
      RECT 16.870000  67.670000 59.825000  67.740000 ;
      RECT 16.870000 171.505000 57.520000 171.575000 ;
      RECT 16.875000  56.505000 57.480000  56.575000 ;
      RECT 16.875000 125.435000 24.540000 125.505000 ;
      RECT 16.875000 125.435000 24.540000 125.505000 ;
      RECT 16.875000 125.435000 57.440000 125.505000 ;
      RECT 16.875000 136.810000 59.690000 136.880000 ;
      RECT 16.875000 136.810000 59.690000 136.880000 ;
      RECT 16.875000 148.505000 57.440000 148.575000 ;
      RECT 16.890000  36.885000 54.390000  36.955000 ;
      RECT 16.890000  36.885000 54.390000  36.955000 ;
      RECT 16.890000  42.940000 60.830000  43.010000 ;
      RECT 16.890000  42.940000 60.830000  43.010000 ;
      RECT 16.900000 182.670000 60.830000 182.740000 ;
      RECT 16.905000  28.010000 57.770000  28.080000 ;
      RECT 16.905000  28.010000 57.770000  28.080000 ;
      RECT 16.905000  90.635000 59.920000  90.705000 ;
      RECT 16.905000  90.635000 59.920000  90.705000 ;
      RECT 16.910000 113.670000 59.795000 113.740000 ;
      RECT 16.910000 113.670000 59.795000 113.740000 ;
      RECT 16.920000  79.575000 24.540000  79.645000 ;
      RECT 16.920000  79.575000 24.540000  79.645000 ;
      RECT 16.920000  79.575000 57.580000  79.645000 ;
      RECT 16.920000 102.575000 24.540000 102.645000 ;
      RECT 16.920000 102.575000 24.540000 102.645000 ;
      RECT 16.920000 102.575000 57.580000 102.645000 ;
      RECT 16.925000 159.670000 59.845000 159.740000 ;
      RECT 16.925000 159.670000 59.845000 159.740000 ;
      RECT 16.940000  67.600000 59.895000  67.670000 ;
      RECT 16.940000  67.600000 59.895000  67.670000 ;
      RECT 16.940000 171.575000 57.590000 171.645000 ;
      RECT 16.945000  56.575000 57.550000  56.645000 ;
      RECT 16.945000 125.505000 24.540000 125.575000 ;
      RECT 16.945000 125.505000 24.540000 125.575000 ;
      RECT 16.945000 125.505000 57.510000 125.575000 ;
      RECT 16.945000 136.740000 59.760000 136.810000 ;
      RECT 16.945000 136.740000 59.760000 136.810000 ;
      RECT 16.945000 148.575000 57.510000 148.645000 ;
      RECT 16.960000  36.955000 54.390000  37.025000 ;
      RECT 16.960000  36.955000 54.390000  37.025000 ;
      RECT 16.960000  42.870000 60.830000  42.940000 ;
      RECT 16.960000  42.870000 60.830000  42.940000 ;
      RECT 16.970000 182.600000 60.830000 182.670000 ;
      RECT 16.975000  27.940000 57.700000  28.010000 ;
      RECT 16.975000  27.940000 57.700000  28.010000 ;
      RECT 16.975000  90.565000 59.990000  90.635000 ;
      RECT 16.975000  90.565000 59.990000  90.635000 ;
      RECT 16.980000 113.600000 59.865000 113.670000 ;
      RECT 16.980000 113.600000 59.865000 113.670000 ;
      RECT 16.990000  79.645000 24.540000  79.715000 ;
      RECT 16.990000  79.645000 24.540000  79.715000 ;
      RECT 16.990000  79.645000 57.650000  79.715000 ;
      RECT 16.990000 102.645000 24.540000 102.715000 ;
      RECT 16.990000 102.645000 24.540000 102.715000 ;
      RECT 16.990000 102.645000 57.650000 102.715000 ;
      RECT 16.995000 159.600000 59.915000 159.670000 ;
      RECT 16.995000 159.600000 59.915000 159.670000 ;
      RECT 17.010000  67.530000 59.965000  67.600000 ;
      RECT 17.010000  67.530000 59.965000  67.600000 ;
      RECT 17.010000 171.645000 57.660000 171.715000 ;
      RECT 17.015000  56.645000 57.620000  56.715000 ;
      RECT 17.015000 125.575000 24.540000 125.645000 ;
      RECT 17.015000 125.575000 24.540000 125.645000 ;
      RECT 17.015000 125.575000 57.580000 125.645000 ;
      RECT 17.015000 136.670000 59.830000 136.740000 ;
      RECT 17.015000 136.670000 59.830000 136.740000 ;
      RECT 17.015000 148.645000 57.580000 148.715000 ;
      RECT 17.030000  37.025000 54.390000  37.095000 ;
      RECT 17.030000  37.025000 54.390000  37.095000 ;
      RECT 17.030000  42.800000 60.830000  42.870000 ;
      RECT 17.030000  42.800000 60.830000  42.870000 ;
      RECT 17.040000 182.530000 60.830000 182.600000 ;
      RECT 17.045000  27.870000 57.630000  27.940000 ;
      RECT 17.045000  27.870000 57.630000  27.940000 ;
      RECT 17.045000  90.495000 60.060000  90.565000 ;
      RECT 17.045000  90.495000 60.060000  90.565000 ;
      RECT 17.050000 113.530000 59.935000 113.600000 ;
      RECT 17.050000 113.530000 59.935000 113.600000 ;
      RECT 17.060000  79.715000 24.540000  79.785000 ;
      RECT 17.060000  79.715000 24.540000  79.785000 ;
      RECT 17.060000  79.715000 57.720000  79.785000 ;
      RECT 17.060000 102.715000 24.540000 102.785000 ;
      RECT 17.060000 102.715000 24.540000 102.785000 ;
      RECT 17.060000 102.715000 57.720000 102.785000 ;
      RECT 17.065000 159.530000 59.985000 159.600000 ;
      RECT 17.065000 159.530000 59.985000 159.600000 ;
      RECT 17.080000  67.460000 60.035000  67.530000 ;
      RECT 17.080000  67.460000 60.035000  67.530000 ;
      RECT 17.080000 171.715000 57.730000 171.785000 ;
      RECT 17.085000  56.715000 57.690000  56.785000 ;
      RECT 17.085000 125.645000 24.540000 125.715000 ;
      RECT 17.085000 125.645000 24.540000 125.715000 ;
      RECT 17.085000 125.645000 57.650000 125.715000 ;
      RECT 17.085000 136.600000 59.900000 136.670000 ;
      RECT 17.085000 136.600000 59.900000 136.670000 ;
      RECT 17.085000 148.715000 57.650000 148.785000 ;
      RECT 17.100000  37.095000 54.390000  37.165000 ;
      RECT 17.100000  37.095000 54.390000  37.165000 ;
      RECT 17.100000  42.730000 60.830000  42.800000 ;
      RECT 17.100000  42.730000 60.830000  42.800000 ;
      RECT 17.110000 182.460000 60.830000 182.530000 ;
      RECT 17.115000  27.800000 57.560000  27.870000 ;
      RECT 17.115000  27.800000 57.560000  27.870000 ;
      RECT 17.115000  90.425000 60.130000  90.495000 ;
      RECT 17.115000  90.425000 60.130000  90.495000 ;
      RECT 17.120000 113.460000 60.005000 113.530000 ;
      RECT 17.120000 113.460000 60.005000 113.530000 ;
      RECT 17.130000  79.785000 24.540000  79.855000 ;
      RECT 17.130000  79.785000 24.540000  79.855000 ;
      RECT 17.130000  79.785000 57.790000  79.855000 ;
      RECT 17.130000 102.785000 24.540000 102.855000 ;
      RECT 17.130000 102.785000 24.540000 102.855000 ;
      RECT 17.130000 102.785000 57.790000 102.855000 ;
      RECT 17.135000 159.460000 60.055000 159.530000 ;
      RECT 17.135000 159.460000 60.055000 159.530000 ;
      RECT 17.150000  67.390000 60.105000  67.460000 ;
      RECT 17.150000  67.390000 60.105000  67.460000 ;
      RECT 17.150000 171.785000 57.800000 171.855000 ;
      RECT 17.155000  56.785000 57.760000  56.855000 ;
      RECT 17.155000 125.715000 24.540000 125.785000 ;
      RECT 17.155000 125.715000 24.540000 125.785000 ;
      RECT 17.155000 125.715000 57.720000 125.785000 ;
      RECT 17.155000 136.530000 59.970000 136.600000 ;
      RECT 17.155000 136.530000 59.970000 136.600000 ;
      RECT 17.155000 148.785000 57.720000 148.855000 ;
      RECT 17.170000  37.165000 54.390000  37.235000 ;
      RECT 17.170000  37.165000 54.390000  37.235000 ;
      RECT 17.170000  42.660000 60.830000  42.730000 ;
      RECT 17.170000  42.660000 60.830000  42.730000 ;
      RECT 17.170000  42.660000 60.970000  43.760000 ;
      RECT 17.180000 182.390000 60.830000 182.460000 ;
      RECT 17.185000  27.730000 57.490000  27.800000 ;
      RECT 17.185000  27.730000 57.490000  27.800000 ;
      RECT 17.185000  90.355000 60.200000  90.425000 ;
      RECT 17.185000  90.355000 60.200000  90.425000 ;
      RECT 17.190000 113.390000 60.075000 113.460000 ;
      RECT 17.190000 113.390000 60.075000 113.460000 ;
      RECT 17.200000  79.855000 24.540000  79.925000 ;
      RECT 17.200000  79.855000 24.540000  79.925000 ;
      RECT 17.200000  79.855000 57.860000  79.925000 ;
      RECT 17.200000 102.855000 24.540000 102.925000 ;
      RECT 17.200000 102.855000 24.540000 102.925000 ;
      RECT 17.200000 102.855000 57.860000 102.925000 ;
      RECT 17.205000 159.390000 60.125000 159.460000 ;
      RECT 17.205000 159.390000 60.125000 159.460000 ;
      RECT 17.220000  67.320000 60.175000  67.390000 ;
      RECT 17.220000  67.320000 60.175000  67.390000 ;
      RECT 17.220000 171.855000 57.870000 171.925000 ;
      RECT 17.225000  56.855000 57.830000  56.925000 ;
      RECT 17.225000 125.785000 24.540000 125.855000 ;
      RECT 17.225000 125.785000 24.540000 125.855000 ;
      RECT 17.225000 125.785000 57.790000 125.855000 ;
      RECT 17.225000 136.460000 60.040000 136.530000 ;
      RECT 17.225000 136.460000 60.040000 136.530000 ;
      RECT 17.225000 148.855000 57.790000 148.925000 ;
      RECT 17.240000  37.235000 54.390000  37.305000 ;
      RECT 17.240000  37.235000 54.390000  37.305000 ;
      RECT 17.250000 182.320000 60.830000 182.390000 ;
      RECT 17.255000  27.660000 57.420000  27.730000 ;
      RECT 17.255000  27.660000 57.420000  27.730000 ;
      RECT 17.255000  90.285000 60.270000  90.355000 ;
      RECT 17.255000  90.285000 60.270000  90.355000 ;
      RECT 17.260000 113.320000 60.145000 113.390000 ;
      RECT 17.260000 113.320000 60.145000 113.390000 ;
      RECT 17.270000  79.925000 24.540000  79.995000 ;
      RECT 17.270000  79.925000 24.540000  79.995000 ;
      RECT 17.270000  79.925000 57.930000  79.995000 ;
      RECT 17.270000 102.925000 24.540000 102.995000 ;
      RECT 17.270000 102.925000 24.540000 102.995000 ;
      RECT 17.270000 102.925000 57.930000 102.995000 ;
      RECT 17.275000 159.320000 60.195000 159.390000 ;
      RECT 17.275000 159.320000 60.195000 159.390000 ;
      RECT 17.290000  67.250000 60.245000  67.320000 ;
      RECT 17.290000  67.250000 60.245000  67.320000 ;
      RECT 17.290000 171.925000 57.940000 171.995000 ;
      RECT 17.295000  56.925000 57.900000  56.995000 ;
      RECT 17.295000 125.855000 24.540000 125.925000 ;
      RECT 17.295000 125.855000 24.540000 125.925000 ;
      RECT 17.295000 125.855000 57.860000 125.925000 ;
      RECT 17.295000 136.390000 60.110000 136.460000 ;
      RECT 17.295000 136.390000 60.110000 136.460000 ;
      RECT 17.295000 148.925000 57.860000 148.995000 ;
      RECT 17.310000  37.305000 54.390000  37.375000 ;
      RECT 17.310000  37.305000 54.390000  37.375000 ;
      RECT 17.320000 182.250000 60.830000 182.320000 ;
      RECT 17.325000  27.590000 57.350000  27.660000 ;
      RECT 17.325000  27.590000 57.350000  27.660000 ;
      RECT 17.325000  90.215000 60.340000  90.285000 ;
      RECT 17.325000  90.215000 60.340000  90.285000 ;
      RECT 17.330000 113.250000 60.215000 113.320000 ;
      RECT 17.330000 113.250000 60.215000 113.320000 ;
      RECT 17.340000  79.995000 24.540000  80.065000 ;
      RECT 17.340000  79.995000 24.540000  80.065000 ;
      RECT 17.340000  79.995000 58.000000  80.065000 ;
      RECT 17.340000 102.995000 24.540000 103.065000 ;
      RECT 17.340000 102.995000 24.540000 103.065000 ;
      RECT 17.340000 102.995000 58.000000 103.065000 ;
      RECT 17.345000 159.250000 60.265000 159.320000 ;
      RECT 17.345000 159.250000 60.265000 159.320000 ;
      RECT 17.360000  67.180000 60.315000  67.250000 ;
      RECT 17.360000  67.180000 60.315000  67.250000 ;
      RECT 17.360000 171.995000 58.010000 172.065000 ;
      RECT 17.365000  56.995000 57.970000  57.065000 ;
      RECT 17.365000 125.925000 24.540000 125.995000 ;
      RECT 17.365000 125.925000 24.540000 125.995000 ;
      RECT 17.365000 125.925000 57.930000 125.995000 ;
      RECT 17.365000 136.320000 60.180000 136.390000 ;
      RECT 17.365000 136.320000 60.180000 136.390000 ;
      RECT 17.365000 148.995000 57.930000 149.065000 ;
      RECT 17.380000  37.375000 54.390000  37.445000 ;
      RECT 17.380000  37.375000 54.390000  37.445000 ;
      RECT 17.390000 182.180000 60.830000 182.250000 ;
      RECT 17.395000  27.520000 57.280000  27.590000 ;
      RECT 17.395000  27.520000 57.280000  27.590000 ;
      RECT 17.395000  90.145000 60.410000  90.215000 ;
      RECT 17.395000  90.145000 60.410000  90.215000 ;
      RECT 17.400000 113.180000 60.285000 113.250000 ;
      RECT 17.400000 113.180000 60.285000 113.250000 ;
      RECT 17.410000  80.065000 24.540000  80.135000 ;
      RECT 17.410000  80.065000 24.540000  80.135000 ;
      RECT 17.410000  80.065000 58.070000  80.135000 ;
      RECT 17.410000 103.065000 24.540000 103.135000 ;
      RECT 17.410000 103.065000 24.540000 103.135000 ;
      RECT 17.410000 103.065000 58.070000 103.135000 ;
      RECT 17.415000 159.180000 60.335000 159.250000 ;
      RECT 17.415000 159.180000 60.335000 159.250000 ;
      RECT 17.430000  67.110000 60.385000  67.180000 ;
      RECT 17.430000  67.110000 60.385000  67.180000 ;
      RECT 17.430000 172.065000 58.080000 172.135000 ;
      RECT 17.435000  57.065000 58.040000  57.135000 ;
      RECT 17.435000 125.995000 24.540000 126.065000 ;
      RECT 17.435000 125.995000 24.540000 126.065000 ;
      RECT 17.435000 125.995000 58.000000 126.065000 ;
      RECT 17.435000 136.250000 60.250000 136.320000 ;
      RECT 17.435000 136.250000 60.250000 136.320000 ;
      RECT 17.435000 149.065000 58.000000 149.135000 ;
      RECT 17.450000  37.445000 54.390000  37.515000 ;
      RECT 17.450000  37.445000 54.390000  37.515000 ;
      RECT 17.460000 182.110000 60.830000 182.180000 ;
      RECT 17.465000  27.450000 57.210000  27.520000 ;
      RECT 17.465000  27.450000 57.210000  27.520000 ;
      RECT 17.465000  90.075000 60.480000  90.145000 ;
      RECT 17.465000  90.075000 60.480000  90.145000 ;
      RECT 17.470000 113.110000 60.355000 113.180000 ;
      RECT 17.470000 113.110000 60.355000 113.180000 ;
      RECT 17.480000  80.135000 24.540000  80.205000 ;
      RECT 17.480000  80.135000 24.540000  80.205000 ;
      RECT 17.480000  80.135000 58.140000  80.205000 ;
      RECT 17.480000 103.135000 24.540000 103.205000 ;
      RECT 17.480000 103.135000 24.540000 103.205000 ;
      RECT 17.480000 103.135000 58.140000 103.205000 ;
      RECT 17.485000 159.110000 60.405000 159.180000 ;
      RECT 17.485000 159.110000 60.405000 159.180000 ;
      RECT 17.500000  67.040000 60.455000  67.110000 ;
      RECT 17.500000  67.040000 60.455000  67.110000 ;
      RECT 17.500000 172.135000 58.150000 172.205000 ;
      RECT 17.505000  57.135000 58.110000  57.205000 ;
      RECT 17.505000 126.065000 24.540000 126.135000 ;
      RECT 17.505000 126.065000 24.540000 126.135000 ;
      RECT 17.505000 126.065000 58.070000 126.135000 ;
      RECT 17.505000 136.180000 60.320000 136.250000 ;
      RECT 17.505000 136.180000 60.320000 136.250000 ;
      RECT 17.505000 149.135000 58.070000 149.205000 ;
      RECT 17.520000  37.515000 54.390000  37.585000 ;
      RECT 17.520000  37.515000 54.390000  37.585000 ;
      RECT 17.530000 182.040000 60.830000 182.110000 ;
      RECT 17.535000  27.380000 57.140000  27.450000 ;
      RECT 17.535000  27.380000 57.140000  27.450000 ;
      RECT 17.535000  90.005000 60.550000  90.075000 ;
      RECT 17.535000  90.005000 60.550000  90.075000 ;
      RECT 17.540000 113.040000 60.425000 113.110000 ;
      RECT 17.540000 113.040000 60.425000 113.110000 ;
      RECT 17.550000  80.205000 24.540000  80.275000 ;
      RECT 17.550000  80.205000 24.540000  80.275000 ;
      RECT 17.550000  80.205000 58.210000  80.275000 ;
      RECT 17.550000 103.205000 24.540000 103.275000 ;
      RECT 17.550000 103.205000 24.540000 103.275000 ;
      RECT 17.550000 103.205000 58.210000 103.275000 ;
      RECT 17.555000 159.040000 60.475000 159.110000 ;
      RECT 17.555000 159.040000 60.475000 159.110000 ;
      RECT 17.570000  66.970000 60.525000  67.040000 ;
      RECT 17.570000  66.970000 60.525000  67.040000 ;
      RECT 17.570000 172.205000 58.220000 172.275000 ;
      RECT 17.575000  57.205000 58.180000  57.275000 ;
      RECT 17.575000 126.135000 24.540000 126.205000 ;
      RECT 17.575000 126.135000 24.540000 126.205000 ;
      RECT 17.575000 126.135000 58.140000 126.205000 ;
      RECT 17.575000 136.110000 60.390000 136.180000 ;
      RECT 17.575000 136.110000 60.390000 136.180000 ;
      RECT 17.575000 149.205000 58.140000 149.275000 ;
      RECT 17.590000  37.585000 54.390000  37.655000 ;
      RECT 17.590000  37.585000 54.390000  37.655000 ;
      RECT 17.600000 181.970000 60.830000 182.040000 ;
      RECT 17.605000  27.310000 57.070000  27.380000 ;
      RECT 17.605000  27.310000 57.070000  27.380000 ;
      RECT 17.605000  89.935000 60.620000  90.005000 ;
      RECT 17.605000  89.935000 60.620000  90.005000 ;
      RECT 17.610000 112.970000 60.495000 113.040000 ;
      RECT 17.610000 112.970000 60.495000 113.040000 ;
      RECT 17.620000  80.275000 24.540000  80.345000 ;
      RECT 17.620000  80.275000 24.540000  80.345000 ;
      RECT 17.620000  80.275000 58.280000  80.345000 ;
      RECT 17.620000 103.275000 24.540000 103.345000 ;
      RECT 17.620000 103.275000 24.540000 103.345000 ;
      RECT 17.620000 103.275000 58.280000 103.345000 ;
      RECT 17.625000 158.970000 60.545000 159.040000 ;
      RECT 17.625000 158.970000 60.545000 159.040000 ;
      RECT 17.640000  66.900000 60.595000  66.970000 ;
      RECT 17.640000  66.900000 60.595000  66.970000 ;
      RECT 17.640000 172.275000 58.290000 172.345000 ;
      RECT 17.645000  57.275000 58.250000  57.345000 ;
      RECT 17.645000 126.205000 24.540000 126.275000 ;
      RECT 17.645000 126.205000 24.540000 126.275000 ;
      RECT 17.645000 126.205000 58.210000 126.275000 ;
      RECT 17.645000 136.040000 60.460000 136.110000 ;
      RECT 17.645000 136.040000 60.460000 136.110000 ;
      RECT 17.645000 149.275000 58.210000 149.345000 ;
      RECT 17.660000  37.655000 54.390000  37.725000 ;
      RECT 17.660000  37.655000 54.390000  37.725000 ;
      RECT 17.670000 181.900000 60.830000 181.970000 ;
      RECT 17.675000  27.240000 57.000000  27.310000 ;
      RECT 17.675000  27.240000 57.000000  27.310000 ;
      RECT 17.675000  89.865000 60.690000  89.935000 ;
      RECT 17.675000  89.865000 60.690000  89.935000 ;
      RECT 17.680000 112.900000 60.565000 112.970000 ;
      RECT 17.680000 112.900000 60.565000 112.970000 ;
      RECT 17.690000  80.345000 24.540000  80.415000 ;
      RECT 17.690000  80.345000 24.540000  80.415000 ;
      RECT 17.690000  80.345000 58.350000  80.415000 ;
      RECT 17.690000  89.850000 57.680000  93.140000 ;
      RECT 17.690000 103.345000 24.540000 103.415000 ;
      RECT 17.690000 103.345000 24.540000 103.415000 ;
      RECT 17.690000 103.345000 58.350000 103.415000 ;
      RECT 17.695000 158.900000 60.615000 158.970000 ;
      RECT 17.695000 158.900000 60.615000 158.970000 ;
      RECT 17.710000  66.830000 60.665000  66.900000 ;
      RECT 17.710000  66.830000 60.665000  66.900000 ;
      RECT 17.710000 172.345000 58.360000 172.415000 ;
      RECT 17.715000  57.345000 58.320000  57.415000 ;
      RECT 17.715000 126.275000 24.540000 126.345000 ;
      RECT 17.715000 126.275000 24.540000 126.345000 ;
      RECT 17.715000 126.275000 58.280000 126.345000 ;
      RECT 17.715000 135.970000 60.530000 136.040000 ;
      RECT 17.715000 135.970000 60.530000 136.040000 ;
      RECT 17.715000 149.345000 58.280000 149.415000 ;
      RECT 17.730000  37.725000 54.390000  37.795000 ;
      RECT 17.730000  37.725000 54.390000  37.795000 ;
      RECT 17.740000 181.830000 60.830000 181.900000 ;
      RECT 17.745000  27.170000 56.930000  27.240000 ;
      RECT 17.745000  27.170000 56.930000  27.240000 ;
      RECT 17.745000  89.795000 60.760000  89.865000 ;
      RECT 17.745000  89.795000 60.760000  89.865000 ;
      RECT 17.750000  66.790000 57.620000  70.140000 ;
      RECT 17.750000  89.790000 60.830000  89.795000 ;
      RECT 17.750000  89.790000 60.830000  89.795000 ;
      RECT 17.750000 112.830000 60.635000 112.900000 ;
      RECT 17.750000 112.830000 60.635000 112.900000 ;
      RECT 17.760000  80.415000 24.540000  80.485000 ;
      RECT 17.760000  80.415000 24.540000  80.485000 ;
      RECT 17.760000  80.415000 58.420000  80.485000 ;
      RECT 17.760000 103.415000 24.540000 103.485000 ;
      RECT 17.760000 103.415000 24.540000 103.485000 ;
      RECT 17.760000 103.415000 58.420000 103.485000 ;
      RECT 17.765000  89.775000 60.830000  89.790000 ;
      RECT 17.765000  89.775000 60.830000  89.790000 ;
      RECT 17.765000 158.830000 60.685000 158.900000 ;
      RECT 17.765000 158.830000 60.685000 158.900000 ;
      RECT 17.775000  80.485000 24.540000  80.500000 ;
      RECT 17.775000  80.485000 24.540000  80.500000 ;
      RECT 17.775000  80.485000 58.490000  80.500000 ;
      RECT 17.775000 103.485000 24.540000 103.500000 ;
      RECT 17.775000 103.485000 24.540000 103.500000 ;
      RECT 17.775000 103.485000 58.490000 103.500000 ;
      RECT 17.780000  66.760000 60.735000  66.830000 ;
      RECT 17.780000  66.760000 60.735000  66.830000 ;
      RECT 17.780000  66.760000 60.970000  66.790000 ;
      RECT 17.780000  89.760000 60.830000  89.775000 ;
      RECT 17.780000  89.760000 60.830000  89.775000 ;
      RECT 17.780000  89.760000 60.970000  89.850000 ;
      RECT 17.780000 172.415000 58.430000 172.485000 ;
      RECT 17.785000  57.415000 58.390000  57.485000 ;
      RECT 17.785000 126.345000 24.540000 126.415000 ;
      RECT 17.785000 126.345000 24.540000 126.415000 ;
      RECT 17.785000 126.345000 58.350000 126.415000 ;
      RECT 17.785000 135.900000 60.600000 135.970000 ;
      RECT 17.785000 135.900000 60.600000 135.970000 ;
      RECT 17.785000 149.415000 58.350000 149.485000 ;
      RECT 17.785000 158.810000 57.585000 162.195000 ;
      RECT 17.795000 172.485000 58.500000 172.500000 ;
      RECT 17.800000  37.795000 54.390000  37.865000 ;
      RECT 17.800000  37.795000 54.390000  37.865000 ;
      RECT 17.800000  57.485000 58.460000  57.500000 ;
      RECT 17.800000 149.485000 58.420000 149.500000 ;
      RECT 17.810000 181.760000 60.830000 181.830000 ;
      RECT 17.810000 181.760000 60.970000 182.820000 ;
      RECT 17.815000  27.100000 56.860000  27.170000 ;
      RECT 17.815000  27.100000 56.860000  27.170000 ;
      RECT 17.820000 112.760000 57.550000 116.180000 ;
      RECT 17.820000 112.760000 60.705000 112.830000 ;
      RECT 17.820000 112.760000 60.705000 112.830000 ;
      RECT 17.820000 112.760000 60.970000 112.760000 ;
      RECT 17.835000 158.760000 60.755000 158.830000 ;
      RECT 17.835000 158.760000 60.755000 158.830000 ;
      RECT 17.835000 158.760000 60.970000 158.810000 ;
      RECT 17.855000 126.415000 24.540000 126.485000 ;
      RECT 17.855000 126.415000 24.540000 126.485000 ;
      RECT 17.855000 126.415000 58.420000 126.485000 ;
      RECT 17.855000 135.830000 60.670000 135.900000 ;
      RECT 17.855000 135.830000 60.670000 135.900000 ;
      RECT 17.870000  37.865000 54.390000  37.935000 ;
      RECT 17.870000  37.865000 54.390000  37.935000 ;
      RECT 17.870000 126.485000 24.540000 126.500000 ;
      RECT 17.870000 126.485000 24.540000 126.500000 ;
      RECT 17.870000 126.485000 58.490000 126.500000 ;
      RECT 17.885000  27.030000 56.790000  27.100000 ;
      RECT 17.885000  27.030000 56.790000  27.100000 ;
      RECT 17.890000 135.795000 57.480000 139.285000 ;
      RECT 17.925000 135.760000 60.740000 135.830000 ;
      RECT 17.925000 135.760000 60.740000 135.830000 ;
      RECT 17.925000 135.760000 60.970000 135.795000 ;
      RECT 17.940000  37.935000 54.390000  38.005000 ;
      RECT 17.940000  37.935000 54.390000  38.005000 ;
      RECT 17.955000  26.960000 56.720000  27.030000 ;
      RECT 17.955000  26.960000 56.720000  27.030000 ;
      RECT 18.010000  38.005000 54.390000  38.075000 ;
      RECT 18.010000  38.005000 54.390000  38.075000 ;
      RECT 18.025000  26.890000 56.650000  26.960000 ;
      RECT 18.025000  26.890000 56.650000  26.960000 ;
      RECT 18.075000  38.075000 54.390000  38.140000 ;
      RECT 18.075000  38.075000 54.390000  38.140000 ;
      RECT 18.095000  26.820000 56.580000  26.890000 ;
      RECT 18.095000  26.820000 56.580000  26.890000 ;
      RECT 18.130000  38.195000 52.655000  40.070000 ;
      RECT 18.145000  38.140000 54.320000  38.210000 ;
      RECT 18.145000  38.140000 54.320000  38.210000 ;
      RECT 18.165000  26.750000 56.510000  26.820000 ;
      RECT 18.165000  26.750000 56.510000  26.820000 ;
      RECT 18.215000  38.210000 54.250000  38.280000 ;
      RECT 18.215000  38.210000 54.250000  38.280000 ;
      RECT 18.235000  26.680000 56.440000  26.750000 ;
      RECT 18.235000  26.680000 56.440000  26.750000 ;
      RECT 18.285000  38.280000 54.180000  38.350000 ;
      RECT 18.285000  38.280000 54.180000  38.350000 ;
      RECT 18.305000  26.610000 56.370000  26.680000 ;
      RECT 18.305000  26.610000 56.370000  26.680000 ;
      RECT 18.355000  38.350000 54.110000  38.420000 ;
      RECT 18.355000  38.350000 54.110000  38.420000 ;
      RECT 18.375000  26.540000 56.300000  26.610000 ;
      RECT 18.375000  26.540000 56.300000  26.610000 ;
      RECT 18.425000  38.420000 54.040000  38.490000 ;
      RECT 18.425000  38.420000 54.040000  38.490000 ;
      RECT 18.445000  26.470000 56.230000  26.540000 ;
      RECT 18.445000  26.470000 56.230000  26.540000 ;
      RECT 18.495000  38.490000 53.970000  38.560000 ;
      RECT 18.495000  38.490000 53.970000  38.560000 ;
      RECT 18.515000  26.400000 56.160000  26.470000 ;
      RECT 18.515000  26.400000 56.160000  26.470000 ;
      RECT 18.565000  38.560000 53.900000  38.630000 ;
      RECT 18.565000  38.560000 53.900000  38.630000 ;
      RECT 18.585000  26.330000 56.090000  26.400000 ;
      RECT 18.585000  26.330000 56.090000  26.400000 ;
      RECT 18.635000  38.630000 53.830000  38.700000 ;
      RECT 18.635000  38.630000 53.830000  38.700000 ;
      RECT 18.655000  26.260000 56.020000  26.330000 ;
      RECT 18.655000  26.260000 56.020000  26.330000 ;
      RECT 18.705000  38.700000 53.760000  38.770000 ;
      RECT 18.705000  38.700000 53.760000  38.770000 ;
      RECT 18.725000  26.190000 55.950000  26.260000 ;
      RECT 18.725000  26.190000 55.950000  26.260000 ;
      RECT 18.775000  38.770000 53.690000  38.840000 ;
      RECT 18.775000  38.770000 53.690000  38.840000 ;
      RECT 18.795000  26.120000 55.880000  26.190000 ;
      RECT 18.795000  26.120000 55.880000  26.190000 ;
      RECT 18.845000  38.840000 53.620000  38.910000 ;
      RECT 18.845000  38.840000 53.620000  38.910000 ;
      RECT 18.865000  26.050000 55.810000  26.120000 ;
      RECT 18.865000  26.050000 55.810000  26.120000 ;
      RECT 18.915000  38.910000 53.550000  38.980000 ;
      RECT 18.915000  38.910000 53.550000  38.980000 ;
      RECT 18.935000  25.980000 55.740000  26.050000 ;
      RECT 18.935000  25.980000 55.740000  26.050000 ;
      RECT 18.935000  25.980000 59.390000  29.430000 ;
      RECT 18.985000  38.980000 53.480000  39.050000 ;
      RECT 18.985000  38.980000 53.480000  39.050000 ;
      RECT 19.055000  39.050000 53.410000  39.120000 ;
      RECT 19.055000  39.050000 53.410000  39.120000 ;
      RECT 19.125000  39.120000 53.340000  39.190000 ;
      RECT 19.125000  39.120000 53.340000  39.190000 ;
      RECT 19.195000  39.190000 53.270000  39.260000 ;
      RECT 19.195000  39.190000 53.270000  39.260000 ;
      RECT 19.265000  39.260000 53.200000  39.330000 ;
      RECT 19.265000  39.260000 53.200000  39.330000 ;
      RECT 19.335000  39.330000 53.130000  39.400000 ;
      RECT 19.335000  39.330000 53.130000  39.400000 ;
      RECT 19.405000  39.400000 53.060000  39.470000 ;
      RECT 19.405000  39.400000 53.060000  39.470000 ;
      RECT 19.475000  39.470000 52.990000  39.540000 ;
      RECT 19.475000  39.470000 52.990000  39.540000 ;
      RECT 19.545000  39.540000 52.920000  39.610000 ;
      RECT 19.545000  39.540000 52.920000  39.610000 ;
      RECT 19.615000  39.610000 52.850000  39.680000 ;
      RECT 19.615000  39.610000 52.850000  39.680000 ;
      RECT 19.685000  39.680000 52.780000  39.750000 ;
      RECT 19.685000  39.680000 52.780000  39.750000 ;
      RECT 19.755000  39.750000 52.710000  39.820000 ;
      RECT 19.755000  39.750000 52.710000  39.820000 ;
      RECT 19.825000  39.820000 52.640000  39.890000 ;
      RECT 19.825000  39.820000 52.640000  39.890000 ;
      RECT 19.895000  39.890000 52.570000  39.960000 ;
      RECT 19.895000  39.890000 52.570000  39.960000 ;
      RECT 19.965000  39.960000 52.500000  40.030000 ;
      RECT 19.965000  39.960000 52.500000  40.030000 ;
      RECT 20.005000  40.030000 52.460000  40.070000 ;
      RECT 20.005000  40.030000 52.460000  40.070000 ;
      RECT 20.400000  40.070000 52.515000  40.210000 ;
      RECT 22.850000  42.520000 60.970000  42.660000 ;
      RECT 24.675000   0.000000 25.615000   0.815000 ;
      RECT 24.675000   0.000000 25.755000   0.675000 ;
      RECT 24.675000   0.675000 50.250000   8.480000 ;
      RECT 24.675000   0.815000 50.110000   8.480000 ;
      RECT 24.675000   8.480000 50.250000   8.565000 ;
      RECT 24.690000   8.480000 50.110000   8.495000 ;
      RECT 24.690000   8.480000 50.110000   8.495000 ;
      RECT 24.705000   8.495000 50.110000   8.510000 ;
      RECT 24.705000   8.495000 50.110000   8.510000 ;
      RECT 24.765000   8.565000 46.695000  12.120000 ;
      RECT 24.775000   8.510000 50.040000   8.580000 ;
      RECT 24.775000   8.510000 50.040000   8.580000 ;
      RECT 24.845000   8.580000 49.970000   8.650000 ;
      RECT 24.845000   8.580000 49.970000   8.650000 ;
      RECT 24.915000   8.650000 49.900000   8.720000 ;
      RECT 24.915000   8.650000 49.900000   8.720000 ;
      RECT 24.985000   8.720000 49.830000   8.790000 ;
      RECT 24.985000   8.720000 49.830000   8.790000 ;
      RECT 25.055000   8.790000 49.760000   8.860000 ;
      RECT 25.055000   8.790000 49.760000   8.860000 ;
      RECT 25.125000   8.860000 49.690000   8.930000 ;
      RECT 25.125000   8.860000 49.690000   8.930000 ;
      RECT 25.195000   8.930000 49.620000   9.000000 ;
      RECT 25.195000   8.930000 49.620000   9.000000 ;
      RECT 25.265000   9.000000 49.550000   9.070000 ;
      RECT 25.265000   9.000000 49.550000   9.070000 ;
      RECT 25.335000   9.070000 49.480000   9.140000 ;
      RECT 25.335000   9.070000 49.480000   9.140000 ;
      RECT 25.405000   9.140000 49.410000   9.210000 ;
      RECT 25.405000   9.140000 49.410000   9.210000 ;
      RECT 25.475000   9.210000 49.340000   9.280000 ;
      RECT 25.475000   9.210000 49.340000   9.280000 ;
      RECT 25.545000   9.280000 49.270000   9.350000 ;
      RECT 25.545000   9.280000 49.270000   9.350000 ;
      RECT 25.615000   9.350000 49.200000   9.420000 ;
      RECT 25.615000   9.350000 49.200000   9.420000 ;
      RECT 25.685000   9.420000 49.130000   9.490000 ;
      RECT 25.685000   9.420000 49.130000   9.490000 ;
      RECT 25.755000   9.490000 49.060000   9.560000 ;
      RECT 25.755000   9.490000 49.060000   9.560000 ;
      RECT 25.825000   9.560000 48.990000   9.630000 ;
      RECT 25.825000   9.560000 48.990000   9.630000 ;
      RECT 25.895000   9.630000 48.920000   9.700000 ;
      RECT 25.895000   9.630000 48.920000   9.700000 ;
      RECT 25.965000   9.700000 48.850000   9.770000 ;
      RECT 25.965000   9.700000 48.850000   9.770000 ;
      RECT 26.035000   9.770000 48.780000   9.840000 ;
      RECT 26.035000   9.770000 48.780000   9.840000 ;
      RECT 26.105000   9.840000 48.710000   9.910000 ;
      RECT 26.105000   9.840000 48.710000   9.910000 ;
      RECT 26.175000   9.910000 48.640000   9.980000 ;
      RECT 26.175000   9.910000 48.640000   9.980000 ;
      RECT 26.245000   9.980000 48.570000  10.050000 ;
      RECT 26.245000   9.980000 48.570000  10.050000 ;
      RECT 26.315000  10.050000 48.500000  10.120000 ;
      RECT 26.315000  10.050000 48.500000  10.120000 ;
      RECT 26.385000  10.120000 48.430000  10.190000 ;
      RECT 26.385000  10.120000 48.430000  10.190000 ;
      RECT 26.455000  10.190000 48.360000  10.260000 ;
      RECT 26.455000  10.190000 48.360000  10.260000 ;
      RECT 26.525000  10.260000 48.290000  10.330000 ;
      RECT 26.525000  10.260000 48.290000  10.330000 ;
      RECT 26.595000  10.330000 48.220000  10.400000 ;
      RECT 26.595000  10.330000 48.220000  10.400000 ;
      RECT 26.665000  10.400000 48.150000  10.470000 ;
      RECT 26.665000  10.400000 48.150000  10.470000 ;
      RECT 26.735000  10.470000 48.080000  10.540000 ;
      RECT 26.735000  10.470000 48.080000  10.540000 ;
      RECT 26.805000  10.540000 48.010000  10.610000 ;
      RECT 26.805000  10.540000 48.010000  10.610000 ;
      RECT 26.875000  10.610000 47.940000  10.680000 ;
      RECT 26.875000  10.610000 47.940000  10.680000 ;
      RECT 26.945000  10.680000 47.870000  10.750000 ;
      RECT 26.945000  10.680000 47.870000  10.750000 ;
      RECT 27.015000  10.750000 47.800000  10.820000 ;
      RECT 27.015000  10.750000 47.800000  10.820000 ;
      RECT 27.085000  10.820000 47.730000  10.890000 ;
      RECT 27.085000  10.820000 47.730000  10.890000 ;
      RECT 27.155000  10.890000 47.660000  10.960000 ;
      RECT 27.155000  10.890000 47.660000  10.960000 ;
      RECT 27.225000  10.960000 47.590000  11.030000 ;
      RECT 27.225000  10.960000 47.590000  11.030000 ;
      RECT 27.295000  11.030000 47.520000  11.100000 ;
      RECT 27.295000  11.030000 47.520000  11.100000 ;
      RECT 27.365000  11.100000 47.450000  11.170000 ;
      RECT 27.365000  11.100000 47.450000  11.170000 ;
      RECT 27.435000  11.170000 47.380000  11.240000 ;
      RECT 27.435000  11.170000 47.380000  11.240000 ;
      RECT 27.505000  11.240000 47.310000  11.310000 ;
      RECT 27.505000  11.240000 47.310000  11.310000 ;
      RECT 27.575000  11.310000 47.240000  11.380000 ;
      RECT 27.575000  11.310000 47.240000  11.380000 ;
      RECT 27.645000  11.380000 47.170000  11.450000 ;
      RECT 27.645000  11.380000 47.170000  11.450000 ;
      RECT 27.715000  11.450000 47.100000  11.520000 ;
      RECT 27.715000  11.450000 47.100000  11.520000 ;
      RECT 27.785000  11.520000 47.030000  11.590000 ;
      RECT 27.785000  11.520000 47.030000  11.590000 ;
      RECT 27.855000  11.590000 46.960000  11.660000 ;
      RECT 27.855000  11.590000 46.960000  11.660000 ;
      RECT 27.925000  11.660000 46.890000  11.730000 ;
      RECT 27.925000  11.660000 46.890000  11.730000 ;
      RECT 27.995000  11.730000 46.820000  11.800000 ;
      RECT 27.995000  11.730000 46.820000  11.800000 ;
      RECT 28.035000   0.000000 50.250000   0.675000 ;
      RECT 28.065000  11.800000 46.750000  11.870000 ;
      RECT 28.065000  11.800000 46.750000  11.870000 ;
      RECT 28.135000  11.870000 46.680000  11.940000 ;
      RECT 28.135000  11.870000 46.680000  11.940000 ;
      RECT 28.175000   0.000000 50.110000   0.815000 ;
      RECT 28.175000   0.000000 50.110000   8.480000 ;
      RECT 28.205000  11.940000 46.610000  12.010000 ;
      RECT 28.205000  11.940000 46.610000  12.010000 ;
      RECT 28.210000  12.010000 46.605000  12.015000 ;
      RECT 28.210000  12.010000 46.605000  12.015000 ;
      RECT 28.260000  12.015000 37.610000  12.065000 ;
      RECT 28.260000  12.015000 37.610000  12.065000 ;
      RECT 28.310000  12.065000 37.610000  12.115000 ;
      RECT 28.310000  12.065000 37.610000  12.115000 ;
      RECT 28.315000  12.115000 37.610000  12.120000 ;
      RECT 28.315000  12.115000 37.610000  12.120000 ;
      RECT 37.175000  12.120000 37.610000  25.940000 ;
      RECT 37.175000  12.120000 46.660000  12.155000 ;
      RECT 37.175000  12.155000 37.750000  25.800000 ;
      RECT 37.175000  25.800000 55.935000  25.980000 ;
      RECT 37.175000  25.940000 55.700000  25.960000 ;
      RECT 37.175000  25.940000 55.700000  25.960000 ;
      RECT 37.175000  25.960000 55.720000  25.980000 ;
      RECT 37.175000  25.960000 55.720000  25.980000 ;
      RECT 54.325000  42.650000 60.830000  42.660000 ;
      RECT 54.325000  42.650000 60.830000  42.660000 ;
      RECT 54.395000  42.580000 60.830000  42.650000 ;
      RECT 54.395000  42.580000 60.830000  42.650000 ;
      RECT 54.465000  42.510000 60.830000  42.580000 ;
      RECT 54.465000  42.510000 60.830000  42.580000 ;
      RECT 54.535000  42.440000 60.830000  42.510000 ;
      RECT 54.535000  42.440000 60.830000  42.510000 ;
      RECT 54.605000  42.370000 60.830000  42.440000 ;
      RECT 54.605000  42.370000 60.830000  42.440000 ;
      RECT 54.675000  42.300000 60.830000  42.370000 ;
      RECT 54.675000  42.300000 60.830000  42.370000 ;
      RECT 54.745000  42.230000 60.830000  42.300000 ;
      RECT 54.745000  42.230000 60.830000  42.300000 ;
      RECT 54.815000  42.160000 60.830000  42.230000 ;
      RECT 54.815000  42.160000 60.830000  42.230000 ;
      RECT 54.885000  42.090000 60.830000  42.160000 ;
      RECT 54.885000  42.090000 60.830000  42.160000 ;
      RECT 54.955000  42.020000 60.830000  42.090000 ;
      RECT 54.955000  42.020000 60.830000  42.090000 ;
      RECT 55.025000  41.950000 60.830000  42.020000 ;
      RECT 55.025000  41.950000 60.830000  42.020000 ;
      RECT 55.095000  41.880000 60.830000  41.950000 ;
      RECT 55.095000  41.880000 60.830000  41.950000 ;
      RECT 55.165000  41.810000 60.830000  41.880000 ;
      RECT 55.165000  41.810000 60.830000  41.880000 ;
      RECT 55.235000  41.740000 60.830000  41.810000 ;
      RECT 55.235000  41.740000 60.830000  41.810000 ;
      RECT 55.305000  41.670000 60.830000  41.740000 ;
      RECT 55.305000  41.670000 60.830000  41.740000 ;
      RECT 55.375000  41.600000 60.830000  41.670000 ;
      RECT 55.375000  41.600000 60.830000  41.670000 ;
      RECT 55.445000  41.530000 60.830000  41.600000 ;
      RECT 55.445000  41.530000 60.830000  41.600000 ;
      RECT 55.515000  41.460000 60.830000  41.530000 ;
      RECT 55.515000  41.460000 60.830000  41.530000 ;
      RECT 55.585000  41.390000 60.830000  41.460000 ;
      RECT 55.585000  41.390000 60.830000  41.460000 ;
      RECT 55.655000  41.320000 60.830000  41.390000 ;
      RECT 55.655000  41.320000 60.830000  41.390000 ;
      RECT 55.725000  41.250000 60.830000  41.320000 ;
      RECT 55.725000  41.250000 60.830000  41.320000 ;
      RECT 55.795000  41.180000 60.830000  41.250000 ;
      RECT 55.795000  41.180000 60.830000  41.250000 ;
      RECT 55.865000  41.110000 60.830000  41.180000 ;
      RECT 55.865000  41.110000 60.830000  41.180000 ;
      RECT 55.935000  41.040000 60.830000  41.110000 ;
      RECT 55.935000  41.040000 60.830000  41.110000 ;
      RECT 56.005000  40.970000 60.830000  41.040000 ;
      RECT 56.005000  40.970000 60.830000  41.040000 ;
      RECT 56.075000  40.900000 60.830000  40.970000 ;
      RECT 56.075000  40.900000 60.830000  40.970000 ;
      RECT 56.145000  40.830000 60.830000  40.900000 ;
      RECT 56.145000  40.830000 60.830000  40.900000 ;
      RECT 56.215000  40.760000 60.830000  40.830000 ;
      RECT 56.215000  40.760000 60.830000  40.830000 ;
      RECT 56.285000  40.690000 60.830000  40.760000 ;
      RECT 56.285000  40.690000 60.830000  40.760000 ;
      RECT 56.355000  40.620000 60.830000  40.690000 ;
      RECT 56.355000  40.620000 60.830000  40.690000 ;
      RECT 56.425000  40.550000 60.830000  40.620000 ;
      RECT 56.425000  40.550000 60.830000  40.620000 ;
      RECT 56.495000  40.480000 60.830000  40.550000 ;
      RECT 56.495000  40.480000 60.830000  40.550000 ;
      RECT 56.565000  40.410000 60.830000  40.480000 ;
      RECT 56.565000  40.410000 60.830000  40.480000 ;
      RECT 56.635000  40.340000 60.830000  40.410000 ;
      RECT 56.635000  40.340000 60.830000  40.410000 ;
      RECT 56.705000  40.270000 60.830000  40.340000 ;
      RECT 56.705000  40.270000 60.830000  40.340000 ;
      RECT 56.775000  40.200000 60.830000  40.270000 ;
      RECT 56.775000  40.200000 60.830000  40.270000 ;
      RECT 56.845000  40.130000 60.830000  40.200000 ;
      RECT 56.845000  40.130000 60.830000  40.200000 ;
      RECT 56.915000  40.060000 60.830000  40.130000 ;
      RECT 56.915000  40.060000 60.830000  40.130000 ;
      RECT 56.985000  39.990000 60.830000  40.060000 ;
      RECT 56.985000  39.990000 60.830000  40.060000 ;
      RECT 56.985000  79.435000 57.440000  79.505000 ;
      RECT 56.985000  79.435000 57.440000  79.505000 ;
      RECT 56.985000  79.505000 57.510000  79.575000 ;
      RECT 56.985000  79.505000 57.510000  79.575000 ;
      RECT 56.985000  79.575000 57.580000  79.645000 ;
      RECT 56.985000  79.575000 57.580000  79.645000 ;
      RECT 56.985000  79.645000 57.650000  79.715000 ;
      RECT 56.985000  79.645000 57.650000  79.715000 ;
      RECT 56.985000  79.715000 57.720000  79.785000 ;
      RECT 56.985000  79.715000 57.720000  79.785000 ;
      RECT 56.985000  79.785000 57.790000  79.855000 ;
      RECT 56.985000  79.785000 57.790000  79.855000 ;
      RECT 56.985000  79.855000 57.860000  79.925000 ;
      RECT 56.985000  79.855000 57.860000  79.925000 ;
      RECT 56.985000  79.925000 57.930000  79.995000 ;
      RECT 56.985000  79.925000 57.930000  79.995000 ;
      RECT 56.985000  79.995000 58.000000  80.065000 ;
      RECT 56.985000  79.995000 58.000000  80.065000 ;
      RECT 56.985000  80.065000 58.070000  80.135000 ;
      RECT 56.985000  80.065000 58.070000  80.135000 ;
      RECT 56.985000  80.135000 58.140000  80.205000 ;
      RECT 56.985000  80.135000 58.140000  80.205000 ;
      RECT 56.985000  80.205000 58.210000  80.275000 ;
      RECT 56.985000  80.205000 58.210000  80.275000 ;
      RECT 56.985000  80.275000 58.280000  80.345000 ;
      RECT 56.985000  80.275000 58.280000  80.345000 ;
      RECT 56.985000  80.345000 58.350000  80.415000 ;
      RECT 56.985000  80.345000 58.350000  80.415000 ;
      RECT 56.985000  80.415000 58.420000  80.485000 ;
      RECT 56.985000  80.415000 58.420000  80.485000 ;
      RECT 56.985000  80.485000 58.490000  80.500000 ;
      RECT 56.985000  80.485000 58.490000  80.500000 ;
      RECT 56.985000  80.500000 58.505000  80.570000 ;
      RECT 56.985000  80.500000 58.505000  80.570000 ;
      RECT 56.985000  80.500000 60.970000  82.770000 ;
      RECT 56.985000  80.570000 58.575000  80.640000 ;
      RECT 56.985000  80.570000 58.575000  80.640000 ;
      RECT 56.985000  80.640000 58.645000  80.710000 ;
      RECT 56.985000  80.640000 58.645000  80.710000 ;
      RECT 56.985000  80.710000 58.715000  80.780000 ;
      RECT 56.985000  80.710000 58.715000  80.780000 ;
      RECT 56.985000  80.780000 58.785000  80.850000 ;
      RECT 56.985000  80.780000 58.785000  80.850000 ;
      RECT 56.985000  80.850000 58.855000  80.920000 ;
      RECT 56.985000  80.850000 58.855000  80.920000 ;
      RECT 56.985000  80.920000 58.925000  80.990000 ;
      RECT 56.985000  80.920000 58.925000  80.990000 ;
      RECT 56.985000  80.990000 58.995000  81.060000 ;
      RECT 56.985000  80.990000 58.995000  81.060000 ;
      RECT 56.985000  81.060000 59.065000  81.130000 ;
      RECT 56.985000  81.060000 59.065000  81.130000 ;
      RECT 56.985000  81.130000 59.135000  81.200000 ;
      RECT 56.985000  81.130000 59.135000  81.200000 ;
      RECT 56.985000  81.200000 59.205000  81.270000 ;
      RECT 56.985000  81.200000 59.205000  81.270000 ;
      RECT 56.985000  81.270000 59.275000  81.340000 ;
      RECT 56.985000  81.270000 59.275000  81.340000 ;
      RECT 56.985000  81.340000 59.345000  81.410000 ;
      RECT 56.985000  81.340000 59.345000  81.410000 ;
      RECT 56.985000  81.410000 59.415000  81.480000 ;
      RECT 56.985000  81.410000 59.415000  81.480000 ;
      RECT 56.985000  81.480000 59.485000  81.550000 ;
      RECT 56.985000  81.480000 59.485000  81.550000 ;
      RECT 56.985000  81.550000 59.555000  81.620000 ;
      RECT 56.985000  81.550000 59.555000  81.620000 ;
      RECT 56.985000  81.620000 59.625000  81.690000 ;
      RECT 56.985000  81.620000 59.625000  81.690000 ;
      RECT 56.985000  81.690000 59.695000  81.760000 ;
      RECT 56.985000  81.690000 59.695000  81.760000 ;
      RECT 56.985000  81.760000 59.765000  81.830000 ;
      RECT 56.985000  81.760000 59.765000  81.830000 ;
      RECT 56.985000  81.830000 59.835000  81.900000 ;
      RECT 56.985000  81.830000 59.835000  81.900000 ;
      RECT 56.985000  81.900000 59.905000  81.970000 ;
      RECT 56.985000  81.900000 59.905000  81.970000 ;
      RECT 56.985000  81.970000 59.975000  82.040000 ;
      RECT 56.985000  81.970000 59.975000  82.040000 ;
      RECT 56.985000  82.040000 60.045000  82.110000 ;
      RECT 56.985000  82.040000 60.045000  82.110000 ;
      RECT 56.985000  82.110000 60.115000  82.180000 ;
      RECT 56.985000  82.110000 60.115000  82.180000 ;
      RECT 56.985000  82.180000 60.185000  82.250000 ;
      RECT 56.985000  82.180000 60.185000  82.250000 ;
      RECT 56.985000  82.250000 60.255000  82.320000 ;
      RECT 56.985000  82.250000 60.255000  82.320000 ;
      RECT 56.985000  82.320000 60.325000  82.390000 ;
      RECT 56.985000  82.320000 60.325000  82.390000 ;
      RECT 56.985000  82.390000 60.395000  82.460000 ;
      RECT 56.985000  82.390000 60.395000  82.460000 ;
      RECT 56.985000  82.460000 60.465000  82.530000 ;
      RECT 56.985000  82.460000 60.465000  82.530000 ;
      RECT 56.985000  82.530000 60.535000  82.600000 ;
      RECT 56.985000  82.530000 60.535000  82.600000 ;
      RECT 56.985000  82.600000 60.605000  82.670000 ;
      RECT 56.985000  82.600000 60.605000  82.670000 ;
      RECT 56.985000  82.670000 60.675000  82.740000 ;
      RECT 56.985000  82.670000 60.675000  82.740000 ;
      RECT 56.985000  82.740000 60.745000  82.810000 ;
      RECT 56.985000  82.740000 60.745000  82.810000 ;
      RECT 56.985000  82.770000 60.970000  89.760000 ;
      RECT 56.985000  82.810000 60.815000  82.825000 ;
      RECT 56.985000  82.810000 60.815000  82.825000 ;
      RECT 56.985000  82.825000 60.830000  89.760000 ;
      RECT 56.985000 102.435000 57.440000 102.505000 ;
      RECT 56.985000 102.435000 57.440000 102.505000 ;
      RECT 56.985000 102.505000 57.510000 102.575000 ;
      RECT 56.985000 102.505000 57.510000 102.575000 ;
      RECT 56.985000 102.575000 57.580000 102.645000 ;
      RECT 56.985000 102.575000 57.580000 102.645000 ;
      RECT 56.985000 102.645000 57.650000 102.715000 ;
      RECT 56.985000 102.645000 57.650000 102.715000 ;
      RECT 56.985000 102.715000 57.720000 102.785000 ;
      RECT 56.985000 102.715000 57.720000 102.785000 ;
      RECT 56.985000 102.785000 57.790000 102.855000 ;
      RECT 56.985000 102.785000 57.790000 102.855000 ;
      RECT 56.985000 102.855000 57.860000 102.925000 ;
      RECT 56.985000 102.855000 57.860000 102.925000 ;
      RECT 56.985000 102.925000 57.930000 102.995000 ;
      RECT 56.985000 102.925000 57.930000 102.995000 ;
      RECT 56.985000 102.995000 58.000000 103.065000 ;
      RECT 56.985000 102.995000 58.000000 103.065000 ;
      RECT 56.985000 103.065000 58.070000 103.135000 ;
      RECT 56.985000 103.065000 58.070000 103.135000 ;
      RECT 56.985000 103.135000 58.140000 103.205000 ;
      RECT 56.985000 103.135000 58.140000 103.205000 ;
      RECT 56.985000 103.205000 58.210000 103.275000 ;
      RECT 56.985000 103.205000 58.210000 103.275000 ;
      RECT 56.985000 103.275000 58.280000 103.345000 ;
      RECT 56.985000 103.275000 58.280000 103.345000 ;
      RECT 56.985000 103.345000 58.350000 103.415000 ;
      RECT 56.985000 103.345000 58.350000 103.415000 ;
      RECT 56.985000 103.415000 58.420000 103.485000 ;
      RECT 56.985000 103.415000 58.420000 103.485000 ;
      RECT 56.985000 103.485000 58.490000 103.500000 ;
      RECT 56.985000 103.485000 58.490000 103.500000 ;
      RECT 56.985000 103.500000 58.505000 103.570000 ;
      RECT 56.985000 103.500000 58.505000 103.570000 ;
      RECT 56.985000 103.500000 60.970000 105.770000 ;
      RECT 56.985000 103.570000 58.575000 103.640000 ;
      RECT 56.985000 103.570000 58.575000 103.640000 ;
      RECT 56.985000 103.640000 58.645000 103.710000 ;
      RECT 56.985000 103.640000 58.645000 103.710000 ;
      RECT 56.985000 103.710000 58.715000 103.780000 ;
      RECT 56.985000 103.710000 58.715000 103.780000 ;
      RECT 56.985000 103.780000 58.785000 103.850000 ;
      RECT 56.985000 103.780000 58.785000 103.850000 ;
      RECT 56.985000 103.850000 58.855000 103.920000 ;
      RECT 56.985000 103.850000 58.855000 103.920000 ;
      RECT 56.985000 103.920000 58.925000 103.990000 ;
      RECT 56.985000 103.920000 58.925000 103.990000 ;
      RECT 56.985000 103.990000 58.995000 104.060000 ;
      RECT 56.985000 103.990000 58.995000 104.060000 ;
      RECT 56.985000 104.060000 59.065000 104.130000 ;
      RECT 56.985000 104.060000 59.065000 104.130000 ;
      RECT 56.985000 104.130000 59.135000 104.200000 ;
      RECT 56.985000 104.130000 59.135000 104.200000 ;
      RECT 56.985000 104.200000 59.205000 104.270000 ;
      RECT 56.985000 104.200000 59.205000 104.270000 ;
      RECT 56.985000 104.270000 59.275000 104.340000 ;
      RECT 56.985000 104.270000 59.275000 104.340000 ;
      RECT 56.985000 104.340000 59.345000 104.410000 ;
      RECT 56.985000 104.340000 59.345000 104.410000 ;
      RECT 56.985000 104.410000 59.415000 104.480000 ;
      RECT 56.985000 104.410000 59.415000 104.480000 ;
      RECT 56.985000 104.480000 59.485000 104.550000 ;
      RECT 56.985000 104.480000 59.485000 104.550000 ;
      RECT 56.985000 104.550000 59.555000 104.620000 ;
      RECT 56.985000 104.550000 59.555000 104.620000 ;
      RECT 56.985000 104.620000 59.625000 104.690000 ;
      RECT 56.985000 104.620000 59.625000 104.690000 ;
      RECT 56.985000 104.690000 59.695000 104.760000 ;
      RECT 56.985000 104.690000 59.695000 104.760000 ;
      RECT 56.985000 104.760000 59.765000 104.830000 ;
      RECT 56.985000 104.760000 59.765000 104.830000 ;
      RECT 56.985000 104.830000 59.835000 104.900000 ;
      RECT 56.985000 104.830000 59.835000 104.900000 ;
      RECT 56.985000 104.900000 59.905000 104.970000 ;
      RECT 56.985000 104.900000 59.905000 104.970000 ;
      RECT 56.985000 104.970000 59.975000 105.040000 ;
      RECT 56.985000 104.970000 59.975000 105.040000 ;
      RECT 56.985000 105.040000 60.045000 105.110000 ;
      RECT 56.985000 105.040000 60.045000 105.110000 ;
      RECT 56.985000 105.110000 60.115000 105.180000 ;
      RECT 56.985000 105.110000 60.115000 105.180000 ;
      RECT 56.985000 105.180000 60.185000 105.250000 ;
      RECT 56.985000 105.180000 60.185000 105.250000 ;
      RECT 56.985000 105.250000 60.255000 105.320000 ;
      RECT 56.985000 105.250000 60.255000 105.320000 ;
      RECT 56.985000 105.320000 60.325000 105.390000 ;
      RECT 56.985000 105.320000 60.325000 105.390000 ;
      RECT 56.985000 105.390000 60.395000 105.460000 ;
      RECT 56.985000 105.390000 60.395000 105.460000 ;
      RECT 56.985000 105.460000 60.465000 105.530000 ;
      RECT 56.985000 105.460000 60.465000 105.530000 ;
      RECT 56.985000 105.530000 60.535000 105.600000 ;
      RECT 56.985000 105.530000 60.535000 105.600000 ;
      RECT 56.985000 105.600000 60.605000 105.670000 ;
      RECT 56.985000 105.600000 60.605000 105.670000 ;
      RECT 56.985000 105.670000 60.675000 105.740000 ;
      RECT 56.985000 105.670000 60.675000 105.740000 ;
      RECT 56.985000 105.740000 60.745000 105.810000 ;
      RECT 56.985000 105.740000 60.745000 105.810000 ;
      RECT 56.985000 105.770000 60.970000 112.760000 ;
      RECT 56.985000 105.810000 60.815000 105.825000 ;
      RECT 56.985000 105.810000 60.815000 105.825000 ;
      RECT 56.985000 105.825000 60.830000 112.705000 ;
      RECT 56.985000 112.705000 60.805000 112.730000 ;
      RECT 56.985000 112.705000 60.805000 112.730000 ;
      RECT 56.985000 112.730000 60.775000 112.760000 ;
      RECT 56.985000 112.730000 60.775000 112.760000 ;
      RECT 56.985000 125.435000 57.440000 125.505000 ;
      RECT 56.985000 125.435000 57.440000 125.505000 ;
      RECT 56.985000 125.505000 57.510000 125.575000 ;
      RECT 56.985000 125.505000 57.510000 125.575000 ;
      RECT 56.985000 125.575000 57.580000 125.645000 ;
      RECT 56.985000 125.575000 57.580000 125.645000 ;
      RECT 56.985000 125.645000 57.650000 125.715000 ;
      RECT 56.985000 125.645000 57.650000 125.715000 ;
      RECT 56.985000 125.715000 57.720000 125.785000 ;
      RECT 56.985000 125.715000 57.720000 125.785000 ;
      RECT 56.985000 125.785000 57.790000 125.855000 ;
      RECT 56.985000 125.785000 57.790000 125.855000 ;
      RECT 56.985000 125.855000 57.860000 125.925000 ;
      RECT 56.985000 125.855000 57.860000 125.925000 ;
      RECT 56.985000 125.925000 57.930000 125.995000 ;
      RECT 56.985000 125.925000 57.930000 125.995000 ;
      RECT 56.985000 125.995000 58.000000 126.065000 ;
      RECT 56.985000 125.995000 58.000000 126.065000 ;
      RECT 56.985000 126.065000 58.070000 126.135000 ;
      RECT 56.985000 126.065000 58.070000 126.135000 ;
      RECT 56.985000 126.135000 58.140000 126.205000 ;
      RECT 56.985000 126.135000 58.140000 126.205000 ;
      RECT 56.985000 126.205000 58.210000 126.275000 ;
      RECT 56.985000 126.205000 58.210000 126.275000 ;
      RECT 56.985000 126.275000 58.280000 126.345000 ;
      RECT 56.985000 126.275000 58.280000 126.345000 ;
      RECT 56.985000 126.345000 58.350000 126.415000 ;
      RECT 56.985000 126.345000 58.350000 126.415000 ;
      RECT 56.985000 126.415000 58.420000 126.485000 ;
      RECT 56.985000 126.415000 58.420000 126.485000 ;
      RECT 56.985000 126.485000 58.490000 126.500000 ;
      RECT 56.985000 126.485000 58.490000 126.500000 ;
      RECT 56.985000 126.500000 58.505000 126.570000 ;
      RECT 56.985000 126.500000 58.505000 126.570000 ;
      RECT 56.985000 126.500000 60.970000 128.770000 ;
      RECT 56.985000 126.570000 58.575000 126.640000 ;
      RECT 56.985000 126.570000 58.575000 126.640000 ;
      RECT 56.985000 126.640000 58.645000 126.710000 ;
      RECT 56.985000 126.640000 58.645000 126.710000 ;
      RECT 56.985000 126.710000 58.715000 126.780000 ;
      RECT 56.985000 126.710000 58.715000 126.780000 ;
      RECT 56.985000 126.780000 58.785000 126.850000 ;
      RECT 56.985000 126.780000 58.785000 126.850000 ;
      RECT 56.985000 126.850000 58.855000 126.920000 ;
      RECT 56.985000 126.850000 58.855000 126.920000 ;
      RECT 56.985000 126.920000 58.925000 126.990000 ;
      RECT 56.985000 126.920000 58.925000 126.990000 ;
      RECT 56.985000 126.990000 58.995000 127.060000 ;
      RECT 56.985000 126.990000 58.995000 127.060000 ;
      RECT 56.985000 127.060000 59.065000 127.130000 ;
      RECT 56.985000 127.060000 59.065000 127.130000 ;
      RECT 56.985000 127.130000 59.135000 127.200000 ;
      RECT 56.985000 127.130000 59.135000 127.200000 ;
      RECT 56.985000 127.200000 59.205000 127.270000 ;
      RECT 56.985000 127.200000 59.205000 127.270000 ;
      RECT 56.985000 127.270000 59.275000 127.340000 ;
      RECT 56.985000 127.270000 59.275000 127.340000 ;
      RECT 56.985000 127.340000 59.345000 127.410000 ;
      RECT 56.985000 127.340000 59.345000 127.410000 ;
      RECT 56.985000 127.410000 59.415000 127.480000 ;
      RECT 56.985000 127.410000 59.415000 127.480000 ;
      RECT 56.985000 127.480000 59.485000 127.550000 ;
      RECT 56.985000 127.480000 59.485000 127.550000 ;
      RECT 56.985000 127.550000 59.555000 127.620000 ;
      RECT 56.985000 127.550000 59.555000 127.620000 ;
      RECT 56.985000 127.620000 59.625000 127.690000 ;
      RECT 56.985000 127.620000 59.625000 127.690000 ;
      RECT 56.985000 127.690000 59.695000 127.760000 ;
      RECT 56.985000 127.690000 59.695000 127.760000 ;
      RECT 56.985000 127.760000 59.765000 127.830000 ;
      RECT 56.985000 127.760000 59.765000 127.830000 ;
      RECT 56.985000 127.830000 59.835000 127.900000 ;
      RECT 56.985000 127.830000 59.835000 127.900000 ;
      RECT 56.985000 127.900000 59.905000 127.970000 ;
      RECT 56.985000 127.900000 59.905000 127.970000 ;
      RECT 56.985000 127.970000 59.975000 128.040000 ;
      RECT 56.985000 127.970000 59.975000 128.040000 ;
      RECT 56.985000 128.040000 60.045000 128.110000 ;
      RECT 56.985000 128.040000 60.045000 128.110000 ;
      RECT 56.985000 128.110000 60.115000 128.180000 ;
      RECT 56.985000 128.110000 60.115000 128.180000 ;
      RECT 56.985000 128.180000 60.185000 128.250000 ;
      RECT 56.985000 128.180000 60.185000 128.250000 ;
      RECT 56.985000 128.250000 60.255000 128.320000 ;
      RECT 56.985000 128.250000 60.255000 128.320000 ;
      RECT 56.985000 128.320000 60.325000 128.390000 ;
      RECT 56.985000 128.320000 60.325000 128.390000 ;
      RECT 56.985000 128.390000 60.395000 128.460000 ;
      RECT 56.985000 128.390000 60.395000 128.460000 ;
      RECT 56.985000 128.460000 60.465000 128.530000 ;
      RECT 56.985000 128.460000 60.465000 128.530000 ;
      RECT 56.985000 128.530000 60.535000 128.600000 ;
      RECT 56.985000 128.530000 60.535000 128.600000 ;
      RECT 56.985000 128.600000 60.605000 128.670000 ;
      RECT 56.985000 128.600000 60.605000 128.670000 ;
      RECT 56.985000 128.670000 60.675000 128.740000 ;
      RECT 56.985000 128.670000 60.675000 128.740000 ;
      RECT 56.985000 128.740000 60.745000 128.810000 ;
      RECT 56.985000 128.740000 60.745000 128.810000 ;
      RECT 56.985000 128.770000 60.970000 135.760000 ;
      RECT 56.985000 128.810000 60.815000 128.825000 ;
      RECT 56.985000 128.810000 60.815000 128.825000 ;
      RECT 56.985000 128.825000 60.830000 135.740000 ;
      RECT 56.985000 135.740000 60.820000 135.750000 ;
      RECT 56.985000 135.740000 60.820000 135.750000 ;
      RECT 56.985000 135.750000 60.810000 135.760000 ;
      RECT 56.985000 135.750000 60.810000 135.760000 ;
      RECT 56.985000 148.435000 57.370000 148.505000 ;
      RECT 56.985000 148.435000 57.370000 148.505000 ;
      RECT 56.985000 148.505000 57.440000 148.575000 ;
      RECT 56.985000 148.505000 57.440000 148.575000 ;
      RECT 56.985000 148.575000 57.510000 148.645000 ;
      RECT 56.985000 148.575000 57.510000 148.645000 ;
      RECT 56.985000 148.645000 57.580000 148.715000 ;
      RECT 56.985000 148.645000 57.580000 148.715000 ;
      RECT 56.985000 148.715000 57.650000 148.785000 ;
      RECT 56.985000 148.715000 57.650000 148.785000 ;
      RECT 56.985000 148.785000 57.720000 148.855000 ;
      RECT 56.985000 148.785000 57.720000 148.855000 ;
      RECT 56.985000 148.855000 57.790000 148.925000 ;
      RECT 56.985000 148.855000 57.790000 148.925000 ;
      RECT 56.985000 148.925000 57.860000 148.995000 ;
      RECT 56.985000 148.925000 57.860000 148.995000 ;
      RECT 56.985000 148.995000 57.930000 149.065000 ;
      RECT 56.985000 148.995000 57.930000 149.065000 ;
      RECT 56.985000 149.065000 58.000000 149.135000 ;
      RECT 56.985000 149.065000 58.000000 149.135000 ;
      RECT 56.985000 149.135000 58.070000 149.205000 ;
      RECT 56.985000 149.135000 58.070000 149.205000 ;
      RECT 56.985000 149.205000 58.140000 149.275000 ;
      RECT 56.985000 149.205000 58.140000 149.275000 ;
      RECT 56.985000 149.275000 58.210000 149.345000 ;
      RECT 56.985000 149.275000 58.210000 149.345000 ;
      RECT 56.985000 149.345000 58.280000 149.415000 ;
      RECT 56.985000 149.345000 58.280000 149.415000 ;
      RECT 56.985000 149.415000 58.350000 149.485000 ;
      RECT 56.985000 149.415000 58.350000 149.485000 ;
      RECT 56.985000 149.485000 58.420000 149.500000 ;
      RECT 56.985000 149.485000 58.420000 149.500000 ;
      RECT 56.985000 149.500000 58.435000 149.570000 ;
      RECT 56.985000 149.500000 58.435000 149.570000 ;
      RECT 56.985000 149.500000 60.970000 151.840000 ;
      RECT 56.985000 149.570000 58.505000 149.640000 ;
      RECT 56.985000 149.570000 58.505000 149.640000 ;
      RECT 56.985000 149.640000 58.575000 149.710000 ;
      RECT 56.985000 149.640000 58.575000 149.710000 ;
      RECT 56.985000 149.710000 58.645000 149.780000 ;
      RECT 56.985000 149.710000 58.645000 149.780000 ;
      RECT 56.985000 149.780000 58.715000 149.850000 ;
      RECT 56.985000 149.780000 58.715000 149.850000 ;
      RECT 56.985000 149.850000 58.785000 149.920000 ;
      RECT 56.985000 149.850000 58.785000 149.920000 ;
      RECT 56.985000 149.920000 58.855000 149.990000 ;
      RECT 56.985000 149.920000 58.855000 149.990000 ;
      RECT 56.985000 149.990000 58.925000 150.060000 ;
      RECT 56.985000 149.990000 58.925000 150.060000 ;
      RECT 56.985000 150.060000 58.995000 150.130000 ;
      RECT 56.985000 150.060000 58.995000 150.130000 ;
      RECT 56.985000 150.130000 59.065000 150.200000 ;
      RECT 56.985000 150.130000 59.065000 150.200000 ;
      RECT 56.985000 150.200000 59.135000 150.270000 ;
      RECT 56.985000 150.200000 59.135000 150.270000 ;
      RECT 56.985000 150.270000 59.205000 150.340000 ;
      RECT 56.985000 150.270000 59.205000 150.340000 ;
      RECT 56.985000 150.340000 59.275000 150.410000 ;
      RECT 56.985000 150.340000 59.275000 150.410000 ;
      RECT 56.985000 150.410000 59.345000 150.480000 ;
      RECT 56.985000 150.410000 59.345000 150.480000 ;
      RECT 56.985000 150.480000 59.415000 150.550000 ;
      RECT 56.985000 150.480000 59.415000 150.550000 ;
      RECT 56.985000 150.550000 59.485000 150.620000 ;
      RECT 56.985000 150.550000 59.485000 150.620000 ;
      RECT 56.985000 150.620000 59.555000 150.690000 ;
      RECT 56.985000 150.620000 59.555000 150.690000 ;
      RECT 56.985000 150.690000 59.625000 150.760000 ;
      RECT 56.985000 150.690000 59.625000 150.760000 ;
      RECT 56.985000 150.760000 59.695000 150.830000 ;
      RECT 56.985000 150.760000 59.695000 150.830000 ;
      RECT 56.985000 150.830000 59.765000 150.900000 ;
      RECT 56.985000 150.830000 59.765000 150.900000 ;
      RECT 56.985000 150.900000 59.835000 150.970000 ;
      RECT 56.985000 150.900000 59.835000 150.970000 ;
      RECT 56.985000 150.970000 59.905000 151.040000 ;
      RECT 56.985000 150.970000 59.905000 151.040000 ;
      RECT 56.985000 151.040000 59.975000 151.110000 ;
      RECT 56.985000 151.040000 59.975000 151.110000 ;
      RECT 56.985000 151.110000 60.045000 151.180000 ;
      RECT 56.985000 151.110000 60.045000 151.180000 ;
      RECT 56.985000 151.180000 60.115000 151.250000 ;
      RECT 56.985000 151.180000 60.115000 151.250000 ;
      RECT 56.985000 151.250000 60.185000 151.320000 ;
      RECT 56.985000 151.250000 60.185000 151.320000 ;
      RECT 56.985000 151.320000 60.255000 151.390000 ;
      RECT 56.985000 151.320000 60.255000 151.390000 ;
      RECT 56.985000 151.390000 60.325000 151.460000 ;
      RECT 56.985000 151.390000 60.325000 151.460000 ;
      RECT 56.985000 151.460000 60.395000 151.530000 ;
      RECT 56.985000 151.460000 60.395000 151.530000 ;
      RECT 56.985000 151.530000 60.465000 151.600000 ;
      RECT 56.985000 151.530000 60.465000 151.600000 ;
      RECT 56.985000 151.600000 60.535000 151.670000 ;
      RECT 56.985000 151.600000 60.535000 151.670000 ;
      RECT 56.985000 151.670000 60.605000 151.740000 ;
      RECT 56.985000 151.670000 60.605000 151.740000 ;
      RECT 56.985000 151.740000 60.675000 151.810000 ;
      RECT 56.985000 151.740000 60.675000 151.810000 ;
      RECT 56.985000 151.810000 60.745000 151.880000 ;
      RECT 56.985000 151.810000 60.745000 151.880000 ;
      RECT 56.985000 151.840000 60.970000 158.760000 ;
      RECT 56.985000 151.880000 60.815000 151.895000 ;
      RECT 56.985000 151.880000 60.815000 151.895000 ;
      RECT 56.985000 151.895000 60.830000 158.755000 ;
      RECT 56.985000 158.755000 60.825000 158.760000 ;
      RECT 56.985000 158.755000 60.825000 158.760000 ;
      RECT 56.990000  56.435000 57.410000  56.505000 ;
      RECT 56.990000  56.435000 57.410000  56.505000 ;
      RECT 56.990000  56.505000 57.480000  56.575000 ;
      RECT 56.990000  56.505000 57.480000  56.575000 ;
      RECT 56.990000  56.575000 57.550000  56.645000 ;
      RECT 56.990000  56.575000 57.550000  56.645000 ;
      RECT 56.990000  56.645000 57.620000  56.715000 ;
      RECT 56.990000  56.645000 57.620000  56.715000 ;
      RECT 56.990000  56.715000 57.690000  56.785000 ;
      RECT 56.990000  56.715000 57.690000  56.785000 ;
      RECT 56.990000  56.785000 57.760000  56.855000 ;
      RECT 56.990000  56.785000 57.760000  56.855000 ;
      RECT 56.990000  56.855000 57.830000  56.925000 ;
      RECT 56.990000  56.855000 57.830000  56.925000 ;
      RECT 56.990000  56.925000 57.900000  56.995000 ;
      RECT 56.990000  56.925000 57.900000  56.995000 ;
      RECT 56.990000  56.995000 57.970000  57.065000 ;
      RECT 56.990000  56.995000 57.970000  57.065000 ;
      RECT 56.990000  57.065000 58.040000  57.135000 ;
      RECT 56.990000  57.065000 58.040000  57.135000 ;
      RECT 56.990000  57.135000 58.110000  57.205000 ;
      RECT 56.990000  57.135000 58.110000  57.205000 ;
      RECT 56.990000  57.205000 58.180000  57.275000 ;
      RECT 56.990000  57.205000 58.180000  57.275000 ;
      RECT 56.990000  57.275000 58.250000  57.345000 ;
      RECT 56.990000  57.275000 58.250000  57.345000 ;
      RECT 56.990000  57.345000 58.320000  57.415000 ;
      RECT 56.990000  57.345000 58.320000  57.415000 ;
      RECT 56.990000  57.415000 58.390000  57.485000 ;
      RECT 56.990000  57.415000 58.390000  57.485000 ;
      RECT 56.990000  57.485000 58.460000  57.500000 ;
      RECT 56.990000  57.485000 58.460000  57.500000 ;
      RECT 56.990000  57.500000 58.475000  57.570000 ;
      RECT 56.990000  57.500000 58.475000  57.570000 ;
      RECT 56.990000  57.500000 60.970000  59.800000 ;
      RECT 56.990000  57.570000 58.545000  57.640000 ;
      RECT 56.990000  57.570000 58.545000  57.640000 ;
      RECT 56.990000  57.640000 58.615000  57.710000 ;
      RECT 56.990000  57.640000 58.615000  57.710000 ;
      RECT 56.990000  57.710000 58.685000  57.780000 ;
      RECT 56.990000  57.710000 58.685000  57.780000 ;
      RECT 56.990000  57.780000 58.755000  57.850000 ;
      RECT 56.990000  57.780000 58.755000  57.850000 ;
      RECT 56.990000  57.850000 58.825000  57.920000 ;
      RECT 56.990000  57.850000 58.825000  57.920000 ;
      RECT 56.990000  57.920000 58.895000  57.990000 ;
      RECT 56.990000  57.920000 58.895000  57.990000 ;
      RECT 56.990000  57.990000 58.965000  58.060000 ;
      RECT 56.990000  57.990000 58.965000  58.060000 ;
      RECT 56.990000  58.060000 59.035000  58.130000 ;
      RECT 56.990000  58.060000 59.035000  58.130000 ;
      RECT 56.990000  58.130000 59.105000  58.200000 ;
      RECT 56.990000  58.130000 59.105000  58.200000 ;
      RECT 56.990000  58.200000 59.175000  58.270000 ;
      RECT 56.990000  58.200000 59.175000  58.270000 ;
      RECT 56.990000  58.270000 59.245000  58.340000 ;
      RECT 56.990000  58.270000 59.245000  58.340000 ;
      RECT 56.990000  58.340000 59.315000  58.410000 ;
      RECT 56.990000  58.340000 59.315000  58.410000 ;
      RECT 56.990000  58.410000 59.385000  58.480000 ;
      RECT 56.990000  58.410000 59.385000  58.480000 ;
      RECT 56.990000  58.480000 59.455000  58.550000 ;
      RECT 56.990000  58.480000 59.455000  58.550000 ;
      RECT 56.990000  58.550000 59.525000  58.620000 ;
      RECT 56.990000  58.550000 59.525000  58.620000 ;
      RECT 56.990000  58.620000 59.595000  58.690000 ;
      RECT 56.990000  58.620000 59.595000  58.690000 ;
      RECT 56.990000  58.690000 59.665000  58.760000 ;
      RECT 56.990000  58.690000 59.665000  58.760000 ;
      RECT 56.990000  58.760000 59.735000  58.830000 ;
      RECT 56.990000  58.760000 59.735000  58.830000 ;
      RECT 56.990000  58.830000 59.805000  58.900000 ;
      RECT 56.990000  58.830000 59.805000  58.900000 ;
      RECT 56.990000  58.900000 59.875000  58.970000 ;
      RECT 56.990000  58.900000 59.875000  58.970000 ;
      RECT 56.990000  58.970000 59.945000  59.040000 ;
      RECT 56.990000  58.970000 59.945000  59.040000 ;
      RECT 56.990000  59.040000 60.015000  59.110000 ;
      RECT 56.990000  59.040000 60.015000  59.110000 ;
      RECT 56.990000  59.110000 60.085000  59.180000 ;
      RECT 56.990000  59.110000 60.085000  59.180000 ;
      RECT 56.990000  59.180000 60.155000  59.250000 ;
      RECT 56.990000  59.180000 60.155000  59.250000 ;
      RECT 56.990000  59.250000 60.225000  59.320000 ;
      RECT 56.990000  59.250000 60.225000  59.320000 ;
      RECT 56.990000  59.320000 60.295000  59.390000 ;
      RECT 56.990000  59.320000 60.295000  59.390000 ;
      RECT 56.990000  59.390000 60.365000  59.460000 ;
      RECT 56.990000  59.390000 60.365000  59.460000 ;
      RECT 56.990000  59.460000 60.435000  59.530000 ;
      RECT 56.990000  59.460000 60.435000  59.530000 ;
      RECT 56.990000  59.530000 60.505000  59.600000 ;
      RECT 56.990000  59.530000 60.505000  59.600000 ;
      RECT 56.990000  59.600000 60.575000  59.670000 ;
      RECT 56.990000  59.600000 60.575000  59.670000 ;
      RECT 56.990000  59.670000 60.645000  59.740000 ;
      RECT 56.990000  59.670000 60.645000  59.740000 ;
      RECT 56.990000  59.740000 60.715000  59.810000 ;
      RECT 56.990000  59.740000 60.715000  59.810000 ;
      RECT 56.990000  59.800000 60.970000  66.760000 ;
      RECT 56.990000  59.810000 60.785000  59.855000 ;
      RECT 56.990000  59.810000 60.785000  59.855000 ;
      RECT 56.990000  59.855000 60.830000  66.735000 ;
      RECT 56.990000  66.735000 60.820000  66.745000 ;
      RECT 56.990000  66.735000 60.820000  66.745000 ;
      RECT 56.990000  66.745000 60.805000  66.760000 ;
      RECT 56.990000  66.745000 60.805000  66.760000 ;
      RECT 57.055000  35.975000 60.970000  39.725000 ;
      RECT 57.055000  39.725000 60.970000  42.520000 ;
      RECT 57.055000  39.920000 60.830000  39.990000 ;
      RECT 57.055000  39.920000 60.830000  39.990000 ;
      RECT 57.125000  39.850000 60.830000  39.920000 ;
      RECT 57.125000  39.850000 60.830000  39.920000 ;
      RECT 57.195000  35.835000 60.830000  39.780000 ;
      RECT 57.195000  39.780000 60.830000  39.850000 ;
      RECT 57.195000  39.780000 60.830000  39.850000 ;
      RECT 58.240000 172.500000 58.515000 172.570000 ;
      RECT 58.240000 172.500000 60.970000 174.760000 ;
      RECT 58.240000 172.570000 58.585000 172.640000 ;
      RECT 58.240000 172.640000 58.655000 172.710000 ;
      RECT 58.240000 172.710000 58.725000 172.780000 ;
      RECT 58.240000 172.780000 58.795000 172.850000 ;
      RECT 58.240000 172.850000 58.865000 172.920000 ;
      RECT 58.240000 172.920000 58.935000 172.990000 ;
      RECT 58.240000 172.990000 59.005000 173.060000 ;
      RECT 58.240000 173.060000 59.075000 173.130000 ;
      RECT 58.240000 173.130000 59.145000 173.200000 ;
      RECT 58.240000 173.200000 59.215000 173.270000 ;
      RECT 58.240000 173.270000 59.285000 173.340000 ;
      RECT 58.240000 173.340000 59.355000 173.410000 ;
      RECT 58.240000 173.410000 59.425000 173.480000 ;
      RECT 58.240000 173.480000 59.495000 173.550000 ;
      RECT 58.240000 173.550000 59.565000 173.620000 ;
      RECT 58.240000 173.620000 59.635000 173.690000 ;
      RECT 58.240000 173.690000 59.705000 173.760000 ;
      RECT 58.240000 173.760000 59.775000 173.830000 ;
      RECT 58.240000 173.830000 59.845000 173.900000 ;
      RECT 58.240000 173.900000 59.915000 173.970000 ;
      RECT 58.240000 173.970000 59.985000 174.040000 ;
      RECT 58.240000 174.040000 60.055000 174.110000 ;
      RECT 58.240000 174.110000 60.125000 174.180000 ;
      RECT 58.240000 174.180000 60.195000 174.250000 ;
      RECT 58.240000 174.250000 60.265000 174.320000 ;
      RECT 58.240000 174.320000 60.335000 174.390000 ;
      RECT 58.240000 174.390000 60.405000 174.460000 ;
      RECT 58.240000 174.460000 60.475000 174.530000 ;
      RECT 58.240000 174.530000 60.545000 174.600000 ;
      RECT 58.240000 174.600000 60.615000 174.670000 ;
      RECT 58.240000 174.670000 60.685000 174.740000 ;
      RECT 58.240000 174.740000 60.755000 174.810000 ;
      RECT 58.240000 174.760000 60.970000 181.760000 ;
      RECT 58.240000 174.810000 60.825000 174.815000 ;
      RECT 58.240000 174.815000 60.830000 181.760000 ;
      RECT 67.480000 190.280000 75.000000 195.355000 ;
      RECT 67.480000 190.295000 75.000000 200.000000 ;
      RECT 70.480000 193.295000 72.000000 197.000000 ;
      RECT 74.430000   0.000000 75.000000 190.155000 ;
      RECT 74.570000   0.000000 75.000000 190.295000 ;
    LAYER met3 ;
      RECT  0.000000   0.000000  0.195000  36.635000 ;
      RECT  0.000000  36.635000  0.670000  37.110000 ;
      RECT  0.000000  36.730000  0.150000  36.880000 ;
      RECT  0.000000  36.880000  0.300000  37.030000 ;
      RECT  0.000000  37.030000  0.450000  37.150000 ;
      RECT  0.000000  37.110000  0.670000  46.360000 ;
      RECT  0.000000  37.150000  0.570000  46.320000 ;
      RECT  0.000000  46.320000  0.420000  46.470000 ;
      RECT  0.000000  46.360000  0.195000  46.835000 ;
      RECT  0.000000  46.470000  0.270000  46.620000 ;
      RECT  0.000000  46.620000  0.120000  46.770000 ;
      RECT  0.000000  46.835000  0.195000 173.455000 ;
      RECT  0.000000 173.455000 13.650000 195.500000 ;
      RECT  0.000000 173.555000 13.650000 195.500000 ;
      RECT  0.000000 173.555000 13.650000 200.000000 ;
      RECT  0.000000 195.500000 75.000000 200.000000 ;
      RECT  0.000000 195.500000 75.000000 200.000000 ;
      RECT 13.800000 101.520000 15.100000 102.035000 ;
      RECT 13.800000 102.035000 15.100000 171.140000 ;
      RECT 13.900000 101.560000 15.425000 101.710000 ;
      RECT 13.900000 101.710000 15.275000 101.860000 ;
      RECT 13.900000 101.860000 15.125000 102.010000 ;
      RECT 13.900000 102.010000 15.100000 102.035000 ;
      RECT 13.900000 102.035000 15.100000 171.140000 ;
      RECT 13.900000 171.140000 14.950000 171.290000 ;
      RECT 13.900000 171.290000 14.800000 171.440000 ;
      RECT 13.900000 171.440000 14.650000 171.590000 ;
      RECT 13.900000 171.590000 14.500000 171.740000 ;
      RECT 13.900000 171.740000 14.350000 171.890000 ;
      RECT 13.900000 171.890000 14.200000 172.040000 ;
      RECT 13.900000 172.040000 14.050000 172.190000 ;
      RECT 14.020000 101.440000 15.575000 101.560000 ;
      RECT 14.170000 101.290000 15.695000 101.440000 ;
      RECT 14.320000 101.140000 15.845000 101.290000 ;
      RECT 14.470000 100.990000 15.995000 101.140000 ;
      RECT 14.620000 100.840000 16.145000 100.990000 ;
      RECT 14.770000 100.690000 16.295000 100.840000 ;
      RECT 14.920000 100.540000 16.445000 100.690000 ;
      RECT 15.070000 100.390000 16.595000 100.540000 ;
      RECT 15.220000 100.240000 16.745000 100.390000 ;
      RECT 15.370000 100.090000 16.895000 100.240000 ;
      RECT 15.520000  99.940000 17.045000 100.090000 ;
      RECT 15.670000  99.790000 17.195000  99.940000 ;
      RECT 15.820000  99.640000 17.345000  99.790000 ;
      RECT 15.970000  99.490000 17.495000  99.640000 ;
      RECT 16.120000  99.340000 17.645000  99.490000 ;
      RECT 16.270000  99.190000 17.795000  99.340000 ;
      RECT 16.420000  99.040000 17.945000  99.190000 ;
      RECT 16.570000  98.890000 18.095000  99.040000 ;
      RECT 16.720000  98.740000 18.245000  98.890000 ;
      RECT 16.870000  98.590000 18.395000  98.740000 ;
      RECT 17.020000  98.440000 18.545000  98.590000 ;
      RECT 17.170000  98.290000 18.695000  98.440000 ;
      RECT 17.320000  98.140000 18.845000  98.290000 ;
      RECT 17.470000  97.990000 18.995000  98.140000 ;
      RECT 17.620000  97.840000 19.145000  97.990000 ;
      RECT 17.770000  97.690000 19.295000  97.840000 ;
      RECT 17.920000  97.540000 19.445000  97.690000 ;
      RECT 18.070000  97.390000 19.595000  97.540000 ;
      RECT 18.220000  97.240000 19.745000  97.390000 ;
      RECT 18.370000  97.090000 19.895000  97.240000 ;
      RECT 18.520000  96.940000 20.045000  97.090000 ;
      RECT 18.670000  96.790000 20.195000  96.940000 ;
      RECT 18.820000  96.640000 20.345000  96.790000 ;
      RECT 18.970000  96.490000 20.495000  96.640000 ;
      RECT 19.120000  96.340000 20.645000  96.490000 ;
      RECT 19.270000  96.190000 20.795000  96.340000 ;
      RECT 19.420000  96.040000 20.945000  96.190000 ;
      RECT 19.570000  95.890000 21.095000  96.040000 ;
      RECT 19.720000  95.740000 21.245000  95.890000 ;
      RECT 19.870000  95.590000 21.395000  95.740000 ;
      RECT 20.020000  95.440000 21.545000  95.590000 ;
      RECT 20.170000  95.290000 21.695000  95.440000 ;
      RECT 20.320000  95.140000 21.845000  95.290000 ;
      RECT 20.470000  94.990000 21.995000  95.140000 ;
      RECT 20.620000  94.840000 22.145000  94.990000 ;
      RECT 20.770000  94.690000 22.295000  94.840000 ;
      RECT 20.920000  94.540000 22.445000  94.690000 ;
      RECT 21.070000  94.390000 22.595000  94.540000 ;
      RECT 21.220000  94.240000 22.745000  94.390000 ;
      RECT 21.370000  94.090000 22.895000  94.240000 ;
      RECT 21.520000  93.940000 23.045000  94.090000 ;
      RECT 21.670000  93.790000 23.195000  93.940000 ;
      RECT 21.695000  93.765000 23.345000  93.790000 ;
      RECT 21.845000  93.615000 23.345000  93.765000 ;
      RECT 21.900000 104.845000 25.530000 168.965000 ;
      RECT 21.900000 104.845000 25.530000 168.965000 ;
      RECT 21.900000 168.965000 25.530000 172.475000 ;
      RECT 21.970000 104.775000 25.530000 104.845000 ;
      RECT 21.995000  93.465000 23.345000  93.615000 ;
      RECT 22.050000 168.965000 25.530000 169.115000 ;
      RECT 22.120000 104.625000 25.530000 104.775000 ;
      RECT 22.145000  93.315000 23.345000  93.465000 ;
      RECT 22.200000 169.115000 25.530000 169.265000 ;
      RECT 22.270000 104.475000 25.530000 104.625000 ;
      RECT 22.295000  93.165000 23.345000  93.315000 ;
      RECT 22.350000 169.265000 25.530000 169.415000 ;
      RECT 22.420000 104.325000 25.530000 104.475000 ;
      RECT 22.445000  93.015000 23.345000  93.165000 ;
      RECT 22.500000 169.415000 25.530000 169.565000 ;
      RECT 22.570000 104.175000 25.530000 104.325000 ;
      RECT 22.595000  92.865000 23.345000  93.015000 ;
      RECT 22.650000 169.565000 25.530000 169.715000 ;
      RECT 22.720000 104.025000 25.530000 104.175000 ;
      RECT 22.745000  92.715000 23.345000  92.865000 ;
      RECT 22.800000 169.715000 25.530000 169.865000 ;
      RECT 22.870000 103.875000 25.530000 104.025000 ;
      RECT 22.895000  92.565000 23.345000  92.715000 ;
      RECT 22.945000  92.375000 23.345000  93.790000 ;
      RECT 22.950000 169.865000 25.530000 170.015000 ;
      RECT 23.020000 103.725000 25.530000 103.875000 ;
      RECT 23.045000  92.415000 23.345000  92.565000 ;
      RECT 23.100000 170.015000 25.530000 170.165000 ;
      RECT 23.170000 103.575000 25.530000 103.725000 ;
      RECT 23.195000  92.265000 23.345000  92.415000 ;
      RECT 23.250000 170.165000 25.530000 170.315000 ;
      RECT 23.320000 103.425000 25.530000 103.575000 ;
      RECT 23.400000 170.315000 25.530000 170.465000 ;
      RECT 23.470000 103.275000 25.530000 103.425000 ;
      RECT 23.550000 170.465000 25.530000 170.615000 ;
      RECT 23.620000 103.125000 25.530000 103.275000 ;
      RECT 23.700000 170.615000 25.530000 170.765000 ;
      RECT 23.770000 102.975000 25.530000 103.125000 ;
      RECT 23.850000 170.765000 25.530000 170.915000 ;
      RECT 23.920000 102.825000 25.530000 102.975000 ;
      RECT 24.000000 170.915000 25.530000 171.065000 ;
      RECT 24.070000 102.675000 25.530000 102.825000 ;
      RECT 24.150000 171.065000 25.530000 171.215000 ;
      RECT 24.220000 102.525000 25.530000 102.675000 ;
      RECT 24.300000 171.215000 25.530000 171.365000 ;
      RECT 24.370000 102.375000 25.530000 102.525000 ;
      RECT 24.450000 171.365000 25.530000 171.515000 ;
      RECT 24.520000 102.225000 25.530000 102.375000 ;
      RECT 24.520000 102.225000 25.530000 104.845000 ;
      RECT 24.525000 102.220000 25.530000 102.225000 ;
      RECT 24.600000 171.515000 25.530000 171.665000 ;
      RECT 24.675000 102.070000 25.535000 102.220000 ;
      RECT 24.695000   0.000000 25.495000  90.225000 ;
      RECT 24.695000  90.225000 25.095000  90.625000 ;
      RECT 24.750000 171.665000 25.530000 171.815000 ;
      RECT 24.795000   0.000000 25.495000  90.225000 ;
      RECT 24.795000  90.225000 25.345000  90.375000 ;
      RECT 24.795000  90.375000 25.195000  90.525000 ;
      RECT 24.795000  90.525000 25.045000  90.675000 ;
      RECT 24.795000  90.675000 24.895000  90.825000 ;
      RECT 24.825000 101.920000 25.685000 102.070000 ;
      RECT 24.900000 171.815000 25.530000 171.965000 ;
      RECT 24.975000 101.770000 25.835000 101.920000 ;
      RECT 25.050000 171.965000 25.530000 172.115000 ;
      RECT 25.125000 101.620000 25.985000 101.770000 ;
      RECT 25.200000 172.115000 25.530000 172.265000 ;
      RECT 25.275000 101.470000 26.135000 101.620000 ;
      RECT 25.350000 172.265000 25.530000 172.415000 ;
      RECT 25.410000 172.475000 25.530000 195.500000 ;
      RECT 25.425000 101.320000 26.285000 101.470000 ;
      RECT 25.500000 172.415000 25.530000 172.565000 ;
      RECT 25.575000 101.170000 26.435000 101.320000 ;
      RECT 25.725000 101.020000 26.585000 101.170000 ;
      RECT 25.875000 100.870000 26.735000 101.020000 ;
      RECT 26.025000 100.720000 26.885000 100.870000 ;
      RECT 26.175000 100.570000 27.035000 100.720000 ;
      RECT 26.325000 100.420000 27.185000 100.570000 ;
      RECT 26.475000 100.270000 27.335000 100.420000 ;
      RECT 26.625000 100.120000 27.485000 100.270000 ;
      RECT 26.775000  99.970000 27.635000 100.120000 ;
      RECT 26.925000  99.820000 27.785000  99.970000 ;
      RECT 27.075000  99.670000 27.935000  99.820000 ;
      RECT 27.225000  99.520000 28.085000  99.670000 ;
      RECT 27.375000  99.370000 28.235000  99.520000 ;
      RECT 27.525000  99.220000 28.385000  99.370000 ;
      RECT 27.675000  99.070000 28.535000  99.220000 ;
      RECT 27.825000  98.920000 28.685000  99.070000 ;
      RECT 27.975000  98.770000 28.835000  98.920000 ;
      RECT 28.125000  98.620000 28.985000  98.770000 ;
      RECT 28.275000  98.470000 29.135000  98.620000 ;
      RECT 28.425000  98.320000 29.285000  98.470000 ;
      RECT 28.575000  98.170000 29.435000  98.320000 ;
      RECT 28.725000  98.020000 29.585000  98.170000 ;
      RECT 28.875000  97.870000 29.735000  98.020000 ;
      RECT 29.025000  97.720000 29.885000  97.870000 ;
      RECT 29.175000  97.570000 30.035000  97.720000 ;
      RECT 29.325000  97.420000 30.185000  97.570000 ;
      RECT 29.475000  97.270000 30.335000  97.420000 ;
      RECT 29.625000  97.120000 30.485000  97.270000 ;
      RECT 29.775000  96.970000 30.635000  97.120000 ;
      RECT 29.925000  93.265000 31.545000  96.210000 ;
      RECT 29.925000  93.265000 31.545000  96.210000 ;
      RECT 29.925000  96.210000 30.935000  96.820000 ;
      RECT 29.925000  96.210000 31.395000  96.360000 ;
      RECT 29.925000  96.360000 31.245000  96.510000 ;
      RECT 29.925000  96.510000 31.095000  96.660000 ;
      RECT 29.925000  96.660000 30.945000  96.810000 ;
      RECT 29.925000  96.810000 30.935000  96.820000 ;
      RECT 29.925000  96.820000 30.785000  96.970000 ;
      RECT 29.950000  93.240000 31.520000  93.265000 ;
      RECT 30.100000  93.090000 31.370000  93.240000 ;
      RECT 30.250000  92.940000 31.220000  93.090000 ;
      RECT 30.400000  92.790000 31.070000  92.940000 ;
      RECT 30.400000  92.790000 31.545000  93.265000 ;
      RECT 32.330000  99.865000 37.490000 110.785000 ;
      RECT 32.330000 105.025000 37.490000 105.820000 ;
      RECT 32.330000 105.025000 37.490000 105.820000 ;
      RECT 32.330000 105.820000 37.490000 105.970000 ;
      RECT 32.330000 105.820000 37.490000 105.970000 ;
      RECT 32.330000 105.820000 42.455000 110.785000 ;
      RECT 32.330000 105.820000 42.455000 175.185000 ;
      RECT 32.330000 105.970000 37.640000 106.120000 ;
      RECT 32.330000 105.970000 37.640000 106.120000 ;
      RECT 32.330000 106.120000 37.790000 106.270000 ;
      RECT 32.330000 106.120000 37.790000 106.270000 ;
      RECT 32.330000 106.270000 37.940000 106.420000 ;
      RECT 32.330000 106.270000 37.940000 106.420000 ;
      RECT 32.330000 106.420000 38.090000 106.570000 ;
      RECT 32.330000 106.420000 38.090000 106.570000 ;
      RECT 32.330000 106.570000 38.240000 106.720000 ;
      RECT 32.330000 106.570000 38.240000 106.720000 ;
      RECT 32.330000 106.720000 38.390000 106.870000 ;
      RECT 32.330000 106.720000 38.390000 106.870000 ;
      RECT 32.330000 106.870000 38.540000 107.020000 ;
      RECT 32.330000 106.870000 38.540000 107.020000 ;
      RECT 32.330000 107.020000 38.690000 107.170000 ;
      RECT 32.330000 107.020000 38.690000 107.170000 ;
      RECT 32.330000 107.170000 38.840000 107.320000 ;
      RECT 32.330000 107.170000 38.840000 107.320000 ;
      RECT 32.330000 107.320000 38.990000 107.470000 ;
      RECT 32.330000 107.320000 38.990000 107.470000 ;
      RECT 32.330000 107.470000 39.140000 107.620000 ;
      RECT 32.330000 107.470000 39.140000 107.620000 ;
      RECT 32.330000 107.620000 39.290000 107.770000 ;
      RECT 32.330000 107.620000 39.290000 107.770000 ;
      RECT 32.330000 107.770000 39.440000 107.920000 ;
      RECT 32.330000 107.770000 39.440000 107.920000 ;
      RECT 32.330000 107.920000 39.590000 108.070000 ;
      RECT 32.330000 107.920000 39.590000 108.070000 ;
      RECT 32.330000 108.070000 39.740000 108.220000 ;
      RECT 32.330000 108.070000 39.740000 108.220000 ;
      RECT 32.330000 108.220000 39.890000 108.370000 ;
      RECT 32.330000 108.220000 39.890000 108.370000 ;
      RECT 32.330000 108.370000 40.040000 108.520000 ;
      RECT 32.330000 108.370000 40.040000 108.520000 ;
      RECT 32.330000 108.520000 40.190000 108.670000 ;
      RECT 32.330000 108.520000 40.190000 108.670000 ;
      RECT 32.330000 108.670000 40.340000 108.820000 ;
      RECT 32.330000 108.670000 40.340000 108.820000 ;
      RECT 32.330000 108.820000 40.490000 108.970000 ;
      RECT 32.330000 108.820000 40.490000 108.970000 ;
      RECT 32.330000 108.970000 40.640000 109.120000 ;
      RECT 32.330000 108.970000 40.640000 109.120000 ;
      RECT 32.330000 109.120000 40.790000 109.270000 ;
      RECT 32.330000 109.120000 40.790000 109.270000 ;
      RECT 32.330000 109.270000 40.940000 109.420000 ;
      RECT 32.330000 109.270000 40.940000 109.420000 ;
      RECT 32.330000 109.420000 41.090000 109.570000 ;
      RECT 32.330000 109.420000 41.090000 109.570000 ;
      RECT 32.330000 109.570000 41.240000 109.720000 ;
      RECT 32.330000 109.570000 41.240000 109.720000 ;
      RECT 32.330000 109.720000 41.390000 109.870000 ;
      RECT 32.330000 109.720000 41.390000 109.870000 ;
      RECT 32.330000 109.870000 41.540000 110.020000 ;
      RECT 32.330000 109.870000 41.540000 110.020000 ;
      RECT 32.330000 110.020000 41.690000 110.170000 ;
      RECT 32.330000 110.020000 41.690000 110.170000 ;
      RECT 32.330000 110.170000 41.840000 110.320000 ;
      RECT 32.330000 110.170000 41.840000 110.320000 ;
      RECT 32.330000 110.320000 41.990000 110.470000 ;
      RECT 32.330000 110.320000 41.990000 110.470000 ;
      RECT 32.330000 110.470000 42.140000 110.620000 ;
      RECT 32.330000 110.470000 42.140000 110.620000 ;
      RECT 32.330000 110.620000 42.290000 110.770000 ;
      RECT 32.330000 110.620000 42.290000 110.770000 ;
      RECT 32.330000 110.770000 42.440000 110.785000 ;
      RECT 32.330000 110.770000 42.440000 110.785000 ;
      RECT 32.330000 110.785000 42.455000 170.295000 ;
      RECT 32.330000 110.785000 42.455000 170.295000 ;
      RECT 32.330000 170.295000 37.565000 175.185000 ;
      RECT 32.390000 104.965000 37.490000 105.025000 ;
      RECT 32.390000 104.965000 37.490000 105.025000 ;
      RECT 32.480000 170.295000 42.305000 170.445000 ;
      RECT 32.480000 170.295000 42.305000 170.445000 ;
      RECT 32.540000 104.815000 37.490000 104.965000 ;
      RECT 32.540000 104.815000 37.490000 104.965000 ;
      RECT 32.630000 170.445000 42.155000 170.595000 ;
      RECT 32.630000 170.445000 42.155000 170.595000 ;
      RECT 32.690000 104.665000 37.490000 104.815000 ;
      RECT 32.690000 104.665000 37.490000 104.815000 ;
      RECT 32.780000 170.595000 42.005000 170.745000 ;
      RECT 32.780000 170.595000 42.005000 170.745000 ;
      RECT 32.840000 104.515000 37.490000 104.665000 ;
      RECT 32.840000 104.515000 37.490000 104.665000 ;
      RECT 32.930000 170.745000 41.855000 170.895000 ;
      RECT 32.930000 170.745000 41.855000 170.895000 ;
      RECT 32.990000 104.365000 37.490000 104.515000 ;
      RECT 32.990000 104.365000 37.490000 104.515000 ;
      RECT 33.080000 170.895000 41.705000 171.045000 ;
      RECT 33.080000 170.895000 41.705000 171.045000 ;
      RECT 33.140000 104.215000 37.490000 104.365000 ;
      RECT 33.140000 104.215000 37.490000 104.365000 ;
      RECT 33.230000 171.045000 41.555000 171.195000 ;
      RECT 33.230000 171.045000 41.555000 171.195000 ;
      RECT 33.290000 104.065000 37.490000 104.215000 ;
      RECT 33.290000 104.065000 37.490000 104.215000 ;
      RECT 33.380000 171.195000 41.405000 171.345000 ;
      RECT 33.380000 171.195000 41.405000 171.345000 ;
      RECT 33.440000 103.915000 37.490000 104.065000 ;
      RECT 33.440000 103.915000 37.490000 104.065000 ;
      RECT 33.530000 171.345000 41.255000 171.495000 ;
      RECT 33.530000 171.345000 41.255000 171.495000 ;
      RECT 33.590000 103.765000 37.490000 103.915000 ;
      RECT 33.590000 103.765000 37.490000 103.915000 ;
      RECT 33.680000 171.495000 41.105000 171.645000 ;
      RECT 33.680000 171.495000 41.105000 171.645000 ;
      RECT 33.740000 103.615000 37.490000 103.765000 ;
      RECT 33.740000 103.615000 37.490000 103.765000 ;
      RECT 33.830000 171.645000 40.955000 171.795000 ;
      RECT 33.830000 171.645000 40.955000 171.795000 ;
      RECT 33.890000 103.465000 37.490000 103.615000 ;
      RECT 33.890000 103.465000 37.490000 103.615000 ;
      RECT 33.980000 171.795000 40.805000 171.945000 ;
      RECT 33.980000 171.795000 40.805000 171.945000 ;
      RECT 34.040000 103.315000 37.490000 103.465000 ;
      RECT 34.040000 103.315000 37.490000 103.465000 ;
      RECT 34.130000 171.945000 40.655000 172.095000 ;
      RECT 34.130000 171.945000 40.655000 172.095000 ;
      RECT 34.190000 103.165000 37.490000 103.315000 ;
      RECT 34.190000 103.165000 37.490000 103.315000 ;
      RECT 34.280000 172.095000 40.505000 172.245000 ;
      RECT 34.280000 172.095000 40.505000 172.245000 ;
      RECT 34.340000 103.015000 37.490000 103.165000 ;
      RECT 34.340000 103.015000 37.490000 103.165000 ;
      RECT 34.430000 172.245000 40.355000 172.395000 ;
      RECT 34.430000 172.245000 40.355000 172.395000 ;
      RECT 34.490000 102.865000 37.490000 103.015000 ;
      RECT 34.490000 102.865000 37.490000 103.015000 ;
      RECT 34.580000 172.395000 40.205000 172.545000 ;
      RECT 34.580000 172.395000 40.205000 172.545000 ;
      RECT 34.640000 102.715000 37.490000 102.865000 ;
      RECT 34.640000 102.715000 37.490000 102.865000 ;
      RECT 34.730000 172.545000 40.055000 172.695000 ;
      RECT 34.730000 172.545000 40.055000 172.695000 ;
      RECT 34.790000 102.565000 37.490000 102.715000 ;
      RECT 34.790000 102.565000 37.490000 102.715000 ;
      RECT 34.880000 172.695000 39.905000 172.845000 ;
      RECT 34.880000 172.695000 39.905000 172.845000 ;
      RECT 34.940000 102.415000 37.490000 102.565000 ;
      RECT 34.940000 102.415000 37.490000 102.565000 ;
      RECT 35.030000 172.845000 39.755000 172.995000 ;
      RECT 35.030000 172.845000 39.755000 172.995000 ;
      RECT 35.090000 102.265000 37.490000 102.415000 ;
      RECT 35.090000 102.265000 37.490000 102.415000 ;
      RECT 35.180000 172.995000 39.605000 173.145000 ;
      RECT 35.180000 172.995000 39.605000 173.145000 ;
      RECT 35.240000 102.115000 37.490000 102.265000 ;
      RECT 35.240000 102.115000 37.490000 102.265000 ;
      RECT 35.330000 173.145000 39.455000 173.295000 ;
      RECT 35.330000 173.145000 39.455000 173.295000 ;
      RECT 35.390000 101.965000 37.490000 102.115000 ;
      RECT 35.390000 101.965000 37.490000 102.115000 ;
      RECT 35.480000 173.295000 39.305000 173.445000 ;
      RECT 35.480000 173.295000 39.305000 173.445000 ;
      RECT 35.540000 101.815000 37.490000 101.965000 ;
      RECT 35.540000 101.815000 37.490000 101.965000 ;
      RECT 35.630000 173.445000 39.155000 173.595000 ;
      RECT 35.630000 173.445000 39.155000 173.595000 ;
      RECT 35.690000 101.665000 37.490000 101.815000 ;
      RECT 35.690000 101.665000 37.490000 101.815000 ;
      RECT 35.780000 173.595000 39.005000 173.745000 ;
      RECT 35.780000 173.595000 39.005000 173.745000 ;
      RECT 35.840000 101.515000 37.490000 101.665000 ;
      RECT 35.840000 101.515000 37.490000 101.665000 ;
      RECT 35.930000 173.745000 38.855000 173.895000 ;
      RECT 35.930000 173.745000 38.855000 173.895000 ;
      RECT 35.990000 101.365000 37.490000 101.515000 ;
      RECT 35.990000 101.365000 37.490000 101.515000 ;
      RECT 36.080000 173.895000 38.705000 174.045000 ;
      RECT 36.080000 173.895000 38.705000 174.045000 ;
      RECT 36.140000 101.215000 37.490000 101.365000 ;
      RECT 36.140000 101.215000 37.490000 101.365000 ;
      RECT 36.230000 174.045000 38.555000 174.195000 ;
      RECT 36.230000 174.045000 38.555000 174.195000 ;
      RECT 36.290000 101.065000 37.490000 101.215000 ;
      RECT 36.290000 101.065000 37.490000 101.215000 ;
      RECT 36.380000 174.195000 38.405000 174.345000 ;
      RECT 36.380000 174.195000 38.405000 174.345000 ;
      RECT 36.440000 100.915000 37.490000 101.065000 ;
      RECT 36.440000 100.915000 37.490000 101.065000 ;
      RECT 36.530000 174.345000 38.255000 174.495000 ;
      RECT 36.530000 174.345000 38.255000 174.495000 ;
      RECT 36.590000 100.765000 37.490000 100.915000 ;
      RECT 36.590000 100.765000 37.490000 100.915000 ;
      RECT 36.680000 174.495000 38.105000 174.645000 ;
      RECT 36.680000 174.495000 38.105000 174.645000 ;
      RECT 36.740000 100.615000 37.490000 100.765000 ;
      RECT 36.740000 100.615000 37.490000 100.765000 ;
      RECT 36.830000 174.645000 37.955000 174.795000 ;
      RECT 36.830000 174.645000 37.955000 174.795000 ;
      RECT 36.890000 100.465000 37.490000 100.615000 ;
      RECT 36.890000 100.465000 37.490000 100.615000 ;
      RECT 36.980000 174.795000 37.805000 174.945000 ;
      RECT 36.980000 174.795000 37.805000 174.945000 ;
      RECT 37.040000 100.315000 37.490000 100.465000 ;
      RECT 37.040000 100.315000 37.490000 100.465000 ;
      RECT 37.130000 174.945000 37.655000 175.095000 ;
      RECT 37.130000 174.945000 37.655000 175.095000 ;
      RECT 37.190000 100.165000 37.490000 100.315000 ;
      RECT 37.190000 100.165000 37.490000 100.315000 ;
      RECT 37.220000 175.185000 37.565000 190.420000 ;
      RECT 37.220000 175.270000 37.305000 175.355000 ;
      RECT 37.220000 175.355000 37.565000 190.420000 ;
      RECT 37.220000 190.420000 49.375000 190.440000 ;
      RECT 37.220000 190.420000 49.375000 190.440000 ;
      RECT 37.220000 190.420000 49.375000 200.000000 ;
      RECT 37.220000 190.440000 75.000000 195.500000 ;
      RECT 37.220000 190.440000 75.000000 195.500000 ;
      RECT 37.220000 190.440000 75.000000 200.000000 ;
      RECT 37.280000 175.095000 37.505000 175.245000 ;
      RECT 37.280000 175.095000 37.505000 175.245000 ;
      RECT 37.295000   0.000000 37.490000 100.060000 ;
      RECT 37.295000 100.060000 37.490000 105.025000 ;
      RECT 37.340000 100.015000 37.490000 100.165000 ;
      RECT 37.340000 100.015000 37.490000 100.165000 ;
      RECT 37.390000 175.245000 37.395000 175.355000 ;
      RECT 37.390000 175.245000 37.395000 175.355000 ;
      RECT 37.480000 175.270000 37.565000 175.355000 ;
      RECT 43.240000 100.380000 44.860000 101.970000 ;
      RECT 43.240000 100.380000 44.860000 101.970000 ;
      RECT 43.240000 101.970000 44.860000 102.580000 ;
      RECT 43.265000 100.355000 44.835000 100.380000 ;
      RECT 43.390000 101.970000 44.860000 102.120000 ;
      RECT 43.415000 100.205000 44.685000 100.355000 ;
      RECT 43.540000 102.120000 44.860000 102.270000 ;
      RECT 43.565000 100.055000 44.535000 100.205000 ;
      RECT 43.690000 102.270000 44.860000 102.420000 ;
      RECT 43.715000  99.905000 44.385000 100.055000 ;
      RECT 43.715000  99.905000 44.860000 100.380000 ;
      RECT 43.840000 102.420000 44.860000 102.570000 ;
      RECT 43.850000 102.570000 44.860000 102.580000 ;
      RECT 43.850000 102.580000 50.265000 107.985000 ;
      RECT 44.000000 102.580000 44.860000 102.730000 ;
      RECT 44.150000 102.730000 45.010000 102.880000 ;
      RECT 44.300000 102.880000 45.160000 103.030000 ;
      RECT 44.450000 103.030000 45.310000 103.180000 ;
      RECT 44.600000 103.180000 45.460000 103.330000 ;
      RECT 44.750000 103.330000 45.610000 103.480000 ;
      RECT 44.900000 103.480000 45.760000 103.630000 ;
      RECT 45.050000 103.630000 45.910000 103.780000 ;
      RECT 45.200000 103.780000 46.060000 103.930000 ;
      RECT 45.350000 103.930000 46.210000 104.080000 ;
      RECT 45.500000 104.080000 46.360000 104.230000 ;
      RECT 45.650000 104.230000 46.510000 104.380000 ;
      RECT 45.800000 104.380000 46.660000 104.530000 ;
      RECT 45.950000 104.530000 46.810000 104.680000 ;
      RECT 46.100000 104.680000 46.960000 104.830000 ;
      RECT 46.250000 104.830000 47.110000 104.980000 ;
      RECT 46.400000 104.980000 47.260000 105.130000 ;
      RECT 46.550000 105.130000 47.410000 105.280000 ;
      RECT 46.700000 105.280000 47.560000 105.430000 ;
      RECT 46.850000 105.430000 47.710000 105.580000 ;
      RECT 47.000000 105.580000 47.860000 105.730000 ;
      RECT 47.150000 105.730000 48.010000 105.880000 ;
      RECT 47.300000 105.880000 48.160000 106.030000 ;
      RECT 47.450000 106.030000 48.310000 106.180000 ;
      RECT 47.600000 106.180000 48.460000 106.330000 ;
      RECT 47.750000 106.330000 48.610000 106.480000 ;
      RECT 47.900000 106.480000 48.760000 106.630000 ;
      RECT 48.050000 106.630000 48.910000 106.780000 ;
      RECT 48.200000 106.780000 49.060000 106.930000 ;
      RECT 48.350000 106.930000 49.210000 107.080000 ;
      RECT 48.500000 107.080000 49.360000 107.230000 ;
      RECT 48.650000 107.230000 49.510000 107.380000 ;
      RECT 48.800000 107.380000 49.660000 107.530000 ;
      RECT 48.950000 107.530000 49.810000 107.680000 ;
      RECT 49.100000 107.680000 49.960000 107.830000 ;
      RECT 49.250000 107.830000 50.110000 107.980000 ;
      RECT 49.255000 107.980000 50.260000 107.985000 ;
      RECT 49.255000 107.985000 50.265000 108.135000 ;
      RECT 49.255000 107.985000 52.885000 110.605000 ;
      RECT 49.255000 108.135000 50.415000 108.285000 ;
      RECT 49.255000 108.285000 50.565000 108.435000 ;
      RECT 49.255000 108.435000 50.715000 108.585000 ;
      RECT 49.255000 108.585000 50.865000 108.735000 ;
      RECT 49.255000 108.735000 51.015000 108.885000 ;
      RECT 49.255000 108.885000 51.165000 109.035000 ;
      RECT 49.255000 109.035000 51.315000 109.185000 ;
      RECT 49.255000 109.185000 51.465000 109.335000 ;
      RECT 49.255000 109.335000 51.615000 109.485000 ;
      RECT 49.255000 109.485000 51.765000 109.635000 ;
      RECT 49.255000 109.635000 51.915000 109.785000 ;
      RECT 49.255000 109.785000 52.065000 109.935000 ;
      RECT 49.255000 109.935000 52.215000 110.085000 ;
      RECT 49.255000 110.085000 52.365000 110.235000 ;
      RECT 49.255000 110.235000 52.515000 110.385000 ;
      RECT 49.255000 110.385000 52.665000 110.535000 ;
      RECT 49.255000 110.535000 52.815000 110.605000 ;
      RECT 49.255000 110.605000 52.885000 168.970000 ;
      RECT 49.255000 110.605000 52.885000 168.970000 ;
      RECT 49.255000 168.970000 49.375000 172.480000 ;
      RECT 49.255000 168.970000 52.735000 169.120000 ;
      RECT 49.255000 169.120000 52.585000 169.270000 ;
      RECT 49.255000 169.270000 52.435000 169.420000 ;
      RECT 49.255000 169.420000 52.285000 169.570000 ;
      RECT 49.255000 169.570000 52.135000 169.720000 ;
      RECT 49.255000 169.720000 51.985000 169.870000 ;
      RECT 49.255000 169.870000 51.835000 170.020000 ;
      RECT 49.255000 170.020000 51.685000 170.170000 ;
      RECT 49.255000 170.170000 51.535000 170.320000 ;
      RECT 49.255000 170.320000 51.385000 170.470000 ;
      RECT 49.255000 170.470000 51.235000 170.620000 ;
      RECT 49.255000 170.620000 51.085000 170.770000 ;
      RECT 49.255000 170.770000 50.935000 170.920000 ;
      RECT 49.255000 170.920000 50.785000 171.070000 ;
      RECT 49.255000 171.070000 50.635000 171.220000 ;
      RECT 49.255000 171.220000 50.485000 171.370000 ;
      RECT 49.255000 171.370000 50.335000 171.520000 ;
      RECT 49.255000 171.520000 50.185000 171.670000 ;
      RECT 49.255000 171.670000 50.035000 171.820000 ;
      RECT 49.255000 171.820000 49.885000 171.970000 ;
      RECT 49.255000 171.970000 49.735000 172.120000 ;
      RECT 49.255000 172.120000 49.585000 172.270000 ;
      RECT 49.255000 172.270000 49.435000 172.420000 ;
      RECT 49.255000 172.420000 49.285000 172.570000 ;
      RECT 49.255000 172.480000 49.375000 190.420000 ;
      RECT 49.290000   0.000000 49.990000  89.650000 ;
      RECT 49.290000   0.000000 50.090000  90.310000 ;
      RECT 49.290000  89.800000 49.440000  89.950000 ;
      RECT 49.290000  89.800000 49.440000  89.950000 ;
      RECT 49.290000  89.950000 49.590000  90.100000 ;
      RECT 49.290000  89.950000 49.590000  90.100000 ;
      RECT 49.290000  90.100000 49.740000  90.250000 ;
      RECT 49.290000  90.100000 49.740000  90.250000 ;
      RECT 49.290000  90.250000 49.890000  90.400000 ;
      RECT 49.290000  90.250000 49.890000  90.400000 ;
      RECT 49.290000  90.310000 55.765000  95.985000 ;
      RECT 49.290000  90.400000 50.040000  90.550000 ;
      RECT 49.290000  90.400000 50.040000  90.550000 ;
      RECT 49.290000  90.550000 50.190000  90.700000 ;
      RECT 49.290000  90.550000 50.190000  90.700000 ;
      RECT 49.290000  90.700000 50.340000  90.850000 ;
      RECT 49.290000  90.700000 50.340000  90.850000 ;
      RECT 49.290000  90.850000 50.490000  91.000000 ;
      RECT 49.290000  90.850000 50.490000  91.000000 ;
      RECT 49.290000  91.000000 50.640000  91.150000 ;
      RECT 49.290000  91.000000 50.640000  91.150000 ;
      RECT 49.290000  91.150000 50.790000  91.300000 ;
      RECT 49.290000  91.150000 50.790000  91.300000 ;
      RECT 49.290000  91.300000 50.940000  91.450000 ;
      RECT 49.290000  91.300000 50.940000  91.450000 ;
      RECT 49.290000  91.450000 51.090000  91.600000 ;
      RECT 49.290000  91.450000 51.090000  91.600000 ;
      RECT 49.290000  91.600000 51.240000  91.750000 ;
      RECT 49.290000  91.600000 51.240000  91.750000 ;
      RECT 49.290000  91.750000 51.390000  91.900000 ;
      RECT 49.290000  91.750000 51.390000  91.900000 ;
      RECT 49.290000  91.900000 51.540000  92.050000 ;
      RECT 49.290000  91.900000 51.540000  92.050000 ;
      RECT 49.290000  92.050000 51.690000  92.200000 ;
      RECT 49.290000  92.050000 51.690000  92.200000 ;
      RECT 49.290000  92.200000 51.840000  92.350000 ;
      RECT 49.290000  92.200000 51.840000  92.350000 ;
      RECT 49.290000  92.350000 51.990000  92.500000 ;
      RECT 49.290000  92.350000 51.990000  92.500000 ;
      RECT 49.290000  92.500000 52.140000  92.650000 ;
      RECT 49.290000  92.500000 52.140000  92.650000 ;
      RECT 49.290000  92.650000 52.290000  92.800000 ;
      RECT 49.290000  92.650000 52.290000  92.800000 ;
      RECT 49.290000  92.800000 52.440000  92.950000 ;
      RECT 49.290000  92.800000 52.440000  92.950000 ;
      RECT 49.290000  92.950000 52.590000  93.100000 ;
      RECT 49.290000  92.950000 52.590000  93.100000 ;
      RECT 49.290000  93.100000 52.740000  93.250000 ;
      RECT 49.290000  93.100000 52.740000  93.250000 ;
      RECT 49.290000  93.250000 52.890000  93.400000 ;
      RECT 49.290000  93.250000 52.890000  93.400000 ;
      RECT 49.290000  93.400000 53.040000  93.550000 ;
      RECT 49.290000  93.400000 53.040000  93.550000 ;
      RECT 49.290000  93.550000 53.190000  93.700000 ;
      RECT 49.290000  93.550000 53.190000  93.700000 ;
      RECT 49.290000  93.700000 53.340000  93.850000 ;
      RECT 49.290000  93.700000 53.340000  93.850000 ;
      RECT 49.290000  93.850000 53.490000  94.000000 ;
      RECT 49.290000  93.850000 53.490000  94.000000 ;
      RECT 49.290000  94.000000 53.640000  94.150000 ;
      RECT 49.290000  94.000000 53.640000  94.150000 ;
      RECT 49.290000  94.150000 53.790000  94.300000 ;
      RECT 49.290000  94.150000 53.790000  94.300000 ;
      RECT 49.290000  94.300000 53.940000  94.450000 ;
      RECT 49.290000  94.300000 53.940000  94.450000 ;
      RECT 49.290000  94.450000 54.090000  94.600000 ;
      RECT 49.290000  94.450000 54.090000  94.600000 ;
      RECT 49.290000  94.600000 54.240000  94.750000 ;
      RECT 49.290000  94.600000 54.240000  94.750000 ;
      RECT 49.290000  94.750000 54.390000  94.900000 ;
      RECT 49.290000  94.750000 54.390000  94.900000 ;
      RECT 49.290000  94.900000 54.540000  95.050000 ;
      RECT 49.290000  94.900000 54.540000  95.050000 ;
      RECT 49.290000  95.050000 54.690000  95.200000 ;
      RECT 49.290000  95.050000 54.690000  95.200000 ;
      RECT 49.290000  95.200000 54.840000  95.350000 ;
      RECT 49.290000  95.200000 54.840000  95.350000 ;
      RECT 49.290000  95.350000 54.990000  95.500000 ;
      RECT 49.290000  95.350000 54.990000  95.500000 ;
      RECT 49.290000  95.500000 55.140000  95.650000 ;
      RECT 49.290000  95.500000 55.140000  95.650000 ;
      RECT 49.290000  95.650000 55.290000  95.800000 ;
      RECT 49.290000  95.650000 55.290000  95.800000 ;
      RECT 49.290000  95.800000 55.440000  95.950000 ;
      RECT 49.290000  95.800000 55.440000  95.950000 ;
      RECT 49.290000  95.950000 55.590000  95.985000 ;
      RECT 49.290000  95.950000 55.590000  95.985000 ;
      RECT 49.290000  95.985000 57.915000  98.135000 ;
      RECT 49.440000  95.985000 55.625000  96.135000 ;
      RECT 49.440000  95.985000 55.625000  96.135000 ;
      RECT 49.590000  96.135000 55.775000  96.285000 ;
      RECT 49.590000  96.135000 55.775000  96.285000 ;
      RECT 49.740000  96.285000 55.925000  96.435000 ;
      RECT 49.740000  96.285000 55.925000  96.435000 ;
      RECT 49.890000  96.435000 56.075000  96.585000 ;
      RECT 49.890000  96.435000 56.075000  96.585000 ;
      RECT 50.040000  96.585000 56.225000  96.735000 ;
      RECT 50.040000  96.585000 56.225000  96.735000 ;
      RECT 50.190000  96.735000 56.375000  96.885000 ;
      RECT 50.190000  96.735000 56.375000  96.885000 ;
      RECT 50.340000  96.885000 56.525000  97.035000 ;
      RECT 50.340000  96.885000 56.525000  97.035000 ;
      RECT 50.490000  97.035000 56.675000  97.185000 ;
      RECT 50.490000  97.035000 56.675000  97.185000 ;
      RECT 50.640000  97.185000 56.825000  97.335000 ;
      RECT 50.640000  97.185000 56.825000  97.335000 ;
      RECT 50.790000  97.335000 56.975000  97.485000 ;
      RECT 50.790000  97.335000 56.975000  97.485000 ;
      RECT 50.940000  97.485000 57.125000  97.635000 ;
      RECT 50.940000  97.485000 57.125000  97.635000 ;
      RECT 51.090000  97.635000 57.275000  97.785000 ;
      RECT 51.090000  97.635000 57.275000  97.785000 ;
      RECT 51.240000  97.785000 57.425000  97.935000 ;
      RECT 51.240000  97.785000 57.425000  97.935000 ;
      RECT 51.390000  97.935000 57.575000  98.085000 ;
      RECT 51.390000  97.935000 57.575000  98.085000 ;
      RECT 51.440000  98.085000 57.725000  98.135000 ;
      RECT 51.440000  98.085000 57.725000  98.135000 ;
      RECT 51.440000  98.135000 57.775000  98.285000 ;
      RECT 51.440000  98.135000 57.775000  98.285000 ;
      RECT 51.440000  98.135000 59.330000  99.550000 ;
      RECT 51.440000  98.285000 57.925000  98.435000 ;
      RECT 51.440000  98.285000 57.925000  98.435000 ;
      RECT 51.440000  98.435000 58.075000  98.585000 ;
      RECT 51.440000  98.435000 58.075000  98.585000 ;
      RECT 51.440000  98.585000 58.225000  98.735000 ;
      RECT 51.440000  98.585000 58.225000  98.735000 ;
      RECT 51.440000  98.735000 58.375000  98.885000 ;
      RECT 51.440000  98.735000 58.375000  98.885000 ;
      RECT 51.440000  98.885000 58.525000  99.035000 ;
      RECT 51.440000  98.885000 58.525000  99.035000 ;
      RECT 51.440000  99.035000 58.675000  99.185000 ;
      RECT 51.440000  99.035000 58.675000  99.185000 ;
      RECT 51.440000  99.185000 58.825000  99.335000 ;
      RECT 51.440000  99.185000 58.825000  99.335000 ;
      RECT 51.440000  99.335000 58.975000  99.485000 ;
      RECT 51.440000  99.335000 58.975000  99.485000 ;
      RECT 51.440000  99.485000 59.125000  99.550000 ;
      RECT 51.440000  99.485000 59.125000  99.550000 ;
      RECT 51.440000  99.550000 61.200000 101.420000 ;
      RECT 51.590000  99.550000 59.190000  99.700000 ;
      RECT 51.590000  99.550000 59.190000  99.700000 ;
      RECT 51.740000  99.700000 59.340000  99.850000 ;
      RECT 51.740000  99.700000 59.340000  99.850000 ;
      RECT 51.890000  99.850000 59.490000 100.000000 ;
      RECT 51.890000  99.850000 59.490000 100.000000 ;
      RECT 52.040000 100.000000 59.640000 100.150000 ;
      RECT 52.040000 100.000000 59.640000 100.150000 ;
      RECT 52.190000 100.150000 59.790000 100.300000 ;
      RECT 52.190000 100.150000 59.790000 100.300000 ;
      RECT 52.340000 100.300000 59.940000 100.450000 ;
      RECT 52.340000 100.300000 59.940000 100.450000 ;
      RECT 52.490000 100.450000 60.090000 100.600000 ;
      RECT 52.490000 100.450000 60.090000 100.600000 ;
      RECT 52.640000 100.600000 60.240000 100.750000 ;
      RECT 52.640000 100.600000 60.240000 100.750000 ;
      RECT 52.790000 100.750000 60.390000 100.900000 ;
      RECT 52.790000 100.750000 60.390000 100.900000 ;
      RECT 52.940000 100.900000 60.540000 101.050000 ;
      RECT 52.940000 100.900000 60.540000 101.050000 ;
      RECT 53.090000 101.050000 60.690000 101.200000 ;
      RECT 53.090000 101.050000 60.690000 101.200000 ;
      RECT 53.240000 101.200000 60.840000 101.350000 ;
      RECT 53.240000 101.200000 60.840000 101.350000 ;
      RECT 53.310000 101.420000 61.200000 107.795000 ;
      RECT 53.350000 101.350000 60.990000 101.460000 ;
      RECT 53.350000 101.350000 60.990000 101.460000 ;
      RECT 53.500000 101.460000 61.100000 101.610000 ;
      RECT 53.500000 101.460000 61.100000 101.610000 ;
      RECT 53.650000 101.610000 61.100000 101.760000 ;
      RECT 53.650000 101.610000 61.100000 101.760000 ;
      RECT 53.800000 101.760000 61.100000 101.910000 ;
      RECT 53.800000 101.760000 61.100000 101.910000 ;
      RECT 53.950000 101.910000 61.100000 102.060000 ;
      RECT 53.950000 101.910000 61.100000 102.060000 ;
      RECT 54.100000 102.060000 61.100000 102.210000 ;
      RECT 54.100000 102.060000 61.100000 102.210000 ;
      RECT 54.250000 102.210000 61.100000 102.360000 ;
      RECT 54.250000 102.210000 61.100000 102.360000 ;
      RECT 54.400000 102.360000 61.100000 102.510000 ;
      RECT 54.400000 102.360000 61.100000 102.510000 ;
      RECT 54.550000 102.510000 61.100000 102.660000 ;
      RECT 54.550000 102.510000 61.100000 102.660000 ;
      RECT 54.700000 102.660000 61.100000 102.810000 ;
      RECT 54.700000 102.660000 61.100000 102.810000 ;
      RECT 54.850000 102.810000 61.100000 102.960000 ;
      RECT 54.850000 102.810000 61.100000 102.960000 ;
      RECT 55.000000 102.960000 61.100000 103.110000 ;
      RECT 55.000000 102.960000 61.100000 103.110000 ;
      RECT 55.150000 103.110000 61.100000 103.260000 ;
      RECT 55.150000 103.110000 61.100000 103.260000 ;
      RECT 55.300000 103.260000 61.100000 103.410000 ;
      RECT 55.300000 103.260000 61.100000 103.410000 ;
      RECT 55.450000 103.410000 61.100000 103.560000 ;
      RECT 55.450000 103.410000 61.100000 103.560000 ;
      RECT 55.600000 103.560000 61.100000 103.710000 ;
      RECT 55.600000 103.560000 61.100000 103.710000 ;
      RECT 55.750000 103.710000 61.100000 103.860000 ;
      RECT 55.750000 103.710000 61.100000 103.860000 ;
      RECT 55.900000 103.860000 61.100000 104.010000 ;
      RECT 55.900000 103.860000 61.100000 104.010000 ;
      RECT 56.050000 104.010000 61.100000 104.160000 ;
      RECT 56.050000 104.010000 61.100000 104.160000 ;
      RECT 56.200000 104.160000 61.100000 104.310000 ;
      RECT 56.200000 104.160000 61.100000 104.310000 ;
      RECT 56.350000 104.310000 61.100000 104.460000 ;
      RECT 56.350000 104.310000 61.100000 104.460000 ;
      RECT 56.500000 104.460000 61.100000 104.610000 ;
      RECT 56.500000 104.460000 61.100000 104.610000 ;
      RECT 56.650000 104.610000 61.100000 104.760000 ;
      RECT 56.650000 104.610000 61.100000 104.760000 ;
      RECT 56.800000 104.760000 61.100000 104.910000 ;
      RECT 56.800000 104.760000 61.100000 104.910000 ;
      RECT 56.950000 104.910000 61.100000 105.060000 ;
      RECT 56.950000 104.910000 61.100000 105.060000 ;
      RECT 57.100000 105.060000 61.100000 105.210000 ;
      RECT 57.100000 105.060000 61.100000 105.210000 ;
      RECT 57.250000 105.210000 61.100000 105.360000 ;
      RECT 57.250000 105.210000 61.100000 105.360000 ;
      RECT 57.400000 105.360000 61.100000 105.510000 ;
      RECT 57.400000 105.360000 61.100000 105.510000 ;
      RECT 57.550000 105.510000 61.100000 105.660000 ;
      RECT 57.550000 105.510000 61.100000 105.660000 ;
      RECT 57.700000 105.660000 61.100000 105.810000 ;
      RECT 57.700000 105.660000 61.100000 105.810000 ;
      RECT 57.850000 105.810000 61.100000 105.960000 ;
      RECT 57.850000 105.810000 61.100000 105.960000 ;
      RECT 58.000000 105.960000 61.100000 106.110000 ;
      RECT 58.000000 105.960000 61.100000 106.110000 ;
      RECT 58.150000 106.110000 61.100000 106.260000 ;
      RECT 58.150000 106.110000 61.100000 106.260000 ;
      RECT 58.300000 106.260000 61.100000 106.410000 ;
      RECT 58.300000 106.260000 61.100000 106.410000 ;
      RECT 58.450000 106.410000 61.100000 106.560000 ;
      RECT 58.450000 106.410000 61.100000 106.560000 ;
      RECT 58.600000 106.560000 61.100000 106.710000 ;
      RECT 58.600000 106.560000 61.100000 106.710000 ;
      RECT 58.750000 106.710000 61.100000 106.860000 ;
      RECT 58.750000 106.710000 61.100000 106.860000 ;
      RECT 58.900000 106.860000 61.100000 107.010000 ;
      RECT 58.900000 106.860000 61.100000 107.010000 ;
      RECT 59.050000 107.010000 61.100000 107.160000 ;
      RECT 59.050000 107.010000 61.100000 107.160000 ;
      RECT 59.200000 107.160000 61.100000 107.310000 ;
      RECT 59.200000 107.160000 61.100000 107.310000 ;
      RECT 59.350000 107.310000 61.100000 107.460000 ;
      RECT 59.350000 107.310000 61.100000 107.460000 ;
      RECT 59.500000 107.460000 61.100000 107.610000 ;
      RECT 59.500000 107.460000 61.100000 107.610000 ;
      RECT 59.650000 107.610000 61.100000 107.760000 ;
      RECT 59.650000 107.610000 61.100000 107.760000 ;
      RECT 59.685000 107.795000 61.200000 172.855000 ;
      RECT 59.685000 107.945000 59.835000 108.095000 ;
      RECT 59.685000 108.095000 59.985000 108.245000 ;
      RECT 59.685000 108.245000 60.135000 108.395000 ;
      RECT 59.685000 108.395000 60.285000 108.545000 ;
      RECT 59.685000 108.545000 60.435000 108.695000 ;
      RECT 59.685000 108.695000 60.585000 108.845000 ;
      RECT 59.685000 108.845000 60.735000 108.995000 ;
      RECT 59.685000 108.995000 60.885000 109.145000 ;
      RECT 59.685000 109.145000 61.035000 109.210000 ;
      RECT 59.685000 109.210000 61.100000 172.855000 ;
      RECT 59.685000 172.855000 61.200000 173.620000 ;
      RECT 59.800000 107.760000 61.100000 107.910000 ;
      RECT 59.800000 107.760000 61.100000 107.910000 ;
      RECT 59.835000 172.855000 61.100000 173.005000 ;
      RECT 59.950000 107.910000 61.100000 108.060000 ;
      RECT 59.950000 107.910000 61.100000 108.060000 ;
      RECT 59.985000 173.005000 61.100000 173.155000 ;
      RECT 60.100000 108.060000 61.100000 108.210000 ;
      RECT 60.100000 108.060000 61.100000 108.210000 ;
      RECT 60.135000 173.155000 61.100000 173.305000 ;
      RECT 60.250000 108.210000 61.100000 108.360000 ;
      RECT 60.250000 108.210000 61.100000 108.360000 ;
      RECT 60.285000 173.305000 61.100000 173.455000 ;
      RECT 60.400000 108.360000 61.100000 108.510000 ;
      RECT 60.400000 108.360000 61.100000 108.510000 ;
      RECT 60.435000 173.455000 61.100000 173.605000 ;
      RECT 60.450000 173.620000 75.000000 174.515000 ;
      RECT 60.550000 108.510000 61.100000 108.660000 ;
      RECT 60.550000 108.510000 61.100000 108.660000 ;
      RECT 60.550000 173.605000 61.100000 173.720000 ;
      RECT 60.700000 108.660000 61.100000 108.810000 ;
      RECT 60.700000 108.660000 61.100000 108.810000 ;
      RECT 60.700000 173.720000 75.000000 173.870000 ;
      RECT 60.850000 108.810000 61.100000 108.960000 ;
      RECT 60.850000 108.810000 61.100000 108.960000 ;
      RECT 60.850000 173.870000 75.000000 174.020000 ;
      RECT 61.000000 108.960000 61.100000 109.110000 ;
      RECT 61.000000 108.960000 61.100000 109.110000 ;
      RECT 61.000000 174.020000 75.000000 174.170000 ;
      RECT 61.150000 174.170000 75.000000 174.320000 ;
      RECT 61.300000 174.320000 75.000000 174.470000 ;
      RECT 61.345000 173.720000 75.000000 190.440000 ;
      RECT 61.345000 173.720000 75.000000 200.000000 ;
      RECT 61.345000 174.470000 75.000000 174.515000 ;
      RECT 61.345000 174.515000 75.000000 190.440000 ;
      RECT 74.590000   0.000000 75.000000 173.620000 ;
      RECT 74.690000   0.000000 75.000000 173.720000 ;
    LAYER met4 ;
      RECT  0.000000   0.000000  1.670000   1.635000 ;
      RECT  0.000000   0.000000 75.000000   1.635000 ;
      RECT  0.000000   7.885000  1.670000   8.485000 ;
      RECT  0.000000   7.885000 75.000000   8.485000 ;
      RECT  0.000000  13.935000  1.365000  14.535000 ;
      RECT  0.000000  13.935000 75.000000  14.535000 ;
      RECT  0.000000  18.785000  1.365000  19.385000 ;
      RECT  0.000000  18.785000 75.000000  19.385000 ;
      RECT  0.000000  24.835000  1.670000  25.435000 ;
      RECT  0.000000  24.835000 75.000000  25.435000 ;
      RECT  0.000000  30.885000  1.670000  31.485000 ;
      RECT  0.000000  30.885000 75.000000  31.485000 ;
      RECT  0.000000  35.735000  1.670000  36.335000 ;
      RECT  0.000000  35.735000 75.000000  36.335000 ;
      RECT  0.000000  40.585000  1.670000  41.185000 ;
      RECT  0.000000  40.585000 75.000000  41.185000 ;
      RECT  0.000000  46.635000  1.670000  47.335000 ;
      RECT  0.000000  46.635000 75.000000  47.435000 ;
      RECT  0.000000  57.035000 75.000000  57.835000 ;
      RECT  0.000000  57.135000  1.670000  57.835000 ;
      RECT  0.000000  63.085000  1.670000  63.685000 ;
      RECT  0.000000  63.085000 75.000000  63.685000 ;
      RECT  0.000000  68.935000  1.670000  69.635000 ;
      RECT  0.000000  68.935000 75.000000  69.635000 ;
      RECT  0.000000  95.400000 75.000000 175.385000 ;
      RECT  1.365000  13.935000 73.635000  19.385000 ;
      RECT  1.570000  47.435000 73.430000  57.035000 ;
      RECT  1.670000   0.000000 73.330000  13.935000 ;
      RECT  1.670000  19.385000 73.330000  95.400000 ;
      RECT  1.670000 175.385000 73.330000 200.000000 ;
      RECT 73.330000   0.000000 75.000000   1.635000 ;
      RECT 73.330000   7.885000 75.000000   8.485000 ;
      RECT 73.330000  24.835000 75.000000  25.435000 ;
      RECT 73.330000  30.885000 75.000000  31.485000 ;
      RECT 73.330000  35.735000 75.000000  36.335000 ;
      RECT 73.330000  40.585000 75.000000  41.185000 ;
      RECT 73.330000  46.635000 75.000000  47.335000 ;
      RECT 73.330000  57.135000 75.000000  57.835000 ;
      RECT 73.330000  63.085000 75.000000  63.685000 ;
      RECT 73.330000  68.935000 75.000000  69.635000 ;
      RECT 73.635000  13.935000 75.000000  14.535000 ;
      RECT 73.635000  18.785000 75.000000  19.385000 ;
    LAYER met5 ;
      RECT  0.000000   0.000000 75.000000   0.535000 ;
      RECT  0.000000  96.585000 75.000000 137.725000 ;
      RECT  0.000000 137.725000 35.045000 147.535000 ;
      RECT  0.000000 147.535000 75.000000 174.185000 ;
      RECT  2.565000  15.035000 72.435000  18.285000 ;
      RECT  2.870000   0.000000 72.130000  15.035000 ;
      RECT  2.870000  18.285000 72.130000  96.585000 ;
      RECT  2.870000 174.185000 72.130000 200.000000 ;
      RECT 39.570000 137.725000 75.000000 147.535000 ;
  END
END sky130_fd_io__top_ground_hvc_wpad
END LIBRARY
