VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram45_256x16
  FOREIGN fakeram45_256x16 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 77.710 BY 40.600 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.485 0.070 2.555 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.905 0.070 2.975 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.325 0.070 3.395 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.745 0.070 3.815 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.165 0.070 4.235 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.585 0.070 4.655 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.005 0.070 5.075 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.425 0.070 5.495 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.845 0.070 5.915 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.265 0.070 6.335 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.685 0.070 6.755 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.105 0.070 7.175 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.525 0.070 7.595 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.945 0.070 8.015 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END w_mask_in[15]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.095 0.070 11.165 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.515 0.070 11.585 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.935 0.070 12.005 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.355 0.070 12.425 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.775 0.070 12.845 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.195 0.070 13.265 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.615 0.070 13.685 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.035 0.070 14.105 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.455 0.070 14.525 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.875 0.070 14.945 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.295 0.070 15.365 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.715 0.070 15.785 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.135 0.070 16.205 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.555 0.070 16.625 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.975 0.070 17.045 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.395 0.070 17.465 ;
    END
  END rd_out[15]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.125 0.070 20.195 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.545 0.070 20.615 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.385 0.070 21.455 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.805 0.070 21.875 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.225 0.070 22.295 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.645 0.070 22.715 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.065 0.070 23.135 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.485 0.070 23.555 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.905 0.070 23.975 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.325 0.070 24.395 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.745 0.070 24.815 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.165 0.070 25.235 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.585 0.070 25.655 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.005 0.070 26.075 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.425 0.070 26.495 ;
    END
  END wd_in[15]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.155 0.070 29.225 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.575 0.070 29.645 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.995 0.070 30.065 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.415 0.070 30.485 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.835 0.070 30.905 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.255 0.070 31.325 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.675 0.070 31.745 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.095 0.070 32.165 ;
    END
  END addr_in[7]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.825 0.070 34.895 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.245 0.070 35.315 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.665 0.070 35.735 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.960 2.100 2.240 38.500 ;
      RECT 5.320 2.100 5.600 38.500 ;
      RECT 8.680 2.100 8.960 38.500 ;
      RECT 12.040 2.100 12.320 38.500 ;
      RECT 15.400 2.100 15.680 38.500 ;
      RECT 18.760 2.100 19.040 38.500 ;
      RECT 22.120 2.100 22.400 38.500 ;
      RECT 25.480 2.100 25.760 38.500 ;
      RECT 28.840 2.100 29.120 38.500 ;
      RECT 32.200 2.100 32.480 38.500 ;
      RECT 35.560 2.100 35.840 38.500 ;
      RECT 38.920 2.100 39.200 38.500 ;
      RECT 42.280 2.100 42.560 38.500 ;
      RECT 45.640 2.100 45.920 38.500 ;
      RECT 49.000 2.100 49.280 38.500 ;
      RECT 52.360 2.100 52.640 38.500 ;
      RECT 55.720 2.100 56.000 38.500 ;
      RECT 59.080 2.100 59.360 38.500 ;
      RECT 62.440 2.100 62.720 38.500 ;
      RECT 65.800 2.100 66.080 38.500 ;
      RECT 69.160 2.100 69.440 38.500 ;
      RECT 72.520 2.100 72.800 38.500 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 3.640 2.100 3.920 38.500 ;
      RECT 7.000 2.100 7.280 38.500 ;
      RECT 10.360 2.100 10.640 38.500 ;
      RECT 13.720 2.100 14.000 38.500 ;
      RECT 17.080 2.100 17.360 38.500 ;
      RECT 20.440 2.100 20.720 38.500 ;
      RECT 23.800 2.100 24.080 38.500 ;
      RECT 27.160 2.100 27.440 38.500 ;
      RECT 30.520 2.100 30.800 38.500 ;
      RECT 33.880 2.100 34.160 38.500 ;
      RECT 37.240 2.100 37.520 38.500 ;
      RECT 40.600 2.100 40.880 38.500 ;
      RECT 43.960 2.100 44.240 38.500 ;
      RECT 47.320 2.100 47.600 38.500 ;
      RECT 50.680 2.100 50.960 38.500 ;
      RECT 54.040 2.100 54.320 38.500 ;
      RECT 57.400 2.100 57.680 38.500 ;
      RECT 60.760 2.100 61.040 38.500 ;
      RECT 64.120 2.100 64.400 38.500 ;
      RECT 67.480 2.100 67.760 38.500 ;
      RECT 70.840 2.100 71.120 38.500 ;
      RECT 74.200 2.100 74.480 38.500 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 77.710 40.600 ;
    LAYER metal2 ;
    RECT 0 0 77.710 40.600 ;
    LAYER metal3 ;
    RECT 0.070 0 77.710 40.600 ;
    RECT 0 0.000 0.070 2.065 ;
    RECT 0 2.135 0.070 2.485 ;
    RECT 0 2.555 0.070 2.905 ;
    RECT 0 2.975 0.070 3.325 ;
    RECT 0 3.395 0.070 3.745 ;
    RECT 0 3.815 0.070 4.165 ;
    RECT 0 4.235 0.070 4.585 ;
    RECT 0 4.655 0.070 5.005 ;
    RECT 0 5.075 0.070 5.425 ;
    RECT 0 5.495 0.070 5.845 ;
    RECT 0 5.915 0.070 6.265 ;
    RECT 0 6.335 0.070 6.685 ;
    RECT 0 6.755 0.070 7.105 ;
    RECT 0 7.175 0.070 7.525 ;
    RECT 0 7.595 0.070 7.945 ;
    RECT 0 8.015 0.070 8.365 ;
    RECT 0 8.435 0.070 11.095 ;
    RECT 0 11.165 0.070 11.515 ;
    RECT 0 11.585 0.070 11.935 ;
    RECT 0 12.005 0.070 12.355 ;
    RECT 0 12.425 0.070 12.775 ;
    RECT 0 12.845 0.070 13.195 ;
    RECT 0 13.265 0.070 13.615 ;
    RECT 0 13.685 0.070 14.035 ;
    RECT 0 14.105 0.070 14.455 ;
    RECT 0 14.525 0.070 14.875 ;
    RECT 0 14.945 0.070 15.295 ;
    RECT 0 15.365 0.070 15.715 ;
    RECT 0 15.785 0.070 16.135 ;
    RECT 0 16.205 0.070 16.555 ;
    RECT 0 16.625 0.070 16.975 ;
    RECT 0 17.045 0.070 17.395 ;
    RECT 0 17.465 0.070 20.125 ;
    RECT 0 20.195 0.070 20.545 ;
    RECT 0 20.615 0.070 20.965 ;
    RECT 0 21.035 0.070 21.385 ;
    RECT 0 21.455 0.070 21.805 ;
    RECT 0 21.875 0.070 22.225 ;
    RECT 0 22.295 0.070 22.645 ;
    RECT 0 22.715 0.070 23.065 ;
    RECT 0 23.135 0.070 23.485 ;
    RECT 0 23.555 0.070 23.905 ;
    RECT 0 23.975 0.070 24.325 ;
    RECT 0 24.395 0.070 24.745 ;
    RECT 0 24.815 0.070 25.165 ;
    RECT 0 25.235 0.070 25.585 ;
    RECT 0 25.655 0.070 26.005 ;
    RECT 0 26.075 0.070 26.425 ;
    RECT 0 26.495 0.070 29.155 ;
    RECT 0 29.225 0.070 29.575 ;
    RECT 0 29.645 0.070 29.995 ;
    RECT 0 30.065 0.070 30.415 ;
    RECT 0 30.485 0.070 30.835 ;
    RECT 0 30.905 0.070 31.255 ;
    RECT 0 31.325 0.070 31.675 ;
    RECT 0 31.745 0.070 32.095 ;
    RECT 0 32.165 0.070 34.825 ;
    RECT 0 34.895 0.070 35.245 ;
    RECT 0 35.315 0.070 35.665 ;
    RECT 0 35.735 0.070 40.600 ;
    LAYER metal4 ;
    RECT 0 0 77.710 2.100 ;
    RECT 0 38.500 77.710 40.600 ;
    RECT 0.000 2.100 1.960 38.500 ;
    RECT 2.240 2.100 3.640 38.500 ;
    RECT 3.920 2.100 5.320 38.500 ;
    RECT 5.600 2.100 7.000 38.500 ;
    RECT 7.280 2.100 8.680 38.500 ;
    RECT 8.960 2.100 10.360 38.500 ;
    RECT 10.640 2.100 12.040 38.500 ;
    RECT 12.320 2.100 13.720 38.500 ;
    RECT 14.000 2.100 15.400 38.500 ;
    RECT 15.680 2.100 17.080 38.500 ;
    RECT 17.360 2.100 18.760 38.500 ;
    RECT 19.040 2.100 20.440 38.500 ;
    RECT 20.720 2.100 22.120 38.500 ;
    RECT 22.400 2.100 23.800 38.500 ;
    RECT 24.080 2.100 25.480 38.500 ;
    RECT 25.760 2.100 27.160 38.500 ;
    RECT 27.440 2.100 28.840 38.500 ;
    RECT 29.120 2.100 30.520 38.500 ;
    RECT 30.800 2.100 32.200 38.500 ;
    RECT 32.480 2.100 33.880 38.500 ;
    RECT 34.160 2.100 35.560 38.500 ;
    RECT 35.840 2.100 37.240 38.500 ;
    RECT 37.520 2.100 38.920 38.500 ;
    RECT 39.200 2.100 40.600 38.500 ;
    RECT 40.880 2.100 42.280 38.500 ;
    RECT 42.560 2.100 43.960 38.500 ;
    RECT 44.240 2.100 45.640 38.500 ;
    RECT 45.920 2.100 47.320 38.500 ;
    RECT 47.600 2.100 49.000 38.500 ;
    RECT 49.280 2.100 50.680 38.500 ;
    RECT 50.960 2.100 52.360 38.500 ;
    RECT 52.640 2.100 54.040 38.500 ;
    RECT 54.320 2.100 55.720 38.500 ;
    RECT 56.000 2.100 57.400 38.500 ;
    RECT 57.680 2.100 59.080 38.500 ;
    RECT 59.360 2.100 60.760 38.500 ;
    RECT 61.040 2.100 62.440 38.500 ;
    RECT 62.720 2.100 64.120 38.500 ;
    RECT 64.400 2.100 65.800 38.500 ;
    RECT 66.080 2.100 67.480 38.500 ;
    RECT 67.760 2.100 69.160 38.500 ;
    RECT 69.440 2.100 70.840 38.500 ;
    RECT 71.120 2.100 72.520 38.500 ;
    RECT 72.800 2.100 74.200 38.500 ;
    RECT 74.480 2.100 77.710 38.500 ;
    LAYER OVERLAP ;
    RECT 0 0 77.710 40.600 ;
  END
END fakeram45_256x16

END LIBRARY
