VERSION 5.7 ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO vref_gen_nmos_with_trim
  CLASS CORE ;
#  CLASS BLOCK ;
  FOREIGN vref_gen_nmos_with_trim ;
  ORIGIN 0.000 0.000 ;
  SIZE 101.280 BY 61.050 ;
  PIN trim9
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 66.300 48.980 66.630 49.310 ;
      LAYER mcon ;
        RECT 66.380 49.060 66.550 49.230 ;
      LAYER met1 ;
        RECT 66.320 49.275 66.610 49.290 ;
        RECT 66.300 49.015 66.620 49.275 ;
        RECT 66.320 49.000 66.610 49.015 ;
      LAYER via ;
        RECT 66.330 49.015 66.590 49.275 ;
      LAYER met2 ;
        RECT 66.395 49.275 66.535 51.560 ;
        RECT 66.300 49.015 66.620 49.275 ;
    END
  END trim9
  PIN trim10
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 73.810 48.980 74.140 49.310 ;
      LAYER mcon ;
        RECT 73.890 49.060 74.060 49.230 ;
      LAYER met1 ;
        RECT 73.830 49.275 74.120 49.290 ;
        RECT 73.810 49.015 74.130 49.275 ;
        RECT 73.830 49.000 74.120 49.015 ;
      LAYER via ;
        RECT 73.840 49.015 74.100 49.275 ;
      LAYER met2 ;
        RECT 73.905 49.275 74.045 51.560 ;
        RECT 73.810 49.015 74.130 49.275 ;
    END
  END trim10
  PIN trim8
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 58.625 48.980 58.955 49.310 ;
      LAYER mcon ;
        RECT 58.705 49.060 58.875 49.230 ;
      LAYER met1 ;
        RECT 58.645 49.275 58.935 49.290 ;
        RECT 58.625 49.015 58.945 49.275 ;
        RECT 58.645 49.000 58.935 49.015 ;
      LAYER via ;
        RECT 58.655 49.015 58.915 49.275 ;
      LAYER met2 ;
        RECT 58.720 49.275 58.860 51.560 ;
        RECT 58.625 49.015 58.945 49.275 ;
    END
  END trim8
  PIN trim7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 51.115 48.980 51.445 49.310 ;
      LAYER mcon ;
        RECT 51.195 49.060 51.365 49.230 ;
      LAYER met1 ;
        RECT 51.135 49.275 51.425 49.290 ;
        RECT 51.115 49.015 51.435 49.275 ;
        RECT 51.135 49.000 51.425 49.015 ;
      LAYER via ;
        RECT 51.145 49.015 51.405 49.275 ;
      LAYER met2 ;
        RECT 51.210 49.275 51.350 51.560 ;
        RECT 51.115 49.015 51.435 49.275 ;
    END
  END trim7
  PIN trim6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 43.305 48.980 43.635 49.310 ;
      LAYER mcon ;
        RECT 43.385 49.060 43.555 49.230 ;
      LAYER met1 ;
        RECT 43.325 49.275 43.615 49.290 ;
        RECT 43.305 49.015 43.625 49.275 ;
        RECT 43.325 49.000 43.615 49.015 ;
      LAYER via ;
        RECT 43.335 49.015 43.595 49.275 ;
      LAYER met2 ;
        RECT 43.400 49.275 43.540 51.560 ;
        RECT 43.305 49.015 43.625 49.275 ;
    END
  END trim6
  PIN trim5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 35.750 48.980 36.080 49.310 ;
      LAYER mcon ;
        RECT 35.830 49.060 36.000 49.230 ;
      LAYER met1 ;
        RECT 35.770 49.275 36.060 49.290 ;
        RECT 35.750 49.015 36.070 49.275 ;
        RECT 35.770 49.000 36.060 49.015 ;
      LAYER via ;
        RECT 35.780 49.015 36.040 49.275 ;
      LAYER met2 ;
        RECT 35.845 49.275 35.985 51.560 ;
        RECT 35.750 49.015 36.070 49.275 ;
    END
  END trim5
  PIN trim4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 28.015 48.980 28.345 49.310 ;
      LAYER mcon ;
        RECT 28.095 49.060 28.265 49.230 ;
      LAYER met1 ;
        RECT 28.035 49.275 28.325 49.290 ;
        RECT 28.015 49.015 28.335 49.275 ;
        RECT 28.035 49.000 28.325 49.015 ;
      LAYER via ;
        RECT 28.045 49.015 28.305 49.275 ;
      LAYER met2 ;
        RECT 28.110 49.275 28.250 51.560 ;
        RECT 28.015 49.015 28.335 49.275 ;
    END
  END trim4
  PIN trim3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 21.025 48.980 21.355 49.310 ;
      LAYER mcon ;
        RECT 21.105 49.060 21.275 49.230 ;
      LAYER met1 ;
        RECT 21.045 49.275 21.335 49.290 ;
        RECT 21.025 49.015 21.345 49.275 ;
        RECT 21.045 49.000 21.335 49.015 ;
      LAYER via ;
        RECT 21.055 49.015 21.315 49.275 ;
      LAYER met2 ;
        RECT 21.115 49.275 21.255 51.560 ;
        RECT 21.025 49.015 21.345 49.275 ;
    END
  END trim3
  PIN trim2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.500 48.980 15.830 49.310 ;
      LAYER mcon ;
        RECT 15.580 49.060 15.750 49.230 ;
      LAYER met1 ;
        RECT 15.520 49.275 15.810 49.290 ;
        RECT 15.500 49.015 15.820 49.275 ;
        RECT 15.520 49.000 15.810 49.015 ;
      LAYER via ;
        RECT 15.530 49.015 15.790 49.275 ;
      LAYER met2 ;
        RECT 15.595 49.275 15.735 51.560 ;
        RECT 15.500 49.015 15.820 49.275 ;
    END
  END trim2
  PIN trim1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.895 48.980 11.225 49.310 ;
      LAYER mcon ;
        RECT 10.975 49.060 11.145 49.230 ;
      LAYER met1 ;
        RECT 10.915 49.275 11.205 49.290 ;
        RECT 10.895 49.015 11.215 49.275 ;
        RECT 10.915 49.000 11.205 49.015 ;
      LAYER via ;
        RECT 10.925 49.015 11.185 49.275 ;
      LAYER met2 ;
        RECT 10.980 49.275 11.120 51.560 ;
        RECT 10.895 49.015 11.215 49.275 ;
    END
  END trim1
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 7.700 50.465 87.545 50.795 ;
        RECT 7.490 49.430 10.200 49.600 ;
        RECT 11.975 49.430 14.685 49.600 ;
        RECT 17.435 49.430 20.145 49.600 ;
        RECT 24.460 49.430 27.170 49.600 ;
        RECT 32.195 49.430 34.905 49.600 ;
        RECT 39.750 49.430 42.460 49.600 ;
        RECT 47.560 49.430 50.270 49.600 ;
        RECT 55.070 49.430 57.780 49.600 ;
        RECT 62.745 49.430 65.455 49.600 ;
        RECT 70.255 49.430 72.965 49.600 ;
        RECT 76.635 47.745 80.295 47.915 ;
        RECT 76.635 42.860 76.805 47.745 ;
        RECT 80.125 42.860 80.295 47.745 ;
        RECT 76.635 42.690 80.295 42.860 ;
        RECT 76.635 37.805 76.805 42.690 ;
        RECT 80.125 37.805 80.295 42.690 ;
        RECT 76.635 37.635 80.295 37.805 ;
        RECT 76.635 32.750 76.805 37.635 ;
        RECT 80.125 32.750 80.295 37.635 ;
        RECT 76.635 32.580 80.295 32.750 ;
        RECT 76.635 27.695 76.805 32.580 ;
        RECT 80.125 27.695 80.295 32.580 ;
        RECT 76.635 27.525 80.295 27.695 ;
        RECT 76.635 22.640 76.805 27.525 ;
        RECT 80.125 22.640 80.295 27.525 ;
        RECT 76.635 22.470 80.295 22.640 ;
        RECT 76.635 17.585 76.805 22.470 ;
        RECT 80.125 17.585 80.295 22.470 ;
        RECT 76.635 17.415 80.295 17.585 ;
        RECT 76.635 12.505 76.805 17.415 ;
        RECT 80.125 12.505 80.295 17.415 ;
        RECT 76.635 12.335 80.295 12.505 ;
        RECT 82.185 47.745 85.845 47.915 ;
        RECT 82.185 42.860 82.355 47.745 ;
        RECT 85.675 42.860 85.845 47.745 ;
        RECT 82.185 42.690 85.845 42.860 ;
        RECT 82.185 37.805 82.355 42.690 ;
        RECT 85.675 37.805 85.845 42.690 ;
        RECT 82.185 37.635 85.845 37.805 ;
        RECT 82.185 32.750 82.355 37.635 ;
        RECT 85.675 32.750 85.845 37.635 ;
        RECT 82.185 32.580 85.845 32.750 ;
        RECT 82.185 27.695 82.355 32.580 ;
        RECT 85.675 27.695 85.845 32.580 ;
        RECT 82.185 27.525 85.845 27.695 ;
        RECT 82.185 22.640 82.355 27.525 ;
        RECT 85.675 22.640 85.845 27.525 ;
        RECT 82.185 22.470 91.515 22.640 ;
        RECT 82.185 17.585 82.355 22.470 ;
        RECT 85.675 17.585 85.845 22.470 ;
        RECT 82.185 17.415 85.845 17.585 ;
        RECT 82.185 12.505 82.355 17.415 ;
        RECT 85.675 12.505 85.845 17.415 ;
        RECT 82.185 12.335 85.845 12.505 ;
        RECT 87.855 17.585 88.025 22.470 ;
        RECT 91.345 17.585 91.515 22.470 ;
        RECT 87.855 17.415 91.515 17.585 ;
        RECT 87.855 12.505 88.025 17.415 ;
        RECT 91.345 12.505 91.515 17.415 ;
        RECT 87.855 12.335 91.515 12.505 ;
      LAYER mcon ;
        RECT 8.090 50.550 8.260 50.720 ;
        RECT 8.450 50.550 8.620 50.720 ;
        RECT 8.810 50.550 8.980 50.720 ;
        RECT 9.170 50.550 9.340 50.720 ;
        RECT 12.580 50.550 12.750 50.720 ;
        RECT 12.940 50.550 13.110 50.720 ;
        RECT 13.300 50.550 13.470 50.720 ;
        RECT 13.660 50.550 13.830 50.720 ;
        RECT 18.040 50.550 18.210 50.720 ;
        RECT 18.400 50.550 18.570 50.720 ;
        RECT 18.760 50.550 18.930 50.720 ;
        RECT 19.120 50.550 19.290 50.720 ;
        RECT 25.065 50.550 25.235 50.720 ;
        RECT 25.425 50.550 25.595 50.720 ;
        RECT 25.785 50.550 25.955 50.720 ;
        RECT 26.145 50.550 26.315 50.720 ;
        RECT 32.800 50.550 32.970 50.720 ;
        RECT 33.160 50.550 33.330 50.720 ;
        RECT 33.520 50.550 33.690 50.720 ;
        RECT 33.880 50.550 34.050 50.720 ;
        RECT 40.355 50.550 40.525 50.720 ;
        RECT 40.715 50.550 40.885 50.720 ;
        RECT 41.075 50.550 41.245 50.720 ;
        RECT 41.435 50.550 41.605 50.720 ;
        RECT 48.165 50.550 48.335 50.720 ;
        RECT 48.525 50.550 48.695 50.720 ;
        RECT 48.885 50.550 49.055 50.720 ;
        RECT 49.245 50.550 49.415 50.720 ;
        RECT 55.675 50.550 55.845 50.720 ;
        RECT 56.035 50.550 56.205 50.720 ;
        RECT 56.395 50.550 56.565 50.720 ;
        RECT 56.755 50.550 56.925 50.720 ;
        RECT 63.350 50.550 63.520 50.720 ;
        RECT 63.710 50.550 63.880 50.720 ;
        RECT 64.070 50.550 64.240 50.720 ;
        RECT 64.430 50.550 64.600 50.720 ;
        RECT 70.860 50.550 71.030 50.720 ;
        RECT 71.220 50.550 71.390 50.720 ;
        RECT 71.580 50.550 71.750 50.720 ;
        RECT 71.940 50.550 72.110 50.720 ;
        RECT 76.825 50.545 76.995 50.715 ;
        RECT 77.185 50.545 77.355 50.715 ;
        RECT 77.545 50.545 77.715 50.715 ;
        RECT 77.905 50.545 78.075 50.715 ;
        RECT 78.265 50.545 78.435 50.715 ;
        RECT 78.625 50.545 78.795 50.715 ;
        RECT 78.985 50.545 79.155 50.715 ;
        RECT 79.345 50.545 79.515 50.715 ;
        RECT 79.705 50.545 79.875 50.715 ;
        RECT 80.065 50.545 80.235 50.715 ;
        RECT 82.375 50.545 82.545 50.715 ;
        RECT 82.735 50.545 82.905 50.715 ;
        RECT 83.095 50.545 83.265 50.715 ;
        RECT 83.455 50.545 83.625 50.715 ;
        RECT 83.815 50.545 83.985 50.715 ;
        RECT 84.175 50.545 84.345 50.715 ;
        RECT 84.535 50.545 84.705 50.715 ;
        RECT 84.895 50.545 85.065 50.715 ;
        RECT 85.255 50.545 85.425 50.715 ;
        RECT 85.615 50.545 85.785 50.715 ;
        RECT 8.095 49.430 8.265 49.600 ;
        RECT 8.455 49.430 8.625 49.600 ;
        RECT 8.815 49.430 8.985 49.600 ;
        RECT 9.175 49.430 9.345 49.600 ;
        RECT 12.580 49.430 12.750 49.600 ;
        RECT 12.940 49.430 13.110 49.600 ;
        RECT 13.300 49.430 13.470 49.600 ;
        RECT 13.660 49.430 13.830 49.600 ;
        RECT 18.040 49.430 18.210 49.600 ;
        RECT 18.400 49.430 18.570 49.600 ;
        RECT 18.760 49.430 18.930 49.600 ;
        RECT 19.120 49.430 19.290 49.600 ;
        RECT 25.065 49.430 25.235 49.600 ;
        RECT 25.425 49.430 25.595 49.600 ;
        RECT 25.785 49.430 25.955 49.600 ;
        RECT 26.145 49.430 26.315 49.600 ;
        RECT 32.800 49.430 32.970 49.600 ;
        RECT 33.160 49.430 33.330 49.600 ;
        RECT 33.520 49.430 33.690 49.600 ;
        RECT 33.880 49.430 34.050 49.600 ;
        RECT 40.355 49.430 40.525 49.600 ;
        RECT 40.715 49.430 40.885 49.600 ;
        RECT 41.075 49.430 41.245 49.600 ;
        RECT 41.435 49.430 41.605 49.600 ;
        RECT 48.165 49.430 48.335 49.600 ;
        RECT 48.525 49.430 48.695 49.600 ;
        RECT 48.885 49.430 49.055 49.600 ;
        RECT 49.245 49.430 49.415 49.600 ;
        RECT 55.675 49.430 55.845 49.600 ;
        RECT 56.035 49.430 56.205 49.600 ;
        RECT 56.395 49.430 56.565 49.600 ;
        RECT 56.755 49.430 56.925 49.600 ;
        RECT 63.350 49.430 63.520 49.600 ;
        RECT 63.710 49.430 63.880 49.600 ;
        RECT 64.070 49.430 64.240 49.600 ;
        RECT 64.430 49.430 64.600 49.600 ;
        RECT 70.860 49.430 71.030 49.600 ;
        RECT 71.220 49.430 71.390 49.600 ;
        RECT 71.580 49.430 71.750 49.600 ;
        RECT 71.940 49.430 72.110 49.600 ;
        RECT 76.825 47.745 76.995 47.915 ;
        RECT 77.185 47.745 77.355 47.915 ;
        RECT 77.545 47.745 77.715 47.915 ;
        RECT 77.905 47.745 78.075 47.915 ;
        RECT 78.265 47.745 78.435 47.915 ;
        RECT 78.625 47.745 78.795 47.915 ;
        RECT 78.985 47.745 79.155 47.915 ;
        RECT 79.345 47.745 79.515 47.915 ;
        RECT 79.705 47.745 79.875 47.915 ;
        RECT 80.065 47.745 80.235 47.915 ;
        RECT 82.375 47.745 82.545 47.915 ;
        RECT 82.735 47.745 82.905 47.915 ;
        RECT 83.095 47.745 83.265 47.915 ;
        RECT 83.455 47.745 83.625 47.915 ;
        RECT 83.815 47.745 83.985 47.915 ;
        RECT 84.175 47.745 84.345 47.915 ;
        RECT 84.535 47.745 84.705 47.915 ;
        RECT 84.895 47.745 85.065 47.915 ;
        RECT 85.255 47.745 85.425 47.915 ;
        RECT 85.615 47.745 85.785 47.915 ;
        RECT 87.895 22.470 88.065 22.640 ;
        RECT 88.255 22.470 88.425 22.640 ;
        RECT 88.615 22.470 88.785 22.640 ;
        RECT 88.975 22.470 89.145 22.640 ;
        RECT 89.335 22.470 89.505 22.640 ;
        RECT 89.695 22.470 89.865 22.640 ;
        RECT 90.055 22.470 90.225 22.640 ;
        RECT 90.415 22.470 90.585 22.640 ;
        RECT 90.775 22.470 90.945 22.640 ;
        RECT 91.135 22.470 91.305 22.640 ;
      LAYER met1 ;
        RECT 0.000 53.165 8.370 53.535 ;
        RECT 7.180 52.655 8.370 53.165 ;
        RECT 83.565 53.165 101.280 53.535 ;
        RECT 83.565 52.655 85.935 53.165 ;
        RECT 0.000 52.285 101.280 52.655 ;
        RECT 7.180 50.295 88.230 52.285 ;
        RECT 8.030 48.965 9.400 50.295 ;
        RECT 12.520 48.965 13.890 50.295 ;
        RECT 17.980 48.965 19.350 50.295 ;
        RECT 25.005 48.965 26.375 50.295 ;
        RECT 32.740 48.965 34.110 50.295 ;
        RECT 40.295 48.965 41.665 50.295 ;
        RECT 48.105 48.965 49.475 50.295 ;
        RECT 55.615 48.965 56.985 50.295 ;
        RECT 63.290 48.965 64.660 50.295 ;
        RECT 70.800 48.965 72.170 50.295 ;
        RECT 76.765 47.715 80.295 50.295 ;
        RECT 82.315 47.715 85.845 50.295 ;
        RECT 87.975 22.670 91.175 22.700 ;
        RECT 87.835 22.440 91.365 22.670 ;
      LAYER via ;
        RECT 76.935 50.490 77.195 50.750 ;
        RECT 77.255 50.490 77.515 50.750 ;
        RECT 77.575 50.490 77.835 50.750 ;
        RECT 77.895 50.490 78.155 50.750 ;
        RECT 78.215 50.490 78.475 50.750 ;
        RECT 78.535 50.490 78.795 50.750 ;
        RECT 78.855 50.490 79.115 50.750 ;
        RECT 79.175 50.490 79.435 50.750 ;
        RECT 79.495 50.490 79.755 50.750 ;
        RECT 79.815 50.490 80.075 50.750 ;
        RECT 82.485 50.490 82.745 50.750 ;
        RECT 82.805 50.490 83.065 50.750 ;
        RECT 83.125 50.490 83.385 50.750 ;
        RECT 83.445 50.490 83.705 50.750 ;
        RECT 83.765 50.490 84.025 50.750 ;
        RECT 84.085 50.490 84.345 50.750 ;
        RECT 84.405 50.490 84.665 50.750 ;
        RECT 84.725 50.490 84.985 50.750 ;
        RECT 85.045 50.490 85.305 50.750 ;
        RECT 85.365 50.490 85.625 50.750 ;
        RECT 76.935 47.715 77.195 47.975 ;
        RECT 77.255 47.715 77.515 47.975 ;
        RECT 77.575 47.715 77.835 47.975 ;
        RECT 77.895 47.715 78.155 47.975 ;
        RECT 78.215 47.715 78.475 47.975 ;
        RECT 78.535 47.715 78.795 47.975 ;
        RECT 78.855 47.715 79.115 47.975 ;
        RECT 79.175 47.715 79.435 47.975 ;
        RECT 79.495 47.715 79.755 47.975 ;
        RECT 79.815 47.715 80.075 47.975 ;
        RECT 82.485 47.715 82.745 47.975 ;
        RECT 82.805 47.715 83.065 47.975 ;
        RECT 83.125 47.715 83.385 47.975 ;
        RECT 83.445 47.715 83.705 47.975 ;
        RECT 83.765 47.715 84.025 47.975 ;
        RECT 84.085 47.715 84.345 47.975 ;
        RECT 84.405 47.715 84.665 47.975 ;
        RECT 84.725 47.715 84.985 47.975 ;
        RECT 85.045 47.715 85.305 47.975 ;
        RECT 85.365 47.715 85.625 47.975 ;
        RECT 88.005 22.440 88.265 22.700 ;
        RECT 88.325 22.440 88.585 22.700 ;
        RECT 88.645 22.440 88.905 22.700 ;
        RECT 88.965 22.440 89.225 22.700 ;
        RECT 89.285 22.440 89.545 22.700 ;
        RECT 89.605 22.440 89.865 22.700 ;
        RECT 89.925 22.440 90.185 22.700 ;
        RECT 90.245 22.440 90.505 22.700 ;
        RECT 90.565 22.440 90.825 22.700 ;
        RECT 90.885 22.440 91.145 22.700 ;
      LAYER met2 ;
        RECT 76.580 12.280 80.330 51.015 ;
        RECT 82.130 12.280 85.880 51.015 ;
        RECT 87.800 12.280 91.550 23.395 ;
    END
  END vpwr
  PIN vref
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 10.105 47.070 11.315 47.580 ;
        RECT 13.475 47.410 15.795 47.580 ;
        RECT 17.600 47.410 21.255 47.580 ;
        RECT 13.475 47.240 15.800 47.410 ;
        RECT 17.600 47.240 21.260 47.410 ;
        RECT 13.485 47.070 15.795 47.240 ;
        RECT 17.600 47.070 21.255 47.240 ;
        RECT 23.185 47.070 29.425 47.580 ;
        RECT 30.920 47.070 37.160 47.580 ;
        RECT 38.475 47.070 44.715 47.580 ;
        RECT 46.285 47.070 52.525 47.580 ;
        RECT 53.795 47.070 60.035 47.580 ;
        RECT 61.470 47.070 67.710 47.580 ;
        RECT 68.980 47.070 75.220 47.580 ;
        RECT 77.515 45.385 77.845 45.465 ;
        RECT 77.515 45.215 78.990 45.385 ;
        RECT 77.515 45.135 77.845 45.215 ;
        RECT 9.825 44.710 11.310 44.880 ;
        RECT 12.560 44.710 15.795 44.880 ;
        RECT 17.600 44.710 21.255 44.880 ;
        RECT 23.185 44.710 28.280 44.880 ;
        RECT 30.920 44.710 36.015 44.880 ;
        RECT 38.475 44.710 43.570 44.880 ;
        RECT 46.285 44.710 51.380 44.880 ;
        RECT 53.795 44.710 58.890 44.880 ;
        RECT 61.470 44.710 66.565 44.880 ;
        RECT 68.980 44.710 74.075 44.880 ;
        RECT 9.825 42.350 11.310 42.520 ;
        RECT 12.560 42.350 15.795 42.520 ;
        RECT 17.600 42.350 21.255 42.520 ;
        RECT 23.185 42.350 28.280 42.520 ;
        RECT 30.920 42.350 36.015 42.520 ;
        RECT 38.475 42.350 43.570 42.520 ;
        RECT 46.285 42.350 51.380 42.520 ;
        RECT 53.795 42.350 58.890 42.520 ;
        RECT 61.470 42.350 66.565 42.520 ;
        RECT 68.980 42.350 74.075 42.520 ;
        RECT 9.825 39.990 11.310 40.160 ;
        RECT 12.560 39.990 15.795 40.160 ;
        RECT 17.600 39.990 21.255 40.160 ;
        RECT 23.185 39.990 28.280 40.160 ;
        RECT 30.920 39.990 36.015 40.160 ;
        RECT 38.475 39.990 43.570 40.160 ;
        RECT 46.285 39.990 51.380 40.160 ;
        RECT 53.795 39.990 58.890 40.160 ;
        RECT 61.470 39.990 66.565 40.160 ;
        RECT 68.980 39.990 74.075 40.160 ;
        RECT 9.825 37.630 11.310 37.800 ;
        RECT 12.560 37.630 15.795 37.800 ;
        RECT 17.600 37.630 21.255 37.800 ;
        RECT 23.185 37.630 28.280 37.800 ;
        RECT 30.920 37.630 36.015 37.800 ;
        RECT 38.475 37.630 43.570 37.800 ;
        RECT 46.285 37.630 51.380 37.800 ;
        RECT 53.795 37.630 58.890 37.800 ;
        RECT 61.470 37.630 66.565 37.800 ;
        RECT 68.980 37.630 74.075 37.800 ;
        RECT 9.825 35.270 11.310 35.440 ;
        RECT 12.560 35.270 15.795 35.440 ;
        RECT 17.600 35.270 21.255 35.440 ;
        RECT 23.185 35.270 28.280 35.440 ;
        RECT 30.920 35.270 36.015 35.440 ;
        RECT 38.475 35.270 43.570 35.440 ;
        RECT 46.285 35.270 51.380 35.440 ;
        RECT 53.795 35.270 58.890 35.440 ;
        RECT 61.470 35.270 66.565 35.440 ;
        RECT 68.980 35.270 74.075 35.440 ;
        RECT 9.825 32.910 11.310 33.080 ;
        RECT 12.560 32.910 15.795 33.080 ;
        RECT 17.600 32.910 21.255 33.080 ;
        RECT 23.185 32.910 28.280 33.080 ;
        RECT 30.920 32.910 36.015 33.080 ;
        RECT 38.475 32.910 43.570 33.080 ;
        RECT 46.285 32.910 51.380 33.080 ;
        RECT 53.795 32.910 58.890 33.080 ;
        RECT 61.470 32.910 66.565 33.080 ;
        RECT 68.980 32.910 74.075 33.080 ;
        RECT 9.825 30.550 11.310 30.720 ;
        RECT 12.560 30.550 15.795 30.720 ;
        RECT 17.600 30.550 21.255 30.720 ;
        RECT 23.185 30.550 28.280 30.720 ;
        RECT 30.920 30.550 36.015 30.720 ;
        RECT 38.475 30.550 43.570 30.720 ;
        RECT 46.285 30.550 51.380 30.720 ;
        RECT 53.795 30.550 58.890 30.720 ;
        RECT 61.470 30.550 66.565 30.720 ;
        RECT 68.980 30.550 74.075 30.720 ;
        RECT 9.825 28.190 11.310 28.360 ;
        RECT 12.560 28.190 15.795 28.360 ;
        RECT 17.600 28.190 21.255 28.360 ;
        RECT 23.185 28.190 28.280 28.360 ;
        RECT 30.920 28.190 36.015 28.360 ;
        RECT 38.475 28.190 43.570 28.360 ;
        RECT 46.285 28.190 51.380 28.360 ;
        RECT 53.795 28.190 58.890 28.360 ;
        RECT 61.470 28.190 66.565 28.360 ;
        RECT 68.980 28.190 74.075 28.360 ;
        RECT 9.825 25.830 11.310 26.000 ;
        RECT 12.560 25.830 15.795 26.000 ;
        RECT 17.600 25.830 21.255 26.000 ;
        RECT 23.185 25.830 28.280 26.000 ;
        RECT 30.920 25.830 36.015 26.000 ;
        RECT 38.475 25.830 43.570 26.000 ;
        RECT 46.285 25.830 51.380 26.000 ;
        RECT 53.795 25.830 58.890 26.000 ;
        RECT 61.470 25.830 66.565 26.000 ;
        RECT 68.980 25.830 74.075 26.000 ;
        RECT 9.825 23.470 11.310 23.640 ;
        RECT 12.560 23.470 15.795 23.640 ;
        RECT 17.600 23.470 21.255 23.640 ;
        RECT 23.185 23.470 28.280 23.640 ;
        RECT 30.920 23.470 36.015 23.640 ;
        RECT 38.475 23.470 43.570 23.640 ;
        RECT 46.285 23.470 51.380 23.640 ;
        RECT 53.795 23.470 58.890 23.640 ;
        RECT 61.470 23.470 66.565 23.640 ;
        RECT 68.980 23.470 74.075 23.640 ;
        RECT 9.825 21.110 11.310 21.280 ;
        RECT 12.560 21.110 15.795 21.280 ;
        RECT 17.600 21.110 21.255 21.280 ;
        RECT 23.185 21.110 28.280 21.280 ;
        RECT 30.920 21.110 36.015 21.280 ;
        RECT 38.475 21.110 43.570 21.280 ;
        RECT 46.285 21.110 51.380 21.280 ;
        RECT 53.795 21.110 58.890 21.280 ;
        RECT 61.470 21.110 66.565 21.280 ;
        RECT 68.980 21.110 74.075 21.280 ;
        RECT 9.825 18.750 11.310 18.920 ;
        RECT 12.560 18.750 15.795 18.920 ;
        RECT 17.600 18.750 21.255 18.920 ;
        RECT 23.185 18.750 28.280 18.920 ;
        RECT 30.920 18.750 36.015 18.920 ;
        RECT 38.475 18.750 43.570 18.920 ;
        RECT 46.285 18.750 51.380 18.920 ;
        RECT 53.795 18.750 58.890 18.920 ;
        RECT 61.470 18.750 66.565 18.920 ;
        RECT 68.980 18.750 74.075 18.920 ;
        RECT 9.825 16.390 11.310 16.560 ;
        RECT 12.560 16.390 15.795 16.560 ;
        RECT 17.600 16.390 21.255 16.560 ;
        RECT 23.185 16.390 28.280 16.560 ;
        RECT 30.920 16.390 36.015 16.560 ;
        RECT 38.475 16.390 43.570 16.560 ;
        RECT 46.285 16.390 51.380 16.560 ;
        RECT 53.795 16.390 58.890 16.560 ;
        RECT 61.470 16.390 66.565 16.560 ;
        RECT 68.980 16.390 74.075 16.560 ;
        RECT 9.825 14.030 11.310 14.200 ;
        RECT 12.560 14.030 15.795 14.200 ;
        RECT 17.600 14.030 21.255 14.200 ;
        RECT 23.185 14.030 28.280 14.200 ;
        RECT 30.920 14.030 36.015 14.200 ;
        RECT 38.475 14.030 43.570 14.200 ;
        RECT 46.285 14.030 51.380 14.200 ;
        RECT 53.795 14.030 58.890 14.200 ;
        RECT 61.470 14.030 66.565 14.200 ;
        RECT 68.980 14.030 74.075 14.200 ;
        RECT 9.825 11.670 11.310 11.840 ;
        RECT 12.560 11.670 15.795 11.840 ;
        RECT 17.600 11.670 21.255 11.840 ;
        RECT 23.185 11.670 28.280 11.840 ;
        RECT 30.920 11.670 36.015 11.840 ;
        RECT 38.475 11.670 43.570 11.840 ;
        RECT 46.285 11.670 51.380 11.840 ;
        RECT 53.795 11.670 58.890 11.840 ;
        RECT 61.470 11.670 66.565 11.840 ;
        RECT 68.980 11.670 74.075 11.840 ;
      LAYER mcon ;
        RECT 10.445 47.105 10.615 47.275 ;
        RECT 10.805 47.105 10.975 47.275 ;
        RECT 14.930 47.105 15.100 47.275 ;
        RECT 15.290 47.105 15.460 47.275 ;
        RECT 20.390 47.105 20.560 47.275 ;
        RECT 20.750 47.105 20.920 47.275 ;
        RECT 27.415 47.105 27.585 47.275 ;
        RECT 27.775 47.105 27.945 47.275 ;
        RECT 28.770 47.270 28.940 47.440 ;
        RECT 29.130 47.270 29.300 47.440 ;
        RECT 35.150 47.105 35.320 47.275 ;
        RECT 35.510 47.105 35.680 47.275 ;
        RECT 36.505 47.270 36.675 47.440 ;
        RECT 36.865 47.270 37.035 47.440 ;
        RECT 42.705 47.105 42.875 47.275 ;
        RECT 43.065 47.105 43.235 47.275 ;
        RECT 44.060 47.270 44.230 47.440 ;
        RECT 44.420 47.270 44.590 47.440 ;
        RECT 50.515 47.105 50.685 47.275 ;
        RECT 50.875 47.105 51.045 47.275 ;
        RECT 51.870 47.270 52.040 47.440 ;
        RECT 52.230 47.270 52.400 47.440 ;
        RECT 58.025 47.105 58.195 47.275 ;
        RECT 58.385 47.105 58.555 47.275 ;
        RECT 59.380 47.270 59.550 47.440 ;
        RECT 59.740 47.270 59.910 47.440 ;
        RECT 65.700 47.105 65.870 47.275 ;
        RECT 66.060 47.105 66.230 47.275 ;
        RECT 67.055 47.270 67.225 47.440 ;
        RECT 67.415 47.270 67.585 47.440 ;
        RECT 73.210 47.105 73.380 47.275 ;
        RECT 73.570 47.105 73.740 47.275 ;
        RECT 74.565 47.270 74.735 47.440 ;
        RECT 74.925 47.270 75.095 47.440 ;
        RECT 77.600 45.215 77.770 45.385 ;
        RECT 78.060 45.215 78.230 45.385 ;
        RECT 78.740 45.215 78.910 45.385 ;
        RECT 10.445 44.710 10.615 44.880 ;
        RECT 10.805 44.710 10.975 44.880 ;
        RECT 14.930 44.710 15.100 44.880 ;
        RECT 15.290 44.710 15.460 44.880 ;
        RECT 20.390 44.710 20.560 44.880 ;
        RECT 20.750 44.710 20.920 44.880 ;
        RECT 27.415 44.710 27.585 44.880 ;
        RECT 27.775 44.710 27.945 44.880 ;
        RECT 35.150 44.710 35.320 44.880 ;
        RECT 35.510 44.710 35.680 44.880 ;
        RECT 42.705 44.710 42.875 44.880 ;
        RECT 43.065 44.710 43.235 44.880 ;
        RECT 50.515 44.710 50.685 44.880 ;
        RECT 50.875 44.710 51.045 44.880 ;
        RECT 58.025 44.710 58.195 44.880 ;
        RECT 58.385 44.710 58.555 44.880 ;
        RECT 65.700 44.710 65.870 44.880 ;
        RECT 66.060 44.710 66.230 44.880 ;
        RECT 73.210 44.710 73.380 44.880 ;
        RECT 73.570 44.710 73.740 44.880 ;
        RECT 10.445 42.350 10.615 42.520 ;
        RECT 10.805 42.350 10.975 42.520 ;
        RECT 14.930 42.350 15.100 42.520 ;
        RECT 15.290 42.350 15.460 42.520 ;
        RECT 20.390 42.350 20.560 42.520 ;
        RECT 20.750 42.350 20.920 42.520 ;
        RECT 27.415 42.350 27.585 42.520 ;
        RECT 27.775 42.350 27.945 42.520 ;
        RECT 35.150 42.350 35.320 42.520 ;
        RECT 35.510 42.350 35.680 42.520 ;
        RECT 42.705 42.350 42.875 42.520 ;
        RECT 43.065 42.350 43.235 42.520 ;
        RECT 50.515 42.350 50.685 42.520 ;
        RECT 50.875 42.350 51.045 42.520 ;
        RECT 58.025 42.350 58.195 42.520 ;
        RECT 58.385 42.350 58.555 42.520 ;
        RECT 65.700 42.350 65.870 42.520 ;
        RECT 66.060 42.350 66.230 42.520 ;
        RECT 73.210 42.350 73.380 42.520 ;
        RECT 73.570 42.350 73.740 42.520 ;
        RECT 10.445 39.990 10.615 40.160 ;
        RECT 10.805 39.990 10.975 40.160 ;
        RECT 14.930 39.990 15.100 40.160 ;
        RECT 15.290 39.990 15.460 40.160 ;
        RECT 20.390 39.990 20.560 40.160 ;
        RECT 20.750 39.990 20.920 40.160 ;
        RECT 27.415 39.990 27.585 40.160 ;
        RECT 27.775 39.990 27.945 40.160 ;
        RECT 35.150 39.990 35.320 40.160 ;
        RECT 35.510 39.990 35.680 40.160 ;
        RECT 42.705 39.990 42.875 40.160 ;
        RECT 43.065 39.990 43.235 40.160 ;
        RECT 50.515 39.990 50.685 40.160 ;
        RECT 50.875 39.990 51.045 40.160 ;
        RECT 58.025 39.990 58.195 40.160 ;
        RECT 58.385 39.990 58.555 40.160 ;
        RECT 65.700 39.990 65.870 40.160 ;
        RECT 66.060 39.990 66.230 40.160 ;
        RECT 73.210 39.990 73.380 40.160 ;
        RECT 73.570 39.990 73.740 40.160 ;
        RECT 10.445 37.630 10.615 37.800 ;
        RECT 10.805 37.630 10.975 37.800 ;
        RECT 14.930 37.630 15.100 37.800 ;
        RECT 15.290 37.630 15.460 37.800 ;
        RECT 20.390 37.630 20.560 37.800 ;
        RECT 20.750 37.630 20.920 37.800 ;
        RECT 27.415 37.630 27.585 37.800 ;
        RECT 27.775 37.630 27.945 37.800 ;
        RECT 35.150 37.630 35.320 37.800 ;
        RECT 35.510 37.630 35.680 37.800 ;
        RECT 42.705 37.630 42.875 37.800 ;
        RECT 43.065 37.630 43.235 37.800 ;
        RECT 50.515 37.630 50.685 37.800 ;
        RECT 50.875 37.630 51.045 37.800 ;
        RECT 58.025 37.630 58.195 37.800 ;
        RECT 58.385 37.630 58.555 37.800 ;
        RECT 65.700 37.630 65.870 37.800 ;
        RECT 66.060 37.630 66.230 37.800 ;
        RECT 73.210 37.630 73.380 37.800 ;
        RECT 73.570 37.630 73.740 37.800 ;
        RECT 10.445 35.270 10.615 35.440 ;
        RECT 10.805 35.270 10.975 35.440 ;
        RECT 14.930 35.270 15.100 35.440 ;
        RECT 15.290 35.270 15.460 35.440 ;
        RECT 20.390 35.270 20.560 35.440 ;
        RECT 20.750 35.270 20.920 35.440 ;
        RECT 27.415 35.270 27.585 35.440 ;
        RECT 27.775 35.270 27.945 35.440 ;
        RECT 35.150 35.270 35.320 35.440 ;
        RECT 35.510 35.270 35.680 35.440 ;
        RECT 42.705 35.270 42.875 35.440 ;
        RECT 43.065 35.270 43.235 35.440 ;
        RECT 50.515 35.270 50.685 35.440 ;
        RECT 50.875 35.270 51.045 35.440 ;
        RECT 58.025 35.270 58.195 35.440 ;
        RECT 58.385 35.270 58.555 35.440 ;
        RECT 65.700 35.270 65.870 35.440 ;
        RECT 66.060 35.270 66.230 35.440 ;
        RECT 73.210 35.270 73.380 35.440 ;
        RECT 73.570 35.270 73.740 35.440 ;
        RECT 10.445 32.910 10.615 33.080 ;
        RECT 10.805 32.910 10.975 33.080 ;
        RECT 14.930 32.910 15.100 33.080 ;
        RECT 15.290 32.910 15.460 33.080 ;
        RECT 20.390 32.910 20.560 33.080 ;
        RECT 20.750 32.910 20.920 33.080 ;
        RECT 27.415 32.910 27.585 33.080 ;
        RECT 27.775 32.910 27.945 33.080 ;
        RECT 35.150 32.910 35.320 33.080 ;
        RECT 35.510 32.910 35.680 33.080 ;
        RECT 42.705 32.910 42.875 33.080 ;
        RECT 43.065 32.910 43.235 33.080 ;
        RECT 50.515 32.910 50.685 33.080 ;
        RECT 50.875 32.910 51.045 33.080 ;
        RECT 58.025 32.910 58.195 33.080 ;
        RECT 58.385 32.910 58.555 33.080 ;
        RECT 65.700 32.910 65.870 33.080 ;
        RECT 66.060 32.910 66.230 33.080 ;
        RECT 73.210 32.910 73.380 33.080 ;
        RECT 73.570 32.910 73.740 33.080 ;
        RECT 10.445 30.550 10.615 30.720 ;
        RECT 10.805 30.550 10.975 30.720 ;
        RECT 14.930 30.550 15.100 30.720 ;
        RECT 15.290 30.550 15.460 30.720 ;
        RECT 20.390 30.550 20.560 30.720 ;
        RECT 20.750 30.550 20.920 30.720 ;
        RECT 27.415 30.550 27.585 30.720 ;
        RECT 27.775 30.550 27.945 30.720 ;
        RECT 35.150 30.550 35.320 30.720 ;
        RECT 35.510 30.550 35.680 30.720 ;
        RECT 42.705 30.550 42.875 30.720 ;
        RECT 43.065 30.550 43.235 30.720 ;
        RECT 50.515 30.550 50.685 30.720 ;
        RECT 50.875 30.550 51.045 30.720 ;
        RECT 58.025 30.550 58.195 30.720 ;
        RECT 58.385 30.550 58.555 30.720 ;
        RECT 65.700 30.550 65.870 30.720 ;
        RECT 66.060 30.550 66.230 30.720 ;
        RECT 73.210 30.550 73.380 30.720 ;
        RECT 73.570 30.550 73.740 30.720 ;
        RECT 10.445 28.190 10.615 28.360 ;
        RECT 10.805 28.190 10.975 28.360 ;
        RECT 14.930 28.190 15.100 28.360 ;
        RECT 15.290 28.190 15.460 28.360 ;
        RECT 20.390 28.190 20.560 28.360 ;
        RECT 20.750 28.190 20.920 28.360 ;
        RECT 27.415 28.190 27.585 28.360 ;
        RECT 27.775 28.190 27.945 28.360 ;
        RECT 35.150 28.190 35.320 28.360 ;
        RECT 35.510 28.190 35.680 28.360 ;
        RECT 42.705 28.190 42.875 28.360 ;
        RECT 43.065 28.190 43.235 28.360 ;
        RECT 50.515 28.190 50.685 28.360 ;
        RECT 50.875 28.190 51.045 28.360 ;
        RECT 58.025 28.190 58.195 28.360 ;
        RECT 58.385 28.190 58.555 28.360 ;
        RECT 65.700 28.190 65.870 28.360 ;
        RECT 66.060 28.190 66.230 28.360 ;
        RECT 73.210 28.190 73.380 28.360 ;
        RECT 73.570 28.190 73.740 28.360 ;
        RECT 10.445 25.830 10.615 26.000 ;
        RECT 10.805 25.830 10.975 26.000 ;
        RECT 14.930 25.830 15.100 26.000 ;
        RECT 15.290 25.830 15.460 26.000 ;
        RECT 20.390 25.830 20.560 26.000 ;
        RECT 20.750 25.830 20.920 26.000 ;
        RECT 27.415 25.830 27.585 26.000 ;
        RECT 27.775 25.830 27.945 26.000 ;
        RECT 35.150 25.830 35.320 26.000 ;
        RECT 35.510 25.830 35.680 26.000 ;
        RECT 42.705 25.830 42.875 26.000 ;
        RECT 43.065 25.830 43.235 26.000 ;
        RECT 50.515 25.830 50.685 26.000 ;
        RECT 50.875 25.830 51.045 26.000 ;
        RECT 58.025 25.830 58.195 26.000 ;
        RECT 58.385 25.830 58.555 26.000 ;
        RECT 65.700 25.830 65.870 26.000 ;
        RECT 66.060 25.830 66.230 26.000 ;
        RECT 73.210 25.830 73.380 26.000 ;
        RECT 73.570 25.830 73.740 26.000 ;
        RECT 10.445 23.470 10.615 23.640 ;
        RECT 10.805 23.470 10.975 23.640 ;
        RECT 14.930 23.470 15.100 23.640 ;
        RECT 15.290 23.470 15.460 23.640 ;
        RECT 20.390 23.470 20.560 23.640 ;
        RECT 20.750 23.470 20.920 23.640 ;
        RECT 27.415 23.470 27.585 23.640 ;
        RECT 27.775 23.470 27.945 23.640 ;
        RECT 35.150 23.470 35.320 23.640 ;
        RECT 35.510 23.470 35.680 23.640 ;
        RECT 42.705 23.470 42.875 23.640 ;
        RECT 43.065 23.470 43.235 23.640 ;
        RECT 50.515 23.470 50.685 23.640 ;
        RECT 50.875 23.470 51.045 23.640 ;
        RECT 58.025 23.470 58.195 23.640 ;
        RECT 58.385 23.470 58.555 23.640 ;
        RECT 65.700 23.470 65.870 23.640 ;
        RECT 66.060 23.470 66.230 23.640 ;
        RECT 73.210 23.470 73.380 23.640 ;
        RECT 73.570 23.470 73.740 23.640 ;
        RECT 10.445 21.110 10.615 21.280 ;
        RECT 10.805 21.110 10.975 21.280 ;
        RECT 14.930 21.110 15.100 21.280 ;
        RECT 15.290 21.110 15.460 21.280 ;
        RECT 20.390 21.110 20.560 21.280 ;
        RECT 20.750 21.110 20.920 21.280 ;
        RECT 27.415 21.110 27.585 21.280 ;
        RECT 27.775 21.110 27.945 21.280 ;
        RECT 35.150 21.110 35.320 21.280 ;
        RECT 35.510 21.110 35.680 21.280 ;
        RECT 42.705 21.110 42.875 21.280 ;
        RECT 43.065 21.110 43.235 21.280 ;
        RECT 50.515 21.110 50.685 21.280 ;
        RECT 50.875 21.110 51.045 21.280 ;
        RECT 58.025 21.110 58.195 21.280 ;
        RECT 58.385 21.110 58.555 21.280 ;
        RECT 65.700 21.110 65.870 21.280 ;
        RECT 66.060 21.110 66.230 21.280 ;
        RECT 73.210 21.110 73.380 21.280 ;
        RECT 73.570 21.110 73.740 21.280 ;
        RECT 10.445 18.750 10.615 18.920 ;
        RECT 10.805 18.750 10.975 18.920 ;
        RECT 14.930 18.750 15.100 18.920 ;
        RECT 15.290 18.750 15.460 18.920 ;
        RECT 20.390 18.750 20.560 18.920 ;
        RECT 20.750 18.750 20.920 18.920 ;
        RECT 27.415 18.750 27.585 18.920 ;
        RECT 27.775 18.750 27.945 18.920 ;
        RECT 35.150 18.750 35.320 18.920 ;
        RECT 35.510 18.750 35.680 18.920 ;
        RECT 42.705 18.750 42.875 18.920 ;
        RECT 43.065 18.750 43.235 18.920 ;
        RECT 50.515 18.750 50.685 18.920 ;
        RECT 50.875 18.750 51.045 18.920 ;
        RECT 58.025 18.750 58.195 18.920 ;
        RECT 58.385 18.750 58.555 18.920 ;
        RECT 65.700 18.750 65.870 18.920 ;
        RECT 66.060 18.750 66.230 18.920 ;
        RECT 73.210 18.750 73.380 18.920 ;
        RECT 73.570 18.750 73.740 18.920 ;
        RECT 10.445 16.390 10.615 16.560 ;
        RECT 10.805 16.390 10.975 16.560 ;
        RECT 14.930 16.390 15.100 16.560 ;
        RECT 15.290 16.390 15.460 16.560 ;
        RECT 20.390 16.390 20.560 16.560 ;
        RECT 20.750 16.390 20.920 16.560 ;
        RECT 27.415 16.390 27.585 16.560 ;
        RECT 27.775 16.390 27.945 16.560 ;
        RECT 35.150 16.390 35.320 16.560 ;
        RECT 35.510 16.390 35.680 16.560 ;
        RECT 42.705 16.390 42.875 16.560 ;
        RECT 43.065 16.390 43.235 16.560 ;
        RECT 50.515 16.390 50.685 16.560 ;
        RECT 50.875 16.390 51.045 16.560 ;
        RECT 58.025 16.390 58.195 16.560 ;
        RECT 58.385 16.390 58.555 16.560 ;
        RECT 65.700 16.390 65.870 16.560 ;
        RECT 66.060 16.390 66.230 16.560 ;
        RECT 73.210 16.390 73.380 16.560 ;
        RECT 73.570 16.390 73.740 16.560 ;
        RECT 10.445 14.030 10.615 14.200 ;
        RECT 10.805 14.030 10.975 14.200 ;
        RECT 14.930 14.030 15.100 14.200 ;
        RECT 15.290 14.030 15.460 14.200 ;
        RECT 20.390 14.030 20.560 14.200 ;
        RECT 20.750 14.030 20.920 14.200 ;
        RECT 27.415 14.030 27.585 14.200 ;
        RECT 27.775 14.030 27.945 14.200 ;
        RECT 35.150 14.030 35.320 14.200 ;
        RECT 35.510 14.030 35.680 14.200 ;
        RECT 42.705 14.030 42.875 14.200 ;
        RECT 43.065 14.030 43.235 14.200 ;
        RECT 50.515 14.030 50.685 14.200 ;
        RECT 50.875 14.030 51.045 14.200 ;
        RECT 58.025 14.030 58.195 14.200 ;
        RECT 58.385 14.030 58.555 14.200 ;
        RECT 65.700 14.030 65.870 14.200 ;
        RECT 66.060 14.030 66.230 14.200 ;
        RECT 73.210 14.030 73.380 14.200 ;
        RECT 73.570 14.030 73.740 14.200 ;
        RECT 10.445 11.670 10.615 11.840 ;
        RECT 10.805 11.670 10.975 11.840 ;
        RECT 14.930 11.670 15.100 11.840 ;
        RECT 15.290 11.670 15.460 11.840 ;
        RECT 20.390 11.670 20.560 11.840 ;
        RECT 20.750 11.670 20.920 11.840 ;
        RECT 27.415 11.670 27.585 11.840 ;
        RECT 27.775 11.670 27.945 11.840 ;
        RECT 35.150 11.670 35.320 11.840 ;
        RECT 35.510 11.670 35.680 11.840 ;
        RECT 42.705 11.670 42.875 11.840 ;
        RECT 43.065 11.670 43.235 11.840 ;
        RECT 50.515 11.670 50.685 11.840 ;
        RECT 50.875 11.670 51.045 11.840 ;
        RECT 58.025 11.670 58.195 11.840 ;
        RECT 58.385 11.670 58.555 11.840 ;
        RECT 65.700 11.670 65.870 11.840 ;
        RECT 66.060 11.670 66.230 11.840 ;
        RECT 73.210 11.670 73.380 11.840 ;
        RECT 73.570 11.670 73.740 11.840 ;
      LAYER met1 ;
        RECT 10.105 46.920 75.990 47.580 ;
        RECT 75.340 45.535 75.990 46.920 ;
        RECT 75.340 45.165 80.840 45.535 ;
        RECT 75.350 45.155 80.840 45.165 ;
        RECT 10.385 44.680 11.035 44.910 ;
        RECT 14.870 44.680 15.520 44.910 ;
        RECT 20.330 44.680 20.980 44.910 ;
        RECT 27.355 44.680 28.005 44.910 ;
        RECT 35.090 44.680 35.740 44.910 ;
        RECT 42.645 44.680 43.295 44.910 ;
        RECT 50.455 44.680 51.105 44.910 ;
        RECT 57.965 44.680 58.615 44.910 ;
        RECT 65.640 44.680 66.290 44.910 ;
        RECT 73.150 44.680 73.800 44.910 ;
        RECT 10.385 44.650 11.025 44.680 ;
        RECT 14.870 44.650 15.510 44.680 ;
        RECT 20.330 44.650 20.970 44.680 ;
        RECT 27.355 44.650 27.995 44.680 ;
        RECT 35.090 44.650 35.730 44.680 ;
        RECT 42.645 44.650 43.285 44.680 ;
        RECT 50.455 44.650 51.095 44.680 ;
        RECT 57.965 44.650 58.605 44.680 ;
        RECT 65.640 44.650 66.280 44.680 ;
        RECT 73.150 44.650 73.790 44.680 ;
        RECT 10.385 42.550 11.025 42.560 ;
        RECT 14.870 42.550 15.510 42.560 ;
        RECT 20.330 42.550 20.970 42.560 ;
        RECT 27.355 42.550 27.995 42.560 ;
        RECT 35.090 42.550 35.730 42.560 ;
        RECT 42.645 42.550 43.285 42.560 ;
        RECT 50.455 42.550 51.095 42.560 ;
        RECT 57.965 42.550 58.605 42.560 ;
        RECT 65.640 42.550 66.280 42.560 ;
        RECT 73.150 42.550 73.790 42.560 ;
        RECT 10.385 42.320 11.035 42.550 ;
        RECT 14.870 42.320 15.520 42.550 ;
        RECT 20.330 42.320 20.980 42.550 ;
        RECT 27.355 42.320 28.005 42.550 ;
        RECT 35.090 42.320 35.740 42.550 ;
        RECT 42.645 42.320 43.295 42.550 ;
        RECT 50.455 42.320 51.105 42.550 ;
        RECT 57.965 42.320 58.615 42.550 ;
        RECT 65.640 42.320 66.290 42.550 ;
        RECT 73.150 42.320 73.800 42.550 ;
        RECT 10.385 42.300 11.025 42.320 ;
        RECT 14.870 42.300 15.510 42.320 ;
        RECT 20.330 42.300 20.970 42.320 ;
        RECT 27.355 42.300 27.995 42.320 ;
        RECT 35.090 42.300 35.730 42.320 ;
        RECT 42.645 42.300 43.285 42.320 ;
        RECT 50.455 42.300 51.095 42.320 ;
        RECT 57.965 42.300 58.605 42.320 ;
        RECT 65.640 42.300 66.280 42.320 ;
        RECT 73.150 42.300 73.790 42.320 ;
        RECT 10.385 40.190 11.025 40.200 ;
        RECT 14.870 40.190 15.510 40.200 ;
        RECT 20.330 40.190 20.970 40.200 ;
        RECT 27.355 40.190 27.995 40.200 ;
        RECT 35.090 40.190 35.730 40.200 ;
        RECT 42.645 40.190 43.285 40.200 ;
        RECT 50.455 40.190 51.095 40.200 ;
        RECT 57.965 40.190 58.605 40.200 ;
        RECT 65.640 40.190 66.280 40.200 ;
        RECT 73.150 40.190 73.790 40.200 ;
        RECT 10.385 39.960 11.035 40.190 ;
        RECT 14.870 39.960 15.520 40.190 ;
        RECT 20.330 39.960 20.980 40.190 ;
        RECT 27.355 39.960 28.005 40.190 ;
        RECT 35.090 39.960 35.740 40.190 ;
        RECT 42.645 39.960 43.295 40.190 ;
        RECT 50.455 39.960 51.105 40.190 ;
        RECT 57.965 39.960 58.615 40.190 ;
        RECT 65.640 39.960 66.290 40.190 ;
        RECT 73.150 39.960 73.800 40.190 ;
        RECT 10.385 39.940 11.025 39.960 ;
        RECT 14.870 39.940 15.510 39.960 ;
        RECT 20.330 39.940 20.970 39.960 ;
        RECT 27.355 39.940 27.995 39.960 ;
        RECT 35.090 39.940 35.730 39.960 ;
        RECT 42.645 39.940 43.285 39.960 ;
        RECT 50.455 39.940 51.095 39.960 ;
        RECT 57.965 39.940 58.605 39.960 ;
        RECT 65.640 39.940 66.280 39.960 ;
        RECT 73.150 39.940 73.790 39.960 ;
        RECT 10.385 37.830 11.025 37.845 ;
        RECT 14.870 37.830 15.510 37.845 ;
        RECT 20.330 37.830 20.970 37.845 ;
        RECT 27.355 37.830 27.995 37.845 ;
        RECT 35.090 37.830 35.730 37.845 ;
        RECT 42.645 37.830 43.285 37.845 ;
        RECT 50.455 37.830 51.095 37.845 ;
        RECT 57.965 37.830 58.605 37.845 ;
        RECT 65.640 37.830 66.280 37.845 ;
        RECT 73.150 37.830 73.790 37.845 ;
        RECT 10.385 37.600 11.035 37.830 ;
        RECT 14.870 37.600 15.520 37.830 ;
        RECT 20.330 37.600 20.980 37.830 ;
        RECT 27.355 37.600 28.005 37.830 ;
        RECT 35.090 37.600 35.740 37.830 ;
        RECT 42.645 37.600 43.295 37.830 ;
        RECT 50.455 37.600 51.105 37.830 ;
        RECT 57.965 37.600 58.615 37.830 ;
        RECT 65.640 37.600 66.290 37.830 ;
        RECT 73.150 37.600 73.800 37.830 ;
        RECT 10.385 37.585 11.025 37.600 ;
        RECT 14.870 37.585 15.510 37.600 ;
        RECT 20.330 37.585 20.970 37.600 ;
        RECT 27.355 37.585 27.995 37.600 ;
        RECT 35.090 37.585 35.730 37.600 ;
        RECT 42.645 37.585 43.285 37.600 ;
        RECT 50.455 37.585 51.095 37.600 ;
        RECT 57.965 37.585 58.605 37.600 ;
        RECT 65.640 37.585 66.280 37.600 ;
        RECT 73.150 37.585 73.790 37.600 ;
        RECT 10.385 35.470 11.025 35.485 ;
        RECT 14.870 35.470 15.510 35.485 ;
        RECT 20.330 35.470 20.970 35.485 ;
        RECT 27.355 35.470 27.995 35.485 ;
        RECT 35.090 35.470 35.730 35.485 ;
        RECT 42.645 35.470 43.285 35.485 ;
        RECT 50.455 35.470 51.095 35.485 ;
        RECT 57.965 35.470 58.605 35.485 ;
        RECT 65.640 35.470 66.280 35.485 ;
        RECT 73.150 35.470 73.790 35.485 ;
        RECT 10.385 35.240 11.035 35.470 ;
        RECT 14.870 35.240 15.520 35.470 ;
        RECT 20.330 35.240 20.980 35.470 ;
        RECT 27.355 35.240 28.005 35.470 ;
        RECT 35.090 35.240 35.740 35.470 ;
        RECT 42.645 35.240 43.295 35.470 ;
        RECT 50.455 35.240 51.105 35.470 ;
        RECT 57.965 35.240 58.615 35.470 ;
        RECT 65.640 35.240 66.290 35.470 ;
        RECT 73.150 35.240 73.800 35.470 ;
        RECT 10.385 35.225 11.025 35.240 ;
        RECT 14.870 35.225 15.510 35.240 ;
        RECT 20.330 35.225 20.970 35.240 ;
        RECT 27.355 35.225 27.995 35.240 ;
        RECT 35.090 35.225 35.730 35.240 ;
        RECT 42.645 35.225 43.285 35.240 ;
        RECT 50.455 35.225 51.095 35.240 ;
        RECT 57.965 35.225 58.605 35.240 ;
        RECT 65.640 35.225 66.280 35.240 ;
        RECT 73.150 35.225 73.790 35.240 ;
        RECT 10.385 33.110 11.025 33.120 ;
        RECT 14.870 33.110 15.510 33.120 ;
        RECT 20.330 33.110 20.970 33.120 ;
        RECT 27.355 33.110 27.995 33.120 ;
        RECT 35.090 33.110 35.730 33.120 ;
        RECT 42.645 33.110 43.285 33.120 ;
        RECT 50.455 33.110 51.095 33.120 ;
        RECT 57.965 33.110 58.605 33.120 ;
        RECT 65.640 33.110 66.280 33.120 ;
        RECT 73.150 33.110 73.790 33.120 ;
        RECT 10.385 32.880 11.035 33.110 ;
        RECT 14.870 32.880 15.520 33.110 ;
        RECT 20.330 32.880 20.980 33.110 ;
        RECT 27.355 32.880 28.005 33.110 ;
        RECT 35.090 32.880 35.740 33.110 ;
        RECT 42.645 32.880 43.295 33.110 ;
        RECT 50.455 32.880 51.105 33.110 ;
        RECT 57.965 32.880 58.615 33.110 ;
        RECT 65.640 32.880 66.290 33.110 ;
        RECT 73.150 32.880 73.800 33.110 ;
        RECT 10.385 32.860 11.025 32.880 ;
        RECT 14.870 32.860 15.510 32.880 ;
        RECT 20.330 32.860 20.970 32.880 ;
        RECT 27.355 32.860 27.995 32.880 ;
        RECT 35.090 32.860 35.730 32.880 ;
        RECT 42.645 32.860 43.285 32.880 ;
        RECT 50.455 32.860 51.095 32.880 ;
        RECT 57.965 32.860 58.605 32.880 ;
        RECT 65.640 32.860 66.280 32.880 ;
        RECT 73.150 32.860 73.790 32.880 ;
        RECT 10.385 30.750 11.025 30.765 ;
        RECT 14.870 30.750 15.510 30.765 ;
        RECT 20.330 30.750 20.970 30.765 ;
        RECT 27.355 30.750 27.995 30.765 ;
        RECT 35.090 30.750 35.730 30.765 ;
        RECT 42.645 30.750 43.285 30.765 ;
        RECT 50.455 30.750 51.095 30.765 ;
        RECT 57.965 30.750 58.605 30.765 ;
        RECT 65.640 30.750 66.280 30.765 ;
        RECT 73.150 30.750 73.790 30.765 ;
        RECT 10.385 30.520 11.035 30.750 ;
        RECT 14.870 30.520 15.520 30.750 ;
        RECT 20.330 30.520 20.980 30.750 ;
        RECT 27.355 30.520 28.005 30.750 ;
        RECT 35.090 30.520 35.740 30.750 ;
        RECT 42.645 30.520 43.295 30.750 ;
        RECT 50.455 30.520 51.105 30.750 ;
        RECT 57.965 30.520 58.615 30.750 ;
        RECT 65.640 30.520 66.290 30.750 ;
        RECT 73.150 30.520 73.800 30.750 ;
        RECT 10.385 30.505 11.025 30.520 ;
        RECT 14.870 30.505 15.510 30.520 ;
        RECT 20.330 30.505 20.970 30.520 ;
        RECT 27.355 30.505 27.995 30.520 ;
        RECT 35.090 30.505 35.730 30.520 ;
        RECT 42.645 30.505 43.285 30.520 ;
        RECT 50.455 30.505 51.095 30.520 ;
        RECT 57.965 30.505 58.605 30.520 ;
        RECT 65.640 30.505 66.280 30.520 ;
        RECT 73.150 30.505 73.790 30.520 ;
        RECT 10.385 28.390 11.025 28.405 ;
        RECT 14.870 28.390 15.510 28.405 ;
        RECT 20.330 28.390 20.970 28.405 ;
        RECT 27.355 28.390 27.995 28.405 ;
        RECT 35.090 28.390 35.730 28.405 ;
        RECT 42.645 28.390 43.285 28.405 ;
        RECT 50.455 28.390 51.095 28.405 ;
        RECT 57.965 28.390 58.605 28.405 ;
        RECT 65.640 28.390 66.280 28.405 ;
        RECT 73.150 28.390 73.790 28.405 ;
        RECT 10.385 28.160 11.035 28.390 ;
        RECT 14.870 28.160 15.520 28.390 ;
        RECT 20.330 28.160 20.980 28.390 ;
        RECT 27.355 28.160 28.005 28.390 ;
        RECT 35.090 28.160 35.740 28.390 ;
        RECT 42.645 28.160 43.295 28.390 ;
        RECT 50.455 28.160 51.105 28.390 ;
        RECT 57.965 28.160 58.615 28.390 ;
        RECT 65.640 28.160 66.290 28.390 ;
        RECT 73.150 28.160 73.800 28.390 ;
        RECT 10.385 28.145 11.025 28.160 ;
        RECT 14.870 28.145 15.510 28.160 ;
        RECT 20.330 28.145 20.970 28.160 ;
        RECT 27.355 28.145 27.995 28.160 ;
        RECT 35.090 28.145 35.730 28.160 ;
        RECT 42.645 28.145 43.285 28.160 ;
        RECT 50.455 28.145 51.095 28.160 ;
        RECT 57.965 28.145 58.605 28.160 ;
        RECT 65.640 28.145 66.280 28.160 ;
        RECT 73.150 28.145 73.790 28.160 ;
        RECT 10.385 26.030 11.025 26.040 ;
        RECT 14.870 26.030 15.510 26.040 ;
        RECT 20.330 26.030 20.970 26.040 ;
        RECT 27.355 26.030 27.995 26.040 ;
        RECT 35.090 26.030 35.730 26.040 ;
        RECT 42.645 26.030 43.285 26.040 ;
        RECT 50.455 26.030 51.095 26.040 ;
        RECT 57.965 26.030 58.605 26.040 ;
        RECT 65.640 26.030 66.280 26.040 ;
        RECT 73.150 26.030 73.790 26.040 ;
        RECT 10.385 25.800 11.035 26.030 ;
        RECT 14.870 25.800 15.520 26.030 ;
        RECT 20.330 25.800 20.980 26.030 ;
        RECT 27.355 25.800 28.005 26.030 ;
        RECT 35.090 25.800 35.740 26.030 ;
        RECT 42.645 25.800 43.295 26.030 ;
        RECT 50.455 25.800 51.105 26.030 ;
        RECT 57.965 25.800 58.615 26.030 ;
        RECT 65.640 25.800 66.290 26.030 ;
        RECT 73.150 25.800 73.800 26.030 ;
        RECT 10.385 25.780 11.025 25.800 ;
        RECT 14.870 25.780 15.510 25.800 ;
        RECT 20.330 25.780 20.970 25.800 ;
        RECT 27.355 25.780 27.995 25.800 ;
        RECT 35.090 25.780 35.730 25.800 ;
        RECT 42.645 25.780 43.285 25.800 ;
        RECT 50.455 25.780 51.095 25.800 ;
        RECT 57.965 25.780 58.605 25.800 ;
        RECT 65.640 25.780 66.280 25.800 ;
        RECT 73.150 25.780 73.790 25.800 ;
        RECT 10.385 23.670 11.025 23.680 ;
        RECT 14.870 23.670 15.510 23.680 ;
        RECT 20.330 23.670 20.970 23.680 ;
        RECT 27.355 23.670 27.995 23.680 ;
        RECT 35.090 23.670 35.730 23.680 ;
        RECT 42.645 23.670 43.285 23.680 ;
        RECT 50.455 23.670 51.095 23.680 ;
        RECT 57.965 23.670 58.605 23.680 ;
        RECT 65.640 23.670 66.280 23.680 ;
        RECT 73.150 23.670 73.790 23.680 ;
        RECT 10.385 23.440 11.035 23.670 ;
        RECT 14.870 23.440 15.520 23.670 ;
        RECT 20.330 23.440 20.980 23.670 ;
        RECT 27.355 23.440 28.005 23.670 ;
        RECT 35.090 23.440 35.740 23.670 ;
        RECT 42.645 23.440 43.295 23.670 ;
        RECT 50.455 23.440 51.105 23.670 ;
        RECT 57.965 23.440 58.615 23.670 ;
        RECT 65.640 23.440 66.290 23.670 ;
        RECT 73.150 23.440 73.800 23.670 ;
        RECT 10.385 23.420 11.025 23.440 ;
        RECT 14.870 23.420 15.510 23.440 ;
        RECT 20.330 23.420 20.970 23.440 ;
        RECT 27.355 23.420 27.995 23.440 ;
        RECT 35.090 23.420 35.730 23.440 ;
        RECT 42.645 23.420 43.285 23.440 ;
        RECT 50.455 23.420 51.095 23.440 ;
        RECT 57.965 23.420 58.605 23.440 ;
        RECT 65.640 23.420 66.280 23.440 ;
        RECT 73.150 23.420 73.790 23.440 ;
        RECT 10.385 21.310 11.025 21.325 ;
        RECT 14.870 21.310 15.510 21.325 ;
        RECT 20.330 21.310 20.970 21.325 ;
        RECT 27.355 21.310 27.995 21.325 ;
        RECT 35.090 21.310 35.730 21.325 ;
        RECT 42.645 21.310 43.285 21.325 ;
        RECT 50.455 21.310 51.095 21.325 ;
        RECT 57.965 21.310 58.605 21.325 ;
        RECT 65.640 21.310 66.280 21.325 ;
        RECT 73.150 21.310 73.790 21.325 ;
        RECT 10.385 21.080 11.035 21.310 ;
        RECT 14.870 21.080 15.520 21.310 ;
        RECT 20.330 21.080 20.980 21.310 ;
        RECT 27.355 21.080 28.005 21.310 ;
        RECT 35.090 21.080 35.740 21.310 ;
        RECT 42.645 21.080 43.295 21.310 ;
        RECT 50.455 21.080 51.105 21.310 ;
        RECT 57.965 21.080 58.615 21.310 ;
        RECT 65.640 21.080 66.290 21.310 ;
        RECT 73.150 21.080 73.800 21.310 ;
        RECT 10.385 21.065 11.025 21.080 ;
        RECT 14.870 21.065 15.510 21.080 ;
        RECT 20.330 21.065 20.970 21.080 ;
        RECT 27.355 21.065 27.995 21.080 ;
        RECT 35.090 21.065 35.730 21.080 ;
        RECT 42.645 21.065 43.285 21.080 ;
        RECT 50.455 21.065 51.095 21.080 ;
        RECT 57.965 21.065 58.605 21.080 ;
        RECT 65.640 21.065 66.280 21.080 ;
        RECT 73.150 21.065 73.790 21.080 ;
        RECT 10.385 18.950 11.025 18.965 ;
        RECT 14.870 18.950 15.510 18.965 ;
        RECT 20.330 18.950 20.970 18.965 ;
        RECT 27.355 18.950 27.995 18.965 ;
        RECT 35.090 18.950 35.730 18.965 ;
        RECT 42.645 18.950 43.285 18.965 ;
        RECT 50.455 18.950 51.095 18.965 ;
        RECT 57.965 18.950 58.605 18.965 ;
        RECT 65.640 18.950 66.280 18.965 ;
        RECT 73.150 18.950 73.790 18.965 ;
        RECT 10.385 18.720 11.035 18.950 ;
        RECT 14.870 18.720 15.520 18.950 ;
        RECT 20.330 18.720 20.980 18.950 ;
        RECT 27.355 18.720 28.005 18.950 ;
        RECT 35.090 18.720 35.740 18.950 ;
        RECT 42.645 18.720 43.295 18.950 ;
        RECT 50.455 18.720 51.105 18.950 ;
        RECT 57.965 18.720 58.615 18.950 ;
        RECT 65.640 18.720 66.290 18.950 ;
        RECT 73.150 18.720 73.800 18.950 ;
        RECT 10.385 18.705 11.025 18.720 ;
        RECT 14.870 18.705 15.510 18.720 ;
        RECT 20.330 18.705 20.970 18.720 ;
        RECT 27.355 18.705 27.995 18.720 ;
        RECT 35.090 18.705 35.730 18.720 ;
        RECT 42.645 18.705 43.285 18.720 ;
        RECT 50.455 18.705 51.095 18.720 ;
        RECT 57.965 18.705 58.605 18.720 ;
        RECT 65.640 18.705 66.280 18.720 ;
        RECT 73.150 18.705 73.790 18.720 ;
        RECT 10.385 16.590 11.025 16.600 ;
        RECT 14.870 16.590 15.510 16.600 ;
        RECT 20.330 16.590 20.970 16.600 ;
        RECT 27.355 16.590 27.995 16.600 ;
        RECT 35.090 16.590 35.730 16.600 ;
        RECT 42.645 16.590 43.285 16.600 ;
        RECT 50.455 16.590 51.095 16.600 ;
        RECT 57.965 16.590 58.605 16.600 ;
        RECT 65.640 16.590 66.280 16.600 ;
        RECT 73.150 16.590 73.790 16.600 ;
        RECT 10.385 16.360 11.035 16.590 ;
        RECT 14.870 16.360 15.520 16.590 ;
        RECT 20.330 16.360 20.980 16.590 ;
        RECT 27.355 16.360 28.005 16.590 ;
        RECT 35.090 16.360 35.740 16.590 ;
        RECT 42.645 16.360 43.295 16.590 ;
        RECT 50.455 16.360 51.105 16.590 ;
        RECT 57.965 16.360 58.615 16.590 ;
        RECT 65.640 16.360 66.290 16.590 ;
        RECT 73.150 16.360 73.800 16.590 ;
        RECT 10.385 16.340 11.025 16.360 ;
        RECT 14.870 16.340 15.510 16.360 ;
        RECT 20.330 16.340 20.970 16.360 ;
        RECT 27.355 16.340 27.995 16.360 ;
        RECT 35.090 16.340 35.730 16.360 ;
        RECT 42.645 16.340 43.285 16.360 ;
        RECT 50.455 16.340 51.095 16.360 ;
        RECT 57.965 16.340 58.605 16.360 ;
        RECT 65.640 16.340 66.280 16.360 ;
        RECT 73.150 16.340 73.790 16.360 ;
        RECT 10.385 14.230 11.025 14.240 ;
        RECT 14.870 14.230 15.510 14.240 ;
        RECT 20.330 14.230 20.970 14.240 ;
        RECT 27.355 14.230 27.995 14.240 ;
        RECT 35.090 14.230 35.730 14.240 ;
        RECT 42.645 14.230 43.285 14.240 ;
        RECT 50.455 14.230 51.095 14.240 ;
        RECT 57.965 14.230 58.605 14.240 ;
        RECT 65.640 14.230 66.280 14.240 ;
        RECT 73.150 14.230 73.790 14.240 ;
        RECT 10.385 14.000 11.035 14.230 ;
        RECT 14.870 14.000 15.520 14.230 ;
        RECT 20.330 14.000 20.980 14.230 ;
        RECT 27.355 14.000 28.005 14.230 ;
        RECT 35.090 14.000 35.740 14.230 ;
        RECT 42.645 14.000 43.295 14.230 ;
        RECT 50.455 14.000 51.105 14.230 ;
        RECT 57.965 14.000 58.615 14.230 ;
        RECT 65.640 14.000 66.290 14.230 ;
        RECT 73.150 14.000 73.800 14.230 ;
        RECT 10.385 13.980 11.025 14.000 ;
        RECT 14.870 13.980 15.510 14.000 ;
        RECT 20.330 13.980 20.970 14.000 ;
        RECT 27.355 13.980 27.995 14.000 ;
        RECT 35.090 13.980 35.730 14.000 ;
        RECT 42.645 13.980 43.285 14.000 ;
        RECT 50.455 13.980 51.095 14.000 ;
        RECT 57.965 13.980 58.605 14.000 ;
        RECT 65.640 13.980 66.280 14.000 ;
        RECT 73.150 13.980 73.790 14.000 ;
        RECT 10.385 11.870 11.025 11.880 ;
        RECT 14.870 11.870 15.510 11.880 ;
        RECT 20.330 11.870 20.970 11.880 ;
        RECT 27.355 11.870 27.995 11.880 ;
        RECT 35.090 11.870 35.730 11.880 ;
        RECT 42.645 11.870 43.285 11.880 ;
        RECT 50.455 11.870 51.095 11.880 ;
        RECT 57.965 11.870 58.605 11.880 ;
        RECT 65.640 11.870 66.280 11.880 ;
        RECT 73.150 11.870 73.790 11.880 ;
        RECT 10.385 11.640 11.035 11.870 ;
        RECT 14.870 11.640 15.520 11.870 ;
        RECT 20.330 11.640 20.980 11.870 ;
        RECT 27.355 11.640 28.005 11.870 ;
        RECT 35.090 11.640 35.740 11.870 ;
        RECT 42.645 11.640 43.295 11.870 ;
        RECT 50.455 11.640 51.105 11.870 ;
        RECT 57.965 11.640 58.615 11.870 ;
        RECT 65.640 11.640 66.290 11.870 ;
        RECT 73.150 11.640 73.800 11.870 ;
        RECT 10.385 11.620 11.025 11.640 ;
        RECT 14.870 11.620 15.510 11.640 ;
        RECT 20.330 11.620 20.970 11.640 ;
        RECT 27.355 11.620 27.995 11.640 ;
        RECT 35.090 11.620 35.730 11.640 ;
        RECT 42.645 11.620 43.285 11.640 ;
        RECT 50.455 11.620 51.095 11.640 ;
        RECT 57.965 11.620 58.605 11.640 ;
        RECT 65.640 11.620 66.280 11.640 ;
        RECT 73.150 11.620 73.790 11.640 ;
      LAYER via ;
        RECT 10.415 47.045 10.675 47.305 ;
        RECT 10.735 47.045 10.995 47.305 ;
        RECT 14.900 47.045 15.160 47.305 ;
        RECT 15.220 47.045 15.480 47.305 ;
        RECT 20.360 47.045 20.620 47.305 ;
        RECT 20.680 47.045 20.940 47.305 ;
        RECT 27.385 47.045 27.645 47.305 ;
        RECT 27.705 47.045 27.965 47.305 ;
        RECT 35.120 47.045 35.380 47.305 ;
        RECT 35.440 47.045 35.700 47.305 ;
        RECT 42.675 47.045 42.935 47.305 ;
        RECT 42.995 47.045 43.255 47.305 ;
        RECT 50.485 47.045 50.745 47.305 ;
        RECT 50.805 47.045 51.065 47.305 ;
        RECT 57.995 47.045 58.255 47.305 ;
        RECT 58.315 47.045 58.575 47.305 ;
        RECT 65.670 47.045 65.930 47.305 ;
        RECT 65.990 47.045 66.250 47.305 ;
        RECT 73.180 47.045 73.440 47.305 ;
        RECT 73.500 47.045 73.760 47.305 ;
        RECT 10.415 44.650 10.675 44.910 ;
        RECT 10.735 44.650 10.995 44.910 ;
        RECT 14.900 44.650 15.160 44.910 ;
        RECT 15.220 44.650 15.480 44.910 ;
        RECT 20.360 44.650 20.620 44.910 ;
        RECT 20.680 44.650 20.940 44.910 ;
        RECT 27.385 44.650 27.645 44.910 ;
        RECT 27.705 44.650 27.965 44.910 ;
        RECT 35.120 44.650 35.380 44.910 ;
        RECT 35.440 44.650 35.700 44.910 ;
        RECT 42.675 44.650 42.935 44.910 ;
        RECT 42.995 44.650 43.255 44.910 ;
        RECT 50.485 44.650 50.745 44.910 ;
        RECT 50.805 44.650 51.065 44.910 ;
        RECT 57.995 44.650 58.255 44.910 ;
        RECT 58.315 44.650 58.575 44.910 ;
        RECT 65.670 44.650 65.930 44.910 ;
        RECT 65.990 44.650 66.250 44.910 ;
        RECT 73.180 44.650 73.440 44.910 ;
        RECT 73.500 44.650 73.760 44.910 ;
        RECT 10.415 42.300 10.675 42.560 ;
        RECT 10.735 42.300 10.995 42.560 ;
        RECT 14.900 42.300 15.160 42.560 ;
        RECT 15.220 42.300 15.480 42.560 ;
        RECT 20.360 42.300 20.620 42.560 ;
        RECT 20.680 42.300 20.940 42.560 ;
        RECT 27.385 42.300 27.645 42.560 ;
        RECT 27.705 42.300 27.965 42.560 ;
        RECT 35.120 42.300 35.380 42.560 ;
        RECT 35.440 42.300 35.700 42.560 ;
        RECT 42.675 42.300 42.935 42.560 ;
        RECT 42.995 42.300 43.255 42.560 ;
        RECT 50.485 42.300 50.745 42.560 ;
        RECT 50.805 42.300 51.065 42.560 ;
        RECT 57.995 42.300 58.255 42.560 ;
        RECT 58.315 42.300 58.575 42.560 ;
        RECT 65.670 42.300 65.930 42.560 ;
        RECT 65.990 42.300 66.250 42.560 ;
        RECT 73.180 42.300 73.440 42.560 ;
        RECT 73.500 42.300 73.760 42.560 ;
        RECT 10.415 39.940 10.675 40.200 ;
        RECT 10.735 39.940 10.995 40.200 ;
        RECT 14.900 39.940 15.160 40.200 ;
        RECT 15.220 39.940 15.480 40.200 ;
        RECT 20.360 39.940 20.620 40.200 ;
        RECT 20.680 39.940 20.940 40.200 ;
        RECT 27.385 39.940 27.645 40.200 ;
        RECT 27.705 39.940 27.965 40.200 ;
        RECT 35.120 39.940 35.380 40.200 ;
        RECT 35.440 39.940 35.700 40.200 ;
        RECT 42.675 39.940 42.935 40.200 ;
        RECT 42.995 39.940 43.255 40.200 ;
        RECT 50.485 39.940 50.745 40.200 ;
        RECT 50.805 39.940 51.065 40.200 ;
        RECT 57.995 39.940 58.255 40.200 ;
        RECT 58.315 39.940 58.575 40.200 ;
        RECT 65.670 39.940 65.930 40.200 ;
        RECT 65.990 39.940 66.250 40.200 ;
        RECT 73.180 39.940 73.440 40.200 ;
        RECT 73.500 39.940 73.760 40.200 ;
        RECT 10.415 37.585 10.675 37.845 ;
        RECT 10.735 37.585 10.995 37.845 ;
        RECT 14.900 37.585 15.160 37.845 ;
        RECT 15.220 37.585 15.480 37.845 ;
        RECT 20.360 37.585 20.620 37.845 ;
        RECT 20.680 37.585 20.940 37.845 ;
        RECT 27.385 37.585 27.645 37.845 ;
        RECT 27.705 37.585 27.965 37.845 ;
        RECT 35.120 37.585 35.380 37.845 ;
        RECT 35.440 37.585 35.700 37.845 ;
        RECT 42.675 37.585 42.935 37.845 ;
        RECT 42.995 37.585 43.255 37.845 ;
        RECT 50.485 37.585 50.745 37.845 ;
        RECT 50.805 37.585 51.065 37.845 ;
        RECT 57.995 37.585 58.255 37.845 ;
        RECT 58.315 37.585 58.575 37.845 ;
        RECT 65.670 37.585 65.930 37.845 ;
        RECT 65.990 37.585 66.250 37.845 ;
        RECT 73.180 37.585 73.440 37.845 ;
        RECT 73.500 37.585 73.760 37.845 ;
        RECT 10.415 35.225 10.675 35.485 ;
        RECT 10.735 35.225 10.995 35.485 ;
        RECT 14.900 35.225 15.160 35.485 ;
        RECT 15.220 35.225 15.480 35.485 ;
        RECT 20.360 35.225 20.620 35.485 ;
        RECT 20.680 35.225 20.940 35.485 ;
        RECT 27.385 35.225 27.645 35.485 ;
        RECT 27.705 35.225 27.965 35.485 ;
        RECT 35.120 35.225 35.380 35.485 ;
        RECT 35.440 35.225 35.700 35.485 ;
        RECT 42.675 35.225 42.935 35.485 ;
        RECT 42.995 35.225 43.255 35.485 ;
        RECT 50.485 35.225 50.745 35.485 ;
        RECT 50.805 35.225 51.065 35.485 ;
        RECT 57.995 35.225 58.255 35.485 ;
        RECT 58.315 35.225 58.575 35.485 ;
        RECT 65.670 35.225 65.930 35.485 ;
        RECT 65.990 35.225 66.250 35.485 ;
        RECT 73.180 35.225 73.440 35.485 ;
        RECT 73.500 35.225 73.760 35.485 ;
        RECT 10.415 32.860 10.675 33.120 ;
        RECT 10.735 32.860 10.995 33.120 ;
        RECT 14.900 32.860 15.160 33.120 ;
        RECT 15.220 32.860 15.480 33.120 ;
        RECT 20.360 32.860 20.620 33.120 ;
        RECT 20.680 32.860 20.940 33.120 ;
        RECT 27.385 32.860 27.645 33.120 ;
        RECT 27.705 32.860 27.965 33.120 ;
        RECT 35.120 32.860 35.380 33.120 ;
        RECT 35.440 32.860 35.700 33.120 ;
        RECT 42.675 32.860 42.935 33.120 ;
        RECT 42.995 32.860 43.255 33.120 ;
        RECT 50.485 32.860 50.745 33.120 ;
        RECT 50.805 32.860 51.065 33.120 ;
        RECT 57.995 32.860 58.255 33.120 ;
        RECT 58.315 32.860 58.575 33.120 ;
        RECT 65.670 32.860 65.930 33.120 ;
        RECT 65.990 32.860 66.250 33.120 ;
        RECT 73.180 32.860 73.440 33.120 ;
        RECT 73.500 32.860 73.760 33.120 ;
        RECT 10.415 30.505 10.675 30.765 ;
        RECT 10.735 30.505 10.995 30.765 ;
        RECT 14.900 30.505 15.160 30.765 ;
        RECT 15.220 30.505 15.480 30.765 ;
        RECT 20.360 30.505 20.620 30.765 ;
        RECT 20.680 30.505 20.940 30.765 ;
        RECT 27.385 30.505 27.645 30.765 ;
        RECT 27.705 30.505 27.965 30.765 ;
        RECT 35.120 30.505 35.380 30.765 ;
        RECT 35.440 30.505 35.700 30.765 ;
        RECT 42.675 30.505 42.935 30.765 ;
        RECT 42.995 30.505 43.255 30.765 ;
        RECT 50.485 30.505 50.745 30.765 ;
        RECT 50.805 30.505 51.065 30.765 ;
        RECT 57.995 30.505 58.255 30.765 ;
        RECT 58.315 30.505 58.575 30.765 ;
        RECT 65.670 30.505 65.930 30.765 ;
        RECT 65.990 30.505 66.250 30.765 ;
        RECT 73.180 30.505 73.440 30.765 ;
        RECT 73.500 30.505 73.760 30.765 ;
        RECT 10.415 28.145 10.675 28.405 ;
        RECT 10.735 28.145 10.995 28.405 ;
        RECT 14.900 28.145 15.160 28.405 ;
        RECT 15.220 28.145 15.480 28.405 ;
        RECT 20.360 28.145 20.620 28.405 ;
        RECT 20.680 28.145 20.940 28.405 ;
        RECT 27.385 28.145 27.645 28.405 ;
        RECT 27.705 28.145 27.965 28.405 ;
        RECT 35.120 28.145 35.380 28.405 ;
        RECT 35.440 28.145 35.700 28.405 ;
        RECT 42.675 28.145 42.935 28.405 ;
        RECT 42.995 28.145 43.255 28.405 ;
        RECT 50.485 28.145 50.745 28.405 ;
        RECT 50.805 28.145 51.065 28.405 ;
        RECT 57.995 28.145 58.255 28.405 ;
        RECT 58.315 28.145 58.575 28.405 ;
        RECT 65.670 28.145 65.930 28.405 ;
        RECT 65.990 28.145 66.250 28.405 ;
        RECT 73.180 28.145 73.440 28.405 ;
        RECT 73.500 28.145 73.760 28.405 ;
        RECT 10.415 25.780 10.675 26.040 ;
        RECT 10.735 25.780 10.995 26.040 ;
        RECT 14.900 25.780 15.160 26.040 ;
        RECT 15.220 25.780 15.480 26.040 ;
        RECT 20.360 25.780 20.620 26.040 ;
        RECT 20.680 25.780 20.940 26.040 ;
        RECT 27.385 25.780 27.645 26.040 ;
        RECT 27.705 25.780 27.965 26.040 ;
        RECT 35.120 25.780 35.380 26.040 ;
        RECT 35.440 25.780 35.700 26.040 ;
        RECT 42.675 25.780 42.935 26.040 ;
        RECT 42.995 25.780 43.255 26.040 ;
        RECT 50.485 25.780 50.745 26.040 ;
        RECT 50.805 25.780 51.065 26.040 ;
        RECT 57.995 25.780 58.255 26.040 ;
        RECT 58.315 25.780 58.575 26.040 ;
        RECT 65.670 25.780 65.930 26.040 ;
        RECT 65.990 25.780 66.250 26.040 ;
        RECT 73.180 25.780 73.440 26.040 ;
        RECT 73.500 25.780 73.760 26.040 ;
        RECT 10.415 23.420 10.675 23.680 ;
        RECT 10.735 23.420 10.995 23.680 ;
        RECT 14.900 23.420 15.160 23.680 ;
        RECT 15.220 23.420 15.480 23.680 ;
        RECT 20.360 23.420 20.620 23.680 ;
        RECT 20.680 23.420 20.940 23.680 ;
        RECT 27.385 23.420 27.645 23.680 ;
        RECT 27.705 23.420 27.965 23.680 ;
        RECT 35.120 23.420 35.380 23.680 ;
        RECT 35.440 23.420 35.700 23.680 ;
        RECT 42.675 23.420 42.935 23.680 ;
        RECT 42.995 23.420 43.255 23.680 ;
        RECT 50.485 23.420 50.745 23.680 ;
        RECT 50.805 23.420 51.065 23.680 ;
        RECT 57.995 23.420 58.255 23.680 ;
        RECT 58.315 23.420 58.575 23.680 ;
        RECT 65.670 23.420 65.930 23.680 ;
        RECT 65.990 23.420 66.250 23.680 ;
        RECT 73.180 23.420 73.440 23.680 ;
        RECT 73.500 23.420 73.760 23.680 ;
        RECT 10.415 21.065 10.675 21.325 ;
        RECT 10.735 21.065 10.995 21.325 ;
        RECT 14.900 21.065 15.160 21.325 ;
        RECT 15.220 21.065 15.480 21.325 ;
        RECT 20.360 21.065 20.620 21.325 ;
        RECT 20.680 21.065 20.940 21.325 ;
        RECT 27.385 21.065 27.645 21.325 ;
        RECT 27.705 21.065 27.965 21.325 ;
        RECT 35.120 21.065 35.380 21.325 ;
        RECT 35.440 21.065 35.700 21.325 ;
        RECT 42.675 21.065 42.935 21.325 ;
        RECT 42.995 21.065 43.255 21.325 ;
        RECT 50.485 21.065 50.745 21.325 ;
        RECT 50.805 21.065 51.065 21.325 ;
        RECT 57.995 21.065 58.255 21.325 ;
        RECT 58.315 21.065 58.575 21.325 ;
        RECT 65.670 21.065 65.930 21.325 ;
        RECT 65.990 21.065 66.250 21.325 ;
        RECT 73.180 21.065 73.440 21.325 ;
        RECT 73.500 21.065 73.760 21.325 ;
        RECT 10.415 18.705 10.675 18.965 ;
        RECT 10.735 18.705 10.995 18.965 ;
        RECT 14.900 18.705 15.160 18.965 ;
        RECT 15.220 18.705 15.480 18.965 ;
        RECT 20.360 18.705 20.620 18.965 ;
        RECT 20.680 18.705 20.940 18.965 ;
        RECT 27.385 18.705 27.645 18.965 ;
        RECT 27.705 18.705 27.965 18.965 ;
        RECT 35.120 18.705 35.380 18.965 ;
        RECT 35.440 18.705 35.700 18.965 ;
        RECT 42.675 18.705 42.935 18.965 ;
        RECT 42.995 18.705 43.255 18.965 ;
        RECT 50.485 18.705 50.745 18.965 ;
        RECT 50.805 18.705 51.065 18.965 ;
        RECT 57.995 18.705 58.255 18.965 ;
        RECT 58.315 18.705 58.575 18.965 ;
        RECT 65.670 18.705 65.930 18.965 ;
        RECT 65.990 18.705 66.250 18.965 ;
        RECT 73.180 18.705 73.440 18.965 ;
        RECT 73.500 18.705 73.760 18.965 ;
        RECT 10.415 16.340 10.675 16.600 ;
        RECT 10.735 16.340 10.995 16.600 ;
        RECT 14.900 16.340 15.160 16.600 ;
        RECT 15.220 16.340 15.480 16.600 ;
        RECT 20.360 16.340 20.620 16.600 ;
        RECT 20.680 16.340 20.940 16.600 ;
        RECT 27.385 16.340 27.645 16.600 ;
        RECT 27.705 16.340 27.965 16.600 ;
        RECT 35.120 16.340 35.380 16.600 ;
        RECT 35.440 16.340 35.700 16.600 ;
        RECT 42.675 16.340 42.935 16.600 ;
        RECT 42.995 16.340 43.255 16.600 ;
        RECT 50.485 16.340 50.745 16.600 ;
        RECT 50.805 16.340 51.065 16.600 ;
        RECT 57.995 16.340 58.255 16.600 ;
        RECT 58.315 16.340 58.575 16.600 ;
        RECT 65.670 16.340 65.930 16.600 ;
        RECT 65.990 16.340 66.250 16.600 ;
        RECT 73.180 16.340 73.440 16.600 ;
        RECT 73.500 16.340 73.760 16.600 ;
        RECT 10.415 13.980 10.675 14.240 ;
        RECT 10.735 13.980 10.995 14.240 ;
        RECT 14.900 13.980 15.160 14.240 ;
        RECT 15.220 13.980 15.480 14.240 ;
        RECT 20.360 13.980 20.620 14.240 ;
        RECT 20.680 13.980 20.940 14.240 ;
        RECT 27.385 13.980 27.645 14.240 ;
        RECT 27.705 13.980 27.965 14.240 ;
        RECT 35.120 13.980 35.380 14.240 ;
        RECT 35.440 13.980 35.700 14.240 ;
        RECT 42.675 13.980 42.935 14.240 ;
        RECT 42.995 13.980 43.255 14.240 ;
        RECT 50.485 13.980 50.745 14.240 ;
        RECT 50.805 13.980 51.065 14.240 ;
        RECT 57.995 13.980 58.255 14.240 ;
        RECT 58.315 13.980 58.575 14.240 ;
        RECT 65.670 13.980 65.930 14.240 ;
        RECT 65.990 13.980 66.250 14.240 ;
        RECT 73.180 13.980 73.440 14.240 ;
        RECT 73.500 13.980 73.760 14.240 ;
        RECT 10.415 11.620 10.675 11.880 ;
        RECT 10.735 11.620 10.995 11.880 ;
        RECT 14.900 11.620 15.160 11.880 ;
        RECT 15.220 11.620 15.480 11.880 ;
        RECT 20.360 11.620 20.620 11.880 ;
        RECT 20.680 11.620 20.940 11.880 ;
        RECT 27.385 11.620 27.645 11.880 ;
        RECT 27.705 11.620 27.965 11.880 ;
        RECT 35.120 11.620 35.380 11.880 ;
        RECT 35.440 11.620 35.700 11.880 ;
        RECT 42.675 11.620 42.935 11.880 ;
        RECT 42.995 11.620 43.255 11.880 ;
        RECT 50.485 11.620 50.745 11.880 ;
        RECT 50.805 11.620 51.065 11.880 ;
        RECT 57.995 11.620 58.255 11.880 ;
        RECT 58.315 11.620 58.575 11.880 ;
        RECT 65.670 11.620 65.930 11.880 ;
        RECT 65.990 11.620 66.250 11.880 ;
        RECT 73.180 11.620 73.440 11.880 ;
        RECT 73.500 11.620 73.760 11.880 ;
      LAYER met2 ;
        RECT 10.385 11.760 11.035 47.305 ;
        RECT 14.870 11.760 15.520 47.305 ;
        RECT 20.330 11.760 20.980 47.305 ;
        RECT 27.355 11.760 28.005 47.305 ;
        RECT 35.090 11.760 35.740 47.305 ;
        RECT 42.645 11.760 43.295 47.305 ;
        RECT 50.455 11.760 51.105 47.305 ;
        RECT 57.965 11.760 58.615 47.305 ;
        RECT 65.640 11.760 66.290 47.305 ;
        RECT 73.150 11.760 73.800 47.305 ;
        RECT 10.385 11.620 11.025 11.760 ;
        RECT 14.870 11.620 15.510 11.760 ;
        RECT 20.330 11.620 20.970 11.760 ;
        RECT 27.355 11.620 27.995 11.760 ;
        RECT 35.090 11.620 35.730 11.760 ;
        RECT 42.645 11.620 43.285 11.760 ;
        RECT 50.455 11.620 51.095 11.760 ;
        RECT 57.965 11.620 58.605 11.760 ;
        RECT 65.640 11.620 66.280 11.760 ;
        RECT 73.150 11.620 73.790 11.760 ;
    END
  END vref
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 7.305 11.065 7.475 47.410 ;
        RECT 16.920 11.065 17.090 47.410 ;
        RECT 22.645 11.065 22.815 47.410 ;
        RECT 30.380 11.065 30.550 47.410 ;
        RECT 37.935 11.065 38.105 47.410 ;
        RECT 45.745 11.065 45.915 47.410 ;
        RECT 53.255 11.065 53.425 47.410 ;
        RECT 60.930 11.065 61.100 47.410 ;
        RECT 68.440 11.065 68.610 47.410 ;
        RECT 89.200 15.665 90.620 15.835 ;
        RECT 90.450 14.275 90.620 15.665 ;
        RECT 89.200 14.105 90.620 14.275 ;
        RECT 89.595 13.600 89.765 14.105 ;
        RECT 88.965 13.270 90.495 13.600 ;
        RECT 7.305 10.735 91.825 11.065 ;
      LAYER mcon ;
        RECT 89.625 13.350 89.795 13.520 ;
        RECT 7.475 10.815 7.645 10.985 ;
        RECT 7.835 10.815 8.005 10.985 ;
        RECT 8.195 10.815 8.365 10.985 ;
        RECT 8.555 10.815 8.725 10.985 ;
        RECT 8.915 10.815 9.085 10.985 ;
        RECT 9.275 10.815 9.445 10.985 ;
        RECT 9.635 10.815 9.805 10.985 ;
        RECT 9.995 10.815 10.165 10.985 ;
        RECT 10.355 10.815 10.525 10.985 ;
        RECT 10.715 10.815 10.885 10.985 ;
        RECT 11.075 10.815 11.245 10.985 ;
        RECT 11.435 10.815 11.605 10.985 ;
        RECT 11.795 10.815 11.965 10.985 ;
        RECT 12.155 10.815 12.325 10.985 ;
        RECT 12.515 10.815 12.685 10.985 ;
        RECT 12.875 10.815 13.045 10.985 ;
        RECT 13.235 10.815 13.405 10.985 ;
        RECT 13.595 10.815 13.765 10.985 ;
        RECT 13.955 10.815 14.125 10.985 ;
        RECT 14.315 10.815 14.485 10.985 ;
        RECT 14.675 10.815 14.845 10.985 ;
        RECT 15.035 10.815 15.205 10.985 ;
        RECT 15.395 10.815 15.565 10.985 ;
        RECT 15.755 10.815 15.925 10.985 ;
        RECT 16.115 10.815 16.285 10.985 ;
        RECT 16.475 10.815 16.645 10.985 ;
        RECT 16.835 10.815 17.005 10.985 ;
        RECT 17.195 10.815 17.365 10.985 ;
        RECT 17.555 10.815 17.725 10.985 ;
        RECT 17.915 10.815 18.085 10.985 ;
        RECT 18.275 10.815 18.445 10.985 ;
        RECT 18.635 10.815 18.805 10.985 ;
        RECT 18.995 10.815 19.165 10.985 ;
        RECT 19.355 10.815 19.525 10.985 ;
        RECT 19.715 10.815 19.885 10.985 ;
        RECT 20.075 10.815 20.245 10.985 ;
        RECT 20.435 10.815 20.605 10.985 ;
        RECT 20.795 10.815 20.965 10.985 ;
        RECT 21.155 10.815 21.325 10.985 ;
        RECT 21.515 10.815 21.685 10.985 ;
        RECT 21.875 10.815 22.045 10.985 ;
        RECT 22.235 10.815 22.405 10.985 ;
        RECT 22.595 10.815 22.765 10.985 ;
        RECT 22.955 10.815 23.125 10.985 ;
        RECT 23.315 10.815 23.485 10.985 ;
        RECT 23.675 10.815 23.845 10.985 ;
        RECT 24.035 10.815 24.205 10.985 ;
        RECT 24.395 10.815 24.565 10.985 ;
        RECT 24.755 10.815 24.925 10.985 ;
        RECT 25.115 10.815 25.285 10.985 ;
        RECT 25.475 10.815 25.645 10.985 ;
        RECT 25.835 10.815 26.005 10.985 ;
        RECT 26.195 10.815 26.365 10.985 ;
        RECT 26.555 10.815 26.725 10.985 ;
        RECT 26.915 10.815 27.085 10.985 ;
        RECT 27.275 10.815 27.445 10.985 ;
        RECT 27.635 10.815 27.805 10.985 ;
        RECT 27.995 10.815 28.165 10.985 ;
        RECT 28.355 10.815 28.525 10.985 ;
        RECT 28.715 10.815 28.885 10.985 ;
        RECT 29.075 10.815 29.245 10.985 ;
        RECT 29.970 10.815 30.140 10.985 ;
        RECT 30.330 10.815 30.500 10.985 ;
        RECT 30.690 10.815 30.860 10.985 ;
        RECT 31.050 10.815 31.220 10.985 ;
        RECT 31.410 10.815 31.580 10.985 ;
        RECT 31.770 10.815 31.940 10.985 ;
        RECT 32.130 10.815 32.300 10.985 ;
        RECT 32.490 10.815 32.660 10.985 ;
        RECT 32.850 10.815 33.020 10.985 ;
        RECT 33.210 10.815 33.380 10.985 ;
        RECT 33.570 10.815 33.740 10.985 ;
        RECT 33.930 10.815 34.100 10.985 ;
        RECT 34.290 10.815 34.460 10.985 ;
        RECT 34.650 10.815 34.820 10.985 ;
        RECT 35.010 10.815 35.180 10.985 ;
        RECT 35.370 10.815 35.540 10.985 ;
        RECT 35.730 10.815 35.900 10.985 ;
        RECT 36.090 10.815 36.260 10.985 ;
        RECT 36.450 10.815 36.620 10.985 ;
        RECT 37.525 10.815 37.695 10.985 ;
        RECT 37.885 10.815 38.055 10.985 ;
        RECT 38.245 10.815 38.415 10.985 ;
        RECT 38.605 10.815 38.775 10.985 ;
        RECT 38.965 10.815 39.135 10.985 ;
        RECT 39.325 10.815 39.495 10.985 ;
        RECT 39.685 10.815 39.855 10.985 ;
        RECT 40.045 10.815 40.215 10.985 ;
        RECT 40.405 10.815 40.575 10.985 ;
        RECT 40.765 10.815 40.935 10.985 ;
        RECT 41.125 10.815 41.295 10.985 ;
        RECT 41.485 10.815 41.655 10.985 ;
        RECT 41.845 10.815 42.015 10.985 ;
        RECT 42.205 10.815 42.375 10.985 ;
        RECT 42.565 10.815 42.735 10.985 ;
        RECT 42.925 10.815 43.095 10.985 ;
        RECT 43.285 10.815 43.455 10.985 ;
        RECT 43.645 10.815 43.815 10.985 ;
        RECT 44.005 10.815 44.175 10.985 ;
        RECT 45.335 10.815 45.505 10.985 ;
        RECT 45.695 10.815 45.865 10.985 ;
        RECT 46.055 10.815 46.225 10.985 ;
        RECT 46.415 10.815 46.585 10.985 ;
        RECT 46.775 10.815 46.945 10.985 ;
        RECT 47.135 10.815 47.305 10.985 ;
        RECT 47.495 10.815 47.665 10.985 ;
        RECT 47.855 10.815 48.025 10.985 ;
        RECT 48.215 10.815 48.385 10.985 ;
        RECT 48.575 10.815 48.745 10.985 ;
        RECT 48.935 10.815 49.105 10.985 ;
        RECT 49.295 10.815 49.465 10.985 ;
        RECT 49.655 10.815 49.825 10.985 ;
        RECT 50.015 10.815 50.185 10.985 ;
        RECT 50.375 10.815 50.545 10.985 ;
        RECT 50.735 10.815 50.905 10.985 ;
        RECT 51.095 10.815 51.265 10.985 ;
        RECT 51.455 10.815 51.625 10.985 ;
        RECT 51.815 10.815 51.985 10.985 ;
        RECT 52.845 10.815 53.015 10.985 ;
        RECT 53.205 10.815 53.375 10.985 ;
        RECT 53.565 10.815 53.735 10.985 ;
        RECT 53.925 10.815 54.095 10.985 ;
        RECT 54.285 10.815 54.455 10.985 ;
        RECT 54.645 10.815 54.815 10.985 ;
        RECT 55.005 10.815 55.175 10.985 ;
        RECT 55.365 10.815 55.535 10.985 ;
        RECT 55.725 10.815 55.895 10.985 ;
        RECT 56.085 10.815 56.255 10.985 ;
        RECT 56.445 10.815 56.615 10.985 ;
        RECT 56.805 10.815 56.975 10.985 ;
        RECT 57.165 10.815 57.335 10.985 ;
        RECT 57.525 10.815 57.695 10.985 ;
        RECT 57.885 10.815 58.055 10.985 ;
        RECT 58.245 10.815 58.415 10.985 ;
        RECT 58.605 10.815 58.775 10.985 ;
        RECT 58.965 10.815 59.135 10.985 ;
        RECT 59.325 10.815 59.495 10.985 ;
        RECT 60.520 10.815 60.690 10.985 ;
        RECT 60.880 10.815 61.050 10.985 ;
        RECT 61.240 10.815 61.410 10.985 ;
        RECT 61.600 10.815 61.770 10.985 ;
        RECT 61.960 10.815 62.130 10.985 ;
        RECT 62.320 10.815 62.490 10.985 ;
        RECT 62.680 10.815 62.850 10.985 ;
        RECT 63.040 10.815 63.210 10.985 ;
        RECT 63.400 10.815 63.570 10.985 ;
        RECT 63.760 10.815 63.930 10.985 ;
        RECT 64.120 10.815 64.290 10.985 ;
        RECT 64.480 10.815 64.650 10.985 ;
        RECT 64.840 10.815 65.010 10.985 ;
        RECT 65.200 10.815 65.370 10.985 ;
        RECT 65.560 10.815 65.730 10.985 ;
        RECT 65.920 10.815 66.090 10.985 ;
        RECT 66.280 10.815 66.450 10.985 ;
        RECT 66.640 10.815 66.810 10.985 ;
        RECT 67.000 10.815 67.170 10.985 ;
        RECT 68.030 10.815 68.200 10.985 ;
        RECT 68.390 10.815 68.560 10.985 ;
        RECT 68.750 10.815 68.920 10.985 ;
        RECT 69.110 10.815 69.280 10.985 ;
        RECT 69.470 10.815 69.640 10.985 ;
        RECT 69.830 10.815 70.000 10.985 ;
        RECT 70.190 10.815 70.360 10.985 ;
        RECT 70.550 10.815 70.720 10.985 ;
        RECT 70.910 10.815 71.080 10.985 ;
        RECT 71.270 10.815 71.440 10.985 ;
        RECT 71.630 10.815 71.800 10.985 ;
        RECT 71.990 10.815 72.160 10.985 ;
        RECT 72.350 10.815 72.520 10.985 ;
        RECT 72.710 10.815 72.880 10.985 ;
        RECT 73.070 10.815 73.240 10.985 ;
        RECT 73.430 10.815 73.600 10.985 ;
        RECT 73.790 10.815 73.960 10.985 ;
        RECT 74.150 10.815 74.320 10.985 ;
        RECT 74.510 10.815 74.680 10.985 ;
        RECT 75.210 10.815 75.380 10.985 ;
        RECT 75.875 10.815 76.045 10.985 ;
        RECT 76.235 10.815 76.405 10.985 ;
        RECT 76.595 10.815 76.765 10.985 ;
        RECT 76.955 10.815 77.125 10.985 ;
        RECT 77.315 10.815 77.485 10.985 ;
        RECT 77.675 10.815 77.845 10.985 ;
        RECT 78.035 10.815 78.205 10.985 ;
        RECT 78.395 10.815 78.565 10.985 ;
        RECT 78.755 10.815 78.925 10.985 ;
        RECT 79.115 10.815 79.285 10.985 ;
        RECT 79.475 10.815 79.645 10.985 ;
        RECT 79.835 10.815 80.005 10.985 ;
        RECT 80.195 10.815 80.365 10.985 ;
        RECT 80.555 10.815 80.725 10.985 ;
        RECT 80.915 10.815 81.085 10.985 ;
        RECT 81.275 10.815 81.445 10.985 ;
        RECT 81.635 10.815 81.805 10.985 ;
        RECT 81.995 10.815 82.165 10.985 ;
        RECT 82.355 10.815 82.525 10.985 ;
        RECT 82.715 10.815 82.885 10.985 ;
        RECT 83.075 10.815 83.245 10.985 ;
        RECT 83.435 10.815 83.605 10.985 ;
        RECT 83.795 10.815 83.965 10.985 ;
        RECT 84.155 10.815 84.325 10.985 ;
        RECT 84.855 10.815 85.025 10.985 ;
        RECT 85.215 10.815 85.385 10.985 ;
        RECT 85.575 10.815 85.745 10.985 ;
        RECT 85.935 10.815 86.105 10.985 ;
        RECT 86.295 10.815 86.465 10.985 ;
        RECT 86.655 10.815 86.825 10.985 ;
        RECT 87.015 10.815 87.185 10.985 ;
        RECT 87.375 10.815 87.545 10.985 ;
        RECT 87.735 10.815 87.905 10.985 ;
        RECT 88.095 10.815 88.265 10.985 ;
        RECT 88.455 10.815 88.625 10.985 ;
        RECT 88.815 10.815 88.985 10.985 ;
        RECT 89.175 10.815 89.345 10.985 ;
        RECT 89.535 10.815 89.705 10.985 ;
        RECT 89.895 10.815 90.065 10.985 ;
        RECT 90.255 10.815 90.425 10.985 ;
        RECT 90.615 10.815 90.785 10.985 ;
        RECT 90.975 10.815 91.145 10.985 ;
        RECT 91.335 10.815 91.505 10.985 ;
      LAYER met1 ;
        RECT 89.565 13.290 89.855 13.580 ;
        RECT 89.640 11.280 89.780 13.290 ;
        RECT 7.180 9.550 92.090 11.280 ;
        RECT 7.180 8.765 8.920 9.550 ;
        RECT 0.000 8.395 8.920 8.765 ;
        RECT 7.180 7.885 8.920 8.395 ;
        RECT 0.000 7.515 8.920 7.885 ;
        RECT 90.350 8.765 92.090 9.550 ;
        RECT 90.350 8.395 101.280 8.765 ;
        RECT 90.350 7.885 92.090 8.395 ;
        RECT 90.350 7.515 101.280 7.885 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 0.000 60.965 101.280 61.135 ;
        RECT 0.000 56.895 101.280 57.065 ;
        RECT 0.000 52.825 3.840 52.995 ;
        RECT 97.440 52.825 101.280 52.995 ;
        RECT 0.000 48.755 3.840 48.925 ;
        RECT 7.490 48.650 10.200 48.820 ;
        RECT 11.975 48.650 14.685 48.820 ;
        RECT 17.435 48.650 20.145 48.820 ;
        RECT 24.460 48.650 27.170 48.820 ;
        RECT 32.195 48.650 34.905 48.820 ;
        RECT 39.750 48.650 42.460 48.820 ;
        RECT 47.560 48.650 50.270 48.820 ;
        RECT 55.070 48.650 57.780 48.820 ;
        RECT 62.745 48.650 65.455 48.820 ;
        RECT 70.255 48.650 72.965 48.820 ;
        RECT 97.440 48.755 101.280 48.925 ;
        RECT 7.965 48.545 9.510 48.650 ;
        RECT 12.480 48.525 13.890 48.650 ;
        RECT 17.980 48.525 19.350 48.650 ;
        RECT 25.005 48.500 26.375 48.650 ;
        RECT 32.740 48.500 34.110 48.650 ;
        RECT 40.295 48.500 41.665 48.650 ;
        RECT 48.105 48.500 49.475 48.650 ;
        RECT 55.615 48.500 56.985 48.650 ;
        RECT 63.290 48.500 64.660 48.650 ;
        RECT 70.800 48.500 72.170 48.650 ;
        RECT 11.525 46.295 11.855 46.625 ;
        RECT 16.010 46.295 16.340 46.625 ;
        RECT 21.470 46.295 21.800 46.625 ;
        RECT 28.495 46.295 28.825 46.625 ;
        RECT 36.230 46.295 36.560 46.625 ;
        RECT 43.785 46.295 44.115 46.625 ;
        RECT 51.595 46.295 51.925 46.625 ;
        RECT 59.105 46.295 59.435 46.625 ;
        RECT 66.780 46.295 67.110 46.625 ;
        RECT 74.290 46.295 74.620 46.625 ;
        RECT 8.045 45.890 11.310 46.060 ;
        RECT 12.530 45.890 15.795 46.060 ;
        RECT 17.645 45.890 21.255 46.060 ;
        RECT 23.360 45.890 28.280 46.060 ;
        RECT 31.095 45.890 36.015 46.060 ;
        RECT 38.650 45.890 43.570 46.060 ;
        RECT 46.460 45.890 51.380 46.060 ;
        RECT 53.970 45.890 58.890 46.060 ;
        RECT 61.645 45.890 66.565 46.060 ;
        RECT 69.155 45.890 74.075 46.060 ;
        RECT 77.980 45.995 79.400 46.165 ;
        RECT 83.530 45.995 84.950 46.165 ;
        RECT 8.095 45.885 9.345 45.890 ;
        RECT 12.580 45.885 13.830 45.890 ;
        RECT 18.040 45.885 19.290 45.890 ;
        RECT 25.065 45.885 26.315 45.890 ;
        RECT 32.800 45.885 34.050 45.890 ;
        RECT 40.355 45.885 41.605 45.890 ;
        RECT 48.165 45.885 49.415 45.890 ;
        RECT 55.675 45.885 56.925 45.890 ;
        RECT 63.350 45.885 64.600 45.890 ;
        RECT 70.860 45.885 72.110 45.890 ;
        RECT 11.525 45.245 11.855 45.575 ;
        RECT 16.010 45.245 16.340 45.575 ;
        RECT 21.470 45.245 21.800 45.575 ;
        RECT 28.495 45.245 28.825 45.575 ;
        RECT 36.230 45.245 36.560 45.575 ;
        RECT 43.785 45.245 44.115 45.575 ;
        RECT 51.595 45.245 51.925 45.575 ;
        RECT 59.105 45.245 59.435 45.575 ;
        RECT 66.780 45.245 67.110 45.575 ;
        RECT 74.290 45.245 74.620 45.575 ;
        RECT 0.000 44.685 3.840 44.855 ;
        RECT 79.230 44.605 79.400 45.995 ;
        RECT 83.065 45.385 83.395 45.465 ;
        RECT 83.065 45.215 84.540 45.385 ;
        RECT 83.065 45.135 83.395 45.215 ;
        RECT 84.780 44.605 84.950 45.995 ;
        RECT 97.440 44.685 101.280 44.855 ;
        RECT 77.980 44.435 79.400 44.605 ;
        RECT 83.530 44.435 84.950 44.605 ;
        RECT 11.525 44.020 11.855 44.350 ;
        RECT 16.010 44.020 16.340 44.350 ;
        RECT 21.470 44.020 21.800 44.350 ;
        RECT 28.495 44.020 28.825 44.350 ;
        RECT 36.230 44.020 36.560 44.350 ;
        RECT 43.785 44.020 44.115 44.350 ;
        RECT 51.595 44.020 51.925 44.350 ;
        RECT 59.105 44.020 59.435 44.350 ;
        RECT 66.780 44.020 67.110 44.350 ;
        RECT 74.290 44.020 74.620 44.350 ;
        RECT 78.375 43.930 78.545 44.435 ;
        RECT 83.925 43.930 84.095 44.435 ;
        RECT 8.045 43.530 11.310 43.700 ;
        RECT 12.530 43.530 15.795 43.700 ;
        RECT 17.645 43.530 21.255 43.700 ;
        RECT 23.360 43.530 28.280 43.700 ;
        RECT 31.095 43.530 36.015 43.700 ;
        RECT 38.650 43.530 43.570 43.700 ;
        RECT 46.460 43.530 51.380 43.700 ;
        RECT 53.970 43.530 58.890 43.700 ;
        RECT 61.645 43.530 66.565 43.700 ;
        RECT 69.155 43.530 74.075 43.700 ;
        RECT 77.745 43.600 79.275 43.930 ;
        RECT 83.295 43.600 84.825 43.930 ;
        RECT 8.095 43.525 9.345 43.530 ;
        RECT 12.580 43.525 13.830 43.530 ;
        RECT 18.040 43.525 19.290 43.530 ;
        RECT 25.065 43.525 26.315 43.530 ;
        RECT 32.800 43.525 34.050 43.530 ;
        RECT 40.355 43.525 41.605 43.530 ;
        RECT 48.165 43.525 49.415 43.530 ;
        RECT 55.675 43.525 56.925 43.530 ;
        RECT 63.350 43.525 64.600 43.530 ;
        RECT 70.860 43.525 72.110 43.530 ;
        RECT 11.525 42.910 11.855 43.240 ;
        RECT 16.010 42.910 16.340 43.240 ;
        RECT 21.470 42.910 21.800 43.240 ;
        RECT 28.495 42.910 28.825 43.240 ;
        RECT 36.230 42.910 36.560 43.240 ;
        RECT 43.785 42.910 44.115 43.240 ;
        RECT 51.595 42.910 51.925 43.240 ;
        RECT 59.105 42.910 59.435 43.240 ;
        RECT 66.780 42.910 67.110 43.240 ;
        RECT 74.290 42.910 74.620 43.240 ;
        RECT 11.525 41.725 11.855 42.055 ;
        RECT 16.010 41.725 16.340 42.055 ;
        RECT 21.470 41.725 21.800 42.055 ;
        RECT 28.495 41.725 28.825 42.055 ;
        RECT 36.230 41.725 36.560 42.055 ;
        RECT 43.785 41.725 44.115 42.055 ;
        RECT 51.595 41.725 51.925 42.055 ;
        RECT 59.105 41.725 59.435 42.055 ;
        RECT 66.780 41.725 67.110 42.055 ;
        RECT 74.290 41.725 74.620 42.055 ;
        RECT 8.045 41.170 11.310 41.340 ;
        RECT 12.530 41.170 15.795 41.340 ;
        RECT 17.645 41.170 21.255 41.340 ;
        RECT 23.360 41.170 28.280 41.340 ;
        RECT 31.095 41.170 36.015 41.340 ;
        RECT 38.650 41.170 43.570 41.340 ;
        RECT 46.460 41.170 51.380 41.340 ;
        RECT 53.970 41.170 58.890 41.340 ;
        RECT 61.645 41.170 66.565 41.340 ;
        RECT 69.155 41.170 74.075 41.340 ;
        RECT 77.980 40.940 79.400 41.110 ;
        RECT 83.530 40.940 84.950 41.110 ;
        RECT 0.000 40.615 3.840 40.785 ;
        RECT 11.525 40.545 11.855 40.875 ;
        RECT 16.010 40.545 16.340 40.875 ;
        RECT 21.470 40.545 21.800 40.875 ;
        RECT 28.495 40.545 28.825 40.875 ;
        RECT 36.230 40.545 36.560 40.875 ;
        RECT 43.785 40.545 44.115 40.875 ;
        RECT 51.595 40.545 51.925 40.875 ;
        RECT 59.105 40.545 59.435 40.875 ;
        RECT 66.780 40.545 67.110 40.875 ;
        RECT 74.290 40.545 74.620 40.875 ;
        RECT 77.515 40.330 77.845 40.410 ;
        RECT 77.515 40.160 78.990 40.330 ;
        RECT 77.515 40.080 77.845 40.160 ;
        RECT 11.525 39.305 11.855 39.635 ;
        RECT 16.010 39.305 16.340 39.635 ;
        RECT 21.470 39.305 21.800 39.635 ;
        RECT 28.495 39.305 28.825 39.635 ;
        RECT 36.230 39.305 36.560 39.635 ;
        RECT 43.785 39.305 44.115 39.635 ;
        RECT 51.595 39.305 51.925 39.635 ;
        RECT 59.105 39.305 59.435 39.635 ;
        RECT 66.780 39.305 67.110 39.635 ;
        RECT 74.290 39.305 74.620 39.635 ;
        RECT 79.230 39.550 79.400 40.940 ;
        RECT 83.065 40.330 83.395 40.410 ;
        RECT 83.065 40.160 84.540 40.330 ;
        RECT 83.065 40.080 83.395 40.160 ;
        RECT 84.780 39.550 84.950 40.940 ;
        RECT 97.440 40.615 101.280 40.785 ;
        RECT 77.980 39.380 79.400 39.550 ;
        RECT 83.530 39.380 84.950 39.550 ;
        RECT 8.045 38.810 11.310 38.980 ;
        RECT 12.530 38.810 15.795 38.980 ;
        RECT 17.645 38.810 21.255 38.980 ;
        RECT 23.360 38.810 28.280 38.980 ;
        RECT 31.095 38.810 36.015 38.980 ;
        RECT 38.650 38.810 43.570 38.980 ;
        RECT 46.460 38.810 51.380 38.980 ;
        RECT 53.970 38.810 58.890 38.980 ;
        RECT 61.645 38.810 66.565 38.980 ;
        RECT 69.155 38.810 74.075 38.980 ;
        RECT 78.375 38.875 78.545 39.380 ;
        RECT 83.925 38.875 84.095 39.380 ;
        RECT 11.525 38.255 11.855 38.585 ;
        RECT 16.010 38.255 16.340 38.585 ;
        RECT 21.470 38.255 21.800 38.585 ;
        RECT 28.495 38.255 28.825 38.585 ;
        RECT 36.230 38.255 36.560 38.585 ;
        RECT 43.785 38.255 44.115 38.585 ;
        RECT 51.595 38.255 51.925 38.585 ;
        RECT 59.105 38.255 59.435 38.585 ;
        RECT 66.780 38.255 67.110 38.585 ;
        RECT 74.290 38.255 74.620 38.585 ;
        RECT 77.745 38.545 79.275 38.875 ;
        RECT 83.295 38.545 84.825 38.875 ;
        RECT 11.525 37.030 11.855 37.360 ;
        RECT 16.010 37.030 16.340 37.360 ;
        RECT 21.470 37.030 21.800 37.360 ;
        RECT 28.495 37.030 28.825 37.360 ;
        RECT 36.230 37.030 36.560 37.360 ;
        RECT 43.785 37.030 44.115 37.360 ;
        RECT 51.595 37.030 51.925 37.360 ;
        RECT 59.105 37.030 59.435 37.360 ;
        RECT 66.780 37.030 67.110 37.360 ;
        RECT 74.290 37.030 74.620 37.360 ;
        RECT 0.000 36.545 3.840 36.715 ;
        RECT 8.045 36.450 11.310 36.620 ;
        RECT 12.530 36.450 15.795 36.620 ;
        RECT 17.645 36.450 21.255 36.620 ;
        RECT 23.360 36.450 28.280 36.620 ;
        RECT 31.095 36.450 36.015 36.620 ;
        RECT 38.650 36.450 43.570 36.620 ;
        RECT 46.460 36.450 51.380 36.620 ;
        RECT 53.970 36.450 58.890 36.620 ;
        RECT 61.645 36.450 66.565 36.620 ;
        RECT 69.155 36.450 74.075 36.620 ;
        RECT 97.440 36.545 101.280 36.715 ;
        RECT 11.525 35.920 11.855 36.250 ;
        RECT 16.010 35.920 16.340 36.250 ;
        RECT 21.470 35.920 21.800 36.250 ;
        RECT 28.495 35.920 28.825 36.250 ;
        RECT 36.230 35.920 36.560 36.250 ;
        RECT 43.785 35.920 44.115 36.250 ;
        RECT 51.595 35.920 51.925 36.250 ;
        RECT 59.105 35.920 59.435 36.250 ;
        RECT 66.780 35.920 67.110 36.250 ;
        RECT 74.290 35.920 74.620 36.250 ;
        RECT 77.980 35.885 79.400 36.055 ;
        RECT 83.530 35.885 84.950 36.055 ;
        RECT 77.515 35.275 77.845 35.355 ;
        RECT 77.515 35.105 78.990 35.275 ;
        RECT 11.525 34.735 11.855 35.065 ;
        RECT 16.010 34.735 16.340 35.065 ;
        RECT 21.470 34.735 21.800 35.065 ;
        RECT 28.495 34.735 28.825 35.065 ;
        RECT 36.230 34.735 36.560 35.065 ;
        RECT 43.785 34.735 44.115 35.065 ;
        RECT 51.595 34.735 51.925 35.065 ;
        RECT 59.105 34.735 59.435 35.065 ;
        RECT 66.780 34.735 67.110 35.065 ;
        RECT 74.290 34.735 74.620 35.065 ;
        RECT 77.515 35.025 77.845 35.105 ;
        RECT 79.230 34.495 79.400 35.885 ;
        RECT 83.065 35.275 83.395 35.355 ;
        RECT 83.065 35.105 84.540 35.275 ;
        RECT 83.065 35.025 83.395 35.105 ;
        RECT 84.780 34.495 84.950 35.885 ;
        RECT 77.980 34.325 79.400 34.495 ;
        RECT 83.530 34.325 84.950 34.495 ;
        RECT 8.045 34.090 11.310 34.260 ;
        RECT 12.530 34.090 15.795 34.260 ;
        RECT 17.645 34.090 21.255 34.260 ;
        RECT 23.360 34.090 28.280 34.260 ;
        RECT 31.095 34.090 36.015 34.260 ;
        RECT 38.650 34.090 43.570 34.260 ;
        RECT 46.460 34.090 51.380 34.260 ;
        RECT 53.970 34.090 58.890 34.260 ;
        RECT 61.645 34.090 66.565 34.260 ;
        RECT 69.155 34.090 74.075 34.260 ;
        RECT 11.525 33.555 11.855 33.885 ;
        RECT 16.010 33.555 16.340 33.885 ;
        RECT 21.470 33.555 21.800 33.885 ;
        RECT 28.495 33.555 28.825 33.885 ;
        RECT 36.230 33.555 36.560 33.885 ;
        RECT 43.785 33.555 44.115 33.885 ;
        RECT 51.595 33.555 51.925 33.885 ;
        RECT 59.105 33.555 59.435 33.885 ;
        RECT 66.780 33.555 67.110 33.885 ;
        RECT 74.290 33.555 74.620 33.885 ;
        RECT 78.375 33.820 78.545 34.325 ;
        RECT 83.925 33.820 84.095 34.325 ;
        RECT 77.745 33.490 79.275 33.820 ;
        RECT 83.295 33.490 84.825 33.820 ;
        RECT 0.000 32.475 3.840 32.645 ;
        RECT 11.525 32.280 11.855 32.610 ;
        RECT 16.010 32.280 16.340 32.610 ;
        RECT 21.470 32.280 21.800 32.610 ;
        RECT 28.495 32.280 28.825 32.610 ;
        RECT 36.230 32.280 36.560 32.610 ;
        RECT 43.785 32.280 44.115 32.610 ;
        RECT 51.595 32.280 51.925 32.610 ;
        RECT 59.105 32.280 59.435 32.610 ;
        RECT 66.780 32.280 67.110 32.610 ;
        RECT 74.290 32.280 74.620 32.610 ;
        RECT 97.440 32.475 101.280 32.645 ;
        RECT 8.045 31.730 11.310 31.900 ;
        RECT 12.530 31.730 15.795 31.900 ;
        RECT 17.645 31.730 21.255 31.900 ;
        RECT 23.360 31.730 28.280 31.900 ;
        RECT 31.095 31.730 36.015 31.900 ;
        RECT 38.650 31.730 43.570 31.900 ;
        RECT 46.460 31.730 51.380 31.900 ;
        RECT 53.970 31.730 58.890 31.900 ;
        RECT 61.645 31.730 66.565 31.900 ;
        RECT 69.155 31.730 74.075 31.900 ;
        RECT 11.525 31.230 11.855 31.560 ;
        RECT 16.010 31.230 16.340 31.560 ;
        RECT 21.470 31.230 21.800 31.560 ;
        RECT 28.495 31.230 28.825 31.560 ;
        RECT 36.230 31.230 36.560 31.560 ;
        RECT 43.785 31.230 44.115 31.560 ;
        RECT 51.595 31.230 51.925 31.560 ;
        RECT 59.105 31.230 59.435 31.560 ;
        RECT 66.780 31.230 67.110 31.560 ;
        RECT 74.290 31.230 74.620 31.560 ;
        RECT 77.980 30.830 79.400 31.000 ;
        RECT 83.530 30.830 84.950 31.000 ;
        RECT 11.525 30.005 11.855 30.335 ;
        RECT 16.010 30.005 16.340 30.335 ;
        RECT 21.470 30.005 21.800 30.335 ;
        RECT 28.495 30.005 28.825 30.335 ;
        RECT 36.230 30.005 36.560 30.335 ;
        RECT 43.785 30.005 44.115 30.335 ;
        RECT 51.595 30.005 51.925 30.335 ;
        RECT 59.105 30.005 59.435 30.335 ;
        RECT 66.780 30.005 67.110 30.335 ;
        RECT 74.290 30.005 74.620 30.335 ;
        RECT 77.515 30.220 77.845 30.300 ;
        RECT 77.515 30.050 78.990 30.220 ;
        RECT 77.515 29.970 77.845 30.050 ;
        RECT 8.045 29.370 11.310 29.540 ;
        RECT 12.530 29.370 15.795 29.540 ;
        RECT 17.645 29.370 21.255 29.540 ;
        RECT 23.360 29.370 28.280 29.540 ;
        RECT 31.095 29.370 36.015 29.540 ;
        RECT 38.650 29.370 43.570 29.540 ;
        RECT 46.460 29.370 51.380 29.540 ;
        RECT 53.970 29.370 58.890 29.540 ;
        RECT 61.645 29.370 66.565 29.540 ;
        RECT 69.155 29.370 74.075 29.540 ;
        RECT 79.230 29.440 79.400 30.830 ;
        RECT 83.065 30.220 83.395 30.300 ;
        RECT 83.065 30.050 84.540 30.220 ;
        RECT 83.065 29.970 83.395 30.050 ;
        RECT 84.780 29.440 84.950 30.830 ;
        RECT 77.980 29.270 79.400 29.440 ;
        RECT 83.530 29.270 84.950 29.440 ;
        RECT 11.525 28.895 11.855 29.225 ;
        RECT 16.010 28.895 16.340 29.225 ;
        RECT 21.470 28.895 21.800 29.225 ;
        RECT 28.495 28.895 28.825 29.225 ;
        RECT 36.230 28.895 36.560 29.225 ;
        RECT 43.785 28.895 44.115 29.225 ;
        RECT 51.595 28.895 51.925 29.225 ;
        RECT 59.105 28.895 59.435 29.225 ;
        RECT 66.780 28.895 67.110 29.225 ;
        RECT 74.290 28.895 74.620 29.225 ;
        RECT 78.375 28.765 78.545 29.270 ;
        RECT 83.925 28.765 84.095 29.270 ;
        RECT 0.000 28.405 3.840 28.575 ;
        RECT 77.745 28.435 79.275 28.765 ;
        RECT 83.295 28.435 84.825 28.765 ;
        RECT 97.440 28.405 101.280 28.575 ;
        RECT 11.525 27.710 11.855 28.040 ;
        RECT 16.010 27.710 16.340 28.040 ;
        RECT 21.470 27.710 21.800 28.040 ;
        RECT 28.495 27.710 28.825 28.040 ;
        RECT 36.230 27.710 36.560 28.040 ;
        RECT 43.785 27.710 44.115 28.040 ;
        RECT 51.595 27.710 51.925 28.040 ;
        RECT 59.105 27.710 59.435 28.040 ;
        RECT 66.780 27.710 67.110 28.040 ;
        RECT 74.290 27.710 74.620 28.040 ;
        RECT 8.045 27.010 11.310 27.180 ;
        RECT 12.530 27.010 15.795 27.180 ;
        RECT 17.645 27.010 21.255 27.180 ;
        RECT 23.360 27.010 28.280 27.180 ;
        RECT 31.095 27.010 36.015 27.180 ;
        RECT 38.650 27.010 43.570 27.180 ;
        RECT 46.460 27.010 51.380 27.180 ;
        RECT 53.970 27.010 58.890 27.180 ;
        RECT 61.645 27.010 66.565 27.180 ;
        RECT 69.155 27.010 74.075 27.180 ;
        RECT 11.525 26.530 11.855 26.860 ;
        RECT 16.010 26.530 16.340 26.860 ;
        RECT 21.470 26.530 21.800 26.860 ;
        RECT 28.495 26.530 28.825 26.860 ;
        RECT 36.230 26.530 36.560 26.860 ;
        RECT 43.785 26.530 44.115 26.860 ;
        RECT 51.595 26.530 51.925 26.860 ;
        RECT 59.105 26.530 59.435 26.860 ;
        RECT 66.780 26.530 67.110 26.860 ;
        RECT 74.290 26.530 74.620 26.860 ;
        RECT 77.980 25.775 79.400 25.945 ;
        RECT 83.530 25.775 84.950 25.945 ;
        RECT 11.525 25.175 11.855 25.505 ;
        RECT 16.010 25.175 16.340 25.505 ;
        RECT 21.470 25.175 21.800 25.505 ;
        RECT 28.495 25.175 28.825 25.505 ;
        RECT 36.230 25.175 36.560 25.505 ;
        RECT 43.785 25.175 44.115 25.505 ;
        RECT 51.595 25.175 51.925 25.505 ;
        RECT 59.105 25.175 59.435 25.505 ;
        RECT 66.780 25.175 67.110 25.505 ;
        RECT 74.290 25.175 74.620 25.505 ;
        RECT 77.515 25.165 77.845 25.245 ;
        RECT 77.515 24.995 78.990 25.165 ;
        RECT 77.515 24.915 77.845 24.995 ;
        RECT 8.045 24.650 11.310 24.820 ;
        RECT 12.530 24.650 15.795 24.820 ;
        RECT 17.645 24.650 21.255 24.820 ;
        RECT 23.360 24.650 28.280 24.820 ;
        RECT 31.095 24.650 36.015 24.820 ;
        RECT 38.650 24.650 43.570 24.820 ;
        RECT 46.460 24.650 51.380 24.820 ;
        RECT 53.970 24.650 58.890 24.820 ;
        RECT 61.645 24.650 66.565 24.820 ;
        RECT 69.155 24.650 74.075 24.820 ;
        RECT 0.000 24.335 3.840 24.505 ;
        RECT 11.525 24.125 11.855 24.455 ;
        RECT 16.010 24.125 16.340 24.455 ;
        RECT 21.470 24.125 21.800 24.455 ;
        RECT 28.495 24.125 28.825 24.455 ;
        RECT 36.230 24.125 36.560 24.455 ;
        RECT 43.785 24.125 44.115 24.455 ;
        RECT 51.595 24.125 51.925 24.455 ;
        RECT 59.105 24.125 59.435 24.455 ;
        RECT 66.780 24.125 67.110 24.455 ;
        RECT 74.290 24.125 74.620 24.455 ;
        RECT 79.230 24.385 79.400 25.775 ;
        RECT 83.065 25.165 83.395 25.245 ;
        RECT 83.065 24.995 84.540 25.165 ;
        RECT 83.065 24.915 83.395 24.995 ;
        RECT 84.780 24.385 84.950 25.775 ;
        RECT 77.980 24.215 79.400 24.385 ;
        RECT 83.530 24.215 84.950 24.385 ;
        RECT 97.440 24.335 101.280 24.505 ;
        RECT 78.375 23.710 78.545 24.215 ;
        RECT 83.925 23.710 84.095 24.215 ;
        RECT 77.745 23.380 79.275 23.710 ;
        RECT 83.295 23.380 84.825 23.710 ;
        RECT 11.525 22.900 11.855 23.230 ;
        RECT 16.010 22.900 16.340 23.230 ;
        RECT 21.470 22.900 21.800 23.230 ;
        RECT 28.495 22.900 28.825 23.230 ;
        RECT 36.230 22.900 36.560 23.230 ;
        RECT 43.785 22.900 44.115 23.230 ;
        RECT 51.595 22.900 51.925 23.230 ;
        RECT 59.105 22.900 59.435 23.230 ;
        RECT 66.780 22.900 67.110 23.230 ;
        RECT 74.290 22.900 74.620 23.230 ;
        RECT 8.045 22.290 11.310 22.460 ;
        RECT 12.530 22.290 15.795 22.460 ;
        RECT 17.645 22.290 21.255 22.460 ;
        RECT 23.360 22.290 28.280 22.460 ;
        RECT 31.095 22.290 36.015 22.460 ;
        RECT 38.650 22.290 43.570 22.460 ;
        RECT 46.460 22.290 51.380 22.460 ;
        RECT 53.970 22.290 58.890 22.460 ;
        RECT 61.645 22.290 66.565 22.460 ;
        RECT 69.155 22.290 74.075 22.460 ;
        RECT 11.525 21.790 11.855 22.120 ;
        RECT 16.010 21.790 16.340 22.120 ;
        RECT 21.470 21.790 21.800 22.120 ;
        RECT 28.495 21.790 28.825 22.120 ;
        RECT 36.230 21.790 36.560 22.120 ;
        RECT 43.785 21.790 44.115 22.120 ;
        RECT 51.595 21.790 51.925 22.120 ;
        RECT 59.105 21.790 59.435 22.120 ;
        RECT 66.780 21.790 67.110 22.120 ;
        RECT 74.290 21.790 74.620 22.120 ;
        RECT 11.525 20.605 11.855 20.935 ;
        RECT 16.010 20.605 16.340 20.935 ;
        RECT 21.470 20.605 21.800 20.935 ;
        RECT 28.495 20.605 28.825 20.935 ;
        RECT 36.230 20.605 36.560 20.935 ;
        RECT 43.785 20.605 44.115 20.935 ;
        RECT 51.595 20.605 51.925 20.935 ;
        RECT 59.105 20.605 59.435 20.935 ;
        RECT 66.780 20.605 67.110 20.935 ;
        RECT 74.290 20.605 74.620 20.935 ;
        RECT 77.980 20.720 79.400 20.890 ;
        RECT 83.530 20.720 84.950 20.890 ;
        RECT 89.200 20.720 90.620 20.890 ;
        RECT 0.000 20.265 3.840 20.435 ;
        RECT 77.515 20.110 77.845 20.190 ;
        RECT 8.045 19.930 11.310 20.100 ;
        RECT 12.530 19.930 15.795 20.100 ;
        RECT 17.645 19.930 21.255 20.100 ;
        RECT 23.360 19.930 28.280 20.100 ;
        RECT 31.095 19.930 36.015 20.100 ;
        RECT 38.650 19.930 43.570 20.100 ;
        RECT 46.460 19.930 51.380 20.100 ;
        RECT 53.970 19.930 58.890 20.100 ;
        RECT 61.645 19.930 66.565 20.100 ;
        RECT 69.155 19.930 74.075 20.100 ;
        RECT 77.515 19.940 78.990 20.110 ;
        RECT 77.515 19.860 77.845 19.940 ;
        RECT 11.525 19.425 11.855 19.755 ;
        RECT 16.010 19.425 16.340 19.755 ;
        RECT 21.470 19.425 21.800 19.755 ;
        RECT 28.495 19.425 28.825 19.755 ;
        RECT 36.230 19.425 36.560 19.755 ;
        RECT 43.785 19.425 44.115 19.755 ;
        RECT 51.595 19.425 51.925 19.755 ;
        RECT 59.105 19.425 59.435 19.755 ;
        RECT 66.780 19.425 67.110 19.755 ;
        RECT 74.290 19.425 74.620 19.755 ;
        RECT 79.230 19.330 79.400 20.720 ;
        RECT 83.065 20.110 83.395 20.190 ;
        RECT 83.065 19.940 84.540 20.110 ;
        RECT 83.065 19.860 83.395 19.940 ;
        RECT 84.780 19.330 84.950 20.720 ;
        RECT 88.735 20.110 89.065 20.190 ;
        RECT 88.735 19.940 90.210 20.110 ;
        RECT 88.735 19.860 89.065 19.940 ;
        RECT 90.450 19.330 90.620 20.720 ;
        RECT 97.440 20.265 101.280 20.435 ;
        RECT 77.980 19.160 79.400 19.330 ;
        RECT 83.530 19.160 84.950 19.330 ;
        RECT 89.200 19.160 90.620 19.330 ;
        RECT 78.375 18.655 78.545 19.160 ;
        RECT 83.925 18.655 84.095 19.160 ;
        RECT 89.595 18.655 89.765 19.160 ;
        RECT 11.525 18.045 11.855 18.375 ;
        RECT 16.010 18.045 16.340 18.375 ;
        RECT 21.470 18.045 21.800 18.375 ;
        RECT 28.495 18.045 28.825 18.375 ;
        RECT 36.230 18.045 36.560 18.375 ;
        RECT 43.785 18.045 44.115 18.375 ;
        RECT 51.595 18.045 51.925 18.375 ;
        RECT 59.105 18.045 59.435 18.375 ;
        RECT 66.780 18.045 67.110 18.375 ;
        RECT 74.290 18.045 74.620 18.375 ;
        RECT 77.745 18.325 79.275 18.655 ;
        RECT 83.295 18.325 84.825 18.655 ;
        RECT 88.965 18.325 90.495 18.655 ;
        RECT 8.045 17.570 11.310 17.740 ;
        RECT 12.530 17.570 15.795 17.740 ;
        RECT 17.645 17.570 21.255 17.740 ;
        RECT 23.360 17.570 28.280 17.740 ;
        RECT 31.095 17.570 36.015 17.740 ;
        RECT 38.650 17.570 43.570 17.740 ;
        RECT 46.460 17.570 51.380 17.740 ;
        RECT 53.970 17.570 58.890 17.740 ;
        RECT 61.645 17.570 66.565 17.740 ;
        RECT 69.155 17.570 74.075 17.740 ;
        RECT 11.525 16.995 11.855 17.325 ;
        RECT 16.010 16.995 16.340 17.325 ;
        RECT 21.470 16.995 21.800 17.325 ;
        RECT 28.495 16.995 28.825 17.325 ;
        RECT 36.230 16.995 36.560 17.325 ;
        RECT 43.785 16.995 44.115 17.325 ;
        RECT 51.595 16.995 51.925 17.325 ;
        RECT 59.105 16.995 59.435 17.325 ;
        RECT 66.780 16.995 67.110 17.325 ;
        RECT 74.290 16.995 74.620 17.325 ;
        RECT 0.000 16.195 3.840 16.365 ;
        RECT 97.440 16.195 101.280 16.365 ;
        RECT 11.525 15.770 11.855 16.100 ;
        RECT 16.010 15.770 16.340 16.100 ;
        RECT 21.470 15.770 21.800 16.100 ;
        RECT 28.495 15.770 28.825 16.100 ;
        RECT 36.230 15.770 36.560 16.100 ;
        RECT 43.785 15.770 44.115 16.100 ;
        RECT 51.595 15.770 51.925 16.100 ;
        RECT 59.105 15.770 59.435 16.100 ;
        RECT 66.780 15.770 67.110 16.100 ;
        RECT 74.290 15.770 74.620 16.100 ;
        RECT 77.980 15.665 79.400 15.835 ;
        RECT 83.530 15.665 84.950 15.835 ;
        RECT 8.045 15.210 11.310 15.380 ;
        RECT 12.530 15.210 15.795 15.380 ;
        RECT 17.645 15.210 21.255 15.380 ;
        RECT 23.360 15.210 28.280 15.380 ;
        RECT 31.095 15.210 36.015 15.380 ;
        RECT 38.650 15.210 43.570 15.380 ;
        RECT 46.460 15.210 51.380 15.380 ;
        RECT 53.970 15.210 58.890 15.380 ;
        RECT 61.645 15.210 66.565 15.380 ;
        RECT 69.155 15.210 74.075 15.380 ;
        RECT 77.515 15.055 77.845 15.135 ;
        RECT 11.525 14.660 11.855 14.990 ;
        RECT 16.010 14.660 16.340 14.990 ;
        RECT 21.470 14.660 21.800 14.990 ;
        RECT 28.495 14.660 28.825 14.990 ;
        RECT 36.230 14.660 36.560 14.990 ;
        RECT 43.785 14.660 44.115 14.990 ;
        RECT 51.595 14.660 51.925 14.990 ;
        RECT 59.105 14.660 59.435 14.990 ;
        RECT 66.780 14.660 67.110 14.990 ;
        RECT 74.290 14.660 74.620 14.990 ;
        RECT 77.515 14.885 78.990 15.055 ;
        RECT 77.515 14.805 77.845 14.885 ;
        RECT 79.230 14.275 79.400 15.665 ;
        RECT 83.065 15.055 83.395 15.135 ;
        RECT 83.065 14.885 84.540 15.055 ;
        RECT 83.065 14.805 83.395 14.885 ;
        RECT 84.780 14.275 84.950 15.665 ;
        RECT 88.735 15.055 89.065 15.135 ;
        RECT 88.735 14.885 90.210 15.055 ;
        RECT 88.735 14.805 89.065 14.885 ;
        RECT 77.980 14.105 79.400 14.275 ;
        RECT 83.530 14.105 84.950 14.275 ;
        RECT 11.525 13.475 11.855 13.805 ;
        RECT 16.010 13.475 16.340 13.805 ;
        RECT 21.470 13.475 21.800 13.805 ;
        RECT 28.495 13.475 28.825 13.805 ;
        RECT 36.230 13.475 36.560 13.805 ;
        RECT 43.785 13.475 44.115 13.805 ;
        RECT 51.595 13.475 51.925 13.805 ;
        RECT 59.105 13.475 59.435 13.805 ;
        RECT 66.780 13.475 67.110 13.805 ;
        RECT 74.290 13.475 74.620 13.805 ;
        RECT 78.375 13.600 78.545 14.105 ;
        RECT 83.925 13.600 84.095 14.105 ;
        RECT 77.745 13.270 79.275 13.600 ;
        RECT 83.295 13.270 84.825 13.600 ;
        RECT 8.045 12.850 11.310 13.020 ;
        RECT 12.530 12.850 15.795 13.020 ;
        RECT 17.645 12.850 21.255 13.020 ;
        RECT 23.360 12.850 28.280 13.020 ;
        RECT 31.095 12.850 36.015 13.020 ;
        RECT 38.650 12.850 43.570 13.020 ;
        RECT 46.460 12.850 51.380 13.020 ;
        RECT 53.970 12.850 58.890 13.020 ;
        RECT 61.645 12.850 66.565 13.020 ;
        RECT 69.155 12.850 74.075 13.020 ;
        RECT 11.525 12.295 11.855 12.625 ;
        RECT 16.010 12.295 16.340 12.625 ;
        RECT 21.470 12.295 21.800 12.625 ;
        RECT 28.495 12.295 28.825 12.625 ;
        RECT 36.230 12.295 36.560 12.625 ;
        RECT 43.785 12.295 44.115 12.625 ;
        RECT 51.595 12.295 51.925 12.625 ;
        RECT 59.105 12.295 59.435 12.625 ;
        RECT 66.780 12.295 67.110 12.625 ;
        RECT 74.290 12.295 74.620 12.625 ;
        RECT 0.000 12.125 3.840 12.295 ;
        RECT 97.440 12.125 101.280 12.295 ;
        RECT 0.000 8.055 3.840 8.225 ;
        RECT 97.440 8.055 101.280 8.225 ;
        RECT 0.000 3.985 101.280 4.155 ;
        RECT 0.000 -0.085 101.280 0.085 ;
      LAYER mcon ;
        RECT 0.155 60.965 0.325 61.135 ;
        RECT 0.635 60.965 0.805 61.135 ;
        RECT 1.115 60.965 1.285 61.135 ;
        RECT 1.595 60.965 1.765 61.135 ;
        RECT 2.075 60.965 2.245 61.135 ;
        RECT 2.555 60.965 2.725 61.135 ;
        RECT 3.035 60.965 3.205 61.135 ;
        RECT 3.515 60.965 3.685 61.135 ;
        RECT 3.995 60.965 4.165 61.135 ;
        RECT 4.475 60.965 4.645 61.135 ;
        RECT 4.955 60.965 5.125 61.135 ;
        RECT 5.435 60.965 5.605 61.135 ;
        RECT 5.915 60.965 6.085 61.135 ;
        RECT 6.395 60.965 6.565 61.135 ;
        RECT 6.875 60.965 7.045 61.135 ;
        RECT 7.355 60.965 7.525 61.135 ;
        RECT 7.835 60.965 8.005 61.135 ;
        RECT 8.315 60.965 8.485 61.135 ;
        RECT 8.795 60.965 8.965 61.135 ;
        RECT 9.275 60.965 9.445 61.135 ;
        RECT 9.755 60.965 9.925 61.135 ;
        RECT 10.235 60.965 10.405 61.135 ;
        RECT 10.715 60.965 10.885 61.135 ;
        RECT 11.195 60.965 11.365 61.135 ;
        RECT 11.675 60.965 11.845 61.135 ;
        RECT 12.155 60.965 12.325 61.135 ;
        RECT 12.635 60.965 12.805 61.135 ;
        RECT 13.115 60.965 13.285 61.135 ;
        RECT 13.595 60.965 13.765 61.135 ;
        RECT 14.075 60.965 14.245 61.135 ;
        RECT 14.555 60.965 14.725 61.135 ;
        RECT 15.035 60.965 15.205 61.135 ;
        RECT 15.515 60.965 15.685 61.135 ;
        RECT 15.995 60.965 16.165 61.135 ;
        RECT 16.475 60.965 16.645 61.135 ;
        RECT 16.955 60.965 17.125 61.135 ;
        RECT 17.435 60.965 17.605 61.135 ;
        RECT 17.915 60.965 18.085 61.135 ;
        RECT 18.395 60.965 18.565 61.135 ;
        RECT 18.875 60.965 19.045 61.135 ;
        RECT 19.355 60.965 19.525 61.135 ;
        RECT 19.835 60.965 20.005 61.135 ;
        RECT 20.315 60.965 20.485 61.135 ;
        RECT 20.795 60.965 20.965 61.135 ;
        RECT 21.275 60.965 21.445 61.135 ;
        RECT 21.755 60.965 21.925 61.135 ;
        RECT 22.235 60.965 22.405 61.135 ;
        RECT 22.715 60.965 22.885 61.135 ;
        RECT 23.195 60.965 23.365 61.135 ;
        RECT 23.675 60.965 23.845 61.135 ;
        RECT 24.155 60.965 24.325 61.135 ;
        RECT 24.635 60.965 24.805 61.135 ;
        RECT 25.115 60.965 25.285 61.135 ;
        RECT 25.595 60.965 25.765 61.135 ;
        RECT 26.075 60.965 26.245 61.135 ;
        RECT 26.555 60.965 26.725 61.135 ;
        RECT 27.035 60.965 27.205 61.135 ;
        RECT 27.515 60.965 27.685 61.135 ;
        RECT 27.995 60.965 28.165 61.135 ;
        RECT 28.475 60.965 28.645 61.135 ;
        RECT 28.955 60.965 29.125 61.135 ;
        RECT 29.435 60.965 29.605 61.135 ;
        RECT 29.915 60.965 30.085 61.135 ;
        RECT 30.395 60.965 30.565 61.135 ;
        RECT 30.875 60.965 31.045 61.135 ;
        RECT 31.355 60.965 31.525 61.135 ;
        RECT 31.835 60.965 32.005 61.135 ;
        RECT 32.315 60.965 32.485 61.135 ;
        RECT 32.795 60.965 32.965 61.135 ;
        RECT 33.275 60.965 33.445 61.135 ;
        RECT 33.755 60.965 33.925 61.135 ;
        RECT 34.235 60.965 34.405 61.135 ;
        RECT 34.715 60.965 34.885 61.135 ;
        RECT 35.195 60.965 35.365 61.135 ;
        RECT 35.675 60.965 35.845 61.135 ;
        RECT 36.155 60.965 36.325 61.135 ;
        RECT 36.635 60.965 36.805 61.135 ;
        RECT 37.115 60.965 37.285 61.135 ;
        RECT 37.595 60.965 37.765 61.135 ;
        RECT 38.075 60.965 38.245 61.135 ;
        RECT 38.555 60.965 38.725 61.135 ;
        RECT 39.035 60.965 39.205 61.135 ;
        RECT 39.515 60.965 39.685 61.135 ;
        RECT 39.995 60.965 40.165 61.135 ;
        RECT 40.475 60.965 40.645 61.135 ;
        RECT 40.955 60.965 41.125 61.135 ;
        RECT 41.435 60.965 41.605 61.135 ;
        RECT 41.915 60.965 42.085 61.135 ;
        RECT 42.395 60.965 42.565 61.135 ;
        RECT 42.875 60.965 43.045 61.135 ;
        RECT 43.355 60.965 43.525 61.135 ;
        RECT 43.835 60.965 44.005 61.135 ;
        RECT 44.315 60.965 44.485 61.135 ;
        RECT 44.795 60.965 44.965 61.135 ;
        RECT 45.275 60.965 45.445 61.135 ;
        RECT 45.755 60.965 45.925 61.135 ;
        RECT 46.235 60.965 46.405 61.135 ;
        RECT 46.715 60.965 46.885 61.135 ;
        RECT 47.195 60.965 47.365 61.135 ;
        RECT 47.675 60.965 47.845 61.135 ;
        RECT 48.155 60.965 48.325 61.135 ;
        RECT 48.635 60.965 48.805 61.135 ;
        RECT 49.115 60.965 49.285 61.135 ;
        RECT 49.595 60.965 49.765 61.135 ;
        RECT 50.075 60.965 50.245 61.135 ;
        RECT 50.555 60.965 50.725 61.135 ;
        RECT 51.035 60.965 51.205 61.135 ;
        RECT 51.515 60.965 51.685 61.135 ;
        RECT 51.995 60.965 52.165 61.135 ;
        RECT 52.475 60.965 52.645 61.135 ;
        RECT 52.955 60.965 53.125 61.135 ;
        RECT 53.435 60.965 53.605 61.135 ;
        RECT 53.915 60.965 54.085 61.135 ;
        RECT 54.395 60.965 54.565 61.135 ;
        RECT 54.875 60.965 55.045 61.135 ;
        RECT 55.355 60.965 55.525 61.135 ;
        RECT 55.835 60.965 56.005 61.135 ;
        RECT 56.315 60.965 56.485 61.135 ;
        RECT 56.795 60.965 56.965 61.135 ;
        RECT 57.275 60.965 57.445 61.135 ;
        RECT 57.755 60.965 57.925 61.135 ;
        RECT 58.235 60.965 58.405 61.135 ;
        RECT 58.715 60.965 58.885 61.135 ;
        RECT 59.195 60.965 59.365 61.135 ;
        RECT 59.675 60.965 59.845 61.135 ;
        RECT 60.155 60.965 60.325 61.135 ;
        RECT 60.635 60.965 60.805 61.135 ;
        RECT 61.115 60.965 61.285 61.135 ;
        RECT 61.595 60.965 61.765 61.135 ;
        RECT 62.075 60.965 62.245 61.135 ;
        RECT 62.555 60.965 62.725 61.135 ;
        RECT 63.035 60.965 63.205 61.135 ;
        RECT 63.515 60.965 63.685 61.135 ;
        RECT 63.995 60.965 64.165 61.135 ;
        RECT 64.475 60.965 64.645 61.135 ;
        RECT 64.955 60.965 65.125 61.135 ;
        RECT 65.435 60.965 65.605 61.135 ;
        RECT 65.915 60.965 66.085 61.135 ;
        RECT 66.395 60.965 66.565 61.135 ;
        RECT 66.875 60.965 67.045 61.135 ;
        RECT 67.355 60.965 67.525 61.135 ;
        RECT 67.835 60.965 68.005 61.135 ;
        RECT 68.315 60.965 68.485 61.135 ;
        RECT 68.795 60.965 68.965 61.135 ;
        RECT 69.275 60.965 69.445 61.135 ;
        RECT 69.755 60.965 69.925 61.135 ;
        RECT 70.235 60.965 70.405 61.135 ;
        RECT 70.715 60.965 70.885 61.135 ;
        RECT 71.195 60.965 71.365 61.135 ;
        RECT 71.675 60.965 71.845 61.135 ;
        RECT 72.155 60.965 72.325 61.135 ;
        RECT 72.635 60.965 72.805 61.135 ;
        RECT 73.115 60.965 73.285 61.135 ;
        RECT 73.595 60.965 73.765 61.135 ;
        RECT 74.075 60.965 74.245 61.135 ;
        RECT 74.555 60.965 74.725 61.135 ;
        RECT 75.035 60.965 75.205 61.135 ;
        RECT 75.515 60.965 75.685 61.135 ;
        RECT 75.995 60.965 76.165 61.135 ;
        RECT 76.475 60.965 76.645 61.135 ;
        RECT 76.955 60.965 77.125 61.135 ;
        RECT 77.435 60.965 77.605 61.135 ;
        RECT 77.915 60.965 78.085 61.135 ;
        RECT 78.395 60.965 78.565 61.135 ;
        RECT 78.875 60.965 79.045 61.135 ;
        RECT 79.355 60.965 79.525 61.135 ;
        RECT 79.835 60.965 80.005 61.135 ;
        RECT 80.315 60.965 80.485 61.135 ;
        RECT 80.795 60.965 80.965 61.135 ;
        RECT 81.275 60.965 81.445 61.135 ;
        RECT 81.755 60.965 81.925 61.135 ;
        RECT 82.235 60.965 82.405 61.135 ;
        RECT 82.715 60.965 82.885 61.135 ;
        RECT 83.195 60.965 83.365 61.135 ;
        RECT 83.675 60.965 83.845 61.135 ;
        RECT 84.155 60.965 84.325 61.135 ;
        RECT 84.635 60.965 84.805 61.135 ;
        RECT 85.115 60.965 85.285 61.135 ;
        RECT 85.595 60.965 85.765 61.135 ;
        RECT 86.075 60.965 86.245 61.135 ;
        RECT 86.555 60.965 86.725 61.135 ;
        RECT 87.035 60.965 87.205 61.135 ;
        RECT 87.515 60.965 87.685 61.135 ;
        RECT 87.995 60.965 88.165 61.135 ;
        RECT 88.475 60.965 88.645 61.135 ;
        RECT 88.955 60.965 89.125 61.135 ;
        RECT 89.435 60.965 89.605 61.135 ;
        RECT 89.915 60.965 90.085 61.135 ;
        RECT 90.395 60.965 90.565 61.135 ;
        RECT 90.875 60.965 91.045 61.135 ;
        RECT 91.355 60.965 91.525 61.135 ;
        RECT 91.835 60.965 92.005 61.135 ;
        RECT 92.315 60.965 92.485 61.135 ;
        RECT 92.795 60.965 92.965 61.135 ;
        RECT 93.275 60.965 93.445 61.135 ;
        RECT 93.755 60.965 93.925 61.135 ;
        RECT 94.235 60.965 94.405 61.135 ;
        RECT 94.715 60.965 94.885 61.135 ;
        RECT 95.195 60.965 95.365 61.135 ;
        RECT 95.675 60.965 95.845 61.135 ;
        RECT 96.155 60.965 96.325 61.135 ;
        RECT 96.635 60.965 96.805 61.135 ;
        RECT 97.115 60.965 97.285 61.135 ;
        RECT 97.595 60.965 97.765 61.135 ;
        RECT 98.075 60.965 98.245 61.135 ;
        RECT 98.555 60.965 98.725 61.135 ;
        RECT 99.035 60.965 99.205 61.135 ;
        RECT 99.515 60.965 99.685 61.135 ;
        RECT 99.995 60.965 100.165 61.135 ;
        RECT 100.475 60.965 100.645 61.135 ;
        RECT 100.955 60.965 101.125 61.135 ;
        RECT 0.155 56.895 0.325 57.065 ;
        RECT 0.635 56.895 0.805 57.065 ;
        RECT 1.115 56.895 1.285 57.065 ;
        RECT 1.595 56.895 1.765 57.065 ;
        RECT 2.075 56.895 2.245 57.065 ;
        RECT 2.555 56.895 2.725 57.065 ;
        RECT 3.035 56.895 3.205 57.065 ;
        RECT 3.515 56.895 3.685 57.065 ;
        RECT 3.995 56.895 4.165 57.065 ;
        RECT 4.475 56.895 4.645 57.065 ;
        RECT 4.955 56.895 5.125 57.065 ;
        RECT 5.435 56.895 5.605 57.065 ;
        RECT 5.915 56.895 6.085 57.065 ;
        RECT 6.395 56.895 6.565 57.065 ;
        RECT 6.875 56.895 7.045 57.065 ;
        RECT 7.355 56.895 7.525 57.065 ;
        RECT 7.835 56.895 8.005 57.065 ;
        RECT 8.315 56.895 8.485 57.065 ;
        RECT 8.795 56.895 8.965 57.065 ;
        RECT 9.275 56.895 9.445 57.065 ;
        RECT 9.755 56.895 9.925 57.065 ;
        RECT 10.235 56.895 10.405 57.065 ;
        RECT 10.715 56.895 10.885 57.065 ;
        RECT 11.195 56.895 11.365 57.065 ;
        RECT 11.675 56.895 11.845 57.065 ;
        RECT 12.155 56.895 12.325 57.065 ;
        RECT 12.635 56.895 12.805 57.065 ;
        RECT 13.115 56.895 13.285 57.065 ;
        RECT 13.595 56.895 13.765 57.065 ;
        RECT 14.075 56.895 14.245 57.065 ;
        RECT 14.555 56.895 14.725 57.065 ;
        RECT 15.035 56.895 15.205 57.065 ;
        RECT 15.515 56.895 15.685 57.065 ;
        RECT 15.995 56.895 16.165 57.065 ;
        RECT 16.475 56.895 16.645 57.065 ;
        RECT 16.955 56.895 17.125 57.065 ;
        RECT 17.435 56.895 17.605 57.065 ;
        RECT 17.915 56.895 18.085 57.065 ;
        RECT 18.395 56.895 18.565 57.065 ;
        RECT 18.875 56.895 19.045 57.065 ;
        RECT 19.355 56.895 19.525 57.065 ;
        RECT 19.835 56.895 20.005 57.065 ;
        RECT 20.315 56.895 20.485 57.065 ;
        RECT 20.795 56.895 20.965 57.065 ;
        RECT 21.275 56.895 21.445 57.065 ;
        RECT 21.755 56.895 21.925 57.065 ;
        RECT 22.235 56.895 22.405 57.065 ;
        RECT 22.715 56.895 22.885 57.065 ;
        RECT 23.195 56.895 23.365 57.065 ;
        RECT 23.675 56.895 23.845 57.065 ;
        RECT 24.155 56.895 24.325 57.065 ;
        RECT 24.635 56.895 24.805 57.065 ;
        RECT 25.115 56.895 25.285 57.065 ;
        RECT 25.595 56.895 25.765 57.065 ;
        RECT 26.075 56.895 26.245 57.065 ;
        RECT 26.555 56.895 26.725 57.065 ;
        RECT 27.035 56.895 27.205 57.065 ;
        RECT 27.515 56.895 27.685 57.065 ;
        RECT 27.995 56.895 28.165 57.065 ;
        RECT 28.475 56.895 28.645 57.065 ;
        RECT 28.955 56.895 29.125 57.065 ;
        RECT 29.435 56.895 29.605 57.065 ;
        RECT 29.915 56.895 30.085 57.065 ;
        RECT 30.395 56.895 30.565 57.065 ;
        RECT 30.875 56.895 31.045 57.065 ;
        RECT 31.355 56.895 31.525 57.065 ;
        RECT 31.835 56.895 32.005 57.065 ;
        RECT 32.315 56.895 32.485 57.065 ;
        RECT 32.795 56.895 32.965 57.065 ;
        RECT 33.275 56.895 33.445 57.065 ;
        RECT 33.755 56.895 33.925 57.065 ;
        RECT 34.235 56.895 34.405 57.065 ;
        RECT 34.715 56.895 34.885 57.065 ;
        RECT 35.195 56.895 35.365 57.065 ;
        RECT 35.675 56.895 35.845 57.065 ;
        RECT 36.155 56.895 36.325 57.065 ;
        RECT 36.635 56.895 36.805 57.065 ;
        RECT 37.115 56.895 37.285 57.065 ;
        RECT 37.595 56.895 37.765 57.065 ;
        RECT 38.075 56.895 38.245 57.065 ;
        RECT 38.555 56.895 38.725 57.065 ;
        RECT 39.035 56.895 39.205 57.065 ;
        RECT 39.515 56.895 39.685 57.065 ;
        RECT 39.995 56.895 40.165 57.065 ;
        RECT 40.475 56.895 40.645 57.065 ;
        RECT 40.955 56.895 41.125 57.065 ;
        RECT 41.435 56.895 41.605 57.065 ;
        RECT 41.915 56.895 42.085 57.065 ;
        RECT 42.395 56.895 42.565 57.065 ;
        RECT 42.875 56.895 43.045 57.065 ;
        RECT 43.355 56.895 43.525 57.065 ;
        RECT 43.835 56.895 44.005 57.065 ;
        RECT 44.315 56.895 44.485 57.065 ;
        RECT 44.795 56.895 44.965 57.065 ;
        RECT 45.275 56.895 45.445 57.065 ;
        RECT 45.755 56.895 45.925 57.065 ;
        RECT 46.235 56.895 46.405 57.065 ;
        RECT 46.715 56.895 46.885 57.065 ;
        RECT 47.195 56.895 47.365 57.065 ;
        RECT 47.675 56.895 47.845 57.065 ;
        RECT 48.155 56.895 48.325 57.065 ;
        RECT 48.635 56.895 48.805 57.065 ;
        RECT 49.115 56.895 49.285 57.065 ;
        RECT 49.595 56.895 49.765 57.065 ;
        RECT 50.075 56.895 50.245 57.065 ;
        RECT 50.555 56.895 50.725 57.065 ;
        RECT 51.035 56.895 51.205 57.065 ;
        RECT 51.515 56.895 51.685 57.065 ;
        RECT 51.995 56.895 52.165 57.065 ;
        RECT 52.475 56.895 52.645 57.065 ;
        RECT 52.955 56.895 53.125 57.065 ;
        RECT 53.435 56.895 53.605 57.065 ;
        RECT 53.915 56.895 54.085 57.065 ;
        RECT 54.395 56.895 54.565 57.065 ;
        RECT 54.875 56.895 55.045 57.065 ;
        RECT 55.355 56.895 55.525 57.065 ;
        RECT 55.835 56.895 56.005 57.065 ;
        RECT 56.315 56.895 56.485 57.065 ;
        RECT 56.795 56.895 56.965 57.065 ;
        RECT 57.275 56.895 57.445 57.065 ;
        RECT 57.755 56.895 57.925 57.065 ;
        RECT 58.235 56.895 58.405 57.065 ;
        RECT 58.715 56.895 58.885 57.065 ;
        RECT 59.195 56.895 59.365 57.065 ;
        RECT 59.675 56.895 59.845 57.065 ;
        RECT 60.155 56.895 60.325 57.065 ;
        RECT 60.635 56.895 60.805 57.065 ;
        RECT 61.115 56.895 61.285 57.065 ;
        RECT 61.595 56.895 61.765 57.065 ;
        RECT 62.075 56.895 62.245 57.065 ;
        RECT 62.555 56.895 62.725 57.065 ;
        RECT 63.035 56.895 63.205 57.065 ;
        RECT 63.515 56.895 63.685 57.065 ;
        RECT 63.995 56.895 64.165 57.065 ;
        RECT 64.475 56.895 64.645 57.065 ;
        RECT 64.955 56.895 65.125 57.065 ;
        RECT 65.435 56.895 65.605 57.065 ;
        RECT 65.915 56.895 66.085 57.065 ;
        RECT 66.395 56.895 66.565 57.065 ;
        RECT 66.875 56.895 67.045 57.065 ;
        RECT 67.355 56.895 67.525 57.065 ;
        RECT 67.835 56.895 68.005 57.065 ;
        RECT 68.315 56.895 68.485 57.065 ;
        RECT 68.795 56.895 68.965 57.065 ;
        RECT 69.275 56.895 69.445 57.065 ;
        RECT 69.755 56.895 69.925 57.065 ;
        RECT 70.235 56.895 70.405 57.065 ;
        RECT 70.715 56.895 70.885 57.065 ;
        RECT 71.195 56.895 71.365 57.065 ;
        RECT 71.675 56.895 71.845 57.065 ;
        RECT 72.155 56.895 72.325 57.065 ;
        RECT 72.635 56.895 72.805 57.065 ;
        RECT 73.115 56.895 73.285 57.065 ;
        RECT 73.595 56.895 73.765 57.065 ;
        RECT 74.075 56.895 74.245 57.065 ;
        RECT 74.555 56.895 74.725 57.065 ;
        RECT 75.035 56.895 75.205 57.065 ;
        RECT 75.515 56.895 75.685 57.065 ;
        RECT 75.995 56.895 76.165 57.065 ;
        RECT 76.475 56.895 76.645 57.065 ;
        RECT 76.955 56.895 77.125 57.065 ;
        RECT 77.435 56.895 77.605 57.065 ;
        RECT 77.915 56.895 78.085 57.065 ;
        RECT 78.395 56.895 78.565 57.065 ;
        RECT 78.875 56.895 79.045 57.065 ;
        RECT 79.355 56.895 79.525 57.065 ;
        RECT 79.835 56.895 80.005 57.065 ;
        RECT 80.315 56.895 80.485 57.065 ;
        RECT 80.795 56.895 80.965 57.065 ;
        RECT 81.275 56.895 81.445 57.065 ;
        RECT 81.755 56.895 81.925 57.065 ;
        RECT 82.235 56.895 82.405 57.065 ;
        RECT 82.715 56.895 82.885 57.065 ;
        RECT 83.195 56.895 83.365 57.065 ;
        RECT 83.675 56.895 83.845 57.065 ;
        RECT 84.155 56.895 84.325 57.065 ;
        RECT 84.635 56.895 84.805 57.065 ;
        RECT 85.115 56.895 85.285 57.065 ;
        RECT 85.595 56.895 85.765 57.065 ;
        RECT 86.075 56.895 86.245 57.065 ;
        RECT 86.555 56.895 86.725 57.065 ;
        RECT 87.035 56.895 87.205 57.065 ;
        RECT 87.515 56.895 87.685 57.065 ;
        RECT 87.995 56.895 88.165 57.065 ;
        RECT 88.475 56.895 88.645 57.065 ;
        RECT 88.955 56.895 89.125 57.065 ;
        RECT 89.435 56.895 89.605 57.065 ;
        RECT 89.915 56.895 90.085 57.065 ;
        RECT 90.395 56.895 90.565 57.065 ;
        RECT 90.875 56.895 91.045 57.065 ;
        RECT 91.355 56.895 91.525 57.065 ;
        RECT 91.835 56.895 92.005 57.065 ;
        RECT 92.315 56.895 92.485 57.065 ;
        RECT 92.795 56.895 92.965 57.065 ;
        RECT 93.275 56.895 93.445 57.065 ;
        RECT 93.755 56.895 93.925 57.065 ;
        RECT 94.235 56.895 94.405 57.065 ;
        RECT 94.715 56.895 94.885 57.065 ;
        RECT 95.195 56.895 95.365 57.065 ;
        RECT 95.675 56.895 95.845 57.065 ;
        RECT 96.155 56.895 96.325 57.065 ;
        RECT 96.635 56.895 96.805 57.065 ;
        RECT 97.115 56.895 97.285 57.065 ;
        RECT 97.595 56.895 97.765 57.065 ;
        RECT 98.075 56.895 98.245 57.065 ;
        RECT 98.555 56.895 98.725 57.065 ;
        RECT 99.035 56.895 99.205 57.065 ;
        RECT 99.515 56.895 99.685 57.065 ;
        RECT 99.995 56.895 100.165 57.065 ;
        RECT 100.475 56.895 100.645 57.065 ;
        RECT 100.955 56.895 101.125 57.065 ;
        RECT 0.155 52.825 0.325 52.995 ;
        RECT 0.635 52.825 0.805 52.995 ;
        RECT 1.115 52.825 1.285 52.995 ;
        RECT 1.595 52.825 1.765 52.995 ;
        RECT 2.075 52.825 2.245 52.995 ;
        RECT 2.555 52.825 2.725 52.995 ;
        RECT 3.035 52.825 3.205 52.995 ;
        RECT 3.515 52.825 3.685 52.995 ;
        RECT 97.595 52.825 97.765 52.995 ;
        RECT 98.075 52.825 98.245 52.995 ;
        RECT 98.555 52.825 98.725 52.995 ;
        RECT 99.035 52.825 99.205 52.995 ;
        RECT 99.515 52.825 99.685 52.995 ;
        RECT 99.995 52.825 100.165 52.995 ;
        RECT 100.475 52.825 100.645 52.995 ;
        RECT 100.955 52.825 101.125 52.995 ;
        RECT 0.155 48.755 0.325 48.925 ;
        RECT 0.635 48.755 0.805 48.925 ;
        RECT 1.115 48.755 1.285 48.925 ;
        RECT 1.595 48.755 1.765 48.925 ;
        RECT 2.075 48.755 2.245 48.925 ;
        RECT 2.555 48.755 2.725 48.925 ;
        RECT 3.035 48.755 3.205 48.925 ;
        RECT 3.515 48.755 3.685 48.925 ;
        RECT 8.095 48.600 8.265 48.770 ;
        RECT 8.455 48.600 8.625 48.770 ;
        RECT 8.815 48.600 8.985 48.770 ;
        RECT 9.175 48.600 9.345 48.770 ;
        RECT 12.580 48.565 12.750 48.735 ;
        RECT 12.940 48.565 13.110 48.735 ;
        RECT 13.300 48.565 13.470 48.735 ;
        RECT 13.660 48.565 13.830 48.735 ;
        RECT 18.040 48.565 18.210 48.735 ;
        RECT 18.400 48.565 18.570 48.735 ;
        RECT 18.760 48.565 18.930 48.735 ;
        RECT 19.120 48.565 19.290 48.735 ;
        RECT 25.065 48.565 25.235 48.735 ;
        RECT 25.425 48.565 25.595 48.735 ;
        RECT 25.785 48.565 25.955 48.735 ;
        RECT 26.145 48.565 26.315 48.735 ;
        RECT 32.800 48.565 32.970 48.735 ;
        RECT 33.160 48.565 33.330 48.735 ;
        RECT 33.520 48.565 33.690 48.735 ;
        RECT 33.880 48.565 34.050 48.735 ;
        RECT 40.355 48.565 40.525 48.735 ;
        RECT 40.715 48.565 40.885 48.735 ;
        RECT 41.075 48.565 41.245 48.735 ;
        RECT 41.435 48.565 41.605 48.735 ;
        RECT 48.165 48.565 48.335 48.735 ;
        RECT 48.525 48.565 48.695 48.735 ;
        RECT 48.885 48.565 49.055 48.735 ;
        RECT 49.245 48.565 49.415 48.735 ;
        RECT 55.675 48.565 55.845 48.735 ;
        RECT 56.035 48.565 56.205 48.735 ;
        RECT 56.395 48.565 56.565 48.735 ;
        RECT 56.755 48.565 56.925 48.735 ;
        RECT 63.350 48.565 63.520 48.735 ;
        RECT 63.710 48.565 63.880 48.735 ;
        RECT 64.070 48.565 64.240 48.735 ;
        RECT 64.430 48.565 64.600 48.735 ;
        RECT 97.595 48.755 97.765 48.925 ;
        RECT 98.075 48.755 98.245 48.925 ;
        RECT 98.555 48.755 98.725 48.925 ;
        RECT 99.035 48.755 99.205 48.925 ;
        RECT 99.515 48.755 99.685 48.925 ;
        RECT 99.995 48.755 100.165 48.925 ;
        RECT 100.475 48.755 100.645 48.925 ;
        RECT 100.955 48.755 101.125 48.925 ;
        RECT 70.860 48.565 71.030 48.735 ;
        RECT 71.220 48.565 71.390 48.735 ;
        RECT 71.580 48.565 71.750 48.735 ;
        RECT 71.940 48.565 72.110 48.735 ;
        RECT 11.605 46.375 11.775 46.545 ;
        RECT 16.090 46.375 16.260 46.545 ;
        RECT 21.550 46.375 21.720 46.545 ;
        RECT 28.575 46.375 28.745 46.545 ;
        RECT 36.310 46.375 36.480 46.545 ;
        RECT 43.865 46.375 44.035 46.545 ;
        RECT 51.675 46.375 51.845 46.545 ;
        RECT 59.185 46.375 59.355 46.545 ;
        RECT 66.860 46.375 67.030 46.545 ;
        RECT 74.370 46.375 74.540 46.545 ;
        RECT 8.455 45.885 8.625 46.055 ;
        RECT 8.815 45.885 8.985 46.055 ;
        RECT 9.175 45.885 9.345 46.055 ;
        RECT 12.940 45.885 13.110 46.055 ;
        RECT 13.300 45.885 13.470 46.055 ;
        RECT 13.660 45.885 13.830 46.055 ;
        RECT 18.400 45.885 18.570 46.055 ;
        RECT 18.760 45.885 18.930 46.055 ;
        RECT 19.120 45.885 19.290 46.055 ;
        RECT 25.425 45.885 25.595 46.055 ;
        RECT 25.785 45.885 25.955 46.055 ;
        RECT 26.145 45.885 26.315 46.055 ;
        RECT 33.160 45.885 33.330 46.055 ;
        RECT 33.520 45.885 33.690 46.055 ;
        RECT 33.880 45.885 34.050 46.055 ;
        RECT 40.715 45.885 40.885 46.055 ;
        RECT 41.075 45.885 41.245 46.055 ;
        RECT 41.435 45.885 41.605 46.055 ;
        RECT 48.525 45.885 48.695 46.055 ;
        RECT 48.885 45.885 49.055 46.055 ;
        RECT 49.245 45.885 49.415 46.055 ;
        RECT 56.035 45.885 56.205 46.055 ;
        RECT 56.395 45.885 56.565 46.055 ;
        RECT 56.755 45.885 56.925 46.055 ;
        RECT 63.710 45.885 63.880 46.055 ;
        RECT 64.070 45.885 64.240 46.055 ;
        RECT 64.430 45.885 64.600 46.055 ;
        RECT 71.220 45.885 71.390 46.055 ;
        RECT 71.580 45.885 71.750 46.055 ;
        RECT 71.940 45.885 72.110 46.055 ;
        RECT 11.605 45.320 11.775 45.490 ;
        RECT 16.090 45.320 16.260 45.490 ;
        RECT 21.550 45.320 21.720 45.490 ;
        RECT 28.575 45.320 28.745 45.490 ;
        RECT 36.310 45.320 36.480 45.490 ;
        RECT 43.865 45.320 44.035 45.490 ;
        RECT 51.675 45.320 51.845 45.490 ;
        RECT 59.185 45.320 59.355 45.490 ;
        RECT 66.860 45.320 67.030 45.490 ;
        RECT 74.370 45.320 74.540 45.490 ;
        RECT 0.155 44.685 0.325 44.855 ;
        RECT 0.635 44.685 0.805 44.855 ;
        RECT 1.115 44.685 1.285 44.855 ;
        RECT 1.595 44.685 1.765 44.855 ;
        RECT 2.075 44.685 2.245 44.855 ;
        RECT 2.555 44.685 2.725 44.855 ;
        RECT 3.035 44.685 3.205 44.855 ;
        RECT 3.515 44.685 3.685 44.855 ;
        RECT 83.150 45.215 83.320 45.385 ;
        RECT 83.610 45.215 83.780 45.385 ;
        RECT 84.290 45.215 84.460 45.385 ;
        RECT 97.595 44.685 97.765 44.855 ;
        RECT 98.075 44.685 98.245 44.855 ;
        RECT 98.555 44.685 98.725 44.855 ;
        RECT 99.035 44.685 99.205 44.855 ;
        RECT 99.515 44.685 99.685 44.855 ;
        RECT 99.995 44.685 100.165 44.855 ;
        RECT 100.475 44.685 100.645 44.855 ;
        RECT 100.955 44.685 101.125 44.855 ;
        RECT 11.605 44.100 11.775 44.270 ;
        RECT 16.090 44.100 16.260 44.270 ;
        RECT 21.550 44.100 21.720 44.270 ;
        RECT 28.575 44.100 28.745 44.270 ;
        RECT 36.310 44.100 36.480 44.270 ;
        RECT 43.865 44.100 44.035 44.270 ;
        RECT 51.675 44.100 51.845 44.270 ;
        RECT 59.185 44.100 59.355 44.270 ;
        RECT 66.860 44.100 67.030 44.270 ;
        RECT 74.370 44.100 74.540 44.270 ;
        RECT 8.455 43.525 8.625 43.695 ;
        RECT 8.815 43.525 8.985 43.695 ;
        RECT 9.175 43.525 9.345 43.695 ;
        RECT 12.940 43.525 13.110 43.695 ;
        RECT 13.300 43.525 13.470 43.695 ;
        RECT 13.660 43.525 13.830 43.695 ;
        RECT 18.400 43.525 18.570 43.695 ;
        RECT 18.760 43.525 18.930 43.695 ;
        RECT 19.120 43.525 19.290 43.695 ;
        RECT 25.425 43.525 25.595 43.695 ;
        RECT 25.785 43.525 25.955 43.695 ;
        RECT 26.145 43.525 26.315 43.695 ;
        RECT 33.160 43.525 33.330 43.695 ;
        RECT 33.520 43.525 33.690 43.695 ;
        RECT 33.880 43.525 34.050 43.695 ;
        RECT 40.715 43.525 40.885 43.695 ;
        RECT 41.075 43.525 41.245 43.695 ;
        RECT 41.435 43.525 41.605 43.695 ;
        RECT 48.525 43.525 48.695 43.695 ;
        RECT 48.885 43.525 49.055 43.695 ;
        RECT 49.245 43.525 49.415 43.695 ;
        RECT 56.035 43.525 56.205 43.695 ;
        RECT 56.395 43.525 56.565 43.695 ;
        RECT 56.755 43.525 56.925 43.695 ;
        RECT 63.710 43.525 63.880 43.695 ;
        RECT 64.070 43.525 64.240 43.695 ;
        RECT 64.430 43.525 64.600 43.695 ;
        RECT 71.220 43.525 71.390 43.695 ;
        RECT 71.580 43.525 71.750 43.695 ;
        RECT 71.940 43.525 72.110 43.695 ;
        RECT 78.405 43.680 78.575 43.850 ;
        RECT 83.955 43.680 84.125 43.850 ;
        RECT 11.605 42.990 11.775 43.160 ;
        RECT 16.090 42.990 16.260 43.160 ;
        RECT 21.550 42.990 21.720 43.160 ;
        RECT 28.575 42.990 28.745 43.160 ;
        RECT 36.310 42.990 36.480 43.160 ;
        RECT 43.865 42.990 44.035 43.160 ;
        RECT 51.675 42.990 51.845 43.160 ;
        RECT 59.185 42.990 59.355 43.160 ;
        RECT 66.860 42.990 67.030 43.160 ;
        RECT 74.370 42.990 74.540 43.160 ;
        RECT 11.605 41.810 11.775 41.980 ;
        RECT 16.090 41.810 16.260 41.980 ;
        RECT 21.550 41.810 21.720 41.980 ;
        RECT 28.575 41.810 28.745 41.980 ;
        RECT 36.310 41.810 36.480 41.980 ;
        RECT 43.865 41.810 44.035 41.980 ;
        RECT 51.675 41.810 51.845 41.980 ;
        RECT 59.185 41.810 59.355 41.980 ;
        RECT 66.860 41.810 67.030 41.980 ;
        RECT 74.370 41.810 74.540 41.980 ;
        RECT 8.095 41.170 8.265 41.340 ;
        RECT 8.455 41.170 8.625 41.340 ;
        RECT 8.815 41.170 8.985 41.340 ;
        RECT 9.175 41.170 9.345 41.340 ;
        RECT 12.580 41.170 12.750 41.340 ;
        RECT 12.940 41.170 13.110 41.340 ;
        RECT 13.300 41.170 13.470 41.340 ;
        RECT 13.660 41.170 13.830 41.340 ;
        RECT 18.040 41.170 18.210 41.340 ;
        RECT 18.400 41.170 18.570 41.340 ;
        RECT 18.760 41.170 18.930 41.340 ;
        RECT 19.120 41.170 19.290 41.340 ;
        RECT 25.065 41.170 25.235 41.340 ;
        RECT 25.425 41.170 25.595 41.340 ;
        RECT 25.785 41.170 25.955 41.340 ;
        RECT 26.145 41.170 26.315 41.340 ;
        RECT 32.800 41.170 32.970 41.340 ;
        RECT 33.160 41.170 33.330 41.340 ;
        RECT 33.520 41.170 33.690 41.340 ;
        RECT 33.880 41.170 34.050 41.340 ;
        RECT 40.355 41.170 40.525 41.340 ;
        RECT 40.715 41.170 40.885 41.340 ;
        RECT 41.075 41.170 41.245 41.340 ;
        RECT 41.435 41.170 41.605 41.340 ;
        RECT 48.165 41.170 48.335 41.340 ;
        RECT 48.525 41.170 48.695 41.340 ;
        RECT 48.885 41.170 49.055 41.340 ;
        RECT 49.245 41.170 49.415 41.340 ;
        RECT 55.675 41.170 55.845 41.340 ;
        RECT 56.035 41.170 56.205 41.340 ;
        RECT 56.395 41.170 56.565 41.340 ;
        RECT 56.755 41.170 56.925 41.340 ;
        RECT 63.350 41.170 63.520 41.340 ;
        RECT 63.710 41.170 63.880 41.340 ;
        RECT 64.070 41.170 64.240 41.340 ;
        RECT 64.430 41.170 64.600 41.340 ;
        RECT 70.860 41.170 71.030 41.340 ;
        RECT 71.220 41.170 71.390 41.340 ;
        RECT 71.580 41.170 71.750 41.340 ;
        RECT 71.940 41.170 72.110 41.340 ;
        RECT 0.155 40.615 0.325 40.785 ;
        RECT 0.635 40.615 0.805 40.785 ;
        RECT 1.115 40.615 1.285 40.785 ;
        RECT 1.595 40.615 1.765 40.785 ;
        RECT 2.075 40.615 2.245 40.785 ;
        RECT 2.555 40.615 2.725 40.785 ;
        RECT 3.035 40.615 3.205 40.785 ;
        RECT 3.515 40.615 3.685 40.785 ;
        RECT 11.605 40.630 11.775 40.800 ;
        RECT 16.090 40.630 16.260 40.800 ;
        RECT 21.550 40.630 21.720 40.800 ;
        RECT 28.575 40.630 28.745 40.800 ;
        RECT 36.310 40.630 36.480 40.800 ;
        RECT 43.865 40.630 44.035 40.800 ;
        RECT 51.675 40.630 51.845 40.800 ;
        RECT 59.185 40.630 59.355 40.800 ;
        RECT 66.860 40.630 67.030 40.800 ;
        RECT 74.370 40.630 74.540 40.800 ;
        RECT 78.055 40.160 78.225 40.330 ;
        RECT 78.750 40.160 78.920 40.330 ;
        RECT 11.605 39.385 11.775 39.555 ;
        RECT 16.090 39.385 16.260 39.555 ;
        RECT 21.550 39.385 21.720 39.555 ;
        RECT 28.575 39.385 28.745 39.555 ;
        RECT 36.310 39.385 36.480 39.555 ;
        RECT 43.865 39.385 44.035 39.555 ;
        RECT 51.675 39.385 51.845 39.555 ;
        RECT 59.185 39.385 59.355 39.555 ;
        RECT 66.860 39.385 67.030 39.555 ;
        RECT 74.370 39.385 74.540 39.555 ;
        RECT 83.950 40.160 84.120 40.330 ;
        RECT 97.595 40.615 97.765 40.785 ;
        RECT 98.075 40.615 98.245 40.785 ;
        RECT 98.555 40.615 98.725 40.785 ;
        RECT 99.035 40.615 99.205 40.785 ;
        RECT 99.515 40.615 99.685 40.785 ;
        RECT 99.995 40.615 100.165 40.785 ;
        RECT 100.475 40.615 100.645 40.785 ;
        RECT 100.955 40.615 101.125 40.785 ;
        RECT 8.095 38.810 8.265 38.980 ;
        RECT 8.455 38.810 8.625 38.980 ;
        RECT 8.815 38.810 8.985 38.980 ;
        RECT 9.175 38.810 9.345 38.980 ;
        RECT 12.580 38.810 12.750 38.980 ;
        RECT 12.940 38.810 13.110 38.980 ;
        RECT 13.300 38.810 13.470 38.980 ;
        RECT 13.660 38.810 13.830 38.980 ;
        RECT 18.040 38.810 18.210 38.980 ;
        RECT 18.400 38.810 18.570 38.980 ;
        RECT 18.760 38.810 18.930 38.980 ;
        RECT 19.120 38.810 19.290 38.980 ;
        RECT 25.065 38.810 25.235 38.980 ;
        RECT 25.425 38.810 25.595 38.980 ;
        RECT 25.785 38.810 25.955 38.980 ;
        RECT 26.145 38.810 26.315 38.980 ;
        RECT 32.800 38.810 32.970 38.980 ;
        RECT 33.160 38.810 33.330 38.980 ;
        RECT 33.520 38.810 33.690 38.980 ;
        RECT 33.880 38.810 34.050 38.980 ;
        RECT 40.355 38.810 40.525 38.980 ;
        RECT 40.715 38.810 40.885 38.980 ;
        RECT 41.075 38.810 41.245 38.980 ;
        RECT 41.435 38.810 41.605 38.980 ;
        RECT 48.165 38.810 48.335 38.980 ;
        RECT 48.525 38.810 48.695 38.980 ;
        RECT 48.885 38.810 49.055 38.980 ;
        RECT 49.245 38.810 49.415 38.980 ;
        RECT 55.675 38.810 55.845 38.980 ;
        RECT 56.035 38.810 56.205 38.980 ;
        RECT 56.395 38.810 56.565 38.980 ;
        RECT 56.755 38.810 56.925 38.980 ;
        RECT 63.350 38.810 63.520 38.980 ;
        RECT 63.710 38.810 63.880 38.980 ;
        RECT 64.070 38.810 64.240 38.980 ;
        RECT 64.430 38.810 64.600 38.980 ;
        RECT 70.860 38.810 71.030 38.980 ;
        RECT 71.220 38.810 71.390 38.980 ;
        RECT 71.580 38.810 71.750 38.980 ;
        RECT 71.940 38.810 72.110 38.980 ;
        RECT 78.405 38.625 78.575 38.795 ;
        RECT 11.605 38.330 11.775 38.500 ;
        RECT 16.090 38.330 16.260 38.500 ;
        RECT 21.550 38.330 21.720 38.500 ;
        RECT 28.575 38.330 28.745 38.500 ;
        RECT 36.310 38.330 36.480 38.500 ;
        RECT 43.865 38.330 44.035 38.500 ;
        RECT 51.675 38.330 51.845 38.500 ;
        RECT 59.185 38.330 59.355 38.500 ;
        RECT 66.860 38.330 67.030 38.500 ;
        RECT 83.955 38.625 84.125 38.795 ;
        RECT 74.370 38.330 74.540 38.500 ;
        RECT 11.605 37.110 11.775 37.280 ;
        RECT 16.090 37.110 16.260 37.280 ;
        RECT 21.550 37.110 21.720 37.280 ;
        RECT 28.575 37.110 28.745 37.280 ;
        RECT 36.310 37.110 36.480 37.280 ;
        RECT 43.865 37.110 44.035 37.280 ;
        RECT 51.675 37.110 51.845 37.280 ;
        RECT 59.185 37.110 59.355 37.280 ;
        RECT 66.860 37.110 67.030 37.280 ;
        RECT 74.370 37.110 74.540 37.280 ;
        RECT 0.155 36.545 0.325 36.715 ;
        RECT 0.635 36.545 0.805 36.715 ;
        RECT 1.115 36.545 1.285 36.715 ;
        RECT 1.595 36.545 1.765 36.715 ;
        RECT 2.075 36.545 2.245 36.715 ;
        RECT 2.555 36.545 2.725 36.715 ;
        RECT 3.035 36.545 3.205 36.715 ;
        RECT 3.515 36.545 3.685 36.715 ;
        RECT 8.095 36.450 8.265 36.620 ;
        RECT 8.455 36.450 8.625 36.620 ;
        RECT 8.815 36.450 8.985 36.620 ;
        RECT 9.175 36.450 9.345 36.620 ;
        RECT 12.580 36.450 12.750 36.620 ;
        RECT 12.940 36.450 13.110 36.620 ;
        RECT 13.300 36.450 13.470 36.620 ;
        RECT 13.660 36.450 13.830 36.620 ;
        RECT 18.040 36.450 18.210 36.620 ;
        RECT 18.400 36.450 18.570 36.620 ;
        RECT 18.760 36.450 18.930 36.620 ;
        RECT 19.120 36.450 19.290 36.620 ;
        RECT 25.065 36.450 25.235 36.620 ;
        RECT 25.425 36.450 25.595 36.620 ;
        RECT 25.785 36.450 25.955 36.620 ;
        RECT 26.145 36.450 26.315 36.620 ;
        RECT 32.800 36.450 32.970 36.620 ;
        RECT 33.160 36.450 33.330 36.620 ;
        RECT 33.520 36.450 33.690 36.620 ;
        RECT 33.880 36.450 34.050 36.620 ;
        RECT 40.355 36.450 40.525 36.620 ;
        RECT 40.715 36.450 40.885 36.620 ;
        RECT 41.075 36.450 41.245 36.620 ;
        RECT 41.435 36.450 41.605 36.620 ;
        RECT 48.165 36.450 48.335 36.620 ;
        RECT 48.525 36.450 48.695 36.620 ;
        RECT 48.885 36.450 49.055 36.620 ;
        RECT 49.245 36.450 49.415 36.620 ;
        RECT 55.675 36.450 55.845 36.620 ;
        RECT 56.035 36.450 56.205 36.620 ;
        RECT 56.395 36.450 56.565 36.620 ;
        RECT 56.755 36.450 56.925 36.620 ;
        RECT 63.350 36.450 63.520 36.620 ;
        RECT 63.710 36.450 63.880 36.620 ;
        RECT 64.070 36.450 64.240 36.620 ;
        RECT 64.430 36.450 64.600 36.620 ;
        RECT 70.860 36.450 71.030 36.620 ;
        RECT 71.220 36.450 71.390 36.620 ;
        RECT 71.580 36.450 71.750 36.620 ;
        RECT 71.940 36.450 72.110 36.620 ;
        RECT 97.595 36.545 97.765 36.715 ;
        RECT 98.075 36.545 98.245 36.715 ;
        RECT 98.555 36.545 98.725 36.715 ;
        RECT 99.035 36.545 99.205 36.715 ;
        RECT 99.515 36.545 99.685 36.715 ;
        RECT 99.995 36.545 100.165 36.715 ;
        RECT 100.475 36.545 100.645 36.715 ;
        RECT 100.955 36.545 101.125 36.715 ;
        RECT 11.605 36.000 11.775 36.170 ;
        RECT 16.090 36.000 16.260 36.170 ;
        RECT 21.550 36.000 21.720 36.170 ;
        RECT 28.575 36.000 28.745 36.170 ;
        RECT 36.310 36.000 36.480 36.170 ;
        RECT 43.865 36.000 44.035 36.170 ;
        RECT 51.675 36.000 51.845 36.170 ;
        RECT 59.185 36.000 59.355 36.170 ;
        RECT 66.860 36.000 67.030 36.170 ;
        RECT 74.370 36.000 74.540 36.170 ;
        RECT 78.405 35.105 78.575 35.275 ;
        RECT 11.605 34.820 11.775 34.990 ;
        RECT 16.090 34.820 16.260 34.990 ;
        RECT 21.550 34.820 21.720 34.990 ;
        RECT 28.575 34.820 28.745 34.990 ;
        RECT 36.310 34.820 36.480 34.990 ;
        RECT 43.865 34.820 44.035 34.990 ;
        RECT 51.675 34.820 51.845 34.990 ;
        RECT 59.185 34.820 59.355 34.990 ;
        RECT 66.860 34.820 67.030 34.990 ;
        RECT 74.370 34.820 74.540 34.990 ;
        RECT 83.955 35.105 84.125 35.275 ;
        RECT 8.095 34.090 8.265 34.260 ;
        RECT 8.455 34.090 8.625 34.260 ;
        RECT 8.815 34.090 8.985 34.260 ;
        RECT 9.175 34.090 9.345 34.260 ;
        RECT 12.580 34.090 12.750 34.260 ;
        RECT 12.940 34.090 13.110 34.260 ;
        RECT 13.300 34.090 13.470 34.260 ;
        RECT 13.660 34.090 13.830 34.260 ;
        RECT 18.040 34.090 18.210 34.260 ;
        RECT 18.400 34.090 18.570 34.260 ;
        RECT 18.760 34.090 18.930 34.260 ;
        RECT 19.120 34.090 19.290 34.260 ;
        RECT 25.065 34.090 25.235 34.260 ;
        RECT 25.425 34.090 25.595 34.260 ;
        RECT 25.785 34.090 25.955 34.260 ;
        RECT 26.145 34.090 26.315 34.260 ;
        RECT 32.800 34.090 32.970 34.260 ;
        RECT 33.160 34.090 33.330 34.260 ;
        RECT 33.520 34.090 33.690 34.260 ;
        RECT 33.880 34.090 34.050 34.260 ;
        RECT 40.355 34.090 40.525 34.260 ;
        RECT 40.715 34.090 40.885 34.260 ;
        RECT 41.075 34.090 41.245 34.260 ;
        RECT 41.435 34.090 41.605 34.260 ;
        RECT 48.165 34.090 48.335 34.260 ;
        RECT 48.525 34.090 48.695 34.260 ;
        RECT 48.885 34.090 49.055 34.260 ;
        RECT 49.245 34.090 49.415 34.260 ;
        RECT 55.675 34.090 55.845 34.260 ;
        RECT 56.035 34.090 56.205 34.260 ;
        RECT 56.395 34.090 56.565 34.260 ;
        RECT 56.755 34.090 56.925 34.260 ;
        RECT 63.350 34.090 63.520 34.260 ;
        RECT 63.710 34.090 63.880 34.260 ;
        RECT 64.070 34.090 64.240 34.260 ;
        RECT 64.430 34.090 64.600 34.260 ;
        RECT 70.860 34.090 71.030 34.260 ;
        RECT 71.220 34.090 71.390 34.260 ;
        RECT 71.580 34.090 71.750 34.260 ;
        RECT 71.940 34.090 72.110 34.260 ;
        RECT 11.605 33.640 11.775 33.810 ;
        RECT 16.090 33.640 16.260 33.810 ;
        RECT 21.550 33.640 21.720 33.810 ;
        RECT 28.575 33.640 28.745 33.810 ;
        RECT 36.310 33.640 36.480 33.810 ;
        RECT 43.865 33.640 44.035 33.810 ;
        RECT 51.675 33.640 51.845 33.810 ;
        RECT 59.185 33.640 59.355 33.810 ;
        RECT 66.860 33.640 67.030 33.810 ;
        RECT 74.370 33.640 74.540 33.810 ;
        RECT 78.405 33.570 78.575 33.740 ;
        RECT 83.955 33.570 84.125 33.740 ;
        RECT 0.155 32.475 0.325 32.645 ;
        RECT 0.635 32.475 0.805 32.645 ;
        RECT 1.115 32.475 1.285 32.645 ;
        RECT 1.595 32.475 1.765 32.645 ;
        RECT 2.075 32.475 2.245 32.645 ;
        RECT 2.555 32.475 2.725 32.645 ;
        RECT 3.035 32.475 3.205 32.645 ;
        RECT 3.515 32.475 3.685 32.645 ;
        RECT 11.605 32.360 11.775 32.530 ;
        RECT 16.090 32.360 16.260 32.530 ;
        RECT 21.550 32.360 21.720 32.530 ;
        RECT 28.575 32.360 28.745 32.530 ;
        RECT 36.310 32.360 36.480 32.530 ;
        RECT 43.865 32.360 44.035 32.530 ;
        RECT 51.675 32.360 51.845 32.530 ;
        RECT 59.185 32.360 59.355 32.530 ;
        RECT 66.860 32.360 67.030 32.530 ;
        RECT 74.370 32.360 74.540 32.530 ;
        RECT 97.595 32.475 97.765 32.645 ;
        RECT 98.075 32.475 98.245 32.645 ;
        RECT 98.555 32.475 98.725 32.645 ;
        RECT 99.035 32.475 99.205 32.645 ;
        RECT 99.515 32.475 99.685 32.645 ;
        RECT 99.995 32.475 100.165 32.645 ;
        RECT 100.475 32.475 100.645 32.645 ;
        RECT 100.955 32.475 101.125 32.645 ;
        RECT 8.095 31.730 8.265 31.900 ;
        RECT 8.455 31.730 8.625 31.900 ;
        RECT 8.815 31.730 8.985 31.900 ;
        RECT 9.175 31.730 9.345 31.900 ;
        RECT 12.580 31.730 12.750 31.900 ;
        RECT 12.940 31.730 13.110 31.900 ;
        RECT 13.300 31.730 13.470 31.900 ;
        RECT 13.660 31.730 13.830 31.900 ;
        RECT 18.040 31.730 18.210 31.900 ;
        RECT 18.400 31.730 18.570 31.900 ;
        RECT 18.760 31.730 18.930 31.900 ;
        RECT 19.120 31.730 19.290 31.900 ;
        RECT 25.065 31.730 25.235 31.900 ;
        RECT 25.425 31.730 25.595 31.900 ;
        RECT 25.785 31.730 25.955 31.900 ;
        RECT 26.145 31.730 26.315 31.900 ;
        RECT 32.800 31.730 32.970 31.900 ;
        RECT 33.160 31.730 33.330 31.900 ;
        RECT 33.520 31.730 33.690 31.900 ;
        RECT 33.880 31.730 34.050 31.900 ;
        RECT 40.355 31.730 40.525 31.900 ;
        RECT 40.715 31.730 40.885 31.900 ;
        RECT 41.075 31.730 41.245 31.900 ;
        RECT 41.435 31.730 41.605 31.900 ;
        RECT 48.165 31.730 48.335 31.900 ;
        RECT 48.525 31.730 48.695 31.900 ;
        RECT 48.885 31.730 49.055 31.900 ;
        RECT 49.245 31.730 49.415 31.900 ;
        RECT 55.675 31.730 55.845 31.900 ;
        RECT 56.035 31.730 56.205 31.900 ;
        RECT 56.395 31.730 56.565 31.900 ;
        RECT 56.755 31.730 56.925 31.900 ;
        RECT 63.350 31.730 63.520 31.900 ;
        RECT 63.710 31.730 63.880 31.900 ;
        RECT 64.070 31.730 64.240 31.900 ;
        RECT 64.430 31.730 64.600 31.900 ;
        RECT 70.860 31.730 71.030 31.900 ;
        RECT 71.220 31.730 71.390 31.900 ;
        RECT 71.580 31.730 71.750 31.900 ;
        RECT 71.940 31.730 72.110 31.900 ;
        RECT 11.605 31.305 11.775 31.475 ;
        RECT 16.090 31.305 16.260 31.475 ;
        RECT 21.550 31.305 21.720 31.475 ;
        RECT 28.575 31.305 28.745 31.475 ;
        RECT 36.310 31.305 36.480 31.475 ;
        RECT 43.865 31.305 44.035 31.475 ;
        RECT 51.675 31.305 51.845 31.475 ;
        RECT 59.185 31.305 59.355 31.475 ;
        RECT 66.860 31.305 67.030 31.475 ;
        RECT 74.370 31.305 74.540 31.475 ;
        RECT 11.605 30.085 11.775 30.255 ;
        RECT 16.090 30.085 16.260 30.255 ;
        RECT 21.550 30.085 21.720 30.255 ;
        RECT 28.575 30.085 28.745 30.255 ;
        RECT 36.310 30.085 36.480 30.255 ;
        RECT 43.865 30.085 44.035 30.255 ;
        RECT 51.675 30.085 51.845 30.255 ;
        RECT 59.185 30.085 59.355 30.255 ;
        RECT 66.860 30.085 67.030 30.255 ;
        RECT 74.370 30.085 74.540 30.255 ;
        RECT 78.405 30.050 78.575 30.220 ;
        RECT 8.095 29.370 8.265 29.540 ;
        RECT 8.455 29.370 8.625 29.540 ;
        RECT 8.815 29.370 8.985 29.540 ;
        RECT 9.175 29.370 9.345 29.540 ;
        RECT 12.580 29.370 12.750 29.540 ;
        RECT 12.940 29.370 13.110 29.540 ;
        RECT 13.300 29.370 13.470 29.540 ;
        RECT 13.660 29.370 13.830 29.540 ;
        RECT 18.040 29.370 18.210 29.540 ;
        RECT 18.400 29.370 18.570 29.540 ;
        RECT 18.760 29.370 18.930 29.540 ;
        RECT 19.120 29.370 19.290 29.540 ;
        RECT 25.065 29.370 25.235 29.540 ;
        RECT 25.425 29.370 25.595 29.540 ;
        RECT 25.785 29.370 25.955 29.540 ;
        RECT 26.145 29.370 26.315 29.540 ;
        RECT 32.800 29.370 32.970 29.540 ;
        RECT 33.160 29.370 33.330 29.540 ;
        RECT 33.520 29.370 33.690 29.540 ;
        RECT 33.880 29.370 34.050 29.540 ;
        RECT 40.355 29.370 40.525 29.540 ;
        RECT 40.715 29.370 40.885 29.540 ;
        RECT 41.075 29.370 41.245 29.540 ;
        RECT 41.435 29.370 41.605 29.540 ;
        RECT 48.165 29.370 48.335 29.540 ;
        RECT 48.525 29.370 48.695 29.540 ;
        RECT 48.885 29.370 49.055 29.540 ;
        RECT 49.245 29.370 49.415 29.540 ;
        RECT 55.675 29.370 55.845 29.540 ;
        RECT 56.035 29.370 56.205 29.540 ;
        RECT 56.395 29.370 56.565 29.540 ;
        RECT 56.755 29.370 56.925 29.540 ;
        RECT 63.350 29.370 63.520 29.540 ;
        RECT 63.710 29.370 63.880 29.540 ;
        RECT 64.070 29.370 64.240 29.540 ;
        RECT 64.430 29.370 64.600 29.540 ;
        RECT 70.860 29.370 71.030 29.540 ;
        RECT 71.220 29.370 71.390 29.540 ;
        RECT 71.580 29.370 71.750 29.540 ;
        RECT 71.940 29.370 72.110 29.540 ;
        RECT 83.955 30.050 84.125 30.220 ;
        RECT 11.605 28.975 11.775 29.145 ;
        RECT 16.090 28.975 16.260 29.145 ;
        RECT 21.550 28.975 21.720 29.145 ;
        RECT 28.575 28.975 28.745 29.145 ;
        RECT 36.310 28.975 36.480 29.145 ;
        RECT 43.865 28.975 44.035 29.145 ;
        RECT 51.675 28.975 51.845 29.145 ;
        RECT 59.185 28.975 59.355 29.145 ;
        RECT 66.860 28.975 67.030 29.145 ;
        RECT 74.370 28.975 74.540 29.145 ;
        RECT 0.155 28.405 0.325 28.575 ;
        RECT 0.635 28.405 0.805 28.575 ;
        RECT 1.115 28.405 1.285 28.575 ;
        RECT 1.595 28.405 1.765 28.575 ;
        RECT 2.075 28.405 2.245 28.575 ;
        RECT 2.555 28.405 2.725 28.575 ;
        RECT 3.035 28.405 3.205 28.575 ;
        RECT 3.515 28.405 3.685 28.575 ;
        RECT 78.405 28.515 78.575 28.685 ;
        RECT 83.955 28.515 84.125 28.685 ;
        RECT 97.595 28.405 97.765 28.575 ;
        RECT 98.075 28.405 98.245 28.575 ;
        RECT 98.555 28.405 98.725 28.575 ;
        RECT 99.035 28.405 99.205 28.575 ;
        RECT 99.515 28.405 99.685 28.575 ;
        RECT 99.995 28.405 100.165 28.575 ;
        RECT 100.475 28.405 100.645 28.575 ;
        RECT 100.955 28.405 101.125 28.575 ;
        RECT 11.605 27.795 11.775 27.965 ;
        RECT 16.090 27.795 16.260 27.965 ;
        RECT 21.550 27.795 21.720 27.965 ;
        RECT 28.575 27.795 28.745 27.965 ;
        RECT 36.310 27.795 36.480 27.965 ;
        RECT 43.865 27.795 44.035 27.965 ;
        RECT 51.675 27.795 51.845 27.965 ;
        RECT 59.185 27.795 59.355 27.965 ;
        RECT 66.860 27.795 67.030 27.965 ;
        RECT 74.370 27.795 74.540 27.965 ;
        RECT 8.095 27.010 8.265 27.180 ;
        RECT 8.455 27.010 8.625 27.180 ;
        RECT 8.815 27.010 8.985 27.180 ;
        RECT 9.175 27.010 9.345 27.180 ;
        RECT 12.580 27.010 12.750 27.180 ;
        RECT 12.940 27.010 13.110 27.180 ;
        RECT 13.300 27.010 13.470 27.180 ;
        RECT 13.660 27.010 13.830 27.180 ;
        RECT 18.040 27.010 18.210 27.180 ;
        RECT 18.400 27.010 18.570 27.180 ;
        RECT 18.760 27.010 18.930 27.180 ;
        RECT 19.120 27.010 19.290 27.180 ;
        RECT 25.065 27.010 25.235 27.180 ;
        RECT 25.425 27.010 25.595 27.180 ;
        RECT 25.785 27.010 25.955 27.180 ;
        RECT 26.145 27.010 26.315 27.180 ;
        RECT 32.800 27.010 32.970 27.180 ;
        RECT 33.160 27.010 33.330 27.180 ;
        RECT 33.520 27.010 33.690 27.180 ;
        RECT 33.880 27.010 34.050 27.180 ;
        RECT 40.355 27.010 40.525 27.180 ;
        RECT 40.715 27.010 40.885 27.180 ;
        RECT 41.075 27.010 41.245 27.180 ;
        RECT 41.435 27.010 41.605 27.180 ;
        RECT 48.165 27.010 48.335 27.180 ;
        RECT 48.525 27.010 48.695 27.180 ;
        RECT 48.885 27.010 49.055 27.180 ;
        RECT 49.245 27.010 49.415 27.180 ;
        RECT 55.675 27.010 55.845 27.180 ;
        RECT 56.035 27.010 56.205 27.180 ;
        RECT 56.395 27.010 56.565 27.180 ;
        RECT 56.755 27.010 56.925 27.180 ;
        RECT 63.350 27.010 63.520 27.180 ;
        RECT 63.710 27.010 63.880 27.180 ;
        RECT 64.070 27.010 64.240 27.180 ;
        RECT 64.430 27.010 64.600 27.180 ;
        RECT 70.860 27.010 71.030 27.180 ;
        RECT 71.220 27.010 71.390 27.180 ;
        RECT 71.580 27.010 71.750 27.180 ;
        RECT 71.940 27.010 72.110 27.180 ;
        RECT 11.605 26.615 11.775 26.785 ;
        RECT 16.090 26.615 16.260 26.785 ;
        RECT 21.550 26.615 21.720 26.785 ;
        RECT 28.575 26.615 28.745 26.785 ;
        RECT 36.310 26.615 36.480 26.785 ;
        RECT 43.865 26.615 44.035 26.785 ;
        RECT 51.675 26.615 51.845 26.785 ;
        RECT 59.185 26.615 59.355 26.785 ;
        RECT 66.860 26.615 67.030 26.785 ;
        RECT 74.370 26.615 74.540 26.785 ;
        RECT 11.605 25.255 11.775 25.425 ;
        RECT 16.090 25.255 16.260 25.425 ;
        RECT 21.550 25.255 21.720 25.425 ;
        RECT 28.575 25.255 28.745 25.425 ;
        RECT 36.310 25.255 36.480 25.425 ;
        RECT 43.865 25.255 44.035 25.425 ;
        RECT 51.675 25.255 51.845 25.425 ;
        RECT 59.185 25.255 59.355 25.425 ;
        RECT 66.860 25.255 67.030 25.425 ;
        RECT 74.370 25.255 74.540 25.425 ;
        RECT 78.405 24.995 78.575 25.165 ;
        RECT 8.095 24.650 8.265 24.820 ;
        RECT 8.455 24.650 8.625 24.820 ;
        RECT 8.815 24.650 8.985 24.820 ;
        RECT 9.175 24.650 9.345 24.820 ;
        RECT 12.580 24.650 12.750 24.820 ;
        RECT 12.940 24.650 13.110 24.820 ;
        RECT 13.300 24.650 13.470 24.820 ;
        RECT 13.660 24.650 13.830 24.820 ;
        RECT 18.040 24.650 18.210 24.820 ;
        RECT 18.400 24.650 18.570 24.820 ;
        RECT 18.760 24.650 18.930 24.820 ;
        RECT 19.120 24.650 19.290 24.820 ;
        RECT 25.065 24.650 25.235 24.820 ;
        RECT 25.425 24.650 25.595 24.820 ;
        RECT 25.785 24.650 25.955 24.820 ;
        RECT 26.145 24.650 26.315 24.820 ;
        RECT 32.800 24.650 32.970 24.820 ;
        RECT 33.160 24.650 33.330 24.820 ;
        RECT 33.520 24.650 33.690 24.820 ;
        RECT 33.880 24.650 34.050 24.820 ;
        RECT 40.355 24.650 40.525 24.820 ;
        RECT 40.715 24.650 40.885 24.820 ;
        RECT 41.075 24.650 41.245 24.820 ;
        RECT 41.435 24.650 41.605 24.820 ;
        RECT 48.165 24.650 48.335 24.820 ;
        RECT 48.525 24.650 48.695 24.820 ;
        RECT 48.885 24.650 49.055 24.820 ;
        RECT 49.245 24.650 49.415 24.820 ;
        RECT 55.675 24.650 55.845 24.820 ;
        RECT 56.035 24.650 56.205 24.820 ;
        RECT 56.395 24.650 56.565 24.820 ;
        RECT 56.755 24.650 56.925 24.820 ;
        RECT 63.350 24.650 63.520 24.820 ;
        RECT 63.710 24.650 63.880 24.820 ;
        RECT 64.070 24.650 64.240 24.820 ;
        RECT 64.430 24.650 64.600 24.820 ;
        RECT 70.860 24.650 71.030 24.820 ;
        RECT 71.220 24.650 71.390 24.820 ;
        RECT 71.580 24.650 71.750 24.820 ;
        RECT 71.940 24.650 72.110 24.820 ;
        RECT 0.155 24.335 0.325 24.505 ;
        RECT 0.635 24.335 0.805 24.505 ;
        RECT 1.115 24.335 1.285 24.505 ;
        RECT 1.595 24.335 1.765 24.505 ;
        RECT 2.075 24.335 2.245 24.505 ;
        RECT 2.555 24.335 2.725 24.505 ;
        RECT 3.035 24.335 3.205 24.505 ;
        RECT 3.515 24.335 3.685 24.505 ;
        RECT 11.605 24.200 11.775 24.370 ;
        RECT 16.090 24.200 16.260 24.370 ;
        RECT 21.550 24.200 21.720 24.370 ;
        RECT 28.575 24.200 28.745 24.370 ;
        RECT 36.310 24.200 36.480 24.370 ;
        RECT 43.865 24.200 44.035 24.370 ;
        RECT 51.675 24.200 51.845 24.370 ;
        RECT 59.185 24.200 59.355 24.370 ;
        RECT 66.860 24.200 67.030 24.370 ;
        RECT 83.955 24.995 84.125 25.165 ;
        RECT 74.370 24.200 74.540 24.370 ;
        RECT 97.595 24.335 97.765 24.505 ;
        RECT 98.075 24.335 98.245 24.505 ;
        RECT 98.555 24.335 98.725 24.505 ;
        RECT 99.035 24.335 99.205 24.505 ;
        RECT 99.515 24.335 99.685 24.505 ;
        RECT 99.995 24.335 100.165 24.505 ;
        RECT 100.475 24.335 100.645 24.505 ;
        RECT 100.955 24.335 101.125 24.505 ;
        RECT 78.405 23.460 78.575 23.630 ;
        RECT 83.955 23.460 84.125 23.630 ;
        RECT 11.605 22.980 11.775 23.150 ;
        RECT 16.090 22.980 16.260 23.150 ;
        RECT 21.550 22.980 21.720 23.150 ;
        RECT 28.575 22.980 28.745 23.150 ;
        RECT 36.310 22.980 36.480 23.150 ;
        RECT 43.865 22.980 44.035 23.150 ;
        RECT 51.675 22.980 51.845 23.150 ;
        RECT 59.185 22.980 59.355 23.150 ;
        RECT 66.860 22.980 67.030 23.150 ;
        RECT 74.370 22.980 74.540 23.150 ;
        RECT 8.095 22.290 8.265 22.460 ;
        RECT 8.455 22.290 8.625 22.460 ;
        RECT 8.815 22.290 8.985 22.460 ;
        RECT 9.175 22.290 9.345 22.460 ;
        RECT 12.580 22.290 12.750 22.460 ;
        RECT 12.940 22.290 13.110 22.460 ;
        RECT 13.300 22.290 13.470 22.460 ;
        RECT 13.660 22.290 13.830 22.460 ;
        RECT 18.040 22.290 18.210 22.460 ;
        RECT 18.400 22.290 18.570 22.460 ;
        RECT 18.760 22.290 18.930 22.460 ;
        RECT 19.120 22.290 19.290 22.460 ;
        RECT 25.065 22.290 25.235 22.460 ;
        RECT 25.425 22.290 25.595 22.460 ;
        RECT 25.785 22.290 25.955 22.460 ;
        RECT 26.145 22.290 26.315 22.460 ;
        RECT 32.800 22.290 32.970 22.460 ;
        RECT 33.160 22.290 33.330 22.460 ;
        RECT 33.520 22.290 33.690 22.460 ;
        RECT 33.880 22.290 34.050 22.460 ;
        RECT 40.355 22.290 40.525 22.460 ;
        RECT 40.715 22.290 40.885 22.460 ;
        RECT 41.075 22.290 41.245 22.460 ;
        RECT 41.435 22.290 41.605 22.460 ;
        RECT 48.165 22.290 48.335 22.460 ;
        RECT 48.525 22.290 48.695 22.460 ;
        RECT 48.885 22.290 49.055 22.460 ;
        RECT 49.245 22.290 49.415 22.460 ;
        RECT 55.675 22.290 55.845 22.460 ;
        RECT 56.035 22.290 56.205 22.460 ;
        RECT 56.395 22.290 56.565 22.460 ;
        RECT 56.755 22.290 56.925 22.460 ;
        RECT 63.350 22.290 63.520 22.460 ;
        RECT 63.710 22.290 63.880 22.460 ;
        RECT 64.070 22.290 64.240 22.460 ;
        RECT 64.430 22.290 64.600 22.460 ;
        RECT 70.860 22.290 71.030 22.460 ;
        RECT 71.220 22.290 71.390 22.460 ;
        RECT 71.580 22.290 71.750 22.460 ;
        RECT 71.940 22.290 72.110 22.460 ;
        RECT 11.605 21.870 11.775 22.040 ;
        RECT 16.090 21.870 16.260 22.040 ;
        RECT 21.550 21.870 21.720 22.040 ;
        RECT 28.575 21.870 28.745 22.040 ;
        RECT 36.310 21.870 36.480 22.040 ;
        RECT 43.865 21.870 44.035 22.040 ;
        RECT 51.675 21.870 51.845 22.040 ;
        RECT 59.185 21.870 59.355 22.040 ;
        RECT 66.860 21.870 67.030 22.040 ;
        RECT 74.370 21.870 74.540 22.040 ;
        RECT 11.605 20.690 11.775 20.860 ;
        RECT 16.090 20.690 16.260 20.860 ;
        RECT 21.550 20.690 21.720 20.860 ;
        RECT 28.575 20.690 28.745 20.860 ;
        RECT 36.310 20.690 36.480 20.860 ;
        RECT 43.865 20.690 44.035 20.860 ;
        RECT 51.675 20.690 51.845 20.860 ;
        RECT 59.185 20.690 59.355 20.860 ;
        RECT 66.860 20.690 67.030 20.860 ;
        RECT 74.370 20.690 74.540 20.860 ;
        RECT 0.155 20.265 0.325 20.435 ;
        RECT 0.635 20.265 0.805 20.435 ;
        RECT 1.115 20.265 1.285 20.435 ;
        RECT 1.595 20.265 1.765 20.435 ;
        RECT 2.075 20.265 2.245 20.435 ;
        RECT 2.555 20.265 2.725 20.435 ;
        RECT 3.035 20.265 3.205 20.435 ;
        RECT 3.515 20.265 3.685 20.435 ;
        RECT 8.095 19.930 8.265 20.100 ;
        RECT 8.455 19.930 8.625 20.100 ;
        RECT 8.815 19.930 8.985 20.100 ;
        RECT 9.175 19.930 9.345 20.100 ;
        RECT 12.580 19.930 12.750 20.100 ;
        RECT 12.940 19.930 13.110 20.100 ;
        RECT 13.300 19.930 13.470 20.100 ;
        RECT 13.660 19.930 13.830 20.100 ;
        RECT 18.040 19.930 18.210 20.100 ;
        RECT 18.400 19.930 18.570 20.100 ;
        RECT 18.760 19.930 18.930 20.100 ;
        RECT 19.120 19.930 19.290 20.100 ;
        RECT 25.065 19.930 25.235 20.100 ;
        RECT 25.425 19.930 25.595 20.100 ;
        RECT 25.785 19.930 25.955 20.100 ;
        RECT 26.145 19.930 26.315 20.100 ;
        RECT 32.800 19.930 32.970 20.100 ;
        RECT 33.160 19.930 33.330 20.100 ;
        RECT 33.520 19.930 33.690 20.100 ;
        RECT 33.880 19.930 34.050 20.100 ;
        RECT 40.355 19.930 40.525 20.100 ;
        RECT 40.715 19.930 40.885 20.100 ;
        RECT 41.075 19.930 41.245 20.100 ;
        RECT 41.435 19.930 41.605 20.100 ;
        RECT 48.165 19.930 48.335 20.100 ;
        RECT 48.525 19.930 48.695 20.100 ;
        RECT 48.885 19.930 49.055 20.100 ;
        RECT 49.245 19.930 49.415 20.100 ;
        RECT 55.675 19.930 55.845 20.100 ;
        RECT 56.035 19.930 56.205 20.100 ;
        RECT 56.395 19.930 56.565 20.100 ;
        RECT 56.755 19.930 56.925 20.100 ;
        RECT 63.350 19.930 63.520 20.100 ;
        RECT 63.710 19.930 63.880 20.100 ;
        RECT 64.070 19.930 64.240 20.100 ;
        RECT 64.430 19.930 64.600 20.100 ;
        RECT 70.860 19.930 71.030 20.100 ;
        RECT 71.220 19.930 71.390 20.100 ;
        RECT 71.580 19.930 71.750 20.100 ;
        RECT 71.940 19.930 72.110 20.100 ;
        RECT 78.405 19.940 78.575 20.110 ;
        RECT 11.605 19.510 11.775 19.680 ;
        RECT 16.090 19.510 16.260 19.680 ;
        RECT 21.550 19.510 21.720 19.680 ;
        RECT 28.575 19.510 28.745 19.680 ;
        RECT 36.310 19.510 36.480 19.680 ;
        RECT 43.865 19.510 44.035 19.680 ;
        RECT 51.675 19.510 51.845 19.680 ;
        RECT 59.185 19.510 59.355 19.680 ;
        RECT 66.860 19.510 67.030 19.680 ;
        RECT 74.370 19.510 74.540 19.680 ;
        RECT 83.955 19.940 84.125 20.110 ;
        RECT 89.625 19.940 89.795 20.110 ;
        RECT 97.595 20.265 97.765 20.435 ;
        RECT 98.075 20.265 98.245 20.435 ;
        RECT 98.555 20.265 98.725 20.435 ;
        RECT 99.035 20.265 99.205 20.435 ;
        RECT 99.515 20.265 99.685 20.435 ;
        RECT 99.995 20.265 100.165 20.435 ;
        RECT 100.475 20.265 100.645 20.435 ;
        RECT 100.955 20.265 101.125 20.435 ;
        RECT 78.405 18.405 78.575 18.575 ;
        RECT 11.605 18.125 11.775 18.295 ;
        RECT 16.090 18.125 16.260 18.295 ;
        RECT 21.550 18.125 21.720 18.295 ;
        RECT 28.575 18.125 28.745 18.295 ;
        RECT 36.310 18.125 36.480 18.295 ;
        RECT 43.865 18.125 44.035 18.295 ;
        RECT 51.675 18.125 51.845 18.295 ;
        RECT 59.185 18.125 59.355 18.295 ;
        RECT 66.860 18.125 67.030 18.295 ;
        RECT 83.955 18.405 84.125 18.575 ;
        RECT 89.625 18.405 89.795 18.575 ;
        RECT 74.370 18.125 74.540 18.295 ;
        RECT 8.095 17.570 8.265 17.740 ;
        RECT 8.455 17.570 8.625 17.740 ;
        RECT 8.815 17.570 8.985 17.740 ;
        RECT 9.175 17.570 9.345 17.740 ;
        RECT 12.580 17.570 12.750 17.740 ;
        RECT 12.940 17.570 13.110 17.740 ;
        RECT 13.300 17.570 13.470 17.740 ;
        RECT 13.660 17.570 13.830 17.740 ;
        RECT 18.040 17.570 18.210 17.740 ;
        RECT 18.400 17.570 18.570 17.740 ;
        RECT 18.760 17.570 18.930 17.740 ;
        RECT 19.120 17.570 19.290 17.740 ;
        RECT 25.065 17.570 25.235 17.740 ;
        RECT 25.425 17.570 25.595 17.740 ;
        RECT 25.785 17.570 25.955 17.740 ;
        RECT 26.145 17.570 26.315 17.740 ;
        RECT 32.800 17.570 32.970 17.740 ;
        RECT 33.160 17.570 33.330 17.740 ;
        RECT 33.520 17.570 33.690 17.740 ;
        RECT 33.880 17.570 34.050 17.740 ;
        RECT 40.355 17.570 40.525 17.740 ;
        RECT 40.715 17.570 40.885 17.740 ;
        RECT 41.075 17.570 41.245 17.740 ;
        RECT 41.435 17.570 41.605 17.740 ;
        RECT 48.165 17.570 48.335 17.740 ;
        RECT 48.525 17.570 48.695 17.740 ;
        RECT 48.885 17.570 49.055 17.740 ;
        RECT 49.245 17.570 49.415 17.740 ;
        RECT 55.675 17.570 55.845 17.740 ;
        RECT 56.035 17.570 56.205 17.740 ;
        RECT 56.395 17.570 56.565 17.740 ;
        RECT 56.755 17.570 56.925 17.740 ;
        RECT 63.350 17.570 63.520 17.740 ;
        RECT 63.710 17.570 63.880 17.740 ;
        RECT 64.070 17.570 64.240 17.740 ;
        RECT 64.430 17.570 64.600 17.740 ;
        RECT 70.860 17.570 71.030 17.740 ;
        RECT 71.220 17.570 71.390 17.740 ;
        RECT 71.580 17.570 71.750 17.740 ;
        RECT 71.940 17.570 72.110 17.740 ;
        RECT 11.605 17.070 11.775 17.240 ;
        RECT 16.090 17.070 16.260 17.240 ;
        RECT 21.550 17.070 21.720 17.240 ;
        RECT 28.575 17.070 28.745 17.240 ;
        RECT 36.310 17.070 36.480 17.240 ;
        RECT 43.865 17.070 44.035 17.240 ;
        RECT 51.675 17.070 51.845 17.240 ;
        RECT 59.185 17.070 59.355 17.240 ;
        RECT 66.860 17.070 67.030 17.240 ;
        RECT 74.370 17.070 74.540 17.240 ;
        RECT 0.155 16.195 0.325 16.365 ;
        RECT 0.635 16.195 0.805 16.365 ;
        RECT 1.115 16.195 1.285 16.365 ;
        RECT 1.595 16.195 1.765 16.365 ;
        RECT 2.075 16.195 2.245 16.365 ;
        RECT 2.555 16.195 2.725 16.365 ;
        RECT 3.035 16.195 3.205 16.365 ;
        RECT 3.515 16.195 3.685 16.365 ;
        RECT 97.595 16.195 97.765 16.365 ;
        RECT 98.075 16.195 98.245 16.365 ;
        RECT 98.555 16.195 98.725 16.365 ;
        RECT 99.035 16.195 99.205 16.365 ;
        RECT 99.515 16.195 99.685 16.365 ;
        RECT 99.995 16.195 100.165 16.365 ;
        RECT 100.475 16.195 100.645 16.365 ;
        RECT 100.955 16.195 101.125 16.365 ;
        RECT 11.605 15.850 11.775 16.020 ;
        RECT 16.090 15.850 16.260 16.020 ;
        RECT 21.550 15.850 21.720 16.020 ;
        RECT 28.575 15.850 28.745 16.020 ;
        RECT 36.310 15.850 36.480 16.020 ;
        RECT 43.865 15.850 44.035 16.020 ;
        RECT 51.675 15.850 51.845 16.020 ;
        RECT 59.185 15.850 59.355 16.020 ;
        RECT 66.860 15.850 67.030 16.020 ;
        RECT 74.370 15.850 74.540 16.020 ;
        RECT 8.095 15.210 8.265 15.380 ;
        RECT 8.455 15.210 8.625 15.380 ;
        RECT 8.815 15.210 8.985 15.380 ;
        RECT 9.175 15.210 9.345 15.380 ;
        RECT 12.580 15.210 12.750 15.380 ;
        RECT 12.940 15.210 13.110 15.380 ;
        RECT 13.300 15.210 13.470 15.380 ;
        RECT 13.660 15.210 13.830 15.380 ;
        RECT 18.040 15.210 18.210 15.380 ;
        RECT 18.400 15.210 18.570 15.380 ;
        RECT 18.760 15.210 18.930 15.380 ;
        RECT 19.120 15.210 19.290 15.380 ;
        RECT 25.065 15.210 25.235 15.380 ;
        RECT 25.425 15.210 25.595 15.380 ;
        RECT 25.785 15.210 25.955 15.380 ;
        RECT 26.145 15.210 26.315 15.380 ;
        RECT 32.800 15.210 32.970 15.380 ;
        RECT 33.160 15.210 33.330 15.380 ;
        RECT 33.520 15.210 33.690 15.380 ;
        RECT 33.880 15.210 34.050 15.380 ;
        RECT 40.355 15.210 40.525 15.380 ;
        RECT 40.715 15.210 40.885 15.380 ;
        RECT 41.075 15.210 41.245 15.380 ;
        RECT 41.435 15.210 41.605 15.380 ;
        RECT 48.165 15.210 48.335 15.380 ;
        RECT 48.525 15.210 48.695 15.380 ;
        RECT 48.885 15.210 49.055 15.380 ;
        RECT 49.245 15.210 49.415 15.380 ;
        RECT 55.675 15.210 55.845 15.380 ;
        RECT 56.035 15.210 56.205 15.380 ;
        RECT 56.395 15.210 56.565 15.380 ;
        RECT 56.755 15.210 56.925 15.380 ;
        RECT 63.350 15.210 63.520 15.380 ;
        RECT 63.710 15.210 63.880 15.380 ;
        RECT 64.070 15.210 64.240 15.380 ;
        RECT 64.430 15.210 64.600 15.380 ;
        RECT 70.860 15.210 71.030 15.380 ;
        RECT 71.220 15.210 71.390 15.380 ;
        RECT 71.580 15.210 71.750 15.380 ;
        RECT 71.940 15.210 72.110 15.380 ;
        RECT 11.605 14.740 11.775 14.910 ;
        RECT 16.090 14.740 16.260 14.910 ;
        RECT 21.550 14.740 21.720 14.910 ;
        RECT 28.575 14.740 28.745 14.910 ;
        RECT 36.310 14.740 36.480 14.910 ;
        RECT 43.865 14.740 44.035 14.910 ;
        RECT 51.675 14.740 51.845 14.910 ;
        RECT 59.185 14.740 59.355 14.910 ;
        RECT 66.860 14.740 67.030 14.910 ;
        RECT 74.370 14.740 74.540 14.910 ;
        RECT 78.405 14.885 78.575 15.055 ;
        RECT 83.955 14.885 84.125 15.055 ;
        RECT 89.625 14.885 89.795 15.055 ;
        RECT 11.605 13.560 11.775 13.730 ;
        RECT 16.090 13.560 16.260 13.730 ;
        RECT 21.550 13.560 21.720 13.730 ;
        RECT 28.575 13.560 28.745 13.730 ;
        RECT 36.310 13.560 36.480 13.730 ;
        RECT 43.865 13.560 44.035 13.730 ;
        RECT 51.675 13.560 51.845 13.730 ;
        RECT 59.185 13.560 59.355 13.730 ;
        RECT 66.860 13.560 67.030 13.730 ;
        RECT 74.370 13.560 74.540 13.730 ;
        RECT 78.405 13.350 78.575 13.520 ;
        RECT 83.955 13.350 84.125 13.520 ;
        RECT 8.095 12.850 8.265 13.020 ;
        RECT 8.455 12.850 8.625 13.020 ;
        RECT 8.815 12.850 8.985 13.020 ;
        RECT 9.175 12.850 9.345 13.020 ;
        RECT 12.580 12.850 12.750 13.020 ;
        RECT 12.940 12.850 13.110 13.020 ;
        RECT 13.300 12.850 13.470 13.020 ;
        RECT 13.660 12.850 13.830 13.020 ;
        RECT 18.040 12.850 18.210 13.020 ;
        RECT 18.400 12.850 18.570 13.020 ;
        RECT 18.760 12.850 18.930 13.020 ;
        RECT 19.120 12.850 19.290 13.020 ;
        RECT 25.065 12.850 25.235 13.020 ;
        RECT 25.425 12.850 25.595 13.020 ;
        RECT 25.785 12.850 25.955 13.020 ;
        RECT 26.145 12.850 26.315 13.020 ;
        RECT 32.800 12.850 32.970 13.020 ;
        RECT 33.160 12.850 33.330 13.020 ;
        RECT 33.520 12.850 33.690 13.020 ;
        RECT 33.880 12.850 34.050 13.020 ;
        RECT 40.355 12.850 40.525 13.020 ;
        RECT 40.715 12.850 40.885 13.020 ;
        RECT 41.075 12.850 41.245 13.020 ;
        RECT 41.435 12.850 41.605 13.020 ;
        RECT 48.165 12.850 48.335 13.020 ;
        RECT 48.525 12.850 48.695 13.020 ;
        RECT 48.885 12.850 49.055 13.020 ;
        RECT 49.245 12.850 49.415 13.020 ;
        RECT 55.675 12.850 55.845 13.020 ;
        RECT 56.035 12.850 56.205 13.020 ;
        RECT 56.395 12.850 56.565 13.020 ;
        RECT 56.755 12.850 56.925 13.020 ;
        RECT 63.350 12.850 63.520 13.020 ;
        RECT 63.710 12.850 63.880 13.020 ;
        RECT 64.070 12.850 64.240 13.020 ;
        RECT 64.430 12.850 64.600 13.020 ;
        RECT 70.860 12.850 71.030 13.020 ;
        RECT 71.220 12.850 71.390 13.020 ;
        RECT 71.580 12.850 71.750 13.020 ;
        RECT 71.940 12.850 72.110 13.020 ;
        RECT 11.605 12.380 11.775 12.550 ;
        RECT 16.090 12.380 16.260 12.550 ;
        RECT 21.550 12.380 21.720 12.550 ;
        RECT 28.575 12.380 28.745 12.550 ;
        RECT 36.310 12.380 36.480 12.550 ;
        RECT 43.865 12.380 44.035 12.550 ;
        RECT 51.675 12.380 51.845 12.550 ;
        RECT 59.185 12.380 59.355 12.550 ;
        RECT 66.860 12.380 67.030 12.550 ;
        RECT 74.370 12.380 74.540 12.550 ;
        RECT 0.155 12.125 0.325 12.295 ;
        RECT 0.635 12.125 0.805 12.295 ;
        RECT 1.115 12.125 1.285 12.295 ;
        RECT 1.595 12.125 1.765 12.295 ;
        RECT 2.075 12.125 2.245 12.295 ;
        RECT 2.555 12.125 2.725 12.295 ;
        RECT 3.035 12.125 3.205 12.295 ;
        RECT 3.515 12.125 3.685 12.295 ;
        RECT 97.595 12.125 97.765 12.295 ;
        RECT 98.075 12.125 98.245 12.295 ;
        RECT 98.555 12.125 98.725 12.295 ;
        RECT 99.035 12.125 99.205 12.295 ;
        RECT 99.515 12.125 99.685 12.295 ;
        RECT 99.995 12.125 100.165 12.295 ;
        RECT 100.475 12.125 100.645 12.295 ;
        RECT 100.955 12.125 101.125 12.295 ;
        RECT 0.155 8.055 0.325 8.225 ;
        RECT 0.635 8.055 0.805 8.225 ;
        RECT 1.115 8.055 1.285 8.225 ;
        RECT 1.595 8.055 1.765 8.225 ;
        RECT 2.075 8.055 2.245 8.225 ;
        RECT 2.555 8.055 2.725 8.225 ;
        RECT 3.035 8.055 3.205 8.225 ;
        RECT 3.515 8.055 3.685 8.225 ;
        RECT 97.595 8.055 97.765 8.225 ;
        RECT 98.075 8.055 98.245 8.225 ;
        RECT 98.555 8.055 98.725 8.225 ;
        RECT 99.035 8.055 99.205 8.225 ;
        RECT 99.515 8.055 99.685 8.225 ;
        RECT 99.995 8.055 100.165 8.225 ;
        RECT 100.475 8.055 100.645 8.225 ;
        RECT 100.955 8.055 101.125 8.225 ;
        RECT 0.155 3.985 0.325 4.155 ;
        RECT 0.635 3.985 0.805 4.155 ;
        RECT 1.115 3.985 1.285 4.155 ;
        RECT 1.595 3.985 1.765 4.155 ;
        RECT 2.075 3.985 2.245 4.155 ;
        RECT 2.555 3.985 2.725 4.155 ;
        RECT 3.035 3.985 3.205 4.155 ;
        RECT 3.515 3.985 3.685 4.155 ;
        RECT 3.995 3.985 4.165 4.155 ;
        RECT 4.475 3.985 4.645 4.155 ;
        RECT 4.955 3.985 5.125 4.155 ;
        RECT 5.435 3.985 5.605 4.155 ;
        RECT 5.915 3.985 6.085 4.155 ;
        RECT 6.395 3.985 6.565 4.155 ;
        RECT 6.875 3.985 7.045 4.155 ;
        RECT 7.355 3.985 7.525 4.155 ;
        RECT 7.835 3.985 8.005 4.155 ;
        RECT 8.315 3.985 8.485 4.155 ;
        RECT 8.795 3.985 8.965 4.155 ;
        RECT 9.275 3.985 9.445 4.155 ;
        RECT 9.755 3.985 9.925 4.155 ;
        RECT 10.235 3.985 10.405 4.155 ;
        RECT 10.715 3.985 10.885 4.155 ;
        RECT 11.195 3.985 11.365 4.155 ;
        RECT 11.675 3.985 11.845 4.155 ;
        RECT 12.155 3.985 12.325 4.155 ;
        RECT 12.635 3.985 12.805 4.155 ;
        RECT 13.115 3.985 13.285 4.155 ;
        RECT 13.595 3.985 13.765 4.155 ;
        RECT 14.075 3.985 14.245 4.155 ;
        RECT 14.555 3.985 14.725 4.155 ;
        RECT 15.035 3.985 15.205 4.155 ;
        RECT 15.515 3.985 15.685 4.155 ;
        RECT 15.995 3.985 16.165 4.155 ;
        RECT 16.475 3.985 16.645 4.155 ;
        RECT 16.955 3.985 17.125 4.155 ;
        RECT 17.435 3.985 17.605 4.155 ;
        RECT 17.915 3.985 18.085 4.155 ;
        RECT 18.395 3.985 18.565 4.155 ;
        RECT 18.875 3.985 19.045 4.155 ;
        RECT 19.355 3.985 19.525 4.155 ;
        RECT 19.835 3.985 20.005 4.155 ;
        RECT 20.315 3.985 20.485 4.155 ;
        RECT 20.795 3.985 20.965 4.155 ;
        RECT 21.275 3.985 21.445 4.155 ;
        RECT 21.755 3.985 21.925 4.155 ;
        RECT 22.235 3.985 22.405 4.155 ;
        RECT 22.715 3.985 22.885 4.155 ;
        RECT 23.195 3.985 23.365 4.155 ;
        RECT 23.675 3.985 23.845 4.155 ;
        RECT 24.155 3.985 24.325 4.155 ;
        RECT 24.635 3.985 24.805 4.155 ;
        RECT 25.115 3.985 25.285 4.155 ;
        RECT 25.595 3.985 25.765 4.155 ;
        RECT 26.075 3.985 26.245 4.155 ;
        RECT 26.555 3.985 26.725 4.155 ;
        RECT 27.035 3.985 27.205 4.155 ;
        RECT 27.515 3.985 27.685 4.155 ;
        RECT 27.995 3.985 28.165 4.155 ;
        RECT 28.475 3.985 28.645 4.155 ;
        RECT 28.955 3.985 29.125 4.155 ;
        RECT 29.435 3.985 29.605 4.155 ;
        RECT 29.915 3.985 30.085 4.155 ;
        RECT 30.395 3.985 30.565 4.155 ;
        RECT 30.875 3.985 31.045 4.155 ;
        RECT 31.355 3.985 31.525 4.155 ;
        RECT 31.835 3.985 32.005 4.155 ;
        RECT 32.315 3.985 32.485 4.155 ;
        RECT 32.795 3.985 32.965 4.155 ;
        RECT 33.275 3.985 33.445 4.155 ;
        RECT 33.755 3.985 33.925 4.155 ;
        RECT 34.235 3.985 34.405 4.155 ;
        RECT 34.715 3.985 34.885 4.155 ;
        RECT 35.195 3.985 35.365 4.155 ;
        RECT 35.675 3.985 35.845 4.155 ;
        RECT 36.155 3.985 36.325 4.155 ;
        RECT 36.635 3.985 36.805 4.155 ;
        RECT 37.115 3.985 37.285 4.155 ;
        RECT 37.595 3.985 37.765 4.155 ;
        RECT 38.075 3.985 38.245 4.155 ;
        RECT 38.555 3.985 38.725 4.155 ;
        RECT 39.035 3.985 39.205 4.155 ;
        RECT 39.515 3.985 39.685 4.155 ;
        RECT 39.995 3.985 40.165 4.155 ;
        RECT 40.475 3.985 40.645 4.155 ;
        RECT 40.955 3.985 41.125 4.155 ;
        RECT 41.435 3.985 41.605 4.155 ;
        RECT 41.915 3.985 42.085 4.155 ;
        RECT 42.395 3.985 42.565 4.155 ;
        RECT 42.875 3.985 43.045 4.155 ;
        RECT 43.355 3.985 43.525 4.155 ;
        RECT 43.835 3.985 44.005 4.155 ;
        RECT 44.315 3.985 44.485 4.155 ;
        RECT 44.795 3.985 44.965 4.155 ;
        RECT 45.275 3.985 45.445 4.155 ;
        RECT 45.755 3.985 45.925 4.155 ;
        RECT 46.235 3.985 46.405 4.155 ;
        RECT 46.715 3.985 46.885 4.155 ;
        RECT 47.195 3.985 47.365 4.155 ;
        RECT 47.675 3.985 47.845 4.155 ;
        RECT 48.155 3.985 48.325 4.155 ;
        RECT 48.635 3.985 48.805 4.155 ;
        RECT 49.115 3.985 49.285 4.155 ;
        RECT 49.595 3.985 49.765 4.155 ;
        RECT 50.075 3.985 50.245 4.155 ;
        RECT 50.555 3.985 50.725 4.155 ;
        RECT 51.035 3.985 51.205 4.155 ;
        RECT 51.515 3.985 51.685 4.155 ;
        RECT 51.995 3.985 52.165 4.155 ;
        RECT 52.475 3.985 52.645 4.155 ;
        RECT 52.955 3.985 53.125 4.155 ;
        RECT 53.435 3.985 53.605 4.155 ;
        RECT 53.915 3.985 54.085 4.155 ;
        RECT 54.395 3.985 54.565 4.155 ;
        RECT 54.875 3.985 55.045 4.155 ;
        RECT 55.355 3.985 55.525 4.155 ;
        RECT 55.835 3.985 56.005 4.155 ;
        RECT 56.315 3.985 56.485 4.155 ;
        RECT 56.795 3.985 56.965 4.155 ;
        RECT 57.275 3.985 57.445 4.155 ;
        RECT 57.755 3.985 57.925 4.155 ;
        RECT 58.235 3.985 58.405 4.155 ;
        RECT 58.715 3.985 58.885 4.155 ;
        RECT 59.195 3.985 59.365 4.155 ;
        RECT 59.675 3.985 59.845 4.155 ;
        RECT 60.155 3.985 60.325 4.155 ;
        RECT 60.635 3.985 60.805 4.155 ;
        RECT 61.115 3.985 61.285 4.155 ;
        RECT 61.595 3.985 61.765 4.155 ;
        RECT 62.075 3.985 62.245 4.155 ;
        RECT 62.555 3.985 62.725 4.155 ;
        RECT 63.035 3.985 63.205 4.155 ;
        RECT 63.515 3.985 63.685 4.155 ;
        RECT 63.995 3.985 64.165 4.155 ;
        RECT 64.475 3.985 64.645 4.155 ;
        RECT 64.955 3.985 65.125 4.155 ;
        RECT 65.435 3.985 65.605 4.155 ;
        RECT 65.915 3.985 66.085 4.155 ;
        RECT 66.395 3.985 66.565 4.155 ;
        RECT 66.875 3.985 67.045 4.155 ;
        RECT 67.355 3.985 67.525 4.155 ;
        RECT 67.835 3.985 68.005 4.155 ;
        RECT 68.315 3.985 68.485 4.155 ;
        RECT 68.795 3.985 68.965 4.155 ;
        RECT 69.275 3.985 69.445 4.155 ;
        RECT 69.755 3.985 69.925 4.155 ;
        RECT 70.235 3.985 70.405 4.155 ;
        RECT 70.715 3.985 70.885 4.155 ;
        RECT 71.195 3.985 71.365 4.155 ;
        RECT 71.675 3.985 71.845 4.155 ;
        RECT 72.155 3.985 72.325 4.155 ;
        RECT 72.635 3.985 72.805 4.155 ;
        RECT 73.115 3.985 73.285 4.155 ;
        RECT 73.595 3.985 73.765 4.155 ;
        RECT 74.075 3.985 74.245 4.155 ;
        RECT 74.555 3.985 74.725 4.155 ;
        RECT 75.035 3.985 75.205 4.155 ;
        RECT 75.515 3.985 75.685 4.155 ;
        RECT 75.995 3.985 76.165 4.155 ;
        RECT 76.475 3.985 76.645 4.155 ;
        RECT 76.955 3.985 77.125 4.155 ;
        RECT 77.435 3.985 77.605 4.155 ;
        RECT 77.915 3.985 78.085 4.155 ;
        RECT 78.395 3.985 78.565 4.155 ;
        RECT 78.875 3.985 79.045 4.155 ;
        RECT 79.355 3.985 79.525 4.155 ;
        RECT 79.835 3.985 80.005 4.155 ;
        RECT 80.315 3.985 80.485 4.155 ;
        RECT 80.795 3.985 80.965 4.155 ;
        RECT 81.275 3.985 81.445 4.155 ;
        RECT 81.755 3.985 81.925 4.155 ;
        RECT 82.235 3.985 82.405 4.155 ;
        RECT 82.715 3.985 82.885 4.155 ;
        RECT 83.195 3.985 83.365 4.155 ;
        RECT 83.675 3.985 83.845 4.155 ;
        RECT 84.155 3.985 84.325 4.155 ;
        RECT 84.635 3.985 84.805 4.155 ;
        RECT 85.115 3.985 85.285 4.155 ;
        RECT 85.595 3.985 85.765 4.155 ;
        RECT 86.075 3.985 86.245 4.155 ;
        RECT 86.555 3.985 86.725 4.155 ;
        RECT 87.035 3.985 87.205 4.155 ;
        RECT 87.515 3.985 87.685 4.155 ;
        RECT 87.995 3.985 88.165 4.155 ;
        RECT 88.475 3.985 88.645 4.155 ;
        RECT 88.955 3.985 89.125 4.155 ;
        RECT 89.435 3.985 89.605 4.155 ;
        RECT 89.915 3.985 90.085 4.155 ;
        RECT 90.395 3.985 90.565 4.155 ;
        RECT 90.875 3.985 91.045 4.155 ;
        RECT 91.355 3.985 91.525 4.155 ;
        RECT 91.835 3.985 92.005 4.155 ;
        RECT 92.315 3.985 92.485 4.155 ;
        RECT 92.795 3.985 92.965 4.155 ;
        RECT 93.275 3.985 93.445 4.155 ;
        RECT 93.755 3.985 93.925 4.155 ;
        RECT 94.235 3.985 94.405 4.155 ;
        RECT 94.715 3.985 94.885 4.155 ;
        RECT 95.195 3.985 95.365 4.155 ;
        RECT 95.675 3.985 95.845 4.155 ;
        RECT 96.155 3.985 96.325 4.155 ;
        RECT 96.635 3.985 96.805 4.155 ;
        RECT 97.115 3.985 97.285 4.155 ;
        RECT 97.595 3.985 97.765 4.155 ;
        RECT 98.075 3.985 98.245 4.155 ;
        RECT 98.555 3.985 98.725 4.155 ;
        RECT 99.035 3.985 99.205 4.155 ;
        RECT 99.515 3.985 99.685 4.155 ;
        RECT 99.995 3.985 100.165 4.155 ;
        RECT 100.475 3.985 100.645 4.155 ;
        RECT 100.955 3.985 101.125 4.155 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
        RECT 13.595 -0.085 13.765 0.085 ;
        RECT 14.075 -0.085 14.245 0.085 ;
        RECT 14.555 -0.085 14.725 0.085 ;
        RECT 15.035 -0.085 15.205 0.085 ;
        RECT 15.515 -0.085 15.685 0.085 ;
        RECT 15.995 -0.085 16.165 0.085 ;
        RECT 16.475 -0.085 16.645 0.085 ;
        RECT 16.955 -0.085 17.125 0.085 ;
        RECT 17.435 -0.085 17.605 0.085 ;
        RECT 17.915 -0.085 18.085 0.085 ;
        RECT 18.395 -0.085 18.565 0.085 ;
        RECT 18.875 -0.085 19.045 0.085 ;
        RECT 19.355 -0.085 19.525 0.085 ;
        RECT 19.835 -0.085 20.005 0.085 ;
        RECT 20.315 -0.085 20.485 0.085 ;
        RECT 20.795 -0.085 20.965 0.085 ;
        RECT 21.275 -0.085 21.445 0.085 ;
        RECT 21.755 -0.085 21.925 0.085 ;
        RECT 22.235 -0.085 22.405 0.085 ;
        RECT 22.715 -0.085 22.885 0.085 ;
        RECT 23.195 -0.085 23.365 0.085 ;
        RECT 23.675 -0.085 23.845 0.085 ;
        RECT 24.155 -0.085 24.325 0.085 ;
        RECT 24.635 -0.085 24.805 0.085 ;
        RECT 25.115 -0.085 25.285 0.085 ;
        RECT 25.595 -0.085 25.765 0.085 ;
        RECT 26.075 -0.085 26.245 0.085 ;
        RECT 26.555 -0.085 26.725 0.085 ;
        RECT 27.035 -0.085 27.205 0.085 ;
        RECT 27.515 -0.085 27.685 0.085 ;
        RECT 27.995 -0.085 28.165 0.085 ;
        RECT 28.475 -0.085 28.645 0.085 ;
        RECT 28.955 -0.085 29.125 0.085 ;
        RECT 29.435 -0.085 29.605 0.085 ;
        RECT 29.915 -0.085 30.085 0.085 ;
        RECT 30.395 -0.085 30.565 0.085 ;
        RECT 30.875 -0.085 31.045 0.085 ;
        RECT 31.355 -0.085 31.525 0.085 ;
        RECT 31.835 -0.085 32.005 0.085 ;
        RECT 32.315 -0.085 32.485 0.085 ;
        RECT 32.795 -0.085 32.965 0.085 ;
        RECT 33.275 -0.085 33.445 0.085 ;
        RECT 33.755 -0.085 33.925 0.085 ;
        RECT 34.235 -0.085 34.405 0.085 ;
        RECT 34.715 -0.085 34.885 0.085 ;
        RECT 35.195 -0.085 35.365 0.085 ;
        RECT 35.675 -0.085 35.845 0.085 ;
        RECT 36.155 -0.085 36.325 0.085 ;
        RECT 36.635 -0.085 36.805 0.085 ;
        RECT 37.115 -0.085 37.285 0.085 ;
        RECT 37.595 -0.085 37.765 0.085 ;
        RECT 38.075 -0.085 38.245 0.085 ;
        RECT 38.555 -0.085 38.725 0.085 ;
        RECT 39.035 -0.085 39.205 0.085 ;
        RECT 39.515 -0.085 39.685 0.085 ;
        RECT 39.995 -0.085 40.165 0.085 ;
        RECT 40.475 -0.085 40.645 0.085 ;
        RECT 40.955 -0.085 41.125 0.085 ;
        RECT 41.435 -0.085 41.605 0.085 ;
        RECT 41.915 -0.085 42.085 0.085 ;
        RECT 42.395 -0.085 42.565 0.085 ;
        RECT 42.875 -0.085 43.045 0.085 ;
        RECT 43.355 -0.085 43.525 0.085 ;
        RECT 43.835 -0.085 44.005 0.085 ;
        RECT 44.315 -0.085 44.485 0.085 ;
        RECT 44.795 -0.085 44.965 0.085 ;
        RECT 45.275 -0.085 45.445 0.085 ;
        RECT 45.755 -0.085 45.925 0.085 ;
        RECT 46.235 -0.085 46.405 0.085 ;
        RECT 46.715 -0.085 46.885 0.085 ;
        RECT 47.195 -0.085 47.365 0.085 ;
        RECT 47.675 -0.085 47.845 0.085 ;
        RECT 48.155 -0.085 48.325 0.085 ;
        RECT 48.635 -0.085 48.805 0.085 ;
        RECT 49.115 -0.085 49.285 0.085 ;
        RECT 49.595 -0.085 49.765 0.085 ;
        RECT 50.075 -0.085 50.245 0.085 ;
        RECT 50.555 -0.085 50.725 0.085 ;
        RECT 51.035 -0.085 51.205 0.085 ;
        RECT 51.515 -0.085 51.685 0.085 ;
        RECT 51.995 -0.085 52.165 0.085 ;
        RECT 52.475 -0.085 52.645 0.085 ;
        RECT 52.955 -0.085 53.125 0.085 ;
        RECT 53.435 -0.085 53.605 0.085 ;
        RECT 53.915 -0.085 54.085 0.085 ;
        RECT 54.395 -0.085 54.565 0.085 ;
        RECT 54.875 -0.085 55.045 0.085 ;
        RECT 55.355 -0.085 55.525 0.085 ;
        RECT 55.835 -0.085 56.005 0.085 ;
        RECT 56.315 -0.085 56.485 0.085 ;
        RECT 56.795 -0.085 56.965 0.085 ;
        RECT 57.275 -0.085 57.445 0.085 ;
        RECT 57.755 -0.085 57.925 0.085 ;
        RECT 58.235 -0.085 58.405 0.085 ;
        RECT 58.715 -0.085 58.885 0.085 ;
        RECT 59.195 -0.085 59.365 0.085 ;
        RECT 59.675 -0.085 59.845 0.085 ;
        RECT 60.155 -0.085 60.325 0.085 ;
        RECT 60.635 -0.085 60.805 0.085 ;
        RECT 61.115 -0.085 61.285 0.085 ;
        RECT 61.595 -0.085 61.765 0.085 ;
        RECT 62.075 -0.085 62.245 0.085 ;
        RECT 62.555 -0.085 62.725 0.085 ;
        RECT 63.035 -0.085 63.205 0.085 ;
        RECT 63.515 -0.085 63.685 0.085 ;
        RECT 63.995 -0.085 64.165 0.085 ;
        RECT 64.475 -0.085 64.645 0.085 ;
        RECT 64.955 -0.085 65.125 0.085 ;
        RECT 65.435 -0.085 65.605 0.085 ;
        RECT 65.915 -0.085 66.085 0.085 ;
        RECT 66.395 -0.085 66.565 0.085 ;
        RECT 66.875 -0.085 67.045 0.085 ;
        RECT 67.355 -0.085 67.525 0.085 ;
        RECT 67.835 -0.085 68.005 0.085 ;
        RECT 68.315 -0.085 68.485 0.085 ;
        RECT 68.795 -0.085 68.965 0.085 ;
        RECT 69.275 -0.085 69.445 0.085 ;
        RECT 69.755 -0.085 69.925 0.085 ;
        RECT 70.235 -0.085 70.405 0.085 ;
        RECT 70.715 -0.085 70.885 0.085 ;
        RECT 71.195 -0.085 71.365 0.085 ;
        RECT 71.675 -0.085 71.845 0.085 ;
        RECT 72.155 -0.085 72.325 0.085 ;
        RECT 72.635 -0.085 72.805 0.085 ;
        RECT 73.115 -0.085 73.285 0.085 ;
        RECT 73.595 -0.085 73.765 0.085 ;
        RECT 74.075 -0.085 74.245 0.085 ;
        RECT 74.555 -0.085 74.725 0.085 ;
        RECT 75.035 -0.085 75.205 0.085 ;
        RECT 75.515 -0.085 75.685 0.085 ;
        RECT 75.995 -0.085 76.165 0.085 ;
        RECT 76.475 -0.085 76.645 0.085 ;
        RECT 76.955 -0.085 77.125 0.085 ;
        RECT 77.435 -0.085 77.605 0.085 ;
        RECT 77.915 -0.085 78.085 0.085 ;
        RECT 78.395 -0.085 78.565 0.085 ;
        RECT 78.875 -0.085 79.045 0.085 ;
        RECT 79.355 -0.085 79.525 0.085 ;
        RECT 79.835 -0.085 80.005 0.085 ;
        RECT 80.315 -0.085 80.485 0.085 ;
        RECT 80.795 -0.085 80.965 0.085 ;
        RECT 81.275 -0.085 81.445 0.085 ;
        RECT 81.755 -0.085 81.925 0.085 ;
        RECT 82.235 -0.085 82.405 0.085 ;
        RECT 82.715 -0.085 82.885 0.085 ;
        RECT 83.195 -0.085 83.365 0.085 ;
        RECT 83.675 -0.085 83.845 0.085 ;
        RECT 84.155 -0.085 84.325 0.085 ;
        RECT 84.635 -0.085 84.805 0.085 ;
        RECT 85.115 -0.085 85.285 0.085 ;
        RECT 85.595 -0.085 85.765 0.085 ;
        RECT 86.075 -0.085 86.245 0.085 ;
        RECT 86.555 -0.085 86.725 0.085 ;
        RECT 87.035 -0.085 87.205 0.085 ;
        RECT 87.515 -0.085 87.685 0.085 ;
        RECT 87.995 -0.085 88.165 0.085 ;
        RECT 88.475 -0.085 88.645 0.085 ;
        RECT 88.955 -0.085 89.125 0.085 ;
        RECT 89.435 -0.085 89.605 0.085 ;
        RECT 89.915 -0.085 90.085 0.085 ;
        RECT 90.395 -0.085 90.565 0.085 ;
        RECT 90.875 -0.085 91.045 0.085 ;
        RECT 91.355 -0.085 91.525 0.085 ;
        RECT 91.835 -0.085 92.005 0.085 ;
        RECT 92.315 -0.085 92.485 0.085 ;
        RECT 92.795 -0.085 92.965 0.085 ;
        RECT 93.275 -0.085 93.445 0.085 ;
        RECT 93.755 -0.085 93.925 0.085 ;
        RECT 94.235 -0.085 94.405 0.085 ;
        RECT 94.715 -0.085 94.885 0.085 ;
        RECT 95.195 -0.085 95.365 0.085 ;
        RECT 95.675 -0.085 95.845 0.085 ;
        RECT 96.155 -0.085 96.325 0.085 ;
        RECT 96.635 -0.085 96.805 0.085 ;
        RECT 97.115 -0.085 97.285 0.085 ;
        RECT 97.595 -0.085 97.765 0.085 ;
        RECT 98.075 -0.085 98.245 0.085 ;
        RECT 98.555 -0.085 98.725 0.085 ;
        RECT 99.035 -0.085 99.205 0.085 ;
        RECT 99.515 -0.085 99.685 0.085 ;
        RECT 99.995 -0.085 100.165 0.085 ;
        RECT 100.475 -0.085 100.645 0.085 ;
        RECT 100.955 -0.085 101.125 0.085 ;
      LAYER met1 ;
        RECT 0.000 60.935 101.280 61.165 ;
        RECT 0.000 60.425 101.280 60.795 ;
        RECT 0.000 57.235 101.280 57.605 ;
        RECT 0.000 56.865 101.280 57.095 ;
        RECT 0.000 56.355 3.840 56.725 ;
        RECT 97.440 56.355 101.280 56.725 ;
        RECT 0.000 52.795 3.840 53.025 ;
        RECT 97.440 52.795 101.280 53.025 ;
        RECT 0.000 49.095 3.840 49.465 ;
        RECT 97.440 49.095 101.280 49.465 ;
        RECT 0.000 48.725 3.840 48.955 ;
        RECT 8.080 48.800 9.360 48.820 ;
        RECT 0.000 48.215 3.840 48.585 ;
        RECT 8.035 48.570 9.405 48.800 ;
        RECT 12.565 48.765 13.845 48.785 ;
        RECT 18.025 48.765 19.305 48.785 ;
        RECT 25.050 48.765 26.330 48.785 ;
        RECT 32.785 48.765 34.065 48.785 ;
        RECT 40.340 48.765 41.620 48.785 ;
        RECT 48.150 48.765 49.430 48.785 ;
        RECT 55.660 48.765 56.940 48.785 ;
        RECT 63.335 48.765 64.615 48.785 ;
        RECT 70.845 48.765 72.125 48.785 ;
        RECT 8.080 48.560 9.360 48.570 ;
        RECT 12.520 48.535 13.890 48.765 ;
        RECT 17.980 48.535 19.350 48.765 ;
        RECT 25.005 48.535 26.375 48.765 ;
        RECT 32.740 48.535 34.110 48.765 ;
        RECT 40.295 48.535 41.665 48.765 ;
        RECT 48.105 48.535 49.475 48.765 ;
        RECT 55.615 48.535 56.985 48.765 ;
        RECT 63.290 48.535 64.660 48.765 ;
        RECT 70.800 48.535 72.170 48.765 ;
        RECT 97.440 48.725 101.280 48.955 ;
        RECT 12.565 48.525 13.845 48.535 ;
        RECT 18.025 48.525 19.305 48.535 ;
        RECT 25.050 48.525 26.330 48.535 ;
        RECT 32.785 48.525 34.065 48.535 ;
        RECT 40.340 48.525 41.620 48.535 ;
        RECT 48.150 48.525 49.430 48.535 ;
        RECT 55.660 48.525 56.940 48.535 ;
        RECT 63.335 48.525 64.615 48.535 ;
        RECT 70.845 48.525 72.125 48.535 ;
        RECT 97.440 48.215 101.280 48.585 ;
        RECT 8.080 46.085 9.360 46.105 ;
        RECT 8.035 45.855 9.405 46.085 ;
        RECT 8.080 45.845 9.360 45.855 ;
        RECT 0.000 45.025 3.840 45.395 ;
        RECT 0.000 44.655 3.840 44.885 ;
        RECT 0.000 44.145 3.840 44.515 ;
        RECT 8.080 43.725 9.360 43.745 ;
        RECT 8.035 43.495 9.405 43.725 ;
        RECT 8.080 43.485 9.360 43.495 ;
        RECT 8.080 41.370 9.360 41.390 ;
        RECT 0.000 40.955 3.840 41.325 ;
        RECT 8.035 41.140 9.405 41.370 ;
        RECT 8.080 41.130 9.360 41.140 ;
        RECT 0.000 40.585 3.840 40.815 ;
        RECT 11.545 40.810 11.835 46.605 ;
        RECT 12.565 46.085 13.845 46.105 ;
        RECT 12.520 45.855 13.890 46.085 ;
        RECT 12.565 45.845 13.845 45.855 ;
        RECT 12.565 43.725 13.845 43.745 ;
        RECT 12.520 43.495 13.890 43.725 ;
        RECT 12.565 43.485 13.845 43.495 ;
        RECT 12.565 41.370 13.845 41.390 ;
        RECT 12.520 41.140 13.890 41.370 ;
        RECT 12.565 41.130 13.845 41.140 ;
        RECT 16.030 40.810 16.320 46.605 ;
        RECT 18.025 46.085 19.305 46.105 ;
        RECT 17.980 45.855 19.350 46.085 ;
        RECT 18.025 45.845 19.305 45.855 ;
        RECT 18.025 43.725 19.305 43.745 ;
        RECT 17.980 43.495 19.350 43.725 ;
        RECT 18.025 43.485 19.305 43.495 ;
        RECT 18.025 41.370 19.305 41.390 ;
        RECT 17.980 41.140 19.350 41.370 ;
        RECT 18.025 41.130 19.305 41.140 ;
        RECT 21.490 40.810 21.780 46.605 ;
        RECT 25.050 46.085 26.330 46.105 ;
        RECT 25.005 45.855 26.375 46.085 ;
        RECT 25.050 45.845 26.330 45.855 ;
        RECT 25.050 43.725 26.330 43.745 ;
        RECT 25.005 43.495 26.375 43.725 ;
        RECT 25.050 43.485 26.330 43.495 ;
        RECT 25.050 41.370 26.330 41.390 ;
        RECT 25.005 41.140 26.375 41.370 ;
        RECT 25.050 41.130 26.330 41.140 ;
        RECT 28.515 40.810 28.805 46.605 ;
        RECT 32.785 46.085 34.065 46.105 ;
        RECT 32.740 45.855 34.110 46.085 ;
        RECT 32.785 45.845 34.065 45.855 ;
        RECT 32.785 43.725 34.065 43.745 ;
        RECT 32.740 43.495 34.110 43.725 ;
        RECT 32.785 43.485 34.065 43.495 ;
        RECT 32.785 41.370 34.065 41.390 ;
        RECT 32.740 41.140 34.110 41.370 ;
        RECT 32.785 41.130 34.065 41.140 ;
        RECT 36.250 40.810 36.540 46.605 ;
        RECT 40.340 46.085 41.620 46.105 ;
        RECT 40.295 45.855 41.665 46.085 ;
        RECT 40.340 45.845 41.620 45.855 ;
        RECT 40.340 43.725 41.620 43.745 ;
        RECT 40.295 43.495 41.665 43.725 ;
        RECT 40.340 43.485 41.620 43.495 ;
        RECT 40.340 41.370 41.620 41.390 ;
        RECT 40.295 41.140 41.665 41.370 ;
        RECT 40.340 41.130 41.620 41.140 ;
        RECT 43.805 40.810 44.095 46.605 ;
        RECT 48.150 46.085 49.430 46.105 ;
        RECT 48.105 45.855 49.475 46.085 ;
        RECT 48.150 45.845 49.430 45.855 ;
        RECT 48.150 43.725 49.430 43.745 ;
        RECT 48.105 43.495 49.475 43.725 ;
        RECT 48.150 43.485 49.430 43.495 ;
        RECT 48.150 41.370 49.430 41.390 ;
        RECT 48.105 41.140 49.475 41.370 ;
        RECT 48.150 41.130 49.430 41.140 ;
        RECT 51.615 40.810 51.905 46.605 ;
        RECT 55.660 46.085 56.940 46.105 ;
        RECT 55.615 45.855 56.985 46.085 ;
        RECT 55.660 45.845 56.940 45.855 ;
        RECT 55.660 43.725 56.940 43.745 ;
        RECT 55.615 43.495 56.985 43.725 ;
        RECT 55.660 43.485 56.940 43.495 ;
        RECT 55.660 41.370 56.940 41.390 ;
        RECT 55.615 41.140 56.985 41.370 ;
        RECT 55.660 41.130 56.940 41.140 ;
        RECT 59.125 40.810 59.415 46.605 ;
        RECT 63.335 46.085 64.615 46.105 ;
        RECT 63.290 45.855 64.660 46.085 ;
        RECT 63.335 45.845 64.615 45.855 ;
        RECT 63.335 43.725 64.615 43.745 ;
        RECT 63.290 43.495 64.660 43.725 ;
        RECT 63.335 43.485 64.615 43.495 ;
        RECT 63.335 41.370 64.615 41.390 ;
        RECT 63.290 41.140 64.660 41.370 ;
        RECT 63.335 41.130 64.615 41.140 ;
        RECT 66.800 40.810 67.090 46.605 ;
        RECT 70.845 46.085 72.125 46.105 ;
        RECT 70.800 45.855 72.170 46.085 ;
        RECT 70.845 45.845 72.125 45.855 ;
        RECT 70.845 43.725 72.125 43.745 ;
        RECT 70.800 43.495 72.170 43.725 ;
        RECT 70.845 43.485 72.125 43.495 ;
        RECT 70.845 41.370 72.125 41.390 ;
        RECT 70.800 41.140 72.170 41.370 ;
        RECT 70.845 41.130 72.125 41.140 ;
        RECT 74.310 40.810 74.600 46.605 ;
        RECT 81.050 45.155 84.610 45.535 ;
        RECT 78.345 43.620 78.635 43.910 ;
        RECT 0.000 40.075 3.840 40.445 ;
        RECT 11.545 40.430 74.605 40.810 ;
        RECT 78.420 40.430 78.560 43.620 ;
        RECT 8.080 39.010 9.360 39.030 ;
        RECT 8.035 38.780 9.405 39.010 ;
        RECT 8.080 38.770 9.360 38.780 ;
        RECT 0.000 36.885 3.840 37.255 ;
        RECT 0.000 36.515 3.840 36.745 ;
        RECT 8.080 36.650 9.360 36.670 ;
        RECT 8.035 36.420 9.405 36.650 ;
        RECT 8.080 36.410 9.360 36.420 ;
        RECT 0.000 36.005 3.840 36.375 ;
        RECT 8.080 34.290 9.360 34.310 ;
        RECT 8.035 34.060 9.405 34.290 ;
        RECT 8.080 34.050 9.360 34.060 ;
        RECT 0.000 32.815 3.840 33.185 ;
        RECT 0.000 32.445 3.840 32.675 ;
        RECT 0.000 31.935 3.840 32.305 ;
        RECT 8.080 31.930 9.360 31.950 ;
        RECT 8.035 31.700 9.405 31.930 ;
        RECT 8.080 31.690 9.360 31.700 ;
        RECT 8.080 29.570 9.360 29.590 ;
        RECT 8.035 29.340 9.405 29.570 ;
        RECT 8.080 29.330 9.360 29.340 ;
        RECT 0.000 28.745 3.840 29.115 ;
        RECT 11.545 29.105 11.835 40.430 ;
        RECT 12.565 39.010 13.845 39.030 ;
        RECT 12.520 38.780 13.890 39.010 ;
        RECT 12.565 38.770 13.845 38.780 ;
        RECT 12.565 36.650 13.845 36.670 ;
        RECT 12.520 36.420 13.890 36.650 ;
        RECT 12.565 36.410 13.845 36.420 ;
        RECT 12.565 34.290 13.845 34.310 ;
        RECT 12.520 34.060 13.890 34.290 ;
        RECT 12.565 34.050 13.845 34.060 ;
        RECT 12.565 31.930 13.845 31.950 ;
        RECT 12.520 31.700 13.890 31.930 ;
        RECT 12.565 31.690 13.845 31.700 ;
        RECT 12.565 29.570 13.845 29.590 ;
        RECT 12.520 29.340 13.890 29.570 ;
        RECT 12.565 29.330 13.845 29.340 ;
        RECT 16.030 29.105 16.320 40.430 ;
        RECT 18.025 39.010 19.305 39.030 ;
        RECT 17.980 38.780 19.350 39.010 ;
        RECT 18.025 38.770 19.305 38.780 ;
        RECT 18.025 36.650 19.305 36.670 ;
        RECT 17.980 36.420 19.350 36.650 ;
        RECT 18.025 36.410 19.305 36.420 ;
        RECT 18.025 34.290 19.305 34.310 ;
        RECT 17.980 34.060 19.350 34.290 ;
        RECT 18.025 34.050 19.305 34.060 ;
        RECT 18.025 31.930 19.305 31.950 ;
        RECT 17.980 31.700 19.350 31.930 ;
        RECT 18.025 31.690 19.305 31.700 ;
        RECT 18.025 29.570 19.305 29.590 ;
        RECT 17.980 29.340 19.350 29.570 ;
        RECT 18.025 29.330 19.305 29.340 ;
        RECT 21.490 29.105 21.780 40.430 ;
        RECT 25.050 39.010 26.330 39.030 ;
        RECT 25.005 38.780 26.375 39.010 ;
        RECT 25.050 38.770 26.330 38.780 ;
        RECT 25.050 36.650 26.330 36.670 ;
        RECT 25.005 36.420 26.375 36.650 ;
        RECT 25.050 36.410 26.330 36.420 ;
        RECT 25.050 34.290 26.330 34.310 ;
        RECT 25.005 34.060 26.375 34.290 ;
        RECT 25.050 34.050 26.330 34.060 ;
        RECT 25.050 31.930 26.330 31.950 ;
        RECT 25.005 31.700 26.375 31.930 ;
        RECT 25.050 31.690 26.330 31.700 ;
        RECT 25.050 29.570 26.330 29.590 ;
        RECT 25.005 29.340 26.375 29.570 ;
        RECT 25.050 29.330 26.330 29.340 ;
        RECT 28.515 29.105 28.805 40.430 ;
        RECT 32.785 39.010 34.065 39.030 ;
        RECT 32.740 38.780 34.110 39.010 ;
        RECT 32.785 38.770 34.065 38.780 ;
        RECT 32.785 36.650 34.065 36.670 ;
        RECT 32.740 36.420 34.110 36.650 ;
        RECT 32.785 36.410 34.065 36.420 ;
        RECT 32.785 34.290 34.065 34.310 ;
        RECT 32.740 34.060 34.110 34.290 ;
        RECT 32.785 34.050 34.065 34.060 ;
        RECT 32.785 31.930 34.065 31.950 ;
        RECT 32.740 31.700 34.110 31.930 ;
        RECT 32.785 31.690 34.065 31.700 ;
        RECT 32.785 29.570 34.065 29.590 ;
        RECT 32.740 29.340 34.110 29.570 ;
        RECT 32.785 29.330 34.065 29.340 ;
        RECT 36.250 29.105 36.540 40.430 ;
        RECT 40.340 39.010 41.620 39.030 ;
        RECT 40.295 38.780 41.665 39.010 ;
        RECT 40.340 38.770 41.620 38.780 ;
        RECT 40.340 36.650 41.620 36.670 ;
        RECT 40.295 36.420 41.665 36.650 ;
        RECT 40.340 36.410 41.620 36.420 ;
        RECT 40.340 34.290 41.620 34.310 ;
        RECT 40.295 34.060 41.665 34.290 ;
        RECT 40.340 34.050 41.620 34.060 ;
        RECT 40.340 31.930 41.620 31.950 ;
        RECT 40.295 31.700 41.665 31.930 ;
        RECT 40.340 31.690 41.620 31.700 ;
        RECT 40.340 29.570 41.620 29.590 ;
        RECT 40.295 29.340 41.665 29.570 ;
        RECT 40.340 29.330 41.620 29.340 ;
        RECT 43.805 29.105 44.095 40.430 ;
        RECT 48.150 39.010 49.430 39.030 ;
        RECT 48.105 38.780 49.475 39.010 ;
        RECT 48.150 38.770 49.430 38.780 ;
        RECT 48.150 36.650 49.430 36.670 ;
        RECT 48.105 36.420 49.475 36.650 ;
        RECT 48.150 36.410 49.430 36.420 ;
        RECT 48.150 34.290 49.430 34.310 ;
        RECT 48.105 34.060 49.475 34.290 ;
        RECT 48.150 34.050 49.430 34.060 ;
        RECT 48.150 31.930 49.430 31.950 ;
        RECT 48.105 31.700 49.475 31.930 ;
        RECT 48.150 31.690 49.430 31.700 ;
        RECT 48.150 29.570 49.430 29.590 ;
        RECT 48.105 29.340 49.475 29.570 ;
        RECT 48.150 29.330 49.430 29.340 ;
        RECT 51.615 29.105 51.905 40.430 ;
        RECT 55.660 39.010 56.940 39.030 ;
        RECT 55.615 38.780 56.985 39.010 ;
        RECT 55.660 38.770 56.940 38.780 ;
        RECT 55.660 36.650 56.940 36.670 ;
        RECT 55.615 36.420 56.985 36.650 ;
        RECT 55.660 36.410 56.940 36.420 ;
        RECT 55.660 34.290 56.940 34.310 ;
        RECT 55.615 34.060 56.985 34.290 ;
        RECT 55.660 34.050 56.940 34.060 ;
        RECT 55.660 31.930 56.940 31.950 ;
        RECT 55.615 31.700 56.985 31.930 ;
        RECT 55.660 31.690 56.940 31.700 ;
        RECT 55.660 29.570 56.940 29.590 ;
        RECT 55.615 29.340 56.985 29.570 ;
        RECT 55.660 29.330 56.940 29.340 ;
        RECT 59.125 29.105 59.415 40.430 ;
        RECT 63.335 39.010 64.615 39.030 ;
        RECT 63.290 38.780 64.660 39.010 ;
        RECT 63.335 38.770 64.615 38.780 ;
        RECT 63.335 36.650 64.615 36.670 ;
        RECT 63.290 36.420 64.660 36.650 ;
        RECT 63.335 36.410 64.615 36.420 ;
        RECT 63.335 34.290 64.615 34.310 ;
        RECT 63.290 34.060 64.660 34.290 ;
        RECT 63.335 34.050 64.615 34.060 ;
        RECT 63.335 31.930 64.615 31.950 ;
        RECT 63.290 31.700 64.660 31.930 ;
        RECT 63.335 31.690 64.615 31.700 ;
        RECT 63.335 29.570 64.615 29.590 ;
        RECT 63.290 29.340 64.660 29.570 ;
        RECT 63.335 29.330 64.615 29.340 ;
        RECT 66.800 29.105 67.090 40.430 ;
        RECT 74.310 40.050 80.540 40.430 ;
        RECT 70.845 39.010 72.125 39.030 ;
        RECT 70.800 38.780 72.170 39.010 ;
        RECT 70.845 38.770 72.125 38.780 ;
        RECT 70.845 36.650 72.125 36.670 ;
        RECT 70.800 36.420 72.170 36.650 ;
        RECT 70.845 36.410 72.125 36.420 ;
        RECT 70.845 34.290 72.125 34.310 ;
        RECT 70.800 34.060 72.170 34.290 ;
        RECT 70.845 34.050 72.125 34.060 ;
        RECT 70.845 31.930 72.125 31.950 ;
        RECT 70.800 31.700 72.170 31.930 ;
        RECT 70.845 31.690 72.125 31.700 ;
        RECT 70.845 29.570 72.125 29.590 ;
        RECT 70.800 29.340 72.170 29.570 ;
        RECT 70.845 29.330 72.125 29.340 ;
        RECT 74.310 29.105 74.600 40.050 ;
        RECT 78.345 38.565 78.635 38.855 ;
        RECT 78.420 35.335 78.560 38.565 ;
        RECT 78.345 35.045 78.635 35.335 ;
        RECT 78.345 33.510 78.635 33.800 ;
        RECT 78.420 30.280 78.560 33.510 ;
        RECT 78.345 29.990 78.635 30.280 ;
        RECT 11.530 28.725 74.605 29.105 ;
        RECT 0.000 28.375 3.840 28.605 ;
        RECT 0.000 27.865 3.840 28.235 ;
        RECT 8.080 27.210 9.360 27.230 ;
        RECT 8.035 26.980 9.405 27.210 ;
        RECT 8.080 26.970 9.360 26.980 ;
        RECT 0.000 24.675 3.840 25.045 ;
        RECT 8.080 24.850 9.360 24.870 ;
        RECT 8.035 24.620 9.405 24.850 ;
        RECT 8.080 24.610 9.360 24.620 ;
        RECT 0.000 24.305 3.840 24.535 ;
        RECT 0.000 23.795 3.840 24.165 ;
        RECT 8.080 22.490 9.360 22.510 ;
        RECT 8.035 22.260 9.405 22.490 ;
        RECT 8.080 22.250 9.360 22.260 ;
        RECT 0.000 20.605 3.840 20.975 ;
        RECT 0.000 20.235 3.840 20.465 ;
        RECT 8.080 20.130 9.360 20.150 ;
        RECT 0.000 19.725 3.840 20.095 ;
        RECT 8.035 19.900 9.405 20.130 ;
        RECT 8.080 19.890 9.360 19.900 ;
        RECT 8.080 17.770 9.360 17.790 ;
        RECT 8.035 17.540 9.405 17.770 ;
        RECT 8.080 17.530 9.360 17.540 ;
        RECT 11.545 17.295 11.835 28.725 ;
        RECT 12.565 27.210 13.845 27.230 ;
        RECT 12.520 26.980 13.890 27.210 ;
        RECT 12.565 26.970 13.845 26.980 ;
        RECT 12.565 24.850 13.845 24.870 ;
        RECT 12.520 24.620 13.890 24.850 ;
        RECT 12.565 24.610 13.845 24.620 ;
        RECT 12.565 22.490 13.845 22.510 ;
        RECT 12.520 22.260 13.890 22.490 ;
        RECT 12.565 22.250 13.845 22.260 ;
        RECT 12.565 20.130 13.845 20.150 ;
        RECT 12.520 19.900 13.890 20.130 ;
        RECT 12.565 19.890 13.845 19.900 ;
        RECT 12.565 17.770 13.845 17.790 ;
        RECT 12.520 17.540 13.890 17.770 ;
        RECT 12.565 17.530 13.845 17.540 ;
        RECT 16.030 17.295 16.320 28.725 ;
        RECT 18.025 27.210 19.305 27.230 ;
        RECT 17.980 26.980 19.350 27.210 ;
        RECT 18.025 26.970 19.305 26.980 ;
        RECT 18.025 24.850 19.305 24.870 ;
        RECT 17.980 24.620 19.350 24.850 ;
        RECT 18.025 24.610 19.305 24.620 ;
        RECT 18.025 22.490 19.305 22.510 ;
        RECT 17.980 22.260 19.350 22.490 ;
        RECT 18.025 22.250 19.305 22.260 ;
        RECT 18.025 20.130 19.305 20.150 ;
        RECT 17.980 19.900 19.350 20.130 ;
        RECT 18.025 19.890 19.305 19.900 ;
        RECT 18.025 17.770 19.305 17.790 ;
        RECT 17.980 17.540 19.350 17.770 ;
        RECT 18.025 17.530 19.305 17.540 ;
        RECT 21.490 17.295 21.780 28.725 ;
        RECT 25.050 27.210 26.330 27.230 ;
        RECT 25.005 26.980 26.375 27.210 ;
        RECT 25.050 26.970 26.330 26.980 ;
        RECT 25.050 24.850 26.330 24.870 ;
        RECT 25.005 24.620 26.375 24.850 ;
        RECT 25.050 24.610 26.330 24.620 ;
        RECT 25.050 22.490 26.330 22.510 ;
        RECT 25.005 22.260 26.375 22.490 ;
        RECT 25.050 22.250 26.330 22.260 ;
        RECT 25.050 20.130 26.330 20.150 ;
        RECT 25.005 19.900 26.375 20.130 ;
        RECT 25.050 19.890 26.330 19.900 ;
        RECT 25.050 17.770 26.330 17.790 ;
        RECT 25.005 17.540 26.375 17.770 ;
        RECT 25.050 17.530 26.330 17.540 ;
        RECT 28.515 17.295 28.805 28.725 ;
        RECT 32.785 27.210 34.065 27.230 ;
        RECT 32.740 26.980 34.110 27.210 ;
        RECT 32.785 26.970 34.065 26.980 ;
        RECT 32.785 24.850 34.065 24.870 ;
        RECT 32.740 24.620 34.110 24.850 ;
        RECT 32.785 24.610 34.065 24.620 ;
        RECT 32.785 22.490 34.065 22.510 ;
        RECT 32.740 22.260 34.110 22.490 ;
        RECT 32.785 22.250 34.065 22.260 ;
        RECT 32.785 20.130 34.065 20.150 ;
        RECT 32.740 19.900 34.110 20.130 ;
        RECT 32.785 19.890 34.065 19.900 ;
        RECT 32.785 17.770 34.065 17.790 ;
        RECT 32.740 17.540 34.110 17.770 ;
        RECT 32.785 17.530 34.065 17.540 ;
        RECT 36.250 17.295 36.540 28.725 ;
        RECT 40.340 27.210 41.620 27.230 ;
        RECT 40.295 26.980 41.665 27.210 ;
        RECT 40.340 26.970 41.620 26.980 ;
        RECT 40.340 24.850 41.620 24.870 ;
        RECT 40.295 24.620 41.665 24.850 ;
        RECT 40.340 24.610 41.620 24.620 ;
        RECT 40.340 22.490 41.620 22.510 ;
        RECT 40.295 22.260 41.665 22.490 ;
        RECT 40.340 22.250 41.620 22.260 ;
        RECT 40.340 20.130 41.620 20.150 ;
        RECT 40.295 19.900 41.665 20.130 ;
        RECT 40.340 19.890 41.620 19.900 ;
        RECT 40.340 17.770 41.620 17.790 ;
        RECT 40.295 17.540 41.665 17.770 ;
        RECT 40.340 17.530 41.620 17.540 ;
        RECT 43.805 17.295 44.095 28.725 ;
        RECT 48.150 27.210 49.430 27.230 ;
        RECT 48.105 26.980 49.475 27.210 ;
        RECT 48.150 26.970 49.430 26.980 ;
        RECT 48.150 24.850 49.430 24.870 ;
        RECT 48.105 24.620 49.475 24.850 ;
        RECT 48.150 24.610 49.430 24.620 ;
        RECT 48.150 22.490 49.430 22.510 ;
        RECT 48.105 22.260 49.475 22.490 ;
        RECT 48.150 22.250 49.430 22.260 ;
        RECT 48.150 20.130 49.430 20.150 ;
        RECT 48.105 19.900 49.475 20.130 ;
        RECT 48.150 19.890 49.430 19.900 ;
        RECT 48.150 17.770 49.430 17.790 ;
        RECT 48.105 17.540 49.475 17.770 ;
        RECT 48.150 17.530 49.430 17.540 ;
        RECT 51.615 17.295 51.905 28.725 ;
        RECT 55.660 27.210 56.940 27.230 ;
        RECT 55.615 26.980 56.985 27.210 ;
        RECT 55.660 26.970 56.940 26.980 ;
        RECT 55.660 24.850 56.940 24.870 ;
        RECT 55.615 24.620 56.985 24.850 ;
        RECT 55.660 24.610 56.940 24.620 ;
        RECT 55.660 22.490 56.940 22.510 ;
        RECT 55.615 22.260 56.985 22.490 ;
        RECT 55.660 22.250 56.940 22.260 ;
        RECT 55.660 20.130 56.940 20.150 ;
        RECT 55.615 19.900 56.985 20.130 ;
        RECT 55.660 19.890 56.940 19.900 ;
        RECT 55.660 17.770 56.940 17.790 ;
        RECT 55.615 17.540 56.985 17.770 ;
        RECT 55.660 17.530 56.940 17.540 ;
        RECT 59.125 17.295 59.415 28.725 ;
        RECT 63.335 27.210 64.615 27.230 ;
        RECT 63.290 26.980 64.660 27.210 ;
        RECT 63.335 26.970 64.615 26.980 ;
        RECT 63.335 24.850 64.615 24.870 ;
        RECT 63.290 24.620 64.660 24.850 ;
        RECT 63.335 24.610 64.615 24.620 ;
        RECT 63.335 22.490 64.615 22.510 ;
        RECT 63.290 22.260 64.660 22.490 ;
        RECT 63.335 22.250 64.615 22.260 ;
        RECT 63.335 20.130 64.615 20.150 ;
        RECT 63.290 19.900 64.660 20.130 ;
        RECT 63.335 19.890 64.615 19.900 ;
        RECT 63.335 17.770 64.615 17.790 ;
        RECT 63.290 17.540 64.660 17.770 ;
        RECT 63.335 17.530 64.615 17.540 ;
        RECT 66.800 17.295 67.090 28.725 ;
        RECT 70.845 27.210 72.125 27.230 ;
        RECT 70.800 26.980 72.170 27.210 ;
        RECT 70.845 26.970 72.125 26.980 ;
        RECT 70.845 24.850 72.125 24.870 ;
        RECT 70.800 24.620 72.170 24.850 ;
        RECT 70.845 24.610 72.125 24.620 ;
        RECT 70.845 22.490 72.125 22.510 ;
        RECT 70.800 22.260 72.170 22.490 ;
        RECT 70.845 22.250 72.125 22.260 ;
        RECT 70.845 20.130 72.125 20.150 ;
        RECT 70.800 19.900 72.170 20.130 ;
        RECT 70.845 19.890 72.125 19.900 ;
        RECT 70.845 17.770 72.125 17.790 ;
        RECT 70.800 17.540 72.170 17.770 ;
        RECT 70.845 17.530 72.125 17.540 ;
        RECT 74.310 17.295 74.600 28.725 ;
        RECT 78.345 28.455 78.635 28.745 ;
        RECT 78.420 25.225 78.560 28.455 ;
        RECT 78.345 24.935 78.635 25.225 ;
        RECT 78.345 23.400 78.635 23.690 ;
        RECT 78.420 20.170 78.560 23.400 ;
        RECT 78.345 19.880 78.635 20.170 ;
        RECT 78.345 18.345 78.635 18.635 ;
        RECT 11.530 16.915 74.605 17.295 ;
        RECT 0.000 16.535 3.840 16.905 ;
        RECT 0.000 16.165 3.840 16.395 ;
        RECT 0.000 15.655 3.840 16.025 ;
        RECT 8.080 15.410 9.360 15.430 ;
        RECT 8.035 15.180 9.405 15.410 ;
        RECT 8.080 15.170 9.360 15.180 ;
        RECT 8.080 13.050 9.360 13.070 ;
        RECT 0.000 12.465 3.840 12.835 ;
        RECT 8.035 12.820 9.405 13.050 ;
        RECT 8.080 12.810 9.360 12.820 ;
        RECT 0.000 12.095 3.840 12.325 ;
        RECT 11.545 12.320 11.835 16.915 ;
        RECT 12.565 15.410 13.845 15.430 ;
        RECT 12.520 15.180 13.890 15.410 ;
        RECT 12.565 15.170 13.845 15.180 ;
        RECT 12.565 13.050 13.845 13.070 ;
        RECT 12.520 12.820 13.890 13.050 ;
        RECT 12.565 12.810 13.845 12.820 ;
        RECT 16.030 12.320 16.320 16.915 ;
        RECT 18.025 15.410 19.305 15.430 ;
        RECT 17.980 15.180 19.350 15.410 ;
        RECT 18.025 15.170 19.305 15.180 ;
        RECT 18.025 13.050 19.305 13.070 ;
        RECT 17.980 12.820 19.350 13.050 ;
        RECT 18.025 12.810 19.305 12.820 ;
        RECT 21.490 12.320 21.780 16.915 ;
        RECT 25.050 15.410 26.330 15.430 ;
        RECT 25.005 15.180 26.375 15.410 ;
        RECT 25.050 15.170 26.330 15.180 ;
        RECT 25.050 13.050 26.330 13.070 ;
        RECT 25.005 12.820 26.375 13.050 ;
        RECT 25.050 12.810 26.330 12.820 ;
        RECT 28.515 12.320 28.805 16.915 ;
        RECT 32.785 15.410 34.065 15.430 ;
        RECT 32.740 15.180 34.110 15.410 ;
        RECT 32.785 15.170 34.065 15.180 ;
        RECT 32.785 13.050 34.065 13.070 ;
        RECT 32.740 12.820 34.110 13.050 ;
        RECT 32.785 12.810 34.065 12.820 ;
        RECT 36.250 12.320 36.540 16.915 ;
        RECT 40.340 15.410 41.620 15.430 ;
        RECT 40.295 15.180 41.665 15.410 ;
        RECT 40.340 15.170 41.620 15.180 ;
        RECT 40.340 13.050 41.620 13.070 ;
        RECT 40.295 12.820 41.665 13.050 ;
        RECT 40.340 12.810 41.620 12.820 ;
        RECT 43.805 12.320 44.095 16.915 ;
        RECT 48.150 15.410 49.430 15.430 ;
        RECT 48.105 15.180 49.475 15.410 ;
        RECT 48.150 15.170 49.430 15.180 ;
        RECT 48.150 13.050 49.430 13.070 ;
        RECT 48.105 12.820 49.475 13.050 ;
        RECT 48.150 12.810 49.430 12.820 ;
        RECT 51.615 12.320 51.905 16.915 ;
        RECT 55.660 15.410 56.940 15.430 ;
        RECT 55.615 15.180 56.985 15.410 ;
        RECT 55.660 15.170 56.940 15.180 ;
        RECT 55.660 13.050 56.940 13.070 ;
        RECT 55.615 12.820 56.985 13.050 ;
        RECT 55.660 12.810 56.940 12.820 ;
        RECT 59.125 12.320 59.415 16.915 ;
        RECT 63.335 15.410 64.615 15.430 ;
        RECT 63.290 15.180 64.660 15.410 ;
        RECT 63.335 15.170 64.615 15.180 ;
        RECT 63.335 13.050 64.615 13.070 ;
        RECT 63.290 12.820 64.660 13.050 ;
        RECT 63.335 12.810 64.615 12.820 ;
        RECT 66.800 12.320 67.090 16.915 ;
        RECT 70.845 15.410 72.125 15.430 ;
        RECT 70.800 15.180 72.170 15.410 ;
        RECT 70.845 15.170 72.125 15.180 ;
        RECT 70.845 13.050 72.125 13.070 ;
        RECT 70.800 12.820 72.170 13.050 ;
        RECT 70.845 12.810 72.125 12.820 ;
        RECT 74.310 12.320 74.600 16.915 ;
        RECT 78.420 15.115 78.560 18.345 ;
        RECT 78.345 14.825 78.635 15.115 ;
        RECT 78.345 13.505 78.635 13.580 ;
        RECT 81.050 13.505 81.245 45.155 ;
        RECT 97.440 45.025 101.280 45.395 ;
        RECT 97.440 44.655 101.280 44.885 ;
        RECT 97.440 44.145 101.280 44.515 ;
        RECT 83.895 43.620 84.185 43.910 ;
        RECT 83.970 40.390 84.110 43.620 ;
        RECT 97.440 40.955 101.280 41.325 ;
        RECT 97.440 40.585 101.280 40.815 ;
        RECT 83.885 40.090 84.185 40.390 ;
        RECT 97.440 40.075 101.280 40.445 ;
        RECT 83.895 38.565 84.185 38.855 ;
        RECT 83.970 35.335 84.110 38.565 ;
        RECT 97.440 36.885 101.280 37.255 ;
        RECT 97.440 36.515 101.280 36.745 ;
        RECT 97.440 36.005 101.280 36.375 ;
        RECT 83.895 35.045 84.185 35.335 ;
        RECT 83.895 33.510 84.185 33.800 ;
        RECT 83.970 30.280 84.110 33.510 ;
        RECT 97.440 32.815 101.280 33.185 ;
        RECT 97.440 32.445 101.280 32.675 ;
        RECT 97.440 31.935 101.280 32.305 ;
        RECT 83.895 29.990 84.185 30.280 ;
        RECT 97.440 28.745 101.280 29.115 ;
        RECT 83.895 28.455 84.185 28.745 ;
        RECT 83.970 25.225 84.110 28.455 ;
        RECT 97.440 28.375 101.280 28.605 ;
        RECT 97.440 27.865 101.280 28.235 ;
        RECT 83.895 24.935 84.185 25.225 ;
        RECT 97.440 24.675 101.280 25.045 ;
        RECT 97.440 24.305 101.280 24.535 ;
        RECT 97.440 23.795 101.280 24.165 ;
        RECT 83.895 23.400 84.185 23.690 ;
        RECT 83.970 20.170 84.110 23.400 ;
        RECT 97.440 20.605 101.280 20.975 ;
        RECT 97.440 20.235 101.280 20.465 ;
        RECT 83.895 19.880 84.185 20.170 ;
        RECT 89.565 20.160 89.855 20.170 ;
        RECT 86.600 19.895 90.260 20.160 ;
        RECT 83.895 18.345 84.185 18.635 ;
        RECT 83.970 15.115 84.110 18.345 ;
        RECT 83.895 14.825 84.185 15.115 ;
        RECT 78.345 13.365 81.245 13.505 ;
        RECT 83.895 13.505 84.185 13.580 ;
        RECT 86.600 13.505 86.795 19.895 ;
        RECT 89.565 19.880 89.855 19.895 ;
        RECT 97.440 19.725 101.280 20.095 ;
        RECT 89.565 18.345 89.855 18.635 ;
        RECT 89.640 15.115 89.780 18.345 ;
        RECT 97.440 16.535 101.280 16.905 ;
        RECT 97.440 16.165 101.280 16.395 ;
        RECT 97.440 15.655 101.280 16.025 ;
        RECT 89.565 14.825 89.855 15.115 ;
        RECT 83.895 13.365 86.795 13.505 ;
        RECT 78.345 13.290 78.635 13.365 ;
        RECT 83.895 13.290 84.185 13.365 ;
        RECT 97.440 12.465 101.280 12.835 ;
        RECT 97.440 12.095 101.280 12.325 ;
        RECT 0.000 11.585 3.840 11.955 ;
        RECT 97.440 11.585 101.280 11.955 ;
        RECT 0.000 8.025 3.840 8.255 ;
        RECT 97.440 8.025 101.280 8.255 ;
        RECT 0.000 4.325 3.840 4.695 ;
        RECT 97.440 4.325 101.280 4.695 ;
        RECT 0.000 3.955 101.280 4.185 ;
        RECT 0.000 3.445 101.280 3.815 ;
        RECT 0.000 0.255 101.280 0.625 ;
        RECT 0.000 -0.115 101.280 0.115 ;
      LAYER via ;
        RECT 8.110 48.560 8.370 48.820 ;
        RECT 8.430 48.560 8.690 48.820 ;
        RECT 8.750 48.560 9.010 48.820 ;
        RECT 9.070 48.560 9.330 48.820 ;
        RECT 12.595 48.525 12.855 48.785 ;
        RECT 12.915 48.525 13.175 48.785 ;
        RECT 13.235 48.525 13.495 48.785 ;
        RECT 13.555 48.525 13.815 48.785 ;
        RECT 18.055 48.525 18.315 48.785 ;
        RECT 18.375 48.525 18.635 48.785 ;
        RECT 18.695 48.525 18.955 48.785 ;
        RECT 19.015 48.525 19.275 48.785 ;
        RECT 25.080 48.525 25.340 48.785 ;
        RECT 25.400 48.525 25.660 48.785 ;
        RECT 25.720 48.525 25.980 48.785 ;
        RECT 26.040 48.525 26.300 48.785 ;
        RECT 32.815 48.525 33.075 48.785 ;
        RECT 33.135 48.525 33.395 48.785 ;
        RECT 33.455 48.525 33.715 48.785 ;
        RECT 33.775 48.525 34.035 48.785 ;
        RECT 40.370 48.525 40.630 48.785 ;
        RECT 40.690 48.525 40.950 48.785 ;
        RECT 41.010 48.525 41.270 48.785 ;
        RECT 41.330 48.525 41.590 48.785 ;
        RECT 48.180 48.525 48.440 48.785 ;
        RECT 48.500 48.525 48.760 48.785 ;
        RECT 48.820 48.525 49.080 48.785 ;
        RECT 49.140 48.525 49.400 48.785 ;
        RECT 55.690 48.525 55.950 48.785 ;
        RECT 56.010 48.525 56.270 48.785 ;
        RECT 56.330 48.525 56.590 48.785 ;
        RECT 56.650 48.525 56.910 48.785 ;
        RECT 63.365 48.525 63.625 48.785 ;
        RECT 63.685 48.525 63.945 48.785 ;
        RECT 64.005 48.525 64.265 48.785 ;
        RECT 64.325 48.525 64.585 48.785 ;
        RECT 70.875 48.525 71.135 48.785 ;
        RECT 71.195 48.525 71.455 48.785 ;
        RECT 71.515 48.525 71.775 48.785 ;
        RECT 71.835 48.525 72.095 48.785 ;
        RECT 8.110 45.845 8.370 46.105 ;
        RECT 8.430 45.845 8.690 46.105 ;
        RECT 8.750 45.845 9.010 46.105 ;
        RECT 9.070 45.845 9.330 46.105 ;
        RECT 8.110 43.485 8.370 43.745 ;
        RECT 8.430 43.485 8.690 43.745 ;
        RECT 8.750 43.485 9.010 43.745 ;
        RECT 9.070 43.485 9.330 43.745 ;
        RECT 8.110 41.130 8.370 41.390 ;
        RECT 8.430 41.130 8.690 41.390 ;
        RECT 8.750 41.130 9.010 41.390 ;
        RECT 9.070 41.130 9.330 41.390 ;
        RECT 12.595 45.845 12.855 46.105 ;
        RECT 12.915 45.845 13.175 46.105 ;
        RECT 13.235 45.845 13.495 46.105 ;
        RECT 13.555 45.845 13.815 46.105 ;
        RECT 12.595 43.485 12.855 43.745 ;
        RECT 12.915 43.485 13.175 43.745 ;
        RECT 13.235 43.485 13.495 43.745 ;
        RECT 13.555 43.485 13.815 43.745 ;
        RECT 12.595 41.130 12.855 41.390 ;
        RECT 12.915 41.130 13.175 41.390 ;
        RECT 13.235 41.130 13.495 41.390 ;
        RECT 13.555 41.130 13.815 41.390 ;
        RECT 18.055 45.845 18.315 46.105 ;
        RECT 18.375 45.845 18.635 46.105 ;
        RECT 18.695 45.845 18.955 46.105 ;
        RECT 19.015 45.845 19.275 46.105 ;
        RECT 18.055 43.485 18.315 43.745 ;
        RECT 18.375 43.485 18.635 43.745 ;
        RECT 18.695 43.485 18.955 43.745 ;
        RECT 19.015 43.485 19.275 43.745 ;
        RECT 18.055 41.130 18.315 41.390 ;
        RECT 18.375 41.130 18.635 41.390 ;
        RECT 18.695 41.130 18.955 41.390 ;
        RECT 19.015 41.130 19.275 41.390 ;
        RECT 25.080 45.845 25.340 46.105 ;
        RECT 25.400 45.845 25.660 46.105 ;
        RECT 25.720 45.845 25.980 46.105 ;
        RECT 26.040 45.845 26.300 46.105 ;
        RECT 25.080 43.485 25.340 43.745 ;
        RECT 25.400 43.485 25.660 43.745 ;
        RECT 25.720 43.485 25.980 43.745 ;
        RECT 26.040 43.485 26.300 43.745 ;
        RECT 25.080 41.130 25.340 41.390 ;
        RECT 25.400 41.130 25.660 41.390 ;
        RECT 25.720 41.130 25.980 41.390 ;
        RECT 26.040 41.130 26.300 41.390 ;
        RECT 32.815 45.845 33.075 46.105 ;
        RECT 33.135 45.845 33.395 46.105 ;
        RECT 33.455 45.845 33.715 46.105 ;
        RECT 33.775 45.845 34.035 46.105 ;
        RECT 32.815 43.485 33.075 43.745 ;
        RECT 33.135 43.485 33.395 43.745 ;
        RECT 33.455 43.485 33.715 43.745 ;
        RECT 33.775 43.485 34.035 43.745 ;
        RECT 32.815 41.130 33.075 41.390 ;
        RECT 33.135 41.130 33.395 41.390 ;
        RECT 33.455 41.130 33.715 41.390 ;
        RECT 33.775 41.130 34.035 41.390 ;
        RECT 40.370 45.845 40.630 46.105 ;
        RECT 40.690 45.845 40.950 46.105 ;
        RECT 41.010 45.845 41.270 46.105 ;
        RECT 41.330 45.845 41.590 46.105 ;
        RECT 40.370 43.485 40.630 43.745 ;
        RECT 40.690 43.485 40.950 43.745 ;
        RECT 41.010 43.485 41.270 43.745 ;
        RECT 41.330 43.485 41.590 43.745 ;
        RECT 40.370 41.130 40.630 41.390 ;
        RECT 40.690 41.130 40.950 41.390 ;
        RECT 41.010 41.130 41.270 41.390 ;
        RECT 41.330 41.130 41.590 41.390 ;
        RECT 48.180 45.845 48.440 46.105 ;
        RECT 48.500 45.845 48.760 46.105 ;
        RECT 48.820 45.845 49.080 46.105 ;
        RECT 49.140 45.845 49.400 46.105 ;
        RECT 48.180 43.485 48.440 43.745 ;
        RECT 48.500 43.485 48.760 43.745 ;
        RECT 48.820 43.485 49.080 43.745 ;
        RECT 49.140 43.485 49.400 43.745 ;
        RECT 48.180 41.130 48.440 41.390 ;
        RECT 48.500 41.130 48.760 41.390 ;
        RECT 48.820 41.130 49.080 41.390 ;
        RECT 49.140 41.130 49.400 41.390 ;
        RECT 55.690 45.845 55.950 46.105 ;
        RECT 56.010 45.845 56.270 46.105 ;
        RECT 56.330 45.845 56.590 46.105 ;
        RECT 56.650 45.845 56.910 46.105 ;
        RECT 55.690 43.485 55.950 43.745 ;
        RECT 56.010 43.485 56.270 43.745 ;
        RECT 56.330 43.485 56.590 43.745 ;
        RECT 56.650 43.485 56.910 43.745 ;
        RECT 55.690 41.130 55.950 41.390 ;
        RECT 56.010 41.130 56.270 41.390 ;
        RECT 56.330 41.130 56.590 41.390 ;
        RECT 56.650 41.130 56.910 41.390 ;
        RECT 63.365 45.845 63.625 46.105 ;
        RECT 63.685 45.845 63.945 46.105 ;
        RECT 64.005 45.845 64.265 46.105 ;
        RECT 64.325 45.845 64.585 46.105 ;
        RECT 63.365 43.485 63.625 43.745 ;
        RECT 63.685 43.485 63.945 43.745 ;
        RECT 64.005 43.485 64.265 43.745 ;
        RECT 64.325 43.485 64.585 43.745 ;
        RECT 63.365 41.130 63.625 41.390 ;
        RECT 63.685 41.130 63.945 41.390 ;
        RECT 64.005 41.130 64.265 41.390 ;
        RECT 64.325 41.130 64.585 41.390 ;
        RECT 70.875 45.845 71.135 46.105 ;
        RECT 71.195 45.845 71.455 46.105 ;
        RECT 71.515 45.845 71.775 46.105 ;
        RECT 71.835 45.845 72.095 46.105 ;
        RECT 70.875 43.485 71.135 43.745 ;
        RECT 71.195 43.485 71.455 43.745 ;
        RECT 71.515 43.485 71.775 43.745 ;
        RECT 71.835 43.485 72.095 43.745 ;
        RECT 70.875 41.130 71.135 41.390 ;
        RECT 71.195 41.130 71.455 41.390 ;
        RECT 71.515 41.130 71.775 41.390 ;
        RECT 71.835 41.130 72.095 41.390 ;
        RECT 8.110 38.770 8.370 39.030 ;
        RECT 8.430 38.770 8.690 39.030 ;
        RECT 8.750 38.770 9.010 39.030 ;
        RECT 9.070 38.770 9.330 39.030 ;
        RECT 8.110 36.410 8.370 36.670 ;
        RECT 8.430 36.410 8.690 36.670 ;
        RECT 8.750 36.410 9.010 36.670 ;
        RECT 9.070 36.410 9.330 36.670 ;
        RECT 8.110 34.050 8.370 34.310 ;
        RECT 8.430 34.050 8.690 34.310 ;
        RECT 8.750 34.050 9.010 34.310 ;
        RECT 9.070 34.050 9.330 34.310 ;
        RECT 8.110 31.690 8.370 31.950 ;
        RECT 8.430 31.690 8.690 31.950 ;
        RECT 8.750 31.690 9.010 31.950 ;
        RECT 9.070 31.690 9.330 31.950 ;
        RECT 8.110 29.330 8.370 29.590 ;
        RECT 8.430 29.330 8.690 29.590 ;
        RECT 8.750 29.330 9.010 29.590 ;
        RECT 9.070 29.330 9.330 29.590 ;
        RECT 12.595 38.770 12.855 39.030 ;
        RECT 12.915 38.770 13.175 39.030 ;
        RECT 13.235 38.770 13.495 39.030 ;
        RECT 13.555 38.770 13.815 39.030 ;
        RECT 12.595 36.410 12.855 36.670 ;
        RECT 12.915 36.410 13.175 36.670 ;
        RECT 13.235 36.410 13.495 36.670 ;
        RECT 13.555 36.410 13.815 36.670 ;
        RECT 12.595 34.050 12.855 34.310 ;
        RECT 12.915 34.050 13.175 34.310 ;
        RECT 13.235 34.050 13.495 34.310 ;
        RECT 13.555 34.050 13.815 34.310 ;
        RECT 12.595 31.690 12.855 31.950 ;
        RECT 12.915 31.690 13.175 31.950 ;
        RECT 13.235 31.690 13.495 31.950 ;
        RECT 13.555 31.690 13.815 31.950 ;
        RECT 12.595 29.330 12.855 29.590 ;
        RECT 12.915 29.330 13.175 29.590 ;
        RECT 13.235 29.330 13.495 29.590 ;
        RECT 13.555 29.330 13.815 29.590 ;
        RECT 18.055 38.770 18.315 39.030 ;
        RECT 18.375 38.770 18.635 39.030 ;
        RECT 18.695 38.770 18.955 39.030 ;
        RECT 19.015 38.770 19.275 39.030 ;
        RECT 18.055 36.410 18.315 36.670 ;
        RECT 18.375 36.410 18.635 36.670 ;
        RECT 18.695 36.410 18.955 36.670 ;
        RECT 19.015 36.410 19.275 36.670 ;
        RECT 18.055 34.050 18.315 34.310 ;
        RECT 18.375 34.050 18.635 34.310 ;
        RECT 18.695 34.050 18.955 34.310 ;
        RECT 19.015 34.050 19.275 34.310 ;
        RECT 18.055 31.690 18.315 31.950 ;
        RECT 18.375 31.690 18.635 31.950 ;
        RECT 18.695 31.690 18.955 31.950 ;
        RECT 19.015 31.690 19.275 31.950 ;
        RECT 18.055 29.330 18.315 29.590 ;
        RECT 18.375 29.330 18.635 29.590 ;
        RECT 18.695 29.330 18.955 29.590 ;
        RECT 19.015 29.330 19.275 29.590 ;
        RECT 25.080 38.770 25.340 39.030 ;
        RECT 25.400 38.770 25.660 39.030 ;
        RECT 25.720 38.770 25.980 39.030 ;
        RECT 26.040 38.770 26.300 39.030 ;
        RECT 25.080 36.410 25.340 36.670 ;
        RECT 25.400 36.410 25.660 36.670 ;
        RECT 25.720 36.410 25.980 36.670 ;
        RECT 26.040 36.410 26.300 36.670 ;
        RECT 25.080 34.050 25.340 34.310 ;
        RECT 25.400 34.050 25.660 34.310 ;
        RECT 25.720 34.050 25.980 34.310 ;
        RECT 26.040 34.050 26.300 34.310 ;
        RECT 25.080 31.690 25.340 31.950 ;
        RECT 25.400 31.690 25.660 31.950 ;
        RECT 25.720 31.690 25.980 31.950 ;
        RECT 26.040 31.690 26.300 31.950 ;
        RECT 25.080 29.330 25.340 29.590 ;
        RECT 25.400 29.330 25.660 29.590 ;
        RECT 25.720 29.330 25.980 29.590 ;
        RECT 26.040 29.330 26.300 29.590 ;
        RECT 32.815 38.770 33.075 39.030 ;
        RECT 33.135 38.770 33.395 39.030 ;
        RECT 33.455 38.770 33.715 39.030 ;
        RECT 33.775 38.770 34.035 39.030 ;
        RECT 32.815 36.410 33.075 36.670 ;
        RECT 33.135 36.410 33.395 36.670 ;
        RECT 33.455 36.410 33.715 36.670 ;
        RECT 33.775 36.410 34.035 36.670 ;
        RECT 32.815 34.050 33.075 34.310 ;
        RECT 33.135 34.050 33.395 34.310 ;
        RECT 33.455 34.050 33.715 34.310 ;
        RECT 33.775 34.050 34.035 34.310 ;
        RECT 32.815 31.690 33.075 31.950 ;
        RECT 33.135 31.690 33.395 31.950 ;
        RECT 33.455 31.690 33.715 31.950 ;
        RECT 33.775 31.690 34.035 31.950 ;
        RECT 32.815 29.330 33.075 29.590 ;
        RECT 33.135 29.330 33.395 29.590 ;
        RECT 33.455 29.330 33.715 29.590 ;
        RECT 33.775 29.330 34.035 29.590 ;
        RECT 40.370 38.770 40.630 39.030 ;
        RECT 40.690 38.770 40.950 39.030 ;
        RECT 41.010 38.770 41.270 39.030 ;
        RECT 41.330 38.770 41.590 39.030 ;
        RECT 40.370 36.410 40.630 36.670 ;
        RECT 40.690 36.410 40.950 36.670 ;
        RECT 41.010 36.410 41.270 36.670 ;
        RECT 41.330 36.410 41.590 36.670 ;
        RECT 40.370 34.050 40.630 34.310 ;
        RECT 40.690 34.050 40.950 34.310 ;
        RECT 41.010 34.050 41.270 34.310 ;
        RECT 41.330 34.050 41.590 34.310 ;
        RECT 40.370 31.690 40.630 31.950 ;
        RECT 40.690 31.690 40.950 31.950 ;
        RECT 41.010 31.690 41.270 31.950 ;
        RECT 41.330 31.690 41.590 31.950 ;
        RECT 40.370 29.330 40.630 29.590 ;
        RECT 40.690 29.330 40.950 29.590 ;
        RECT 41.010 29.330 41.270 29.590 ;
        RECT 41.330 29.330 41.590 29.590 ;
        RECT 48.180 38.770 48.440 39.030 ;
        RECT 48.500 38.770 48.760 39.030 ;
        RECT 48.820 38.770 49.080 39.030 ;
        RECT 49.140 38.770 49.400 39.030 ;
        RECT 48.180 36.410 48.440 36.670 ;
        RECT 48.500 36.410 48.760 36.670 ;
        RECT 48.820 36.410 49.080 36.670 ;
        RECT 49.140 36.410 49.400 36.670 ;
        RECT 48.180 34.050 48.440 34.310 ;
        RECT 48.500 34.050 48.760 34.310 ;
        RECT 48.820 34.050 49.080 34.310 ;
        RECT 49.140 34.050 49.400 34.310 ;
        RECT 48.180 31.690 48.440 31.950 ;
        RECT 48.500 31.690 48.760 31.950 ;
        RECT 48.820 31.690 49.080 31.950 ;
        RECT 49.140 31.690 49.400 31.950 ;
        RECT 48.180 29.330 48.440 29.590 ;
        RECT 48.500 29.330 48.760 29.590 ;
        RECT 48.820 29.330 49.080 29.590 ;
        RECT 49.140 29.330 49.400 29.590 ;
        RECT 55.690 38.770 55.950 39.030 ;
        RECT 56.010 38.770 56.270 39.030 ;
        RECT 56.330 38.770 56.590 39.030 ;
        RECT 56.650 38.770 56.910 39.030 ;
        RECT 55.690 36.410 55.950 36.670 ;
        RECT 56.010 36.410 56.270 36.670 ;
        RECT 56.330 36.410 56.590 36.670 ;
        RECT 56.650 36.410 56.910 36.670 ;
        RECT 55.690 34.050 55.950 34.310 ;
        RECT 56.010 34.050 56.270 34.310 ;
        RECT 56.330 34.050 56.590 34.310 ;
        RECT 56.650 34.050 56.910 34.310 ;
        RECT 55.690 31.690 55.950 31.950 ;
        RECT 56.010 31.690 56.270 31.950 ;
        RECT 56.330 31.690 56.590 31.950 ;
        RECT 56.650 31.690 56.910 31.950 ;
        RECT 55.690 29.330 55.950 29.590 ;
        RECT 56.010 29.330 56.270 29.590 ;
        RECT 56.330 29.330 56.590 29.590 ;
        RECT 56.650 29.330 56.910 29.590 ;
        RECT 63.365 38.770 63.625 39.030 ;
        RECT 63.685 38.770 63.945 39.030 ;
        RECT 64.005 38.770 64.265 39.030 ;
        RECT 64.325 38.770 64.585 39.030 ;
        RECT 63.365 36.410 63.625 36.670 ;
        RECT 63.685 36.410 63.945 36.670 ;
        RECT 64.005 36.410 64.265 36.670 ;
        RECT 64.325 36.410 64.585 36.670 ;
        RECT 63.365 34.050 63.625 34.310 ;
        RECT 63.685 34.050 63.945 34.310 ;
        RECT 64.005 34.050 64.265 34.310 ;
        RECT 64.325 34.050 64.585 34.310 ;
        RECT 63.365 31.690 63.625 31.950 ;
        RECT 63.685 31.690 63.945 31.950 ;
        RECT 64.005 31.690 64.265 31.950 ;
        RECT 64.325 31.690 64.585 31.950 ;
        RECT 63.365 29.330 63.625 29.590 ;
        RECT 63.685 29.330 63.945 29.590 ;
        RECT 64.005 29.330 64.265 29.590 ;
        RECT 64.325 29.330 64.585 29.590 ;
        RECT 70.875 38.770 71.135 39.030 ;
        RECT 71.195 38.770 71.455 39.030 ;
        RECT 71.515 38.770 71.775 39.030 ;
        RECT 71.835 38.770 72.095 39.030 ;
        RECT 70.875 36.410 71.135 36.670 ;
        RECT 71.195 36.410 71.455 36.670 ;
        RECT 71.515 36.410 71.775 36.670 ;
        RECT 71.835 36.410 72.095 36.670 ;
        RECT 70.875 34.050 71.135 34.310 ;
        RECT 71.195 34.050 71.455 34.310 ;
        RECT 71.515 34.050 71.775 34.310 ;
        RECT 71.835 34.050 72.095 34.310 ;
        RECT 70.875 31.690 71.135 31.950 ;
        RECT 71.195 31.690 71.455 31.950 ;
        RECT 71.515 31.690 71.775 31.950 ;
        RECT 71.835 31.690 72.095 31.950 ;
        RECT 70.875 29.330 71.135 29.590 ;
        RECT 71.195 29.330 71.455 29.590 ;
        RECT 71.515 29.330 71.775 29.590 ;
        RECT 71.835 29.330 72.095 29.590 ;
        RECT 8.110 26.970 8.370 27.230 ;
        RECT 8.430 26.970 8.690 27.230 ;
        RECT 8.750 26.970 9.010 27.230 ;
        RECT 9.070 26.970 9.330 27.230 ;
        RECT 8.110 24.610 8.370 24.870 ;
        RECT 8.430 24.610 8.690 24.870 ;
        RECT 8.750 24.610 9.010 24.870 ;
        RECT 9.070 24.610 9.330 24.870 ;
        RECT 8.110 22.250 8.370 22.510 ;
        RECT 8.430 22.250 8.690 22.510 ;
        RECT 8.750 22.250 9.010 22.510 ;
        RECT 9.070 22.250 9.330 22.510 ;
        RECT 8.110 19.890 8.370 20.150 ;
        RECT 8.430 19.890 8.690 20.150 ;
        RECT 8.750 19.890 9.010 20.150 ;
        RECT 9.070 19.890 9.330 20.150 ;
        RECT 8.110 17.530 8.370 17.790 ;
        RECT 8.430 17.530 8.690 17.790 ;
        RECT 8.750 17.530 9.010 17.790 ;
        RECT 9.070 17.530 9.330 17.790 ;
        RECT 12.595 26.970 12.855 27.230 ;
        RECT 12.915 26.970 13.175 27.230 ;
        RECT 13.235 26.970 13.495 27.230 ;
        RECT 13.555 26.970 13.815 27.230 ;
        RECT 12.595 24.610 12.855 24.870 ;
        RECT 12.915 24.610 13.175 24.870 ;
        RECT 13.235 24.610 13.495 24.870 ;
        RECT 13.555 24.610 13.815 24.870 ;
        RECT 12.595 22.250 12.855 22.510 ;
        RECT 12.915 22.250 13.175 22.510 ;
        RECT 13.235 22.250 13.495 22.510 ;
        RECT 13.555 22.250 13.815 22.510 ;
        RECT 12.595 19.890 12.855 20.150 ;
        RECT 12.915 19.890 13.175 20.150 ;
        RECT 13.235 19.890 13.495 20.150 ;
        RECT 13.555 19.890 13.815 20.150 ;
        RECT 12.595 17.530 12.855 17.790 ;
        RECT 12.915 17.530 13.175 17.790 ;
        RECT 13.235 17.530 13.495 17.790 ;
        RECT 13.555 17.530 13.815 17.790 ;
        RECT 18.055 26.970 18.315 27.230 ;
        RECT 18.375 26.970 18.635 27.230 ;
        RECT 18.695 26.970 18.955 27.230 ;
        RECT 19.015 26.970 19.275 27.230 ;
        RECT 18.055 24.610 18.315 24.870 ;
        RECT 18.375 24.610 18.635 24.870 ;
        RECT 18.695 24.610 18.955 24.870 ;
        RECT 19.015 24.610 19.275 24.870 ;
        RECT 18.055 22.250 18.315 22.510 ;
        RECT 18.375 22.250 18.635 22.510 ;
        RECT 18.695 22.250 18.955 22.510 ;
        RECT 19.015 22.250 19.275 22.510 ;
        RECT 18.055 19.890 18.315 20.150 ;
        RECT 18.375 19.890 18.635 20.150 ;
        RECT 18.695 19.890 18.955 20.150 ;
        RECT 19.015 19.890 19.275 20.150 ;
        RECT 18.055 17.530 18.315 17.790 ;
        RECT 18.375 17.530 18.635 17.790 ;
        RECT 18.695 17.530 18.955 17.790 ;
        RECT 19.015 17.530 19.275 17.790 ;
        RECT 25.080 26.970 25.340 27.230 ;
        RECT 25.400 26.970 25.660 27.230 ;
        RECT 25.720 26.970 25.980 27.230 ;
        RECT 26.040 26.970 26.300 27.230 ;
        RECT 25.080 24.610 25.340 24.870 ;
        RECT 25.400 24.610 25.660 24.870 ;
        RECT 25.720 24.610 25.980 24.870 ;
        RECT 26.040 24.610 26.300 24.870 ;
        RECT 25.080 22.250 25.340 22.510 ;
        RECT 25.400 22.250 25.660 22.510 ;
        RECT 25.720 22.250 25.980 22.510 ;
        RECT 26.040 22.250 26.300 22.510 ;
        RECT 25.080 19.890 25.340 20.150 ;
        RECT 25.400 19.890 25.660 20.150 ;
        RECT 25.720 19.890 25.980 20.150 ;
        RECT 26.040 19.890 26.300 20.150 ;
        RECT 25.080 17.530 25.340 17.790 ;
        RECT 25.400 17.530 25.660 17.790 ;
        RECT 25.720 17.530 25.980 17.790 ;
        RECT 26.040 17.530 26.300 17.790 ;
        RECT 32.815 26.970 33.075 27.230 ;
        RECT 33.135 26.970 33.395 27.230 ;
        RECT 33.455 26.970 33.715 27.230 ;
        RECT 33.775 26.970 34.035 27.230 ;
        RECT 32.815 24.610 33.075 24.870 ;
        RECT 33.135 24.610 33.395 24.870 ;
        RECT 33.455 24.610 33.715 24.870 ;
        RECT 33.775 24.610 34.035 24.870 ;
        RECT 32.815 22.250 33.075 22.510 ;
        RECT 33.135 22.250 33.395 22.510 ;
        RECT 33.455 22.250 33.715 22.510 ;
        RECT 33.775 22.250 34.035 22.510 ;
        RECT 32.815 19.890 33.075 20.150 ;
        RECT 33.135 19.890 33.395 20.150 ;
        RECT 33.455 19.890 33.715 20.150 ;
        RECT 33.775 19.890 34.035 20.150 ;
        RECT 32.815 17.530 33.075 17.790 ;
        RECT 33.135 17.530 33.395 17.790 ;
        RECT 33.455 17.530 33.715 17.790 ;
        RECT 33.775 17.530 34.035 17.790 ;
        RECT 40.370 26.970 40.630 27.230 ;
        RECT 40.690 26.970 40.950 27.230 ;
        RECT 41.010 26.970 41.270 27.230 ;
        RECT 41.330 26.970 41.590 27.230 ;
        RECT 40.370 24.610 40.630 24.870 ;
        RECT 40.690 24.610 40.950 24.870 ;
        RECT 41.010 24.610 41.270 24.870 ;
        RECT 41.330 24.610 41.590 24.870 ;
        RECT 40.370 22.250 40.630 22.510 ;
        RECT 40.690 22.250 40.950 22.510 ;
        RECT 41.010 22.250 41.270 22.510 ;
        RECT 41.330 22.250 41.590 22.510 ;
        RECT 40.370 19.890 40.630 20.150 ;
        RECT 40.690 19.890 40.950 20.150 ;
        RECT 41.010 19.890 41.270 20.150 ;
        RECT 41.330 19.890 41.590 20.150 ;
        RECT 40.370 17.530 40.630 17.790 ;
        RECT 40.690 17.530 40.950 17.790 ;
        RECT 41.010 17.530 41.270 17.790 ;
        RECT 41.330 17.530 41.590 17.790 ;
        RECT 48.180 26.970 48.440 27.230 ;
        RECT 48.500 26.970 48.760 27.230 ;
        RECT 48.820 26.970 49.080 27.230 ;
        RECT 49.140 26.970 49.400 27.230 ;
        RECT 48.180 24.610 48.440 24.870 ;
        RECT 48.500 24.610 48.760 24.870 ;
        RECT 48.820 24.610 49.080 24.870 ;
        RECT 49.140 24.610 49.400 24.870 ;
        RECT 48.180 22.250 48.440 22.510 ;
        RECT 48.500 22.250 48.760 22.510 ;
        RECT 48.820 22.250 49.080 22.510 ;
        RECT 49.140 22.250 49.400 22.510 ;
        RECT 48.180 19.890 48.440 20.150 ;
        RECT 48.500 19.890 48.760 20.150 ;
        RECT 48.820 19.890 49.080 20.150 ;
        RECT 49.140 19.890 49.400 20.150 ;
        RECT 48.180 17.530 48.440 17.790 ;
        RECT 48.500 17.530 48.760 17.790 ;
        RECT 48.820 17.530 49.080 17.790 ;
        RECT 49.140 17.530 49.400 17.790 ;
        RECT 55.690 26.970 55.950 27.230 ;
        RECT 56.010 26.970 56.270 27.230 ;
        RECT 56.330 26.970 56.590 27.230 ;
        RECT 56.650 26.970 56.910 27.230 ;
        RECT 55.690 24.610 55.950 24.870 ;
        RECT 56.010 24.610 56.270 24.870 ;
        RECT 56.330 24.610 56.590 24.870 ;
        RECT 56.650 24.610 56.910 24.870 ;
        RECT 55.690 22.250 55.950 22.510 ;
        RECT 56.010 22.250 56.270 22.510 ;
        RECT 56.330 22.250 56.590 22.510 ;
        RECT 56.650 22.250 56.910 22.510 ;
        RECT 55.690 19.890 55.950 20.150 ;
        RECT 56.010 19.890 56.270 20.150 ;
        RECT 56.330 19.890 56.590 20.150 ;
        RECT 56.650 19.890 56.910 20.150 ;
        RECT 55.690 17.530 55.950 17.790 ;
        RECT 56.010 17.530 56.270 17.790 ;
        RECT 56.330 17.530 56.590 17.790 ;
        RECT 56.650 17.530 56.910 17.790 ;
        RECT 63.365 26.970 63.625 27.230 ;
        RECT 63.685 26.970 63.945 27.230 ;
        RECT 64.005 26.970 64.265 27.230 ;
        RECT 64.325 26.970 64.585 27.230 ;
        RECT 63.365 24.610 63.625 24.870 ;
        RECT 63.685 24.610 63.945 24.870 ;
        RECT 64.005 24.610 64.265 24.870 ;
        RECT 64.325 24.610 64.585 24.870 ;
        RECT 63.365 22.250 63.625 22.510 ;
        RECT 63.685 22.250 63.945 22.510 ;
        RECT 64.005 22.250 64.265 22.510 ;
        RECT 64.325 22.250 64.585 22.510 ;
        RECT 63.365 19.890 63.625 20.150 ;
        RECT 63.685 19.890 63.945 20.150 ;
        RECT 64.005 19.890 64.265 20.150 ;
        RECT 64.325 19.890 64.585 20.150 ;
        RECT 63.365 17.530 63.625 17.790 ;
        RECT 63.685 17.530 63.945 17.790 ;
        RECT 64.005 17.530 64.265 17.790 ;
        RECT 64.325 17.530 64.585 17.790 ;
        RECT 70.875 26.970 71.135 27.230 ;
        RECT 71.195 26.970 71.455 27.230 ;
        RECT 71.515 26.970 71.775 27.230 ;
        RECT 71.835 26.970 72.095 27.230 ;
        RECT 70.875 24.610 71.135 24.870 ;
        RECT 71.195 24.610 71.455 24.870 ;
        RECT 71.515 24.610 71.775 24.870 ;
        RECT 71.835 24.610 72.095 24.870 ;
        RECT 70.875 22.250 71.135 22.510 ;
        RECT 71.195 22.250 71.455 22.510 ;
        RECT 71.515 22.250 71.775 22.510 ;
        RECT 71.835 22.250 72.095 22.510 ;
        RECT 70.875 19.890 71.135 20.150 ;
        RECT 71.195 19.890 71.455 20.150 ;
        RECT 71.515 19.890 71.775 20.150 ;
        RECT 71.835 19.890 72.095 20.150 ;
        RECT 70.875 17.530 71.135 17.790 ;
        RECT 71.195 17.530 71.455 17.790 ;
        RECT 71.515 17.530 71.775 17.790 ;
        RECT 71.835 17.530 72.095 17.790 ;
        RECT 8.110 15.170 8.370 15.430 ;
        RECT 8.430 15.170 8.690 15.430 ;
        RECT 8.750 15.170 9.010 15.430 ;
        RECT 9.070 15.170 9.330 15.430 ;
        RECT 8.110 12.810 8.370 13.070 ;
        RECT 8.430 12.810 8.690 13.070 ;
        RECT 8.750 12.810 9.010 13.070 ;
        RECT 9.070 12.810 9.330 13.070 ;
        RECT 12.595 15.170 12.855 15.430 ;
        RECT 12.915 15.170 13.175 15.430 ;
        RECT 13.235 15.170 13.495 15.430 ;
        RECT 13.555 15.170 13.815 15.430 ;
        RECT 12.595 12.810 12.855 13.070 ;
        RECT 12.915 12.810 13.175 13.070 ;
        RECT 13.235 12.810 13.495 13.070 ;
        RECT 13.555 12.810 13.815 13.070 ;
        RECT 18.055 15.170 18.315 15.430 ;
        RECT 18.375 15.170 18.635 15.430 ;
        RECT 18.695 15.170 18.955 15.430 ;
        RECT 19.015 15.170 19.275 15.430 ;
        RECT 18.055 12.810 18.315 13.070 ;
        RECT 18.375 12.810 18.635 13.070 ;
        RECT 18.695 12.810 18.955 13.070 ;
        RECT 19.015 12.810 19.275 13.070 ;
        RECT 25.080 15.170 25.340 15.430 ;
        RECT 25.400 15.170 25.660 15.430 ;
        RECT 25.720 15.170 25.980 15.430 ;
        RECT 26.040 15.170 26.300 15.430 ;
        RECT 25.080 12.810 25.340 13.070 ;
        RECT 25.400 12.810 25.660 13.070 ;
        RECT 25.720 12.810 25.980 13.070 ;
        RECT 26.040 12.810 26.300 13.070 ;
        RECT 32.815 15.170 33.075 15.430 ;
        RECT 33.135 15.170 33.395 15.430 ;
        RECT 33.455 15.170 33.715 15.430 ;
        RECT 33.775 15.170 34.035 15.430 ;
        RECT 32.815 12.810 33.075 13.070 ;
        RECT 33.135 12.810 33.395 13.070 ;
        RECT 33.455 12.810 33.715 13.070 ;
        RECT 33.775 12.810 34.035 13.070 ;
        RECT 40.370 15.170 40.630 15.430 ;
        RECT 40.690 15.170 40.950 15.430 ;
        RECT 41.010 15.170 41.270 15.430 ;
        RECT 41.330 15.170 41.590 15.430 ;
        RECT 40.370 12.810 40.630 13.070 ;
        RECT 40.690 12.810 40.950 13.070 ;
        RECT 41.010 12.810 41.270 13.070 ;
        RECT 41.330 12.810 41.590 13.070 ;
        RECT 48.180 15.170 48.440 15.430 ;
        RECT 48.500 15.170 48.760 15.430 ;
        RECT 48.820 15.170 49.080 15.430 ;
        RECT 49.140 15.170 49.400 15.430 ;
        RECT 48.180 12.810 48.440 13.070 ;
        RECT 48.500 12.810 48.760 13.070 ;
        RECT 48.820 12.810 49.080 13.070 ;
        RECT 49.140 12.810 49.400 13.070 ;
        RECT 55.690 15.170 55.950 15.430 ;
        RECT 56.010 15.170 56.270 15.430 ;
        RECT 56.330 15.170 56.590 15.430 ;
        RECT 56.650 15.170 56.910 15.430 ;
        RECT 55.690 12.810 55.950 13.070 ;
        RECT 56.010 12.810 56.270 13.070 ;
        RECT 56.330 12.810 56.590 13.070 ;
        RECT 56.650 12.810 56.910 13.070 ;
        RECT 63.365 15.170 63.625 15.430 ;
        RECT 63.685 15.170 63.945 15.430 ;
        RECT 64.005 15.170 64.265 15.430 ;
        RECT 64.325 15.170 64.585 15.430 ;
        RECT 63.365 12.810 63.625 13.070 ;
        RECT 63.685 12.810 63.945 13.070 ;
        RECT 64.005 12.810 64.265 13.070 ;
        RECT 64.325 12.810 64.585 13.070 ;
        RECT 70.875 15.170 71.135 15.430 ;
        RECT 71.195 15.170 71.455 15.430 ;
        RECT 71.515 15.170 71.775 15.430 ;
        RECT 71.835 15.170 72.095 15.430 ;
        RECT 70.875 12.810 71.135 13.070 ;
        RECT 71.195 12.810 71.455 13.070 ;
        RECT 71.515 12.810 71.775 13.070 ;
        RECT 71.835 12.810 72.095 13.070 ;
      LAYER met2 ;
        RECT 8.080 12.810 9.360 48.820 ;
        RECT 12.565 12.810 13.845 48.785 ;
        RECT 18.025 12.810 19.305 48.785 ;
        RECT 25.050 12.810 26.330 48.785 ;
        RECT 32.785 12.810 34.065 48.785 ;
        RECT 40.340 12.810 41.620 48.785 ;
        RECT 48.150 12.810 49.430 48.785 ;
        RECT 55.660 12.810 56.940 48.785 ;
        RECT 63.335 12.810 64.615 48.785 ;
        RECT 70.845 12.810 72.125 48.785 ;
  END
END vref_gen_nmos_with_trim
END LIBRARY

