../sky130_temp_sensor/SLC.lef