../../../../test/Nangate45/Nangate45_tech.lef