VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

VIA Element_via1_2_41040_18_1_1140_36_36
  VIARULE M2_M1 ;
  CUTSIZE 0.018 0.018 ;
  LAYERS M1 V1 M2 ;
  CUTSPACING 0.018 0.018 ;
  ENCLOSURE 0 0 0.002 0 ;
  ROWCOL 1 1140 ;
END Element_via1_2_41040_18_1_1140_36_36

VIA Element_VIA23_1_3_36_36
    LAYER M2 ;
      RECT  -0.05 -0.009 0.05 0.009 ;
    LAYER M3 ;
      RECT  -0.045 -0.014 0.045 0.014 ;
    LAYER V2 ;
      RECT  0.027 -0.009 0.045 0.009 ;
      RECT  -0.009 -0.009 0.009 0.009 ;
      RECT  -0.045 -0.009 -0.027 0.009 ;
END Element_VIA23_1_3_36_36

VIA Element_VIA34_1_2_58_52
    LAYER M3 ;
      RECT  -0.04 -0.017 0.04 0.017 ;
    LAYER M4 ;
      RECT  -0.046 -0.012 0.046 0.012 ;
    LAYER V3 ;
      RECT  0.017 -0.012 0.035 0.012 ;
      RECT  -0.035 -0.012 -0.017 0.012 ;
END Element_VIA34_1_2_58_52

VIA Element_VIA45_1_2_58_58
    LAYER M4 ;
      RECT  -0.052 -0.012 0.052 0.012 ;
    LAYER M5 ;
      RECT  -0.06 -0.023 0.06 0.023 ;
    LAYER V4 ;
      RECT  0.017 -0.012 0.041 0.012 ;
      RECT  -0.041 -0.012 -0.017 0.012 ;
END Element_VIA45_1_2_58_58

VIA Element_VIA45_2_2_58_58
    LAYER M4 ;
      RECT  -0.052 -0.06 0.052 0.06 ;
    LAYER M5 ;
      RECT  -0.06 -0.052 0.06 0.052 ;
    LAYER V4 ;
      RECT  0.017 0.017 0.041 0.041 ;
      RECT  -0.041 0.017 -0.017 0.041 ;
      RECT  0.017 -0.041 0.041 -0.017 ;
      RECT  -0.041 -0.041 -0.017 -0.017 ;
END Element_VIA45_2_2_58_58

MACRO Element
  FOREIGN Element 0 0 ;
  CLASS BLOCK ;
  SIZE 43.2 BY 43.2 ;
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER M5 ;
        RECT  41.4 0.684 41.52 42.516 ;
        RECT  38.424 0.684 38.544 42.516 ;
        RECT  35.448 0.684 35.568 42.516 ;
        RECT  32.472 0.684 32.592 42.516 ;
        RECT  29.496 0.684 29.616 42.516 ;
        RECT  26.52 0.684 26.64 42.516 ;
        RECT  23.544 0.684 23.664 42.516 ;
        RECT  20.568 0.684 20.688 42.516 ;
        RECT  17.592 0.684 17.712 42.516 ;
        RECT  14.616 0.684 14.736 42.516 ;
        RECT  11.64 0.684 11.76 42.516 ;
        RECT  8.664 0.684 8.784 42.516 ;
        RECT  5.688 0.684 5.808 42.516 ;
        RECT  2.712 0.684 2.832 42.516 ;
      LAYER M2 ;
        RECT  1.08 41.841 42.12 41.859 ;
        RECT  1.08 41.301 42.12 41.319 ;
        RECT  1.08 40.761 42.12 40.779 ;
        RECT  1.08 40.221 42.12 40.239 ;
        RECT  1.08 39.681 42.12 39.699 ;
        RECT  1.08 39.141 42.12 39.159 ;
        RECT  1.08 38.601 42.12 38.619 ;
        RECT  1.08 38.061 42.12 38.079 ;
        RECT  1.08 37.521 42.12 37.539 ;
        RECT  1.08 36.981 42.12 36.999 ;
        RECT  1.08 36.441 42.12 36.459 ;
        RECT  1.08 35.901 42.12 35.919 ;
        RECT  1.08 35.361 42.12 35.379 ;
        RECT  1.08 34.821 42.12 34.839 ;
        RECT  1.08 34.281 42.12 34.299 ;
        RECT  1.08 33.741 42.12 33.759 ;
        RECT  1.08 33.201 42.12 33.219 ;
        RECT  1.08 32.661 42.12 32.679 ;
        RECT  1.08 32.121 42.12 32.139 ;
        RECT  1.08 31.581 42.12 31.599 ;
        RECT  1.08 31.041 42.12 31.059 ;
        RECT  1.08 30.501 42.12 30.519 ;
        RECT  1.08 29.961 42.12 29.979 ;
        RECT  1.08 29.421 42.12 29.439 ;
        RECT  1.08 28.881 42.12 28.899 ;
        RECT  1.08 28.341 42.12 28.359 ;
        RECT  1.08 27.801 42.12 27.819 ;
        RECT  1.08 27.261 42.12 27.279 ;
        RECT  1.08 26.721 42.12 26.739 ;
        RECT  1.08 26.181 42.12 26.199 ;
        RECT  1.08 25.641 42.12 25.659 ;
        RECT  1.08 25.101 42.12 25.119 ;
        RECT  1.08 24.561 42.12 24.579 ;
        RECT  1.08 24.021 42.12 24.039 ;
        RECT  1.08 23.481 42.12 23.499 ;
        RECT  1.08 22.941 42.12 22.959 ;
        RECT  1.08 22.401 42.12 22.419 ;
        RECT  1.08 21.861 42.12 21.879 ;
        RECT  1.08 21.321 42.12 21.339 ;
        RECT  1.08 20.781 42.12 20.799 ;
        RECT  1.08 20.241 42.12 20.259 ;
        RECT  1.08 19.701 42.12 19.719 ;
        RECT  1.08 19.161 42.12 19.179 ;
        RECT  1.08 18.621 42.12 18.639 ;
        RECT  1.08 18.081 42.12 18.099 ;
        RECT  1.08 17.541 42.12 17.559 ;
        RECT  1.08 17.001 42.12 17.019 ;
        RECT  1.08 16.461 42.12 16.479 ;
        RECT  1.08 15.921 42.12 15.939 ;
        RECT  1.08 15.381 42.12 15.399 ;
        RECT  1.08 14.841 42.12 14.859 ;
        RECT  1.08 14.301 42.12 14.319 ;
        RECT  1.08 13.761 42.12 13.779 ;
        RECT  1.08 13.221 42.12 13.239 ;
        RECT  1.08 12.681 42.12 12.699 ;
        RECT  1.08 12.141 42.12 12.159 ;
        RECT  1.08 11.601 42.12 11.619 ;
        RECT  1.08 11.061 42.12 11.079 ;
        RECT  1.08 10.521 42.12 10.539 ;
        RECT  1.08 9.981 42.12 9.999 ;
        RECT  1.08 9.441 42.12 9.459 ;
        RECT  1.08 8.901 42.12 8.919 ;
        RECT  1.08 8.361 42.12 8.379 ;
        RECT  1.08 7.821 42.12 7.839 ;
        RECT  1.08 7.281 42.12 7.299 ;
        RECT  1.08 6.741 42.12 6.759 ;
        RECT  1.08 6.201 42.12 6.219 ;
        RECT  1.08 5.661 42.12 5.679 ;
        RECT  1.08 5.121 42.12 5.139 ;
        RECT  1.08 4.581 42.12 4.599 ;
        RECT  1.08 4.041 42.12 4.059 ;
        RECT  1.08 3.501 42.12 3.519 ;
        RECT  1.08 2.961 42.12 2.979 ;
        RECT  1.08 2.421 42.12 2.439 ;
        RECT  1.08 1.881 42.12 1.899 ;
        RECT  1.08 1.341 42.12 1.359 ;
      LAYER M1 ;
        RECT  1.08 41.841 42.12 41.859 ;
        RECT  1.08 41.301 42.12 41.319 ;
        RECT  1.08 40.761 42.12 40.779 ;
        RECT  1.08 40.221 42.12 40.239 ;
        RECT  1.08 39.681 42.12 39.699 ;
        RECT  1.08 39.141 42.12 39.159 ;
        RECT  1.08 38.601 42.12 38.619 ;
        RECT  1.08 38.061 42.12 38.079 ;
        RECT  1.08 37.521 42.12 37.539 ;
        RECT  1.08 36.981 42.12 36.999 ;
        RECT  1.08 36.441 42.12 36.459 ;
        RECT  1.08 35.901 42.12 35.919 ;
        RECT  1.08 35.361 42.12 35.379 ;
        RECT  1.08 34.821 42.12 34.839 ;
        RECT  1.08 34.281 42.12 34.299 ;
        RECT  1.08 33.741 42.12 33.759 ;
        RECT  1.08 33.201 42.12 33.219 ;
        RECT  1.08 32.661 42.12 32.679 ;
        RECT  1.08 32.121 42.12 32.139 ;
        RECT  1.08 31.581 42.12 31.599 ;
        RECT  1.08 31.041 42.12 31.059 ;
        RECT  1.08 30.501 42.12 30.519 ;
        RECT  1.08 29.961 42.12 29.979 ;
        RECT  1.08 29.421 42.12 29.439 ;
        RECT  1.08 28.881 42.12 28.899 ;
        RECT  1.08 28.341 42.12 28.359 ;
        RECT  1.08 27.801 42.12 27.819 ;
        RECT  1.08 27.261 42.12 27.279 ;
        RECT  1.08 26.721 42.12 26.739 ;
        RECT  1.08 26.181 42.12 26.199 ;
        RECT  1.08 25.641 42.12 25.659 ;
        RECT  1.08 25.101 42.12 25.119 ;
        RECT  1.08 24.561 42.12 24.579 ;
        RECT  1.08 24.021 42.12 24.039 ;
        RECT  1.08 23.481 42.12 23.499 ;
        RECT  1.08 22.941 42.12 22.959 ;
        RECT  1.08 22.401 42.12 22.419 ;
        RECT  1.08 21.861 42.12 21.879 ;
        RECT  1.08 21.321 42.12 21.339 ;
        RECT  1.08 20.781 42.12 20.799 ;
        RECT  1.08 20.241 42.12 20.259 ;
        RECT  1.08 19.701 42.12 19.719 ;
        RECT  1.08 19.161 42.12 19.179 ;
        RECT  1.08 18.621 42.12 18.639 ;
        RECT  1.08 18.081 42.12 18.099 ;
        RECT  1.08 17.541 42.12 17.559 ;
        RECT  1.08 17.001 42.12 17.019 ;
        RECT  1.08 16.461 42.12 16.479 ;
        RECT  1.08 15.921 42.12 15.939 ;
        RECT  1.08 15.381 42.12 15.399 ;
        RECT  1.08 14.841 42.12 14.859 ;
        RECT  1.08 14.301 42.12 14.319 ;
        RECT  1.08 13.761 42.12 13.779 ;
        RECT  1.08 13.221 42.12 13.239 ;
        RECT  1.08 12.681 42.12 12.699 ;
        RECT  1.08 12.141 42.12 12.159 ;
        RECT  1.08 11.601 42.12 11.619 ;
        RECT  1.08 11.061 42.12 11.079 ;
        RECT  1.08 10.521 42.12 10.539 ;
        RECT  1.08 9.981 42.12 9.999 ;
        RECT  1.08 9.441 42.12 9.459 ;
        RECT  1.08 8.901 42.12 8.919 ;
        RECT  1.08 8.361 42.12 8.379 ;
        RECT  1.08 7.821 42.12 7.839 ;
        RECT  1.08 7.281 42.12 7.299 ;
        RECT  1.08 6.741 42.12 6.759 ;
        RECT  1.08 6.201 42.12 6.219 ;
        RECT  1.08 5.661 42.12 5.679 ;
        RECT  1.08 5.121 42.12 5.139 ;
        RECT  1.08 4.581 42.12 4.599 ;
        RECT  1.08 4.041 42.12 4.059 ;
        RECT  1.08 3.501 42.12 3.519 ;
        RECT  1.08 2.961 42.12 2.979 ;
        RECT  1.08 2.421 42.12 2.439 ;
        RECT  1.08 1.881 42.12 1.899 ;
        RECT  1.08 1.341 42.12 1.359 ;
      LAYER M5 ;
        RECT  42.396 0.684 42.516 42.516 ;
      LAYER M4 ;
        RECT  0.684 42.396 42.516 42.516 ;
        RECT  0.684 0.684 42.516 0.804 ;
      LAYER M5 ;
        RECT  0.684 0.684 0.804 42.516 ;
      VIA 42.456 42.456 Element_VIA45_2_2_58_58 ;
      VIA 42.456 0.744 Element_VIA45_2_2_58_58 ;
      VIA 41.46 42.456 Element_VIA45_2_2_58_58 ;
      VIA 41.46 0.744 Element_VIA45_2_2_58_58 ;
      VIA 38.484 42.456 Element_VIA45_2_2_58_58 ;
      VIA 38.484 0.744 Element_VIA45_2_2_58_58 ;
      VIA 35.508 42.456 Element_VIA45_2_2_58_58 ;
      VIA 35.508 0.744 Element_VIA45_2_2_58_58 ;
      VIA 32.532 42.456 Element_VIA45_2_2_58_58 ;
      VIA 32.532 0.744 Element_VIA45_2_2_58_58 ;
      VIA 29.556 42.456 Element_VIA45_2_2_58_58 ;
      VIA 29.556 0.744 Element_VIA45_2_2_58_58 ;
      VIA 26.58 42.456 Element_VIA45_2_2_58_58 ;
      VIA 26.58 0.744 Element_VIA45_2_2_58_58 ;
      VIA 23.604 42.456 Element_VIA45_2_2_58_58 ;
      VIA 23.604 0.744 Element_VIA45_2_2_58_58 ;
      VIA 20.628 42.456 Element_VIA45_2_2_58_58 ;
      VIA 20.628 0.744 Element_VIA45_2_2_58_58 ;
      VIA 17.652 42.456 Element_VIA45_2_2_58_58 ;
      VIA 17.652 0.744 Element_VIA45_2_2_58_58 ;
      VIA 14.676 42.456 Element_VIA45_2_2_58_58 ;
      VIA 14.676 0.744 Element_VIA45_2_2_58_58 ;
      VIA 11.7 42.456 Element_VIA45_2_2_58_58 ;
      VIA 11.7 0.744 Element_VIA45_2_2_58_58 ;
      VIA 8.724 42.456 Element_VIA45_2_2_58_58 ;
      VIA 8.724 0.744 Element_VIA45_2_2_58_58 ;
      VIA 5.748 42.456 Element_VIA45_2_2_58_58 ;
      VIA 5.748 0.744 Element_VIA45_2_2_58_58 ;
      VIA 2.772 42.456 Element_VIA45_2_2_58_58 ;
      VIA 2.772 0.744 Element_VIA45_2_2_58_58 ;
      VIA 0.744 42.456 Element_VIA45_2_2_58_58 ;
      VIA 0.744 0.744 Element_VIA45_2_2_58_58 ;
      VIA 41.46 41.85 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 41.833 41.505 41.867 ;
      VIA 41.46 41.85 Element_VIA34_1_2_58_52 ;
      VIA 41.46 41.85 Element_VIA23_1_3_36_36 ;
      VIA 41.46 41.31 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 41.293 41.505 41.327 ;
      VIA 41.46 41.31 Element_VIA34_1_2_58_52 ;
      VIA 41.46 41.31 Element_VIA23_1_3_36_36 ;
      VIA 41.46 40.77 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 40.753 41.505 40.787 ;
      VIA 41.46 40.77 Element_VIA34_1_2_58_52 ;
      VIA 41.46 40.77 Element_VIA23_1_3_36_36 ;
      VIA 41.46 40.23 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 40.213 41.505 40.247 ;
      VIA 41.46 40.23 Element_VIA34_1_2_58_52 ;
      VIA 41.46 40.23 Element_VIA23_1_3_36_36 ;
      VIA 41.46 39.69 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 39.673 41.505 39.707 ;
      VIA 41.46 39.69 Element_VIA34_1_2_58_52 ;
      VIA 41.46 39.69 Element_VIA23_1_3_36_36 ;
      VIA 41.46 39.15 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 39.133 41.505 39.167 ;
      VIA 41.46 39.15 Element_VIA34_1_2_58_52 ;
      VIA 41.46 39.15 Element_VIA23_1_3_36_36 ;
      VIA 41.46 38.61 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 38.593 41.505 38.627 ;
      VIA 41.46 38.61 Element_VIA34_1_2_58_52 ;
      VIA 41.46 38.61 Element_VIA23_1_3_36_36 ;
      VIA 41.46 38.07 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 38.053 41.505 38.087 ;
      VIA 41.46 38.07 Element_VIA34_1_2_58_52 ;
      VIA 41.46 38.07 Element_VIA23_1_3_36_36 ;
      VIA 41.46 37.53 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 37.513 41.505 37.547 ;
      VIA 41.46 37.53 Element_VIA34_1_2_58_52 ;
      VIA 41.46 37.53 Element_VIA23_1_3_36_36 ;
      VIA 41.46 36.99 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 36.973 41.505 37.007 ;
      VIA 41.46 36.99 Element_VIA34_1_2_58_52 ;
      VIA 41.46 36.99 Element_VIA23_1_3_36_36 ;
      VIA 41.46 36.45 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 36.433 41.505 36.467 ;
      VIA 41.46 36.45 Element_VIA34_1_2_58_52 ;
      VIA 41.46 36.45 Element_VIA23_1_3_36_36 ;
      VIA 41.46 35.91 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 35.893 41.505 35.927 ;
      VIA 41.46 35.91 Element_VIA34_1_2_58_52 ;
      VIA 41.46 35.91 Element_VIA23_1_3_36_36 ;
      VIA 41.46 35.37 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 35.353 41.505 35.387 ;
      VIA 41.46 35.37 Element_VIA34_1_2_58_52 ;
      VIA 41.46 35.37 Element_VIA23_1_3_36_36 ;
      VIA 41.46 34.83 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 34.813 41.505 34.847 ;
      VIA 41.46 34.83 Element_VIA34_1_2_58_52 ;
      VIA 41.46 34.83 Element_VIA23_1_3_36_36 ;
      VIA 41.46 34.29 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 34.273 41.505 34.307 ;
      VIA 41.46 34.29 Element_VIA34_1_2_58_52 ;
      VIA 41.46 34.29 Element_VIA23_1_3_36_36 ;
      VIA 41.46 33.75 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 33.733 41.505 33.767 ;
      VIA 41.46 33.75 Element_VIA34_1_2_58_52 ;
      VIA 41.46 33.75 Element_VIA23_1_3_36_36 ;
      VIA 41.46 33.21 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 33.193 41.505 33.227 ;
      VIA 41.46 33.21 Element_VIA34_1_2_58_52 ;
      VIA 41.46 33.21 Element_VIA23_1_3_36_36 ;
      VIA 41.46 32.67 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 32.653 41.505 32.687 ;
      VIA 41.46 32.67 Element_VIA34_1_2_58_52 ;
      VIA 41.46 32.67 Element_VIA23_1_3_36_36 ;
      VIA 41.46 32.13 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 32.113 41.505 32.147 ;
      VIA 41.46 32.13 Element_VIA34_1_2_58_52 ;
      VIA 41.46 32.13 Element_VIA23_1_3_36_36 ;
      VIA 41.46 31.59 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 31.573 41.505 31.607 ;
      VIA 41.46 31.59 Element_VIA34_1_2_58_52 ;
      VIA 41.46 31.59 Element_VIA23_1_3_36_36 ;
      VIA 41.46 31.05 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 31.033 41.505 31.067 ;
      VIA 41.46 31.05 Element_VIA34_1_2_58_52 ;
      VIA 41.46 31.05 Element_VIA23_1_3_36_36 ;
      VIA 41.46 30.51 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 30.493 41.505 30.527 ;
      VIA 41.46 30.51 Element_VIA34_1_2_58_52 ;
      VIA 41.46 30.51 Element_VIA23_1_3_36_36 ;
      VIA 41.46 29.97 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 29.953 41.505 29.987 ;
      VIA 41.46 29.97 Element_VIA34_1_2_58_52 ;
      VIA 41.46 29.97 Element_VIA23_1_3_36_36 ;
      VIA 41.46 29.43 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 29.413 41.505 29.447 ;
      VIA 41.46 29.43 Element_VIA34_1_2_58_52 ;
      VIA 41.46 29.43 Element_VIA23_1_3_36_36 ;
      VIA 41.46 28.89 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 28.873 41.505 28.907 ;
      VIA 41.46 28.89 Element_VIA34_1_2_58_52 ;
      VIA 41.46 28.89 Element_VIA23_1_3_36_36 ;
      VIA 41.46 28.35 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 28.333 41.505 28.367 ;
      VIA 41.46 28.35 Element_VIA34_1_2_58_52 ;
      VIA 41.46 28.35 Element_VIA23_1_3_36_36 ;
      VIA 41.46 27.81 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 27.793 41.505 27.827 ;
      VIA 41.46 27.81 Element_VIA34_1_2_58_52 ;
      VIA 41.46 27.81 Element_VIA23_1_3_36_36 ;
      VIA 41.46 27.27 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 27.253 41.505 27.287 ;
      VIA 41.46 27.27 Element_VIA34_1_2_58_52 ;
      VIA 41.46 27.27 Element_VIA23_1_3_36_36 ;
      VIA 41.46 26.73 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 26.713 41.505 26.747 ;
      VIA 41.46 26.73 Element_VIA34_1_2_58_52 ;
      VIA 41.46 26.73 Element_VIA23_1_3_36_36 ;
      VIA 41.46 26.19 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 26.173 41.505 26.207 ;
      VIA 41.46 26.19 Element_VIA34_1_2_58_52 ;
      VIA 41.46 26.19 Element_VIA23_1_3_36_36 ;
      VIA 41.46 25.65 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 25.633 41.505 25.667 ;
      VIA 41.46 25.65 Element_VIA34_1_2_58_52 ;
      VIA 41.46 25.65 Element_VIA23_1_3_36_36 ;
      VIA 41.46 25.11 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 25.093 41.505 25.127 ;
      VIA 41.46 25.11 Element_VIA34_1_2_58_52 ;
      VIA 41.46 25.11 Element_VIA23_1_3_36_36 ;
      VIA 41.46 24.57 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 24.553 41.505 24.587 ;
      VIA 41.46 24.57 Element_VIA34_1_2_58_52 ;
      VIA 41.46 24.57 Element_VIA23_1_3_36_36 ;
      VIA 41.46 24.03 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 24.013 41.505 24.047 ;
      VIA 41.46 24.03 Element_VIA34_1_2_58_52 ;
      VIA 41.46 24.03 Element_VIA23_1_3_36_36 ;
      VIA 41.46 23.49 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 23.473 41.505 23.507 ;
      VIA 41.46 23.49 Element_VIA34_1_2_58_52 ;
      VIA 41.46 23.49 Element_VIA23_1_3_36_36 ;
      VIA 41.46 22.95 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 22.933 41.505 22.967 ;
      VIA 41.46 22.95 Element_VIA34_1_2_58_52 ;
      VIA 41.46 22.95 Element_VIA23_1_3_36_36 ;
      VIA 41.46 22.41 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 22.393 41.505 22.427 ;
      VIA 41.46 22.41 Element_VIA34_1_2_58_52 ;
      VIA 41.46 22.41 Element_VIA23_1_3_36_36 ;
      VIA 41.46 21.87 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 21.853 41.505 21.887 ;
      VIA 41.46 21.87 Element_VIA34_1_2_58_52 ;
      VIA 41.46 21.87 Element_VIA23_1_3_36_36 ;
      VIA 41.46 21.33 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 21.313 41.505 21.347 ;
      VIA 41.46 21.33 Element_VIA34_1_2_58_52 ;
      VIA 41.46 21.33 Element_VIA23_1_3_36_36 ;
      VIA 41.46 20.79 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 20.773 41.505 20.807 ;
      VIA 41.46 20.79 Element_VIA34_1_2_58_52 ;
      VIA 41.46 20.79 Element_VIA23_1_3_36_36 ;
      VIA 41.46 20.25 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 20.233 41.505 20.267 ;
      VIA 41.46 20.25 Element_VIA34_1_2_58_52 ;
      VIA 41.46 20.25 Element_VIA23_1_3_36_36 ;
      VIA 41.46 19.71 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 19.693 41.505 19.727 ;
      VIA 41.46 19.71 Element_VIA34_1_2_58_52 ;
      VIA 41.46 19.71 Element_VIA23_1_3_36_36 ;
      VIA 41.46 19.17 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 19.153 41.505 19.187 ;
      VIA 41.46 19.17 Element_VIA34_1_2_58_52 ;
      VIA 41.46 19.17 Element_VIA23_1_3_36_36 ;
      VIA 41.46 18.63 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 18.613 41.505 18.647 ;
      VIA 41.46 18.63 Element_VIA34_1_2_58_52 ;
      VIA 41.46 18.63 Element_VIA23_1_3_36_36 ;
      VIA 41.46 18.09 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 18.073 41.505 18.107 ;
      VIA 41.46 18.09 Element_VIA34_1_2_58_52 ;
      VIA 41.46 18.09 Element_VIA23_1_3_36_36 ;
      VIA 41.46 17.55 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 17.533 41.505 17.567 ;
      VIA 41.46 17.55 Element_VIA34_1_2_58_52 ;
      VIA 41.46 17.55 Element_VIA23_1_3_36_36 ;
      VIA 41.46 17.01 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 16.993 41.505 17.027 ;
      VIA 41.46 17.01 Element_VIA34_1_2_58_52 ;
      VIA 41.46 17.01 Element_VIA23_1_3_36_36 ;
      VIA 41.46 16.47 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 16.453 41.505 16.487 ;
      VIA 41.46 16.47 Element_VIA34_1_2_58_52 ;
      VIA 41.46 16.47 Element_VIA23_1_3_36_36 ;
      VIA 41.46 15.93 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 15.913 41.505 15.947 ;
      VIA 41.46 15.93 Element_VIA34_1_2_58_52 ;
      VIA 41.46 15.93 Element_VIA23_1_3_36_36 ;
      VIA 41.46 15.39 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 15.373 41.505 15.407 ;
      VIA 41.46 15.39 Element_VIA34_1_2_58_52 ;
      VIA 41.46 15.39 Element_VIA23_1_3_36_36 ;
      VIA 41.46 14.85 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 14.833 41.505 14.867 ;
      VIA 41.46 14.85 Element_VIA34_1_2_58_52 ;
      VIA 41.46 14.85 Element_VIA23_1_3_36_36 ;
      VIA 41.46 14.31 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 14.293 41.505 14.327 ;
      VIA 41.46 14.31 Element_VIA34_1_2_58_52 ;
      VIA 41.46 14.31 Element_VIA23_1_3_36_36 ;
      VIA 41.46 13.77 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 13.753 41.505 13.787 ;
      VIA 41.46 13.77 Element_VIA34_1_2_58_52 ;
      VIA 41.46 13.77 Element_VIA23_1_3_36_36 ;
      VIA 41.46 13.23 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 13.213 41.505 13.247 ;
      VIA 41.46 13.23 Element_VIA34_1_2_58_52 ;
      VIA 41.46 13.23 Element_VIA23_1_3_36_36 ;
      VIA 41.46 12.69 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 12.673 41.505 12.707 ;
      VIA 41.46 12.69 Element_VIA34_1_2_58_52 ;
      VIA 41.46 12.69 Element_VIA23_1_3_36_36 ;
      VIA 41.46 12.15 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 12.133 41.505 12.167 ;
      VIA 41.46 12.15 Element_VIA34_1_2_58_52 ;
      VIA 41.46 12.15 Element_VIA23_1_3_36_36 ;
      VIA 41.46 11.61 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 11.593 41.505 11.627 ;
      VIA 41.46 11.61 Element_VIA34_1_2_58_52 ;
      VIA 41.46 11.61 Element_VIA23_1_3_36_36 ;
      VIA 41.46 11.07 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 11.053 41.505 11.087 ;
      VIA 41.46 11.07 Element_VIA34_1_2_58_52 ;
      VIA 41.46 11.07 Element_VIA23_1_3_36_36 ;
      VIA 41.46 10.53 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 10.513 41.505 10.547 ;
      VIA 41.46 10.53 Element_VIA34_1_2_58_52 ;
      VIA 41.46 10.53 Element_VIA23_1_3_36_36 ;
      VIA 41.46 9.99 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 9.973 41.505 10.007 ;
      VIA 41.46 9.99 Element_VIA34_1_2_58_52 ;
      VIA 41.46 9.99 Element_VIA23_1_3_36_36 ;
      VIA 41.46 9.45 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 9.433 41.505 9.467 ;
      VIA 41.46 9.45 Element_VIA34_1_2_58_52 ;
      VIA 41.46 9.45 Element_VIA23_1_3_36_36 ;
      VIA 41.46 8.91 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 8.893 41.505 8.927 ;
      VIA 41.46 8.91 Element_VIA34_1_2_58_52 ;
      VIA 41.46 8.91 Element_VIA23_1_3_36_36 ;
      VIA 41.46 8.37 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 8.353 41.505 8.387 ;
      VIA 41.46 8.37 Element_VIA34_1_2_58_52 ;
      VIA 41.46 8.37 Element_VIA23_1_3_36_36 ;
      VIA 41.46 7.83 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 7.813 41.505 7.847 ;
      VIA 41.46 7.83 Element_VIA34_1_2_58_52 ;
      VIA 41.46 7.83 Element_VIA23_1_3_36_36 ;
      VIA 41.46 7.29 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 7.273 41.505 7.307 ;
      VIA 41.46 7.29 Element_VIA34_1_2_58_52 ;
      VIA 41.46 7.29 Element_VIA23_1_3_36_36 ;
      VIA 41.46 6.75 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 6.733 41.505 6.767 ;
      VIA 41.46 6.75 Element_VIA34_1_2_58_52 ;
      VIA 41.46 6.75 Element_VIA23_1_3_36_36 ;
      VIA 41.46 6.21 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 6.193 41.505 6.227 ;
      VIA 41.46 6.21 Element_VIA34_1_2_58_52 ;
      VIA 41.46 6.21 Element_VIA23_1_3_36_36 ;
      VIA 41.46 5.67 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 5.653 41.505 5.687 ;
      VIA 41.46 5.67 Element_VIA34_1_2_58_52 ;
      VIA 41.46 5.67 Element_VIA23_1_3_36_36 ;
      VIA 41.46 5.13 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 5.113 41.505 5.147 ;
      VIA 41.46 5.13 Element_VIA34_1_2_58_52 ;
      VIA 41.46 5.13 Element_VIA23_1_3_36_36 ;
      VIA 41.46 4.59 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 4.573 41.505 4.607 ;
      VIA 41.46 4.59 Element_VIA34_1_2_58_52 ;
      VIA 41.46 4.59 Element_VIA23_1_3_36_36 ;
      VIA 41.46 4.05 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 4.033 41.505 4.067 ;
      VIA 41.46 4.05 Element_VIA34_1_2_58_52 ;
      VIA 41.46 4.05 Element_VIA23_1_3_36_36 ;
      VIA 41.46 3.51 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 3.493 41.505 3.527 ;
      VIA 41.46 3.51 Element_VIA34_1_2_58_52 ;
      VIA 41.46 3.51 Element_VIA23_1_3_36_36 ;
      VIA 41.46 2.97 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 2.953 41.505 2.987 ;
      VIA 41.46 2.97 Element_VIA34_1_2_58_52 ;
      VIA 41.46 2.97 Element_VIA23_1_3_36_36 ;
      VIA 41.46 2.43 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 2.413 41.505 2.447 ;
      VIA 41.46 2.43 Element_VIA34_1_2_58_52 ;
      VIA 41.46 2.43 Element_VIA23_1_3_36_36 ;
      VIA 41.46 1.89 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 1.873 41.505 1.907 ;
      VIA 41.46 1.89 Element_VIA34_1_2_58_52 ;
      VIA 41.46 1.89 Element_VIA23_1_3_36_36 ;
      VIA 41.46 1.35 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.415 1.333 41.505 1.367 ;
      VIA 41.46 1.35 Element_VIA34_1_2_58_52 ;
      VIA 41.46 1.35 Element_VIA23_1_3_36_36 ;
      VIA 38.484 41.85 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 41.833 38.529 41.867 ;
      VIA 38.484 41.85 Element_VIA34_1_2_58_52 ;
      VIA 38.484 41.85 Element_VIA23_1_3_36_36 ;
      VIA 38.484 41.31 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 41.293 38.529 41.327 ;
      VIA 38.484 41.31 Element_VIA34_1_2_58_52 ;
      VIA 38.484 41.31 Element_VIA23_1_3_36_36 ;
      VIA 38.484 40.77 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 40.753 38.529 40.787 ;
      VIA 38.484 40.77 Element_VIA34_1_2_58_52 ;
      VIA 38.484 40.77 Element_VIA23_1_3_36_36 ;
      VIA 38.484 40.23 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 40.213 38.529 40.247 ;
      VIA 38.484 40.23 Element_VIA34_1_2_58_52 ;
      VIA 38.484 40.23 Element_VIA23_1_3_36_36 ;
      VIA 38.484 39.69 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 39.673 38.529 39.707 ;
      VIA 38.484 39.69 Element_VIA34_1_2_58_52 ;
      VIA 38.484 39.69 Element_VIA23_1_3_36_36 ;
      VIA 38.484 39.15 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 39.133 38.529 39.167 ;
      VIA 38.484 39.15 Element_VIA34_1_2_58_52 ;
      VIA 38.484 39.15 Element_VIA23_1_3_36_36 ;
      VIA 38.484 38.61 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 38.593 38.529 38.627 ;
      VIA 38.484 38.61 Element_VIA34_1_2_58_52 ;
      VIA 38.484 38.61 Element_VIA23_1_3_36_36 ;
      VIA 38.484 38.07 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 38.053 38.529 38.087 ;
      VIA 38.484 38.07 Element_VIA34_1_2_58_52 ;
      VIA 38.484 38.07 Element_VIA23_1_3_36_36 ;
      VIA 38.484 37.53 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 37.513 38.529 37.547 ;
      VIA 38.484 37.53 Element_VIA34_1_2_58_52 ;
      VIA 38.484 37.53 Element_VIA23_1_3_36_36 ;
      VIA 38.484 36.99 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 36.973 38.529 37.007 ;
      VIA 38.484 36.99 Element_VIA34_1_2_58_52 ;
      VIA 38.484 36.99 Element_VIA23_1_3_36_36 ;
      VIA 38.484 36.45 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 36.433 38.529 36.467 ;
      VIA 38.484 36.45 Element_VIA34_1_2_58_52 ;
      VIA 38.484 36.45 Element_VIA23_1_3_36_36 ;
      VIA 38.484 35.91 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 35.893 38.529 35.927 ;
      VIA 38.484 35.91 Element_VIA34_1_2_58_52 ;
      VIA 38.484 35.91 Element_VIA23_1_3_36_36 ;
      VIA 38.484 35.37 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 35.353 38.529 35.387 ;
      VIA 38.484 35.37 Element_VIA34_1_2_58_52 ;
      VIA 38.484 35.37 Element_VIA23_1_3_36_36 ;
      VIA 38.484 34.83 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 34.813 38.529 34.847 ;
      VIA 38.484 34.83 Element_VIA34_1_2_58_52 ;
      VIA 38.484 34.83 Element_VIA23_1_3_36_36 ;
      VIA 38.484 34.29 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 34.273 38.529 34.307 ;
      VIA 38.484 34.29 Element_VIA34_1_2_58_52 ;
      VIA 38.484 34.29 Element_VIA23_1_3_36_36 ;
      VIA 38.484 33.75 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 33.733 38.529 33.767 ;
      VIA 38.484 33.75 Element_VIA34_1_2_58_52 ;
      VIA 38.484 33.75 Element_VIA23_1_3_36_36 ;
      VIA 38.484 33.21 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 33.193 38.529 33.227 ;
      VIA 38.484 33.21 Element_VIA34_1_2_58_52 ;
      VIA 38.484 33.21 Element_VIA23_1_3_36_36 ;
      VIA 38.484 32.67 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 32.653 38.529 32.687 ;
      VIA 38.484 32.67 Element_VIA34_1_2_58_52 ;
      VIA 38.484 32.67 Element_VIA23_1_3_36_36 ;
      VIA 38.484 32.13 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 32.113 38.529 32.147 ;
      VIA 38.484 32.13 Element_VIA34_1_2_58_52 ;
      VIA 38.484 32.13 Element_VIA23_1_3_36_36 ;
      VIA 38.484 31.59 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 31.573 38.529 31.607 ;
      VIA 38.484 31.59 Element_VIA34_1_2_58_52 ;
      VIA 38.484 31.59 Element_VIA23_1_3_36_36 ;
      VIA 38.484 31.05 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 31.033 38.529 31.067 ;
      VIA 38.484 31.05 Element_VIA34_1_2_58_52 ;
      VIA 38.484 31.05 Element_VIA23_1_3_36_36 ;
      VIA 38.484 30.51 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 30.493 38.529 30.527 ;
      VIA 38.484 30.51 Element_VIA34_1_2_58_52 ;
      VIA 38.484 30.51 Element_VIA23_1_3_36_36 ;
      VIA 38.484 29.97 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 29.953 38.529 29.987 ;
      VIA 38.484 29.97 Element_VIA34_1_2_58_52 ;
      VIA 38.484 29.97 Element_VIA23_1_3_36_36 ;
      VIA 38.484 29.43 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 29.413 38.529 29.447 ;
      VIA 38.484 29.43 Element_VIA34_1_2_58_52 ;
      VIA 38.484 29.43 Element_VIA23_1_3_36_36 ;
      VIA 38.484 28.89 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 28.873 38.529 28.907 ;
      VIA 38.484 28.89 Element_VIA34_1_2_58_52 ;
      VIA 38.484 28.89 Element_VIA23_1_3_36_36 ;
      VIA 38.484 28.35 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 28.333 38.529 28.367 ;
      VIA 38.484 28.35 Element_VIA34_1_2_58_52 ;
      VIA 38.484 28.35 Element_VIA23_1_3_36_36 ;
      VIA 38.484 27.81 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 27.793 38.529 27.827 ;
      VIA 38.484 27.81 Element_VIA34_1_2_58_52 ;
      VIA 38.484 27.81 Element_VIA23_1_3_36_36 ;
      VIA 38.484 27.27 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 27.253 38.529 27.287 ;
      VIA 38.484 27.27 Element_VIA34_1_2_58_52 ;
      VIA 38.484 27.27 Element_VIA23_1_3_36_36 ;
      VIA 38.484 26.73 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 26.713 38.529 26.747 ;
      VIA 38.484 26.73 Element_VIA34_1_2_58_52 ;
      VIA 38.484 26.73 Element_VIA23_1_3_36_36 ;
      VIA 38.484 26.19 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 26.173 38.529 26.207 ;
      VIA 38.484 26.19 Element_VIA34_1_2_58_52 ;
      VIA 38.484 26.19 Element_VIA23_1_3_36_36 ;
      VIA 38.484 25.65 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 25.633 38.529 25.667 ;
      VIA 38.484 25.65 Element_VIA34_1_2_58_52 ;
      VIA 38.484 25.65 Element_VIA23_1_3_36_36 ;
      VIA 38.484 25.11 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 25.093 38.529 25.127 ;
      VIA 38.484 25.11 Element_VIA34_1_2_58_52 ;
      VIA 38.484 25.11 Element_VIA23_1_3_36_36 ;
      VIA 38.484 24.57 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 24.553 38.529 24.587 ;
      VIA 38.484 24.57 Element_VIA34_1_2_58_52 ;
      VIA 38.484 24.57 Element_VIA23_1_3_36_36 ;
      VIA 38.484 24.03 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 24.013 38.529 24.047 ;
      VIA 38.484 24.03 Element_VIA34_1_2_58_52 ;
      VIA 38.484 24.03 Element_VIA23_1_3_36_36 ;
      VIA 38.484 23.49 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 23.473 38.529 23.507 ;
      VIA 38.484 23.49 Element_VIA34_1_2_58_52 ;
      VIA 38.484 23.49 Element_VIA23_1_3_36_36 ;
      VIA 38.484 22.95 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 22.933 38.529 22.967 ;
      VIA 38.484 22.95 Element_VIA34_1_2_58_52 ;
      VIA 38.484 22.95 Element_VIA23_1_3_36_36 ;
      VIA 38.484 22.41 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 22.393 38.529 22.427 ;
      VIA 38.484 22.41 Element_VIA34_1_2_58_52 ;
      VIA 38.484 22.41 Element_VIA23_1_3_36_36 ;
      VIA 38.484 21.87 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 21.853 38.529 21.887 ;
      VIA 38.484 21.87 Element_VIA34_1_2_58_52 ;
      VIA 38.484 21.87 Element_VIA23_1_3_36_36 ;
      VIA 38.484 21.33 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 21.313 38.529 21.347 ;
      VIA 38.484 21.33 Element_VIA34_1_2_58_52 ;
      VIA 38.484 21.33 Element_VIA23_1_3_36_36 ;
      VIA 38.484 20.79 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 20.773 38.529 20.807 ;
      VIA 38.484 20.79 Element_VIA34_1_2_58_52 ;
      VIA 38.484 20.79 Element_VIA23_1_3_36_36 ;
      VIA 38.484 20.25 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 20.233 38.529 20.267 ;
      VIA 38.484 20.25 Element_VIA34_1_2_58_52 ;
      VIA 38.484 20.25 Element_VIA23_1_3_36_36 ;
      VIA 38.484 19.71 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 19.693 38.529 19.727 ;
      VIA 38.484 19.71 Element_VIA34_1_2_58_52 ;
      VIA 38.484 19.71 Element_VIA23_1_3_36_36 ;
      VIA 38.484 19.17 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 19.153 38.529 19.187 ;
      VIA 38.484 19.17 Element_VIA34_1_2_58_52 ;
      VIA 38.484 19.17 Element_VIA23_1_3_36_36 ;
      VIA 38.484 18.63 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 18.613 38.529 18.647 ;
      VIA 38.484 18.63 Element_VIA34_1_2_58_52 ;
      VIA 38.484 18.63 Element_VIA23_1_3_36_36 ;
      VIA 38.484 18.09 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 18.073 38.529 18.107 ;
      VIA 38.484 18.09 Element_VIA34_1_2_58_52 ;
      VIA 38.484 18.09 Element_VIA23_1_3_36_36 ;
      VIA 38.484 17.55 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 17.533 38.529 17.567 ;
      VIA 38.484 17.55 Element_VIA34_1_2_58_52 ;
      VIA 38.484 17.55 Element_VIA23_1_3_36_36 ;
      VIA 38.484 17.01 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 16.993 38.529 17.027 ;
      VIA 38.484 17.01 Element_VIA34_1_2_58_52 ;
      VIA 38.484 17.01 Element_VIA23_1_3_36_36 ;
      VIA 38.484 16.47 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 16.453 38.529 16.487 ;
      VIA 38.484 16.47 Element_VIA34_1_2_58_52 ;
      VIA 38.484 16.47 Element_VIA23_1_3_36_36 ;
      VIA 38.484 15.93 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 15.913 38.529 15.947 ;
      VIA 38.484 15.93 Element_VIA34_1_2_58_52 ;
      VIA 38.484 15.93 Element_VIA23_1_3_36_36 ;
      VIA 38.484 15.39 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 15.373 38.529 15.407 ;
      VIA 38.484 15.39 Element_VIA34_1_2_58_52 ;
      VIA 38.484 15.39 Element_VIA23_1_3_36_36 ;
      VIA 38.484 14.85 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 14.833 38.529 14.867 ;
      VIA 38.484 14.85 Element_VIA34_1_2_58_52 ;
      VIA 38.484 14.85 Element_VIA23_1_3_36_36 ;
      VIA 38.484 14.31 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 14.293 38.529 14.327 ;
      VIA 38.484 14.31 Element_VIA34_1_2_58_52 ;
      VIA 38.484 14.31 Element_VIA23_1_3_36_36 ;
      VIA 38.484 13.77 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 13.753 38.529 13.787 ;
      VIA 38.484 13.77 Element_VIA34_1_2_58_52 ;
      VIA 38.484 13.77 Element_VIA23_1_3_36_36 ;
      VIA 38.484 13.23 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 13.213 38.529 13.247 ;
      VIA 38.484 13.23 Element_VIA34_1_2_58_52 ;
      VIA 38.484 13.23 Element_VIA23_1_3_36_36 ;
      VIA 38.484 12.69 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 12.673 38.529 12.707 ;
      VIA 38.484 12.69 Element_VIA34_1_2_58_52 ;
      VIA 38.484 12.69 Element_VIA23_1_3_36_36 ;
      VIA 38.484 12.15 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 12.133 38.529 12.167 ;
      VIA 38.484 12.15 Element_VIA34_1_2_58_52 ;
      VIA 38.484 12.15 Element_VIA23_1_3_36_36 ;
      VIA 38.484 11.61 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 11.593 38.529 11.627 ;
      VIA 38.484 11.61 Element_VIA34_1_2_58_52 ;
      VIA 38.484 11.61 Element_VIA23_1_3_36_36 ;
      VIA 38.484 11.07 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 11.053 38.529 11.087 ;
      VIA 38.484 11.07 Element_VIA34_1_2_58_52 ;
      VIA 38.484 11.07 Element_VIA23_1_3_36_36 ;
      VIA 38.484 10.53 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 10.513 38.529 10.547 ;
      VIA 38.484 10.53 Element_VIA34_1_2_58_52 ;
      VIA 38.484 10.53 Element_VIA23_1_3_36_36 ;
      VIA 38.484 9.99 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 9.973 38.529 10.007 ;
      VIA 38.484 9.99 Element_VIA34_1_2_58_52 ;
      VIA 38.484 9.99 Element_VIA23_1_3_36_36 ;
      VIA 38.484 9.45 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 9.433 38.529 9.467 ;
      VIA 38.484 9.45 Element_VIA34_1_2_58_52 ;
      VIA 38.484 9.45 Element_VIA23_1_3_36_36 ;
      VIA 38.484 8.91 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 8.893 38.529 8.927 ;
      VIA 38.484 8.91 Element_VIA34_1_2_58_52 ;
      VIA 38.484 8.91 Element_VIA23_1_3_36_36 ;
      VIA 38.484 8.37 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 8.353 38.529 8.387 ;
      VIA 38.484 8.37 Element_VIA34_1_2_58_52 ;
      VIA 38.484 8.37 Element_VIA23_1_3_36_36 ;
      VIA 38.484 7.83 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 7.813 38.529 7.847 ;
      VIA 38.484 7.83 Element_VIA34_1_2_58_52 ;
      VIA 38.484 7.83 Element_VIA23_1_3_36_36 ;
      VIA 38.484 7.29 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 7.273 38.529 7.307 ;
      VIA 38.484 7.29 Element_VIA34_1_2_58_52 ;
      VIA 38.484 7.29 Element_VIA23_1_3_36_36 ;
      VIA 38.484 6.75 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 6.733 38.529 6.767 ;
      VIA 38.484 6.75 Element_VIA34_1_2_58_52 ;
      VIA 38.484 6.75 Element_VIA23_1_3_36_36 ;
      VIA 38.484 6.21 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 6.193 38.529 6.227 ;
      VIA 38.484 6.21 Element_VIA34_1_2_58_52 ;
      VIA 38.484 6.21 Element_VIA23_1_3_36_36 ;
      VIA 38.484 5.67 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 5.653 38.529 5.687 ;
      VIA 38.484 5.67 Element_VIA34_1_2_58_52 ;
      VIA 38.484 5.67 Element_VIA23_1_3_36_36 ;
      VIA 38.484 5.13 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 5.113 38.529 5.147 ;
      VIA 38.484 5.13 Element_VIA34_1_2_58_52 ;
      VIA 38.484 5.13 Element_VIA23_1_3_36_36 ;
      VIA 38.484 4.59 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 4.573 38.529 4.607 ;
      VIA 38.484 4.59 Element_VIA34_1_2_58_52 ;
      VIA 38.484 4.59 Element_VIA23_1_3_36_36 ;
      VIA 38.484 4.05 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 4.033 38.529 4.067 ;
      VIA 38.484 4.05 Element_VIA34_1_2_58_52 ;
      VIA 38.484 4.05 Element_VIA23_1_3_36_36 ;
      VIA 38.484 3.51 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 3.493 38.529 3.527 ;
      VIA 38.484 3.51 Element_VIA34_1_2_58_52 ;
      VIA 38.484 3.51 Element_VIA23_1_3_36_36 ;
      VIA 38.484 2.97 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 2.953 38.529 2.987 ;
      VIA 38.484 2.97 Element_VIA34_1_2_58_52 ;
      VIA 38.484 2.97 Element_VIA23_1_3_36_36 ;
      VIA 38.484 2.43 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 2.413 38.529 2.447 ;
      VIA 38.484 2.43 Element_VIA34_1_2_58_52 ;
      VIA 38.484 2.43 Element_VIA23_1_3_36_36 ;
      VIA 38.484 1.89 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 1.873 38.529 1.907 ;
      VIA 38.484 1.89 Element_VIA34_1_2_58_52 ;
      VIA 38.484 1.89 Element_VIA23_1_3_36_36 ;
      VIA 38.484 1.35 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.439 1.333 38.529 1.367 ;
      VIA 38.484 1.35 Element_VIA34_1_2_58_52 ;
      VIA 38.484 1.35 Element_VIA23_1_3_36_36 ;
      VIA 35.508 41.85 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 41.833 35.553 41.867 ;
      VIA 35.508 41.85 Element_VIA34_1_2_58_52 ;
      VIA 35.508 41.85 Element_VIA23_1_3_36_36 ;
      VIA 35.508 41.31 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 41.293 35.553 41.327 ;
      VIA 35.508 41.31 Element_VIA34_1_2_58_52 ;
      VIA 35.508 41.31 Element_VIA23_1_3_36_36 ;
      VIA 35.508 40.77 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 40.753 35.553 40.787 ;
      VIA 35.508 40.77 Element_VIA34_1_2_58_52 ;
      VIA 35.508 40.77 Element_VIA23_1_3_36_36 ;
      VIA 35.508 40.23 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 40.213 35.553 40.247 ;
      VIA 35.508 40.23 Element_VIA34_1_2_58_52 ;
      VIA 35.508 40.23 Element_VIA23_1_3_36_36 ;
      VIA 35.508 39.69 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 39.673 35.553 39.707 ;
      VIA 35.508 39.69 Element_VIA34_1_2_58_52 ;
      VIA 35.508 39.69 Element_VIA23_1_3_36_36 ;
      VIA 35.508 39.15 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 39.133 35.553 39.167 ;
      VIA 35.508 39.15 Element_VIA34_1_2_58_52 ;
      VIA 35.508 39.15 Element_VIA23_1_3_36_36 ;
      VIA 35.508 38.61 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 38.593 35.553 38.627 ;
      VIA 35.508 38.61 Element_VIA34_1_2_58_52 ;
      VIA 35.508 38.61 Element_VIA23_1_3_36_36 ;
      VIA 35.508 38.07 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 38.053 35.553 38.087 ;
      VIA 35.508 38.07 Element_VIA34_1_2_58_52 ;
      VIA 35.508 38.07 Element_VIA23_1_3_36_36 ;
      VIA 35.508 37.53 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 37.513 35.553 37.547 ;
      VIA 35.508 37.53 Element_VIA34_1_2_58_52 ;
      VIA 35.508 37.53 Element_VIA23_1_3_36_36 ;
      VIA 35.508 36.99 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 36.973 35.553 37.007 ;
      VIA 35.508 36.99 Element_VIA34_1_2_58_52 ;
      VIA 35.508 36.99 Element_VIA23_1_3_36_36 ;
      VIA 35.508 36.45 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 36.433 35.553 36.467 ;
      VIA 35.508 36.45 Element_VIA34_1_2_58_52 ;
      VIA 35.508 36.45 Element_VIA23_1_3_36_36 ;
      VIA 35.508 35.91 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 35.893 35.553 35.927 ;
      VIA 35.508 35.91 Element_VIA34_1_2_58_52 ;
      VIA 35.508 35.91 Element_VIA23_1_3_36_36 ;
      VIA 35.508 35.37 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 35.353 35.553 35.387 ;
      VIA 35.508 35.37 Element_VIA34_1_2_58_52 ;
      VIA 35.508 35.37 Element_VIA23_1_3_36_36 ;
      VIA 35.508 34.83 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 34.813 35.553 34.847 ;
      VIA 35.508 34.83 Element_VIA34_1_2_58_52 ;
      VIA 35.508 34.83 Element_VIA23_1_3_36_36 ;
      VIA 35.508 34.29 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 34.273 35.553 34.307 ;
      VIA 35.508 34.29 Element_VIA34_1_2_58_52 ;
      VIA 35.508 34.29 Element_VIA23_1_3_36_36 ;
      VIA 35.508 33.75 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 33.733 35.553 33.767 ;
      VIA 35.508 33.75 Element_VIA34_1_2_58_52 ;
      VIA 35.508 33.75 Element_VIA23_1_3_36_36 ;
      VIA 35.508 33.21 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 33.193 35.553 33.227 ;
      VIA 35.508 33.21 Element_VIA34_1_2_58_52 ;
      VIA 35.508 33.21 Element_VIA23_1_3_36_36 ;
      VIA 35.508 32.67 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 32.653 35.553 32.687 ;
      VIA 35.508 32.67 Element_VIA34_1_2_58_52 ;
      VIA 35.508 32.67 Element_VIA23_1_3_36_36 ;
      VIA 35.508 32.13 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 32.113 35.553 32.147 ;
      VIA 35.508 32.13 Element_VIA34_1_2_58_52 ;
      VIA 35.508 32.13 Element_VIA23_1_3_36_36 ;
      VIA 35.508 31.59 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 31.573 35.553 31.607 ;
      VIA 35.508 31.59 Element_VIA34_1_2_58_52 ;
      VIA 35.508 31.59 Element_VIA23_1_3_36_36 ;
      VIA 35.508 31.05 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 31.033 35.553 31.067 ;
      VIA 35.508 31.05 Element_VIA34_1_2_58_52 ;
      VIA 35.508 31.05 Element_VIA23_1_3_36_36 ;
      VIA 35.508 30.51 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 30.493 35.553 30.527 ;
      VIA 35.508 30.51 Element_VIA34_1_2_58_52 ;
      VIA 35.508 30.51 Element_VIA23_1_3_36_36 ;
      VIA 35.508 29.97 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 29.953 35.553 29.987 ;
      VIA 35.508 29.97 Element_VIA34_1_2_58_52 ;
      VIA 35.508 29.97 Element_VIA23_1_3_36_36 ;
      VIA 35.508 29.43 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 29.413 35.553 29.447 ;
      VIA 35.508 29.43 Element_VIA34_1_2_58_52 ;
      VIA 35.508 29.43 Element_VIA23_1_3_36_36 ;
      VIA 35.508 28.89 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 28.873 35.553 28.907 ;
      VIA 35.508 28.89 Element_VIA34_1_2_58_52 ;
      VIA 35.508 28.89 Element_VIA23_1_3_36_36 ;
      VIA 35.508 28.35 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 28.333 35.553 28.367 ;
      VIA 35.508 28.35 Element_VIA34_1_2_58_52 ;
      VIA 35.508 28.35 Element_VIA23_1_3_36_36 ;
      VIA 35.508 27.81 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 27.793 35.553 27.827 ;
      VIA 35.508 27.81 Element_VIA34_1_2_58_52 ;
      VIA 35.508 27.81 Element_VIA23_1_3_36_36 ;
      VIA 35.508 27.27 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 27.253 35.553 27.287 ;
      VIA 35.508 27.27 Element_VIA34_1_2_58_52 ;
      VIA 35.508 27.27 Element_VIA23_1_3_36_36 ;
      VIA 35.508 26.73 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 26.713 35.553 26.747 ;
      VIA 35.508 26.73 Element_VIA34_1_2_58_52 ;
      VIA 35.508 26.73 Element_VIA23_1_3_36_36 ;
      VIA 35.508 26.19 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 26.173 35.553 26.207 ;
      VIA 35.508 26.19 Element_VIA34_1_2_58_52 ;
      VIA 35.508 26.19 Element_VIA23_1_3_36_36 ;
      VIA 35.508 25.65 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 25.633 35.553 25.667 ;
      VIA 35.508 25.65 Element_VIA34_1_2_58_52 ;
      VIA 35.508 25.65 Element_VIA23_1_3_36_36 ;
      VIA 35.508 25.11 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 25.093 35.553 25.127 ;
      VIA 35.508 25.11 Element_VIA34_1_2_58_52 ;
      VIA 35.508 25.11 Element_VIA23_1_3_36_36 ;
      VIA 35.508 24.57 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 24.553 35.553 24.587 ;
      VIA 35.508 24.57 Element_VIA34_1_2_58_52 ;
      VIA 35.508 24.57 Element_VIA23_1_3_36_36 ;
      VIA 35.508 24.03 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 24.013 35.553 24.047 ;
      VIA 35.508 24.03 Element_VIA34_1_2_58_52 ;
      VIA 35.508 24.03 Element_VIA23_1_3_36_36 ;
      VIA 35.508 23.49 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 23.473 35.553 23.507 ;
      VIA 35.508 23.49 Element_VIA34_1_2_58_52 ;
      VIA 35.508 23.49 Element_VIA23_1_3_36_36 ;
      VIA 35.508 22.95 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 22.933 35.553 22.967 ;
      VIA 35.508 22.95 Element_VIA34_1_2_58_52 ;
      VIA 35.508 22.95 Element_VIA23_1_3_36_36 ;
      VIA 35.508 22.41 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 22.393 35.553 22.427 ;
      VIA 35.508 22.41 Element_VIA34_1_2_58_52 ;
      VIA 35.508 22.41 Element_VIA23_1_3_36_36 ;
      VIA 35.508 21.87 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 21.853 35.553 21.887 ;
      VIA 35.508 21.87 Element_VIA34_1_2_58_52 ;
      VIA 35.508 21.87 Element_VIA23_1_3_36_36 ;
      VIA 35.508 21.33 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 21.313 35.553 21.347 ;
      VIA 35.508 21.33 Element_VIA34_1_2_58_52 ;
      VIA 35.508 21.33 Element_VIA23_1_3_36_36 ;
      VIA 35.508 20.79 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 20.773 35.553 20.807 ;
      VIA 35.508 20.79 Element_VIA34_1_2_58_52 ;
      VIA 35.508 20.79 Element_VIA23_1_3_36_36 ;
      VIA 35.508 20.25 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 20.233 35.553 20.267 ;
      VIA 35.508 20.25 Element_VIA34_1_2_58_52 ;
      VIA 35.508 20.25 Element_VIA23_1_3_36_36 ;
      VIA 35.508 19.71 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 19.693 35.553 19.727 ;
      VIA 35.508 19.71 Element_VIA34_1_2_58_52 ;
      VIA 35.508 19.71 Element_VIA23_1_3_36_36 ;
      VIA 35.508 19.17 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 19.153 35.553 19.187 ;
      VIA 35.508 19.17 Element_VIA34_1_2_58_52 ;
      VIA 35.508 19.17 Element_VIA23_1_3_36_36 ;
      VIA 35.508 18.63 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 18.613 35.553 18.647 ;
      VIA 35.508 18.63 Element_VIA34_1_2_58_52 ;
      VIA 35.508 18.63 Element_VIA23_1_3_36_36 ;
      VIA 35.508 18.09 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 18.073 35.553 18.107 ;
      VIA 35.508 18.09 Element_VIA34_1_2_58_52 ;
      VIA 35.508 18.09 Element_VIA23_1_3_36_36 ;
      VIA 35.508 17.55 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 17.533 35.553 17.567 ;
      VIA 35.508 17.55 Element_VIA34_1_2_58_52 ;
      VIA 35.508 17.55 Element_VIA23_1_3_36_36 ;
      VIA 35.508 17.01 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 16.993 35.553 17.027 ;
      VIA 35.508 17.01 Element_VIA34_1_2_58_52 ;
      VIA 35.508 17.01 Element_VIA23_1_3_36_36 ;
      VIA 35.508 16.47 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 16.453 35.553 16.487 ;
      VIA 35.508 16.47 Element_VIA34_1_2_58_52 ;
      VIA 35.508 16.47 Element_VIA23_1_3_36_36 ;
      VIA 35.508 15.93 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 15.913 35.553 15.947 ;
      VIA 35.508 15.93 Element_VIA34_1_2_58_52 ;
      VIA 35.508 15.93 Element_VIA23_1_3_36_36 ;
      VIA 35.508 15.39 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 15.373 35.553 15.407 ;
      VIA 35.508 15.39 Element_VIA34_1_2_58_52 ;
      VIA 35.508 15.39 Element_VIA23_1_3_36_36 ;
      VIA 35.508 14.85 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 14.833 35.553 14.867 ;
      VIA 35.508 14.85 Element_VIA34_1_2_58_52 ;
      VIA 35.508 14.85 Element_VIA23_1_3_36_36 ;
      VIA 35.508 14.31 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 14.293 35.553 14.327 ;
      VIA 35.508 14.31 Element_VIA34_1_2_58_52 ;
      VIA 35.508 14.31 Element_VIA23_1_3_36_36 ;
      VIA 35.508 13.77 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 13.753 35.553 13.787 ;
      VIA 35.508 13.77 Element_VIA34_1_2_58_52 ;
      VIA 35.508 13.77 Element_VIA23_1_3_36_36 ;
      VIA 35.508 13.23 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 13.213 35.553 13.247 ;
      VIA 35.508 13.23 Element_VIA34_1_2_58_52 ;
      VIA 35.508 13.23 Element_VIA23_1_3_36_36 ;
      VIA 35.508 12.69 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 12.673 35.553 12.707 ;
      VIA 35.508 12.69 Element_VIA34_1_2_58_52 ;
      VIA 35.508 12.69 Element_VIA23_1_3_36_36 ;
      VIA 35.508 12.15 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 12.133 35.553 12.167 ;
      VIA 35.508 12.15 Element_VIA34_1_2_58_52 ;
      VIA 35.508 12.15 Element_VIA23_1_3_36_36 ;
      VIA 35.508 11.61 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 11.593 35.553 11.627 ;
      VIA 35.508 11.61 Element_VIA34_1_2_58_52 ;
      VIA 35.508 11.61 Element_VIA23_1_3_36_36 ;
      VIA 35.508 11.07 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 11.053 35.553 11.087 ;
      VIA 35.508 11.07 Element_VIA34_1_2_58_52 ;
      VIA 35.508 11.07 Element_VIA23_1_3_36_36 ;
      VIA 35.508 10.53 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 10.513 35.553 10.547 ;
      VIA 35.508 10.53 Element_VIA34_1_2_58_52 ;
      VIA 35.508 10.53 Element_VIA23_1_3_36_36 ;
      VIA 35.508 9.99 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 9.973 35.553 10.007 ;
      VIA 35.508 9.99 Element_VIA34_1_2_58_52 ;
      VIA 35.508 9.99 Element_VIA23_1_3_36_36 ;
      VIA 35.508 9.45 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 9.433 35.553 9.467 ;
      VIA 35.508 9.45 Element_VIA34_1_2_58_52 ;
      VIA 35.508 9.45 Element_VIA23_1_3_36_36 ;
      VIA 35.508 8.91 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 8.893 35.553 8.927 ;
      VIA 35.508 8.91 Element_VIA34_1_2_58_52 ;
      VIA 35.508 8.91 Element_VIA23_1_3_36_36 ;
      VIA 35.508 8.37 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 8.353 35.553 8.387 ;
      VIA 35.508 8.37 Element_VIA34_1_2_58_52 ;
      VIA 35.508 8.37 Element_VIA23_1_3_36_36 ;
      VIA 35.508 7.83 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 7.813 35.553 7.847 ;
      VIA 35.508 7.83 Element_VIA34_1_2_58_52 ;
      VIA 35.508 7.83 Element_VIA23_1_3_36_36 ;
      VIA 35.508 7.29 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 7.273 35.553 7.307 ;
      VIA 35.508 7.29 Element_VIA34_1_2_58_52 ;
      VIA 35.508 7.29 Element_VIA23_1_3_36_36 ;
      VIA 35.508 6.75 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 6.733 35.553 6.767 ;
      VIA 35.508 6.75 Element_VIA34_1_2_58_52 ;
      VIA 35.508 6.75 Element_VIA23_1_3_36_36 ;
      VIA 35.508 6.21 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 6.193 35.553 6.227 ;
      VIA 35.508 6.21 Element_VIA34_1_2_58_52 ;
      VIA 35.508 6.21 Element_VIA23_1_3_36_36 ;
      VIA 35.508 5.67 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 5.653 35.553 5.687 ;
      VIA 35.508 5.67 Element_VIA34_1_2_58_52 ;
      VIA 35.508 5.67 Element_VIA23_1_3_36_36 ;
      VIA 35.508 5.13 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 5.113 35.553 5.147 ;
      VIA 35.508 5.13 Element_VIA34_1_2_58_52 ;
      VIA 35.508 5.13 Element_VIA23_1_3_36_36 ;
      VIA 35.508 4.59 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 4.573 35.553 4.607 ;
      VIA 35.508 4.59 Element_VIA34_1_2_58_52 ;
      VIA 35.508 4.59 Element_VIA23_1_3_36_36 ;
      VIA 35.508 4.05 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 4.033 35.553 4.067 ;
      VIA 35.508 4.05 Element_VIA34_1_2_58_52 ;
      VIA 35.508 4.05 Element_VIA23_1_3_36_36 ;
      VIA 35.508 3.51 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 3.493 35.553 3.527 ;
      VIA 35.508 3.51 Element_VIA34_1_2_58_52 ;
      VIA 35.508 3.51 Element_VIA23_1_3_36_36 ;
      VIA 35.508 2.97 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 2.953 35.553 2.987 ;
      VIA 35.508 2.97 Element_VIA34_1_2_58_52 ;
      VIA 35.508 2.97 Element_VIA23_1_3_36_36 ;
      VIA 35.508 2.43 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 2.413 35.553 2.447 ;
      VIA 35.508 2.43 Element_VIA34_1_2_58_52 ;
      VIA 35.508 2.43 Element_VIA23_1_3_36_36 ;
      VIA 35.508 1.89 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 1.873 35.553 1.907 ;
      VIA 35.508 1.89 Element_VIA34_1_2_58_52 ;
      VIA 35.508 1.89 Element_VIA23_1_3_36_36 ;
      VIA 35.508 1.35 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.463 1.333 35.553 1.367 ;
      VIA 35.508 1.35 Element_VIA34_1_2_58_52 ;
      VIA 35.508 1.35 Element_VIA23_1_3_36_36 ;
      VIA 32.532 41.85 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 41.833 32.577 41.867 ;
      VIA 32.532 41.85 Element_VIA34_1_2_58_52 ;
      VIA 32.532 41.85 Element_VIA23_1_3_36_36 ;
      VIA 32.532 41.31 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 41.293 32.577 41.327 ;
      VIA 32.532 41.31 Element_VIA34_1_2_58_52 ;
      VIA 32.532 41.31 Element_VIA23_1_3_36_36 ;
      VIA 32.532 40.77 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 40.753 32.577 40.787 ;
      VIA 32.532 40.77 Element_VIA34_1_2_58_52 ;
      VIA 32.532 40.77 Element_VIA23_1_3_36_36 ;
      VIA 32.532 40.23 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 40.213 32.577 40.247 ;
      VIA 32.532 40.23 Element_VIA34_1_2_58_52 ;
      VIA 32.532 40.23 Element_VIA23_1_3_36_36 ;
      VIA 32.532 39.69 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 39.673 32.577 39.707 ;
      VIA 32.532 39.69 Element_VIA34_1_2_58_52 ;
      VIA 32.532 39.69 Element_VIA23_1_3_36_36 ;
      VIA 32.532 39.15 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 39.133 32.577 39.167 ;
      VIA 32.532 39.15 Element_VIA34_1_2_58_52 ;
      VIA 32.532 39.15 Element_VIA23_1_3_36_36 ;
      VIA 32.532 38.61 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 38.593 32.577 38.627 ;
      VIA 32.532 38.61 Element_VIA34_1_2_58_52 ;
      VIA 32.532 38.61 Element_VIA23_1_3_36_36 ;
      VIA 32.532 38.07 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 38.053 32.577 38.087 ;
      VIA 32.532 38.07 Element_VIA34_1_2_58_52 ;
      VIA 32.532 38.07 Element_VIA23_1_3_36_36 ;
      VIA 32.532 37.53 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 37.513 32.577 37.547 ;
      VIA 32.532 37.53 Element_VIA34_1_2_58_52 ;
      VIA 32.532 37.53 Element_VIA23_1_3_36_36 ;
      VIA 32.532 36.99 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 36.973 32.577 37.007 ;
      VIA 32.532 36.99 Element_VIA34_1_2_58_52 ;
      VIA 32.532 36.99 Element_VIA23_1_3_36_36 ;
      VIA 32.532 36.45 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 36.433 32.577 36.467 ;
      VIA 32.532 36.45 Element_VIA34_1_2_58_52 ;
      VIA 32.532 36.45 Element_VIA23_1_3_36_36 ;
      VIA 32.532 35.91 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 35.893 32.577 35.927 ;
      VIA 32.532 35.91 Element_VIA34_1_2_58_52 ;
      VIA 32.532 35.91 Element_VIA23_1_3_36_36 ;
      VIA 32.532 35.37 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 35.353 32.577 35.387 ;
      VIA 32.532 35.37 Element_VIA34_1_2_58_52 ;
      VIA 32.532 35.37 Element_VIA23_1_3_36_36 ;
      VIA 32.532 34.83 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 34.813 32.577 34.847 ;
      VIA 32.532 34.83 Element_VIA34_1_2_58_52 ;
      VIA 32.532 34.83 Element_VIA23_1_3_36_36 ;
      VIA 32.532 34.29 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 34.273 32.577 34.307 ;
      VIA 32.532 34.29 Element_VIA34_1_2_58_52 ;
      VIA 32.532 34.29 Element_VIA23_1_3_36_36 ;
      VIA 32.532 33.75 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 33.733 32.577 33.767 ;
      VIA 32.532 33.75 Element_VIA34_1_2_58_52 ;
      VIA 32.532 33.75 Element_VIA23_1_3_36_36 ;
      VIA 32.532 33.21 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 33.193 32.577 33.227 ;
      VIA 32.532 33.21 Element_VIA34_1_2_58_52 ;
      VIA 32.532 33.21 Element_VIA23_1_3_36_36 ;
      VIA 32.532 32.67 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 32.653 32.577 32.687 ;
      VIA 32.532 32.67 Element_VIA34_1_2_58_52 ;
      VIA 32.532 32.67 Element_VIA23_1_3_36_36 ;
      VIA 32.532 32.13 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 32.113 32.577 32.147 ;
      VIA 32.532 32.13 Element_VIA34_1_2_58_52 ;
      VIA 32.532 32.13 Element_VIA23_1_3_36_36 ;
      VIA 32.532 31.59 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 31.573 32.577 31.607 ;
      VIA 32.532 31.59 Element_VIA34_1_2_58_52 ;
      VIA 32.532 31.59 Element_VIA23_1_3_36_36 ;
      VIA 32.532 31.05 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 31.033 32.577 31.067 ;
      VIA 32.532 31.05 Element_VIA34_1_2_58_52 ;
      VIA 32.532 31.05 Element_VIA23_1_3_36_36 ;
      VIA 32.532 30.51 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 30.493 32.577 30.527 ;
      VIA 32.532 30.51 Element_VIA34_1_2_58_52 ;
      VIA 32.532 30.51 Element_VIA23_1_3_36_36 ;
      VIA 32.532 29.97 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 29.953 32.577 29.987 ;
      VIA 32.532 29.97 Element_VIA34_1_2_58_52 ;
      VIA 32.532 29.97 Element_VIA23_1_3_36_36 ;
      VIA 32.532 29.43 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 29.413 32.577 29.447 ;
      VIA 32.532 29.43 Element_VIA34_1_2_58_52 ;
      VIA 32.532 29.43 Element_VIA23_1_3_36_36 ;
      VIA 32.532 28.89 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 28.873 32.577 28.907 ;
      VIA 32.532 28.89 Element_VIA34_1_2_58_52 ;
      VIA 32.532 28.89 Element_VIA23_1_3_36_36 ;
      VIA 32.532 28.35 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 28.333 32.577 28.367 ;
      VIA 32.532 28.35 Element_VIA34_1_2_58_52 ;
      VIA 32.532 28.35 Element_VIA23_1_3_36_36 ;
      VIA 32.532 27.81 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 27.793 32.577 27.827 ;
      VIA 32.532 27.81 Element_VIA34_1_2_58_52 ;
      VIA 32.532 27.81 Element_VIA23_1_3_36_36 ;
      VIA 32.532 27.27 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 27.253 32.577 27.287 ;
      VIA 32.532 27.27 Element_VIA34_1_2_58_52 ;
      VIA 32.532 27.27 Element_VIA23_1_3_36_36 ;
      VIA 32.532 26.73 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 26.713 32.577 26.747 ;
      VIA 32.532 26.73 Element_VIA34_1_2_58_52 ;
      VIA 32.532 26.73 Element_VIA23_1_3_36_36 ;
      VIA 32.532 26.19 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 26.173 32.577 26.207 ;
      VIA 32.532 26.19 Element_VIA34_1_2_58_52 ;
      VIA 32.532 26.19 Element_VIA23_1_3_36_36 ;
      VIA 32.532 25.65 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 25.633 32.577 25.667 ;
      VIA 32.532 25.65 Element_VIA34_1_2_58_52 ;
      VIA 32.532 25.65 Element_VIA23_1_3_36_36 ;
      VIA 32.532 25.11 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 25.093 32.577 25.127 ;
      VIA 32.532 25.11 Element_VIA34_1_2_58_52 ;
      VIA 32.532 25.11 Element_VIA23_1_3_36_36 ;
      VIA 32.532 24.57 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 24.553 32.577 24.587 ;
      VIA 32.532 24.57 Element_VIA34_1_2_58_52 ;
      VIA 32.532 24.57 Element_VIA23_1_3_36_36 ;
      VIA 32.532 24.03 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 24.013 32.577 24.047 ;
      VIA 32.532 24.03 Element_VIA34_1_2_58_52 ;
      VIA 32.532 24.03 Element_VIA23_1_3_36_36 ;
      VIA 32.532 23.49 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 23.473 32.577 23.507 ;
      VIA 32.532 23.49 Element_VIA34_1_2_58_52 ;
      VIA 32.532 23.49 Element_VIA23_1_3_36_36 ;
      VIA 32.532 22.95 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 22.933 32.577 22.967 ;
      VIA 32.532 22.95 Element_VIA34_1_2_58_52 ;
      VIA 32.532 22.95 Element_VIA23_1_3_36_36 ;
      VIA 32.532 22.41 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 22.393 32.577 22.427 ;
      VIA 32.532 22.41 Element_VIA34_1_2_58_52 ;
      VIA 32.532 22.41 Element_VIA23_1_3_36_36 ;
      VIA 32.532 21.87 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 21.853 32.577 21.887 ;
      VIA 32.532 21.87 Element_VIA34_1_2_58_52 ;
      VIA 32.532 21.87 Element_VIA23_1_3_36_36 ;
      VIA 32.532 21.33 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 21.313 32.577 21.347 ;
      VIA 32.532 21.33 Element_VIA34_1_2_58_52 ;
      VIA 32.532 21.33 Element_VIA23_1_3_36_36 ;
      VIA 32.532 20.79 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 20.773 32.577 20.807 ;
      VIA 32.532 20.79 Element_VIA34_1_2_58_52 ;
      VIA 32.532 20.79 Element_VIA23_1_3_36_36 ;
      VIA 32.532 20.25 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 20.233 32.577 20.267 ;
      VIA 32.532 20.25 Element_VIA34_1_2_58_52 ;
      VIA 32.532 20.25 Element_VIA23_1_3_36_36 ;
      VIA 32.532 19.71 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 19.693 32.577 19.727 ;
      VIA 32.532 19.71 Element_VIA34_1_2_58_52 ;
      VIA 32.532 19.71 Element_VIA23_1_3_36_36 ;
      VIA 32.532 19.17 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 19.153 32.577 19.187 ;
      VIA 32.532 19.17 Element_VIA34_1_2_58_52 ;
      VIA 32.532 19.17 Element_VIA23_1_3_36_36 ;
      VIA 32.532 18.63 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 18.613 32.577 18.647 ;
      VIA 32.532 18.63 Element_VIA34_1_2_58_52 ;
      VIA 32.532 18.63 Element_VIA23_1_3_36_36 ;
      VIA 32.532 18.09 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 18.073 32.577 18.107 ;
      VIA 32.532 18.09 Element_VIA34_1_2_58_52 ;
      VIA 32.532 18.09 Element_VIA23_1_3_36_36 ;
      VIA 32.532 17.55 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 17.533 32.577 17.567 ;
      VIA 32.532 17.55 Element_VIA34_1_2_58_52 ;
      VIA 32.532 17.55 Element_VIA23_1_3_36_36 ;
      VIA 32.532 17.01 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 16.993 32.577 17.027 ;
      VIA 32.532 17.01 Element_VIA34_1_2_58_52 ;
      VIA 32.532 17.01 Element_VIA23_1_3_36_36 ;
      VIA 32.532 16.47 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 16.453 32.577 16.487 ;
      VIA 32.532 16.47 Element_VIA34_1_2_58_52 ;
      VIA 32.532 16.47 Element_VIA23_1_3_36_36 ;
      VIA 32.532 15.93 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 15.913 32.577 15.947 ;
      VIA 32.532 15.93 Element_VIA34_1_2_58_52 ;
      VIA 32.532 15.93 Element_VIA23_1_3_36_36 ;
      VIA 32.532 15.39 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 15.373 32.577 15.407 ;
      VIA 32.532 15.39 Element_VIA34_1_2_58_52 ;
      VIA 32.532 15.39 Element_VIA23_1_3_36_36 ;
      VIA 32.532 14.85 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 14.833 32.577 14.867 ;
      VIA 32.532 14.85 Element_VIA34_1_2_58_52 ;
      VIA 32.532 14.85 Element_VIA23_1_3_36_36 ;
      VIA 32.532 14.31 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 14.293 32.577 14.327 ;
      VIA 32.532 14.31 Element_VIA34_1_2_58_52 ;
      VIA 32.532 14.31 Element_VIA23_1_3_36_36 ;
      VIA 32.532 13.77 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 13.753 32.577 13.787 ;
      VIA 32.532 13.77 Element_VIA34_1_2_58_52 ;
      VIA 32.532 13.77 Element_VIA23_1_3_36_36 ;
      VIA 32.532 13.23 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 13.213 32.577 13.247 ;
      VIA 32.532 13.23 Element_VIA34_1_2_58_52 ;
      VIA 32.532 13.23 Element_VIA23_1_3_36_36 ;
      VIA 32.532 12.69 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 12.673 32.577 12.707 ;
      VIA 32.532 12.69 Element_VIA34_1_2_58_52 ;
      VIA 32.532 12.69 Element_VIA23_1_3_36_36 ;
      VIA 32.532 12.15 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 12.133 32.577 12.167 ;
      VIA 32.532 12.15 Element_VIA34_1_2_58_52 ;
      VIA 32.532 12.15 Element_VIA23_1_3_36_36 ;
      VIA 32.532 11.61 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 11.593 32.577 11.627 ;
      VIA 32.532 11.61 Element_VIA34_1_2_58_52 ;
      VIA 32.532 11.61 Element_VIA23_1_3_36_36 ;
      VIA 32.532 11.07 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 11.053 32.577 11.087 ;
      VIA 32.532 11.07 Element_VIA34_1_2_58_52 ;
      VIA 32.532 11.07 Element_VIA23_1_3_36_36 ;
      VIA 32.532 10.53 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 10.513 32.577 10.547 ;
      VIA 32.532 10.53 Element_VIA34_1_2_58_52 ;
      VIA 32.532 10.53 Element_VIA23_1_3_36_36 ;
      VIA 32.532 9.99 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 9.973 32.577 10.007 ;
      VIA 32.532 9.99 Element_VIA34_1_2_58_52 ;
      VIA 32.532 9.99 Element_VIA23_1_3_36_36 ;
      VIA 32.532 9.45 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 9.433 32.577 9.467 ;
      VIA 32.532 9.45 Element_VIA34_1_2_58_52 ;
      VIA 32.532 9.45 Element_VIA23_1_3_36_36 ;
      VIA 32.532 8.91 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 8.893 32.577 8.927 ;
      VIA 32.532 8.91 Element_VIA34_1_2_58_52 ;
      VIA 32.532 8.91 Element_VIA23_1_3_36_36 ;
      VIA 32.532 8.37 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 8.353 32.577 8.387 ;
      VIA 32.532 8.37 Element_VIA34_1_2_58_52 ;
      VIA 32.532 8.37 Element_VIA23_1_3_36_36 ;
      VIA 32.532 7.83 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 7.813 32.577 7.847 ;
      VIA 32.532 7.83 Element_VIA34_1_2_58_52 ;
      VIA 32.532 7.83 Element_VIA23_1_3_36_36 ;
      VIA 32.532 7.29 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 7.273 32.577 7.307 ;
      VIA 32.532 7.29 Element_VIA34_1_2_58_52 ;
      VIA 32.532 7.29 Element_VIA23_1_3_36_36 ;
      VIA 32.532 6.75 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 6.733 32.577 6.767 ;
      VIA 32.532 6.75 Element_VIA34_1_2_58_52 ;
      VIA 32.532 6.75 Element_VIA23_1_3_36_36 ;
      VIA 32.532 6.21 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 6.193 32.577 6.227 ;
      VIA 32.532 6.21 Element_VIA34_1_2_58_52 ;
      VIA 32.532 6.21 Element_VIA23_1_3_36_36 ;
      VIA 32.532 5.67 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 5.653 32.577 5.687 ;
      VIA 32.532 5.67 Element_VIA34_1_2_58_52 ;
      VIA 32.532 5.67 Element_VIA23_1_3_36_36 ;
      VIA 32.532 5.13 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 5.113 32.577 5.147 ;
      VIA 32.532 5.13 Element_VIA34_1_2_58_52 ;
      VIA 32.532 5.13 Element_VIA23_1_3_36_36 ;
      VIA 32.532 4.59 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 4.573 32.577 4.607 ;
      VIA 32.532 4.59 Element_VIA34_1_2_58_52 ;
      VIA 32.532 4.59 Element_VIA23_1_3_36_36 ;
      VIA 32.532 4.05 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 4.033 32.577 4.067 ;
      VIA 32.532 4.05 Element_VIA34_1_2_58_52 ;
      VIA 32.532 4.05 Element_VIA23_1_3_36_36 ;
      VIA 32.532 3.51 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 3.493 32.577 3.527 ;
      VIA 32.532 3.51 Element_VIA34_1_2_58_52 ;
      VIA 32.532 3.51 Element_VIA23_1_3_36_36 ;
      VIA 32.532 2.97 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 2.953 32.577 2.987 ;
      VIA 32.532 2.97 Element_VIA34_1_2_58_52 ;
      VIA 32.532 2.97 Element_VIA23_1_3_36_36 ;
      VIA 32.532 2.43 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 2.413 32.577 2.447 ;
      VIA 32.532 2.43 Element_VIA34_1_2_58_52 ;
      VIA 32.532 2.43 Element_VIA23_1_3_36_36 ;
      VIA 32.532 1.89 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 1.873 32.577 1.907 ;
      VIA 32.532 1.89 Element_VIA34_1_2_58_52 ;
      VIA 32.532 1.89 Element_VIA23_1_3_36_36 ;
      VIA 32.532 1.35 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.487 1.333 32.577 1.367 ;
      VIA 32.532 1.35 Element_VIA34_1_2_58_52 ;
      VIA 32.532 1.35 Element_VIA23_1_3_36_36 ;
      VIA 29.556 41.85 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 41.833 29.601 41.867 ;
      VIA 29.556 41.85 Element_VIA34_1_2_58_52 ;
      VIA 29.556 41.85 Element_VIA23_1_3_36_36 ;
      VIA 29.556 41.31 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 41.293 29.601 41.327 ;
      VIA 29.556 41.31 Element_VIA34_1_2_58_52 ;
      VIA 29.556 41.31 Element_VIA23_1_3_36_36 ;
      VIA 29.556 40.77 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 40.753 29.601 40.787 ;
      VIA 29.556 40.77 Element_VIA34_1_2_58_52 ;
      VIA 29.556 40.77 Element_VIA23_1_3_36_36 ;
      VIA 29.556 40.23 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 40.213 29.601 40.247 ;
      VIA 29.556 40.23 Element_VIA34_1_2_58_52 ;
      VIA 29.556 40.23 Element_VIA23_1_3_36_36 ;
      VIA 29.556 39.69 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 39.673 29.601 39.707 ;
      VIA 29.556 39.69 Element_VIA34_1_2_58_52 ;
      VIA 29.556 39.69 Element_VIA23_1_3_36_36 ;
      VIA 29.556 39.15 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 39.133 29.601 39.167 ;
      VIA 29.556 39.15 Element_VIA34_1_2_58_52 ;
      VIA 29.556 39.15 Element_VIA23_1_3_36_36 ;
      VIA 29.556 38.61 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 38.593 29.601 38.627 ;
      VIA 29.556 38.61 Element_VIA34_1_2_58_52 ;
      VIA 29.556 38.61 Element_VIA23_1_3_36_36 ;
      VIA 29.556 38.07 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 38.053 29.601 38.087 ;
      VIA 29.556 38.07 Element_VIA34_1_2_58_52 ;
      VIA 29.556 38.07 Element_VIA23_1_3_36_36 ;
      VIA 29.556 37.53 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 37.513 29.601 37.547 ;
      VIA 29.556 37.53 Element_VIA34_1_2_58_52 ;
      VIA 29.556 37.53 Element_VIA23_1_3_36_36 ;
      VIA 29.556 36.99 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 36.973 29.601 37.007 ;
      VIA 29.556 36.99 Element_VIA34_1_2_58_52 ;
      VIA 29.556 36.99 Element_VIA23_1_3_36_36 ;
      VIA 29.556 36.45 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 36.433 29.601 36.467 ;
      VIA 29.556 36.45 Element_VIA34_1_2_58_52 ;
      VIA 29.556 36.45 Element_VIA23_1_3_36_36 ;
      VIA 29.556 35.91 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 35.893 29.601 35.927 ;
      VIA 29.556 35.91 Element_VIA34_1_2_58_52 ;
      VIA 29.556 35.91 Element_VIA23_1_3_36_36 ;
      VIA 29.556 35.37 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 35.353 29.601 35.387 ;
      VIA 29.556 35.37 Element_VIA34_1_2_58_52 ;
      VIA 29.556 35.37 Element_VIA23_1_3_36_36 ;
      VIA 29.556 34.83 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 34.813 29.601 34.847 ;
      VIA 29.556 34.83 Element_VIA34_1_2_58_52 ;
      VIA 29.556 34.83 Element_VIA23_1_3_36_36 ;
      VIA 29.556 34.29 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 34.273 29.601 34.307 ;
      VIA 29.556 34.29 Element_VIA34_1_2_58_52 ;
      VIA 29.556 34.29 Element_VIA23_1_3_36_36 ;
      VIA 29.556 33.75 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 33.733 29.601 33.767 ;
      VIA 29.556 33.75 Element_VIA34_1_2_58_52 ;
      VIA 29.556 33.75 Element_VIA23_1_3_36_36 ;
      VIA 29.556 33.21 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 33.193 29.601 33.227 ;
      VIA 29.556 33.21 Element_VIA34_1_2_58_52 ;
      VIA 29.556 33.21 Element_VIA23_1_3_36_36 ;
      VIA 29.556 32.67 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 32.653 29.601 32.687 ;
      VIA 29.556 32.67 Element_VIA34_1_2_58_52 ;
      VIA 29.556 32.67 Element_VIA23_1_3_36_36 ;
      VIA 29.556 32.13 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 32.113 29.601 32.147 ;
      VIA 29.556 32.13 Element_VIA34_1_2_58_52 ;
      VIA 29.556 32.13 Element_VIA23_1_3_36_36 ;
      VIA 29.556 31.59 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 31.573 29.601 31.607 ;
      VIA 29.556 31.59 Element_VIA34_1_2_58_52 ;
      VIA 29.556 31.59 Element_VIA23_1_3_36_36 ;
      VIA 29.556 31.05 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 31.033 29.601 31.067 ;
      VIA 29.556 31.05 Element_VIA34_1_2_58_52 ;
      VIA 29.556 31.05 Element_VIA23_1_3_36_36 ;
      VIA 29.556 30.51 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 30.493 29.601 30.527 ;
      VIA 29.556 30.51 Element_VIA34_1_2_58_52 ;
      VIA 29.556 30.51 Element_VIA23_1_3_36_36 ;
      VIA 29.556 29.97 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 29.953 29.601 29.987 ;
      VIA 29.556 29.97 Element_VIA34_1_2_58_52 ;
      VIA 29.556 29.97 Element_VIA23_1_3_36_36 ;
      VIA 29.556 29.43 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 29.413 29.601 29.447 ;
      VIA 29.556 29.43 Element_VIA34_1_2_58_52 ;
      VIA 29.556 29.43 Element_VIA23_1_3_36_36 ;
      VIA 29.556 28.89 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 28.873 29.601 28.907 ;
      VIA 29.556 28.89 Element_VIA34_1_2_58_52 ;
      VIA 29.556 28.89 Element_VIA23_1_3_36_36 ;
      VIA 29.556 28.35 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 28.333 29.601 28.367 ;
      VIA 29.556 28.35 Element_VIA34_1_2_58_52 ;
      VIA 29.556 28.35 Element_VIA23_1_3_36_36 ;
      VIA 29.556 27.81 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 27.793 29.601 27.827 ;
      VIA 29.556 27.81 Element_VIA34_1_2_58_52 ;
      VIA 29.556 27.81 Element_VIA23_1_3_36_36 ;
      VIA 29.556 27.27 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 27.253 29.601 27.287 ;
      VIA 29.556 27.27 Element_VIA34_1_2_58_52 ;
      VIA 29.556 27.27 Element_VIA23_1_3_36_36 ;
      VIA 29.556 26.73 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 26.713 29.601 26.747 ;
      VIA 29.556 26.73 Element_VIA34_1_2_58_52 ;
      VIA 29.556 26.73 Element_VIA23_1_3_36_36 ;
      VIA 29.556 26.19 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 26.173 29.601 26.207 ;
      VIA 29.556 26.19 Element_VIA34_1_2_58_52 ;
      VIA 29.556 26.19 Element_VIA23_1_3_36_36 ;
      VIA 29.556 25.65 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 25.633 29.601 25.667 ;
      VIA 29.556 25.65 Element_VIA34_1_2_58_52 ;
      VIA 29.556 25.65 Element_VIA23_1_3_36_36 ;
      VIA 29.556 25.11 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 25.093 29.601 25.127 ;
      VIA 29.556 25.11 Element_VIA34_1_2_58_52 ;
      VIA 29.556 25.11 Element_VIA23_1_3_36_36 ;
      VIA 29.556 24.57 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 24.553 29.601 24.587 ;
      VIA 29.556 24.57 Element_VIA34_1_2_58_52 ;
      VIA 29.556 24.57 Element_VIA23_1_3_36_36 ;
      VIA 29.556 24.03 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 24.013 29.601 24.047 ;
      VIA 29.556 24.03 Element_VIA34_1_2_58_52 ;
      VIA 29.556 24.03 Element_VIA23_1_3_36_36 ;
      VIA 29.556 23.49 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 23.473 29.601 23.507 ;
      VIA 29.556 23.49 Element_VIA34_1_2_58_52 ;
      VIA 29.556 23.49 Element_VIA23_1_3_36_36 ;
      VIA 29.556 22.95 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 22.933 29.601 22.967 ;
      VIA 29.556 22.95 Element_VIA34_1_2_58_52 ;
      VIA 29.556 22.95 Element_VIA23_1_3_36_36 ;
      VIA 29.556 22.41 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 22.393 29.601 22.427 ;
      VIA 29.556 22.41 Element_VIA34_1_2_58_52 ;
      VIA 29.556 22.41 Element_VIA23_1_3_36_36 ;
      VIA 29.556 21.87 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 21.853 29.601 21.887 ;
      VIA 29.556 21.87 Element_VIA34_1_2_58_52 ;
      VIA 29.556 21.87 Element_VIA23_1_3_36_36 ;
      VIA 29.556 21.33 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 21.313 29.601 21.347 ;
      VIA 29.556 21.33 Element_VIA34_1_2_58_52 ;
      VIA 29.556 21.33 Element_VIA23_1_3_36_36 ;
      VIA 29.556 20.79 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 20.773 29.601 20.807 ;
      VIA 29.556 20.79 Element_VIA34_1_2_58_52 ;
      VIA 29.556 20.79 Element_VIA23_1_3_36_36 ;
      VIA 29.556 20.25 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 20.233 29.601 20.267 ;
      VIA 29.556 20.25 Element_VIA34_1_2_58_52 ;
      VIA 29.556 20.25 Element_VIA23_1_3_36_36 ;
      VIA 29.556 19.71 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 19.693 29.601 19.727 ;
      VIA 29.556 19.71 Element_VIA34_1_2_58_52 ;
      VIA 29.556 19.71 Element_VIA23_1_3_36_36 ;
      VIA 29.556 19.17 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 19.153 29.601 19.187 ;
      VIA 29.556 19.17 Element_VIA34_1_2_58_52 ;
      VIA 29.556 19.17 Element_VIA23_1_3_36_36 ;
      VIA 29.556 18.63 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 18.613 29.601 18.647 ;
      VIA 29.556 18.63 Element_VIA34_1_2_58_52 ;
      VIA 29.556 18.63 Element_VIA23_1_3_36_36 ;
      VIA 29.556 18.09 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 18.073 29.601 18.107 ;
      VIA 29.556 18.09 Element_VIA34_1_2_58_52 ;
      VIA 29.556 18.09 Element_VIA23_1_3_36_36 ;
      VIA 29.556 17.55 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 17.533 29.601 17.567 ;
      VIA 29.556 17.55 Element_VIA34_1_2_58_52 ;
      VIA 29.556 17.55 Element_VIA23_1_3_36_36 ;
      VIA 29.556 17.01 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 16.993 29.601 17.027 ;
      VIA 29.556 17.01 Element_VIA34_1_2_58_52 ;
      VIA 29.556 17.01 Element_VIA23_1_3_36_36 ;
      VIA 29.556 16.47 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 16.453 29.601 16.487 ;
      VIA 29.556 16.47 Element_VIA34_1_2_58_52 ;
      VIA 29.556 16.47 Element_VIA23_1_3_36_36 ;
      VIA 29.556 15.93 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 15.913 29.601 15.947 ;
      VIA 29.556 15.93 Element_VIA34_1_2_58_52 ;
      VIA 29.556 15.93 Element_VIA23_1_3_36_36 ;
      VIA 29.556 15.39 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 15.373 29.601 15.407 ;
      VIA 29.556 15.39 Element_VIA34_1_2_58_52 ;
      VIA 29.556 15.39 Element_VIA23_1_3_36_36 ;
      VIA 29.556 14.85 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 14.833 29.601 14.867 ;
      VIA 29.556 14.85 Element_VIA34_1_2_58_52 ;
      VIA 29.556 14.85 Element_VIA23_1_3_36_36 ;
      VIA 29.556 14.31 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 14.293 29.601 14.327 ;
      VIA 29.556 14.31 Element_VIA34_1_2_58_52 ;
      VIA 29.556 14.31 Element_VIA23_1_3_36_36 ;
      VIA 29.556 13.77 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 13.753 29.601 13.787 ;
      VIA 29.556 13.77 Element_VIA34_1_2_58_52 ;
      VIA 29.556 13.77 Element_VIA23_1_3_36_36 ;
      VIA 29.556 13.23 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 13.213 29.601 13.247 ;
      VIA 29.556 13.23 Element_VIA34_1_2_58_52 ;
      VIA 29.556 13.23 Element_VIA23_1_3_36_36 ;
      VIA 29.556 12.69 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 12.673 29.601 12.707 ;
      VIA 29.556 12.69 Element_VIA34_1_2_58_52 ;
      VIA 29.556 12.69 Element_VIA23_1_3_36_36 ;
      VIA 29.556 12.15 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 12.133 29.601 12.167 ;
      VIA 29.556 12.15 Element_VIA34_1_2_58_52 ;
      VIA 29.556 12.15 Element_VIA23_1_3_36_36 ;
      VIA 29.556 11.61 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 11.593 29.601 11.627 ;
      VIA 29.556 11.61 Element_VIA34_1_2_58_52 ;
      VIA 29.556 11.61 Element_VIA23_1_3_36_36 ;
      VIA 29.556 11.07 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 11.053 29.601 11.087 ;
      VIA 29.556 11.07 Element_VIA34_1_2_58_52 ;
      VIA 29.556 11.07 Element_VIA23_1_3_36_36 ;
      VIA 29.556 10.53 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 10.513 29.601 10.547 ;
      VIA 29.556 10.53 Element_VIA34_1_2_58_52 ;
      VIA 29.556 10.53 Element_VIA23_1_3_36_36 ;
      VIA 29.556 9.99 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 9.973 29.601 10.007 ;
      VIA 29.556 9.99 Element_VIA34_1_2_58_52 ;
      VIA 29.556 9.99 Element_VIA23_1_3_36_36 ;
      VIA 29.556 9.45 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 9.433 29.601 9.467 ;
      VIA 29.556 9.45 Element_VIA34_1_2_58_52 ;
      VIA 29.556 9.45 Element_VIA23_1_3_36_36 ;
      VIA 29.556 8.91 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 8.893 29.601 8.927 ;
      VIA 29.556 8.91 Element_VIA34_1_2_58_52 ;
      VIA 29.556 8.91 Element_VIA23_1_3_36_36 ;
      VIA 29.556 8.37 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 8.353 29.601 8.387 ;
      VIA 29.556 8.37 Element_VIA34_1_2_58_52 ;
      VIA 29.556 8.37 Element_VIA23_1_3_36_36 ;
      VIA 29.556 7.83 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 7.813 29.601 7.847 ;
      VIA 29.556 7.83 Element_VIA34_1_2_58_52 ;
      VIA 29.556 7.83 Element_VIA23_1_3_36_36 ;
      VIA 29.556 7.29 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 7.273 29.601 7.307 ;
      VIA 29.556 7.29 Element_VIA34_1_2_58_52 ;
      VIA 29.556 7.29 Element_VIA23_1_3_36_36 ;
      VIA 29.556 6.75 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 6.733 29.601 6.767 ;
      VIA 29.556 6.75 Element_VIA34_1_2_58_52 ;
      VIA 29.556 6.75 Element_VIA23_1_3_36_36 ;
      VIA 29.556 6.21 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 6.193 29.601 6.227 ;
      VIA 29.556 6.21 Element_VIA34_1_2_58_52 ;
      VIA 29.556 6.21 Element_VIA23_1_3_36_36 ;
      VIA 29.556 5.67 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 5.653 29.601 5.687 ;
      VIA 29.556 5.67 Element_VIA34_1_2_58_52 ;
      VIA 29.556 5.67 Element_VIA23_1_3_36_36 ;
      VIA 29.556 5.13 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 5.113 29.601 5.147 ;
      VIA 29.556 5.13 Element_VIA34_1_2_58_52 ;
      VIA 29.556 5.13 Element_VIA23_1_3_36_36 ;
      VIA 29.556 4.59 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 4.573 29.601 4.607 ;
      VIA 29.556 4.59 Element_VIA34_1_2_58_52 ;
      VIA 29.556 4.59 Element_VIA23_1_3_36_36 ;
      VIA 29.556 4.05 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 4.033 29.601 4.067 ;
      VIA 29.556 4.05 Element_VIA34_1_2_58_52 ;
      VIA 29.556 4.05 Element_VIA23_1_3_36_36 ;
      VIA 29.556 3.51 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 3.493 29.601 3.527 ;
      VIA 29.556 3.51 Element_VIA34_1_2_58_52 ;
      VIA 29.556 3.51 Element_VIA23_1_3_36_36 ;
      VIA 29.556 2.97 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 2.953 29.601 2.987 ;
      VIA 29.556 2.97 Element_VIA34_1_2_58_52 ;
      VIA 29.556 2.97 Element_VIA23_1_3_36_36 ;
      VIA 29.556 2.43 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 2.413 29.601 2.447 ;
      VIA 29.556 2.43 Element_VIA34_1_2_58_52 ;
      VIA 29.556 2.43 Element_VIA23_1_3_36_36 ;
      VIA 29.556 1.89 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 1.873 29.601 1.907 ;
      VIA 29.556 1.89 Element_VIA34_1_2_58_52 ;
      VIA 29.556 1.89 Element_VIA23_1_3_36_36 ;
      VIA 29.556 1.35 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.511 1.333 29.601 1.367 ;
      VIA 29.556 1.35 Element_VIA34_1_2_58_52 ;
      VIA 29.556 1.35 Element_VIA23_1_3_36_36 ;
      VIA 26.58 41.85 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 41.833 26.625 41.867 ;
      VIA 26.58 41.85 Element_VIA34_1_2_58_52 ;
      VIA 26.58 41.85 Element_VIA23_1_3_36_36 ;
      VIA 26.58 41.31 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 41.293 26.625 41.327 ;
      VIA 26.58 41.31 Element_VIA34_1_2_58_52 ;
      VIA 26.58 41.31 Element_VIA23_1_3_36_36 ;
      VIA 26.58 40.77 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 40.753 26.625 40.787 ;
      VIA 26.58 40.77 Element_VIA34_1_2_58_52 ;
      VIA 26.58 40.77 Element_VIA23_1_3_36_36 ;
      VIA 26.58 40.23 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 40.213 26.625 40.247 ;
      VIA 26.58 40.23 Element_VIA34_1_2_58_52 ;
      VIA 26.58 40.23 Element_VIA23_1_3_36_36 ;
      VIA 26.58 39.69 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 39.673 26.625 39.707 ;
      VIA 26.58 39.69 Element_VIA34_1_2_58_52 ;
      VIA 26.58 39.69 Element_VIA23_1_3_36_36 ;
      VIA 26.58 39.15 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 39.133 26.625 39.167 ;
      VIA 26.58 39.15 Element_VIA34_1_2_58_52 ;
      VIA 26.58 39.15 Element_VIA23_1_3_36_36 ;
      VIA 26.58 38.61 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 38.593 26.625 38.627 ;
      VIA 26.58 38.61 Element_VIA34_1_2_58_52 ;
      VIA 26.58 38.61 Element_VIA23_1_3_36_36 ;
      VIA 26.58 38.07 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 38.053 26.625 38.087 ;
      VIA 26.58 38.07 Element_VIA34_1_2_58_52 ;
      VIA 26.58 38.07 Element_VIA23_1_3_36_36 ;
      VIA 26.58 37.53 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 37.513 26.625 37.547 ;
      VIA 26.58 37.53 Element_VIA34_1_2_58_52 ;
      VIA 26.58 37.53 Element_VIA23_1_3_36_36 ;
      VIA 26.58 36.99 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 36.973 26.625 37.007 ;
      VIA 26.58 36.99 Element_VIA34_1_2_58_52 ;
      VIA 26.58 36.99 Element_VIA23_1_3_36_36 ;
      VIA 26.58 36.45 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 36.433 26.625 36.467 ;
      VIA 26.58 36.45 Element_VIA34_1_2_58_52 ;
      VIA 26.58 36.45 Element_VIA23_1_3_36_36 ;
      VIA 26.58 35.91 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 35.893 26.625 35.927 ;
      VIA 26.58 35.91 Element_VIA34_1_2_58_52 ;
      VIA 26.58 35.91 Element_VIA23_1_3_36_36 ;
      VIA 26.58 35.37 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 35.353 26.625 35.387 ;
      VIA 26.58 35.37 Element_VIA34_1_2_58_52 ;
      VIA 26.58 35.37 Element_VIA23_1_3_36_36 ;
      VIA 26.58 34.83 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 34.813 26.625 34.847 ;
      VIA 26.58 34.83 Element_VIA34_1_2_58_52 ;
      VIA 26.58 34.83 Element_VIA23_1_3_36_36 ;
      VIA 26.58 34.29 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 34.273 26.625 34.307 ;
      VIA 26.58 34.29 Element_VIA34_1_2_58_52 ;
      VIA 26.58 34.29 Element_VIA23_1_3_36_36 ;
      VIA 26.58 33.75 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 33.733 26.625 33.767 ;
      VIA 26.58 33.75 Element_VIA34_1_2_58_52 ;
      VIA 26.58 33.75 Element_VIA23_1_3_36_36 ;
      VIA 26.58 33.21 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 33.193 26.625 33.227 ;
      VIA 26.58 33.21 Element_VIA34_1_2_58_52 ;
      VIA 26.58 33.21 Element_VIA23_1_3_36_36 ;
      VIA 26.58 32.67 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 32.653 26.625 32.687 ;
      VIA 26.58 32.67 Element_VIA34_1_2_58_52 ;
      VIA 26.58 32.67 Element_VIA23_1_3_36_36 ;
      VIA 26.58 32.13 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 32.113 26.625 32.147 ;
      VIA 26.58 32.13 Element_VIA34_1_2_58_52 ;
      VIA 26.58 32.13 Element_VIA23_1_3_36_36 ;
      VIA 26.58 31.59 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 31.573 26.625 31.607 ;
      VIA 26.58 31.59 Element_VIA34_1_2_58_52 ;
      VIA 26.58 31.59 Element_VIA23_1_3_36_36 ;
      VIA 26.58 31.05 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 31.033 26.625 31.067 ;
      VIA 26.58 31.05 Element_VIA34_1_2_58_52 ;
      VIA 26.58 31.05 Element_VIA23_1_3_36_36 ;
      VIA 26.58 30.51 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 30.493 26.625 30.527 ;
      VIA 26.58 30.51 Element_VIA34_1_2_58_52 ;
      VIA 26.58 30.51 Element_VIA23_1_3_36_36 ;
      VIA 26.58 29.97 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 29.953 26.625 29.987 ;
      VIA 26.58 29.97 Element_VIA34_1_2_58_52 ;
      VIA 26.58 29.97 Element_VIA23_1_3_36_36 ;
      VIA 26.58 29.43 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 29.413 26.625 29.447 ;
      VIA 26.58 29.43 Element_VIA34_1_2_58_52 ;
      VIA 26.58 29.43 Element_VIA23_1_3_36_36 ;
      VIA 26.58 28.89 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 28.873 26.625 28.907 ;
      VIA 26.58 28.89 Element_VIA34_1_2_58_52 ;
      VIA 26.58 28.89 Element_VIA23_1_3_36_36 ;
      VIA 26.58 28.35 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 28.333 26.625 28.367 ;
      VIA 26.58 28.35 Element_VIA34_1_2_58_52 ;
      VIA 26.58 28.35 Element_VIA23_1_3_36_36 ;
      VIA 26.58 27.81 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 27.793 26.625 27.827 ;
      VIA 26.58 27.81 Element_VIA34_1_2_58_52 ;
      VIA 26.58 27.81 Element_VIA23_1_3_36_36 ;
      VIA 26.58 27.27 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 27.253 26.625 27.287 ;
      VIA 26.58 27.27 Element_VIA34_1_2_58_52 ;
      VIA 26.58 27.27 Element_VIA23_1_3_36_36 ;
      VIA 26.58 26.73 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 26.713 26.625 26.747 ;
      VIA 26.58 26.73 Element_VIA34_1_2_58_52 ;
      VIA 26.58 26.73 Element_VIA23_1_3_36_36 ;
      VIA 26.58 26.19 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 26.173 26.625 26.207 ;
      VIA 26.58 26.19 Element_VIA34_1_2_58_52 ;
      VIA 26.58 26.19 Element_VIA23_1_3_36_36 ;
      VIA 26.58 25.65 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 25.633 26.625 25.667 ;
      VIA 26.58 25.65 Element_VIA34_1_2_58_52 ;
      VIA 26.58 25.65 Element_VIA23_1_3_36_36 ;
      VIA 26.58 25.11 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 25.093 26.625 25.127 ;
      VIA 26.58 25.11 Element_VIA34_1_2_58_52 ;
      VIA 26.58 25.11 Element_VIA23_1_3_36_36 ;
      VIA 26.58 24.57 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 24.553 26.625 24.587 ;
      VIA 26.58 24.57 Element_VIA34_1_2_58_52 ;
      VIA 26.58 24.57 Element_VIA23_1_3_36_36 ;
      VIA 26.58 24.03 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 24.013 26.625 24.047 ;
      VIA 26.58 24.03 Element_VIA34_1_2_58_52 ;
      VIA 26.58 24.03 Element_VIA23_1_3_36_36 ;
      VIA 26.58 23.49 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 23.473 26.625 23.507 ;
      VIA 26.58 23.49 Element_VIA34_1_2_58_52 ;
      VIA 26.58 23.49 Element_VIA23_1_3_36_36 ;
      VIA 26.58 22.95 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 22.933 26.625 22.967 ;
      VIA 26.58 22.95 Element_VIA34_1_2_58_52 ;
      VIA 26.58 22.95 Element_VIA23_1_3_36_36 ;
      VIA 26.58 22.41 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 22.393 26.625 22.427 ;
      VIA 26.58 22.41 Element_VIA34_1_2_58_52 ;
      VIA 26.58 22.41 Element_VIA23_1_3_36_36 ;
      VIA 26.58 21.87 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 21.853 26.625 21.887 ;
      VIA 26.58 21.87 Element_VIA34_1_2_58_52 ;
      VIA 26.58 21.87 Element_VIA23_1_3_36_36 ;
      VIA 26.58 21.33 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 21.313 26.625 21.347 ;
      VIA 26.58 21.33 Element_VIA34_1_2_58_52 ;
      VIA 26.58 21.33 Element_VIA23_1_3_36_36 ;
      VIA 26.58 20.79 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 20.773 26.625 20.807 ;
      VIA 26.58 20.79 Element_VIA34_1_2_58_52 ;
      VIA 26.58 20.79 Element_VIA23_1_3_36_36 ;
      VIA 26.58 20.25 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 20.233 26.625 20.267 ;
      VIA 26.58 20.25 Element_VIA34_1_2_58_52 ;
      VIA 26.58 20.25 Element_VIA23_1_3_36_36 ;
      VIA 26.58 19.71 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 19.693 26.625 19.727 ;
      VIA 26.58 19.71 Element_VIA34_1_2_58_52 ;
      VIA 26.58 19.71 Element_VIA23_1_3_36_36 ;
      VIA 26.58 19.17 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 19.153 26.625 19.187 ;
      VIA 26.58 19.17 Element_VIA34_1_2_58_52 ;
      VIA 26.58 19.17 Element_VIA23_1_3_36_36 ;
      VIA 26.58 18.63 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 18.613 26.625 18.647 ;
      VIA 26.58 18.63 Element_VIA34_1_2_58_52 ;
      VIA 26.58 18.63 Element_VIA23_1_3_36_36 ;
      VIA 26.58 18.09 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 18.073 26.625 18.107 ;
      VIA 26.58 18.09 Element_VIA34_1_2_58_52 ;
      VIA 26.58 18.09 Element_VIA23_1_3_36_36 ;
      VIA 26.58 17.55 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 17.533 26.625 17.567 ;
      VIA 26.58 17.55 Element_VIA34_1_2_58_52 ;
      VIA 26.58 17.55 Element_VIA23_1_3_36_36 ;
      VIA 26.58 17.01 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 16.993 26.625 17.027 ;
      VIA 26.58 17.01 Element_VIA34_1_2_58_52 ;
      VIA 26.58 17.01 Element_VIA23_1_3_36_36 ;
      VIA 26.58 16.47 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 16.453 26.625 16.487 ;
      VIA 26.58 16.47 Element_VIA34_1_2_58_52 ;
      VIA 26.58 16.47 Element_VIA23_1_3_36_36 ;
      VIA 26.58 15.93 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 15.913 26.625 15.947 ;
      VIA 26.58 15.93 Element_VIA34_1_2_58_52 ;
      VIA 26.58 15.93 Element_VIA23_1_3_36_36 ;
      VIA 26.58 15.39 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 15.373 26.625 15.407 ;
      VIA 26.58 15.39 Element_VIA34_1_2_58_52 ;
      VIA 26.58 15.39 Element_VIA23_1_3_36_36 ;
      VIA 26.58 14.85 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 14.833 26.625 14.867 ;
      VIA 26.58 14.85 Element_VIA34_1_2_58_52 ;
      VIA 26.58 14.85 Element_VIA23_1_3_36_36 ;
      VIA 26.58 14.31 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 14.293 26.625 14.327 ;
      VIA 26.58 14.31 Element_VIA34_1_2_58_52 ;
      VIA 26.58 14.31 Element_VIA23_1_3_36_36 ;
      VIA 26.58 13.77 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 13.753 26.625 13.787 ;
      VIA 26.58 13.77 Element_VIA34_1_2_58_52 ;
      VIA 26.58 13.77 Element_VIA23_1_3_36_36 ;
      VIA 26.58 13.23 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 13.213 26.625 13.247 ;
      VIA 26.58 13.23 Element_VIA34_1_2_58_52 ;
      VIA 26.58 13.23 Element_VIA23_1_3_36_36 ;
      VIA 26.58 12.69 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 12.673 26.625 12.707 ;
      VIA 26.58 12.69 Element_VIA34_1_2_58_52 ;
      VIA 26.58 12.69 Element_VIA23_1_3_36_36 ;
      VIA 26.58 12.15 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 12.133 26.625 12.167 ;
      VIA 26.58 12.15 Element_VIA34_1_2_58_52 ;
      VIA 26.58 12.15 Element_VIA23_1_3_36_36 ;
      VIA 26.58 11.61 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 11.593 26.625 11.627 ;
      VIA 26.58 11.61 Element_VIA34_1_2_58_52 ;
      VIA 26.58 11.61 Element_VIA23_1_3_36_36 ;
      VIA 26.58 11.07 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 11.053 26.625 11.087 ;
      VIA 26.58 11.07 Element_VIA34_1_2_58_52 ;
      VIA 26.58 11.07 Element_VIA23_1_3_36_36 ;
      VIA 26.58 10.53 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 10.513 26.625 10.547 ;
      VIA 26.58 10.53 Element_VIA34_1_2_58_52 ;
      VIA 26.58 10.53 Element_VIA23_1_3_36_36 ;
      VIA 26.58 9.99 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 9.973 26.625 10.007 ;
      VIA 26.58 9.99 Element_VIA34_1_2_58_52 ;
      VIA 26.58 9.99 Element_VIA23_1_3_36_36 ;
      VIA 26.58 9.45 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 9.433 26.625 9.467 ;
      VIA 26.58 9.45 Element_VIA34_1_2_58_52 ;
      VIA 26.58 9.45 Element_VIA23_1_3_36_36 ;
      VIA 26.58 8.91 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 8.893 26.625 8.927 ;
      VIA 26.58 8.91 Element_VIA34_1_2_58_52 ;
      VIA 26.58 8.91 Element_VIA23_1_3_36_36 ;
      VIA 26.58 8.37 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 8.353 26.625 8.387 ;
      VIA 26.58 8.37 Element_VIA34_1_2_58_52 ;
      VIA 26.58 8.37 Element_VIA23_1_3_36_36 ;
      VIA 26.58 7.83 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 7.813 26.625 7.847 ;
      VIA 26.58 7.83 Element_VIA34_1_2_58_52 ;
      VIA 26.58 7.83 Element_VIA23_1_3_36_36 ;
      VIA 26.58 7.29 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 7.273 26.625 7.307 ;
      VIA 26.58 7.29 Element_VIA34_1_2_58_52 ;
      VIA 26.58 7.29 Element_VIA23_1_3_36_36 ;
      VIA 26.58 6.75 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 6.733 26.625 6.767 ;
      VIA 26.58 6.75 Element_VIA34_1_2_58_52 ;
      VIA 26.58 6.75 Element_VIA23_1_3_36_36 ;
      VIA 26.58 6.21 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 6.193 26.625 6.227 ;
      VIA 26.58 6.21 Element_VIA34_1_2_58_52 ;
      VIA 26.58 6.21 Element_VIA23_1_3_36_36 ;
      VIA 26.58 5.67 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 5.653 26.625 5.687 ;
      VIA 26.58 5.67 Element_VIA34_1_2_58_52 ;
      VIA 26.58 5.67 Element_VIA23_1_3_36_36 ;
      VIA 26.58 5.13 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 5.113 26.625 5.147 ;
      VIA 26.58 5.13 Element_VIA34_1_2_58_52 ;
      VIA 26.58 5.13 Element_VIA23_1_3_36_36 ;
      VIA 26.58 4.59 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 4.573 26.625 4.607 ;
      VIA 26.58 4.59 Element_VIA34_1_2_58_52 ;
      VIA 26.58 4.59 Element_VIA23_1_3_36_36 ;
      VIA 26.58 4.05 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 4.033 26.625 4.067 ;
      VIA 26.58 4.05 Element_VIA34_1_2_58_52 ;
      VIA 26.58 4.05 Element_VIA23_1_3_36_36 ;
      VIA 26.58 3.51 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 3.493 26.625 3.527 ;
      VIA 26.58 3.51 Element_VIA34_1_2_58_52 ;
      VIA 26.58 3.51 Element_VIA23_1_3_36_36 ;
      VIA 26.58 2.97 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 2.953 26.625 2.987 ;
      VIA 26.58 2.97 Element_VIA34_1_2_58_52 ;
      VIA 26.58 2.97 Element_VIA23_1_3_36_36 ;
      VIA 26.58 2.43 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 2.413 26.625 2.447 ;
      VIA 26.58 2.43 Element_VIA34_1_2_58_52 ;
      VIA 26.58 2.43 Element_VIA23_1_3_36_36 ;
      VIA 26.58 1.89 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 1.873 26.625 1.907 ;
      VIA 26.58 1.89 Element_VIA34_1_2_58_52 ;
      VIA 26.58 1.89 Element_VIA23_1_3_36_36 ;
      VIA 26.58 1.35 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.535 1.333 26.625 1.367 ;
      VIA 26.58 1.35 Element_VIA34_1_2_58_52 ;
      VIA 26.58 1.35 Element_VIA23_1_3_36_36 ;
      VIA 23.604 41.85 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 41.833 23.649 41.867 ;
      VIA 23.604 41.85 Element_VIA34_1_2_58_52 ;
      VIA 23.604 41.85 Element_VIA23_1_3_36_36 ;
      VIA 23.604 41.31 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 41.293 23.649 41.327 ;
      VIA 23.604 41.31 Element_VIA34_1_2_58_52 ;
      VIA 23.604 41.31 Element_VIA23_1_3_36_36 ;
      VIA 23.604 40.77 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 40.753 23.649 40.787 ;
      VIA 23.604 40.77 Element_VIA34_1_2_58_52 ;
      VIA 23.604 40.77 Element_VIA23_1_3_36_36 ;
      VIA 23.604 40.23 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 40.213 23.649 40.247 ;
      VIA 23.604 40.23 Element_VIA34_1_2_58_52 ;
      VIA 23.604 40.23 Element_VIA23_1_3_36_36 ;
      VIA 23.604 39.69 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 39.673 23.649 39.707 ;
      VIA 23.604 39.69 Element_VIA34_1_2_58_52 ;
      VIA 23.604 39.69 Element_VIA23_1_3_36_36 ;
      VIA 23.604 39.15 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 39.133 23.649 39.167 ;
      VIA 23.604 39.15 Element_VIA34_1_2_58_52 ;
      VIA 23.604 39.15 Element_VIA23_1_3_36_36 ;
      VIA 23.604 38.61 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 38.593 23.649 38.627 ;
      VIA 23.604 38.61 Element_VIA34_1_2_58_52 ;
      VIA 23.604 38.61 Element_VIA23_1_3_36_36 ;
      VIA 23.604 38.07 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 38.053 23.649 38.087 ;
      VIA 23.604 38.07 Element_VIA34_1_2_58_52 ;
      VIA 23.604 38.07 Element_VIA23_1_3_36_36 ;
      VIA 23.604 37.53 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 37.513 23.649 37.547 ;
      VIA 23.604 37.53 Element_VIA34_1_2_58_52 ;
      VIA 23.604 37.53 Element_VIA23_1_3_36_36 ;
      VIA 23.604 36.99 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 36.973 23.649 37.007 ;
      VIA 23.604 36.99 Element_VIA34_1_2_58_52 ;
      VIA 23.604 36.99 Element_VIA23_1_3_36_36 ;
      VIA 23.604 36.45 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 36.433 23.649 36.467 ;
      VIA 23.604 36.45 Element_VIA34_1_2_58_52 ;
      VIA 23.604 36.45 Element_VIA23_1_3_36_36 ;
      VIA 23.604 35.91 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 35.893 23.649 35.927 ;
      VIA 23.604 35.91 Element_VIA34_1_2_58_52 ;
      VIA 23.604 35.91 Element_VIA23_1_3_36_36 ;
      VIA 23.604 35.37 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 35.353 23.649 35.387 ;
      VIA 23.604 35.37 Element_VIA34_1_2_58_52 ;
      VIA 23.604 35.37 Element_VIA23_1_3_36_36 ;
      VIA 23.604 34.83 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 34.813 23.649 34.847 ;
      VIA 23.604 34.83 Element_VIA34_1_2_58_52 ;
      VIA 23.604 34.83 Element_VIA23_1_3_36_36 ;
      VIA 23.604 34.29 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 34.273 23.649 34.307 ;
      VIA 23.604 34.29 Element_VIA34_1_2_58_52 ;
      VIA 23.604 34.29 Element_VIA23_1_3_36_36 ;
      VIA 23.604 33.75 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 33.733 23.649 33.767 ;
      VIA 23.604 33.75 Element_VIA34_1_2_58_52 ;
      VIA 23.604 33.75 Element_VIA23_1_3_36_36 ;
      VIA 23.604 33.21 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 33.193 23.649 33.227 ;
      VIA 23.604 33.21 Element_VIA34_1_2_58_52 ;
      VIA 23.604 33.21 Element_VIA23_1_3_36_36 ;
      VIA 23.604 32.67 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 32.653 23.649 32.687 ;
      VIA 23.604 32.67 Element_VIA34_1_2_58_52 ;
      VIA 23.604 32.67 Element_VIA23_1_3_36_36 ;
      VIA 23.604 32.13 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 32.113 23.649 32.147 ;
      VIA 23.604 32.13 Element_VIA34_1_2_58_52 ;
      VIA 23.604 32.13 Element_VIA23_1_3_36_36 ;
      VIA 23.604 31.59 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 31.573 23.649 31.607 ;
      VIA 23.604 31.59 Element_VIA34_1_2_58_52 ;
      VIA 23.604 31.59 Element_VIA23_1_3_36_36 ;
      VIA 23.604 31.05 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 31.033 23.649 31.067 ;
      VIA 23.604 31.05 Element_VIA34_1_2_58_52 ;
      VIA 23.604 31.05 Element_VIA23_1_3_36_36 ;
      VIA 23.604 30.51 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 30.493 23.649 30.527 ;
      VIA 23.604 30.51 Element_VIA34_1_2_58_52 ;
      VIA 23.604 30.51 Element_VIA23_1_3_36_36 ;
      VIA 23.604 29.97 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 29.953 23.649 29.987 ;
      VIA 23.604 29.97 Element_VIA34_1_2_58_52 ;
      VIA 23.604 29.97 Element_VIA23_1_3_36_36 ;
      VIA 23.604 29.43 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 29.413 23.649 29.447 ;
      VIA 23.604 29.43 Element_VIA34_1_2_58_52 ;
      VIA 23.604 29.43 Element_VIA23_1_3_36_36 ;
      VIA 23.604 28.89 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 28.873 23.649 28.907 ;
      VIA 23.604 28.89 Element_VIA34_1_2_58_52 ;
      VIA 23.604 28.89 Element_VIA23_1_3_36_36 ;
      VIA 23.604 28.35 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 28.333 23.649 28.367 ;
      VIA 23.604 28.35 Element_VIA34_1_2_58_52 ;
      VIA 23.604 28.35 Element_VIA23_1_3_36_36 ;
      VIA 23.604 27.81 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 27.793 23.649 27.827 ;
      VIA 23.604 27.81 Element_VIA34_1_2_58_52 ;
      VIA 23.604 27.81 Element_VIA23_1_3_36_36 ;
      VIA 23.604 27.27 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 27.253 23.649 27.287 ;
      VIA 23.604 27.27 Element_VIA34_1_2_58_52 ;
      VIA 23.604 27.27 Element_VIA23_1_3_36_36 ;
      VIA 23.604 26.73 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 26.713 23.649 26.747 ;
      VIA 23.604 26.73 Element_VIA34_1_2_58_52 ;
      VIA 23.604 26.73 Element_VIA23_1_3_36_36 ;
      VIA 23.604 26.19 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 26.173 23.649 26.207 ;
      VIA 23.604 26.19 Element_VIA34_1_2_58_52 ;
      VIA 23.604 26.19 Element_VIA23_1_3_36_36 ;
      VIA 23.604 25.65 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 25.633 23.649 25.667 ;
      VIA 23.604 25.65 Element_VIA34_1_2_58_52 ;
      VIA 23.604 25.65 Element_VIA23_1_3_36_36 ;
      VIA 23.604 25.11 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 25.093 23.649 25.127 ;
      VIA 23.604 25.11 Element_VIA34_1_2_58_52 ;
      VIA 23.604 25.11 Element_VIA23_1_3_36_36 ;
      VIA 23.604 24.57 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 24.553 23.649 24.587 ;
      VIA 23.604 24.57 Element_VIA34_1_2_58_52 ;
      VIA 23.604 24.57 Element_VIA23_1_3_36_36 ;
      VIA 23.604 24.03 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 24.013 23.649 24.047 ;
      VIA 23.604 24.03 Element_VIA34_1_2_58_52 ;
      VIA 23.604 24.03 Element_VIA23_1_3_36_36 ;
      VIA 23.604 23.49 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 23.473 23.649 23.507 ;
      VIA 23.604 23.49 Element_VIA34_1_2_58_52 ;
      VIA 23.604 23.49 Element_VIA23_1_3_36_36 ;
      VIA 23.604 22.95 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 22.933 23.649 22.967 ;
      VIA 23.604 22.95 Element_VIA34_1_2_58_52 ;
      VIA 23.604 22.95 Element_VIA23_1_3_36_36 ;
      VIA 23.604 22.41 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 22.393 23.649 22.427 ;
      VIA 23.604 22.41 Element_VIA34_1_2_58_52 ;
      VIA 23.604 22.41 Element_VIA23_1_3_36_36 ;
      VIA 23.604 21.87 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 21.853 23.649 21.887 ;
      VIA 23.604 21.87 Element_VIA34_1_2_58_52 ;
      VIA 23.604 21.87 Element_VIA23_1_3_36_36 ;
      VIA 23.604 21.33 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 21.313 23.649 21.347 ;
      VIA 23.604 21.33 Element_VIA34_1_2_58_52 ;
      VIA 23.604 21.33 Element_VIA23_1_3_36_36 ;
      VIA 23.604 20.79 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 20.773 23.649 20.807 ;
      VIA 23.604 20.79 Element_VIA34_1_2_58_52 ;
      VIA 23.604 20.79 Element_VIA23_1_3_36_36 ;
      VIA 23.604 20.25 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 20.233 23.649 20.267 ;
      VIA 23.604 20.25 Element_VIA34_1_2_58_52 ;
      VIA 23.604 20.25 Element_VIA23_1_3_36_36 ;
      VIA 23.604 19.71 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 19.693 23.649 19.727 ;
      VIA 23.604 19.71 Element_VIA34_1_2_58_52 ;
      VIA 23.604 19.71 Element_VIA23_1_3_36_36 ;
      VIA 23.604 19.17 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 19.153 23.649 19.187 ;
      VIA 23.604 19.17 Element_VIA34_1_2_58_52 ;
      VIA 23.604 19.17 Element_VIA23_1_3_36_36 ;
      VIA 23.604 18.63 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 18.613 23.649 18.647 ;
      VIA 23.604 18.63 Element_VIA34_1_2_58_52 ;
      VIA 23.604 18.63 Element_VIA23_1_3_36_36 ;
      VIA 23.604 18.09 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 18.073 23.649 18.107 ;
      VIA 23.604 18.09 Element_VIA34_1_2_58_52 ;
      VIA 23.604 18.09 Element_VIA23_1_3_36_36 ;
      VIA 23.604 17.55 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 17.533 23.649 17.567 ;
      VIA 23.604 17.55 Element_VIA34_1_2_58_52 ;
      VIA 23.604 17.55 Element_VIA23_1_3_36_36 ;
      VIA 23.604 17.01 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 16.993 23.649 17.027 ;
      VIA 23.604 17.01 Element_VIA34_1_2_58_52 ;
      VIA 23.604 17.01 Element_VIA23_1_3_36_36 ;
      VIA 23.604 16.47 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 16.453 23.649 16.487 ;
      VIA 23.604 16.47 Element_VIA34_1_2_58_52 ;
      VIA 23.604 16.47 Element_VIA23_1_3_36_36 ;
      VIA 23.604 15.93 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 15.913 23.649 15.947 ;
      VIA 23.604 15.93 Element_VIA34_1_2_58_52 ;
      VIA 23.604 15.93 Element_VIA23_1_3_36_36 ;
      VIA 23.604 15.39 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 15.373 23.649 15.407 ;
      VIA 23.604 15.39 Element_VIA34_1_2_58_52 ;
      VIA 23.604 15.39 Element_VIA23_1_3_36_36 ;
      VIA 23.604 14.85 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 14.833 23.649 14.867 ;
      VIA 23.604 14.85 Element_VIA34_1_2_58_52 ;
      VIA 23.604 14.85 Element_VIA23_1_3_36_36 ;
      VIA 23.604 14.31 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 14.293 23.649 14.327 ;
      VIA 23.604 14.31 Element_VIA34_1_2_58_52 ;
      VIA 23.604 14.31 Element_VIA23_1_3_36_36 ;
      VIA 23.604 13.77 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 13.753 23.649 13.787 ;
      VIA 23.604 13.77 Element_VIA34_1_2_58_52 ;
      VIA 23.604 13.77 Element_VIA23_1_3_36_36 ;
      VIA 23.604 13.23 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 13.213 23.649 13.247 ;
      VIA 23.604 13.23 Element_VIA34_1_2_58_52 ;
      VIA 23.604 13.23 Element_VIA23_1_3_36_36 ;
      VIA 23.604 12.69 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 12.673 23.649 12.707 ;
      VIA 23.604 12.69 Element_VIA34_1_2_58_52 ;
      VIA 23.604 12.69 Element_VIA23_1_3_36_36 ;
      VIA 23.604 12.15 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 12.133 23.649 12.167 ;
      VIA 23.604 12.15 Element_VIA34_1_2_58_52 ;
      VIA 23.604 12.15 Element_VIA23_1_3_36_36 ;
      VIA 23.604 11.61 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 11.593 23.649 11.627 ;
      VIA 23.604 11.61 Element_VIA34_1_2_58_52 ;
      VIA 23.604 11.61 Element_VIA23_1_3_36_36 ;
      VIA 23.604 11.07 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 11.053 23.649 11.087 ;
      VIA 23.604 11.07 Element_VIA34_1_2_58_52 ;
      VIA 23.604 11.07 Element_VIA23_1_3_36_36 ;
      VIA 23.604 10.53 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 10.513 23.649 10.547 ;
      VIA 23.604 10.53 Element_VIA34_1_2_58_52 ;
      VIA 23.604 10.53 Element_VIA23_1_3_36_36 ;
      VIA 23.604 9.99 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 9.973 23.649 10.007 ;
      VIA 23.604 9.99 Element_VIA34_1_2_58_52 ;
      VIA 23.604 9.99 Element_VIA23_1_3_36_36 ;
      VIA 23.604 9.45 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 9.433 23.649 9.467 ;
      VIA 23.604 9.45 Element_VIA34_1_2_58_52 ;
      VIA 23.604 9.45 Element_VIA23_1_3_36_36 ;
      VIA 23.604 8.91 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 8.893 23.649 8.927 ;
      VIA 23.604 8.91 Element_VIA34_1_2_58_52 ;
      VIA 23.604 8.91 Element_VIA23_1_3_36_36 ;
      VIA 23.604 8.37 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 8.353 23.649 8.387 ;
      VIA 23.604 8.37 Element_VIA34_1_2_58_52 ;
      VIA 23.604 8.37 Element_VIA23_1_3_36_36 ;
      VIA 23.604 7.83 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 7.813 23.649 7.847 ;
      VIA 23.604 7.83 Element_VIA34_1_2_58_52 ;
      VIA 23.604 7.83 Element_VIA23_1_3_36_36 ;
      VIA 23.604 7.29 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 7.273 23.649 7.307 ;
      VIA 23.604 7.29 Element_VIA34_1_2_58_52 ;
      VIA 23.604 7.29 Element_VIA23_1_3_36_36 ;
      VIA 23.604 6.75 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 6.733 23.649 6.767 ;
      VIA 23.604 6.75 Element_VIA34_1_2_58_52 ;
      VIA 23.604 6.75 Element_VIA23_1_3_36_36 ;
      VIA 23.604 6.21 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 6.193 23.649 6.227 ;
      VIA 23.604 6.21 Element_VIA34_1_2_58_52 ;
      VIA 23.604 6.21 Element_VIA23_1_3_36_36 ;
      VIA 23.604 5.67 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 5.653 23.649 5.687 ;
      VIA 23.604 5.67 Element_VIA34_1_2_58_52 ;
      VIA 23.604 5.67 Element_VIA23_1_3_36_36 ;
      VIA 23.604 5.13 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 5.113 23.649 5.147 ;
      VIA 23.604 5.13 Element_VIA34_1_2_58_52 ;
      VIA 23.604 5.13 Element_VIA23_1_3_36_36 ;
      VIA 23.604 4.59 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 4.573 23.649 4.607 ;
      VIA 23.604 4.59 Element_VIA34_1_2_58_52 ;
      VIA 23.604 4.59 Element_VIA23_1_3_36_36 ;
      VIA 23.604 4.05 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 4.033 23.649 4.067 ;
      VIA 23.604 4.05 Element_VIA34_1_2_58_52 ;
      VIA 23.604 4.05 Element_VIA23_1_3_36_36 ;
      VIA 23.604 3.51 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 3.493 23.649 3.527 ;
      VIA 23.604 3.51 Element_VIA34_1_2_58_52 ;
      VIA 23.604 3.51 Element_VIA23_1_3_36_36 ;
      VIA 23.604 2.97 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 2.953 23.649 2.987 ;
      VIA 23.604 2.97 Element_VIA34_1_2_58_52 ;
      VIA 23.604 2.97 Element_VIA23_1_3_36_36 ;
      VIA 23.604 2.43 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 2.413 23.649 2.447 ;
      VIA 23.604 2.43 Element_VIA34_1_2_58_52 ;
      VIA 23.604 2.43 Element_VIA23_1_3_36_36 ;
      VIA 23.604 1.89 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 1.873 23.649 1.907 ;
      VIA 23.604 1.89 Element_VIA34_1_2_58_52 ;
      VIA 23.604 1.89 Element_VIA23_1_3_36_36 ;
      VIA 23.604 1.35 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.559 1.333 23.649 1.367 ;
      VIA 23.604 1.35 Element_VIA34_1_2_58_52 ;
      VIA 23.604 1.35 Element_VIA23_1_3_36_36 ;
      VIA 20.628 41.85 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 41.833 20.673 41.867 ;
      VIA 20.628 41.85 Element_VIA34_1_2_58_52 ;
      VIA 20.628 41.85 Element_VIA23_1_3_36_36 ;
      VIA 20.628 41.31 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 41.293 20.673 41.327 ;
      VIA 20.628 41.31 Element_VIA34_1_2_58_52 ;
      VIA 20.628 41.31 Element_VIA23_1_3_36_36 ;
      VIA 20.628 40.77 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 40.753 20.673 40.787 ;
      VIA 20.628 40.77 Element_VIA34_1_2_58_52 ;
      VIA 20.628 40.77 Element_VIA23_1_3_36_36 ;
      VIA 20.628 40.23 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 40.213 20.673 40.247 ;
      VIA 20.628 40.23 Element_VIA34_1_2_58_52 ;
      VIA 20.628 40.23 Element_VIA23_1_3_36_36 ;
      VIA 20.628 39.69 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 39.673 20.673 39.707 ;
      VIA 20.628 39.69 Element_VIA34_1_2_58_52 ;
      VIA 20.628 39.69 Element_VIA23_1_3_36_36 ;
      VIA 20.628 39.15 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 39.133 20.673 39.167 ;
      VIA 20.628 39.15 Element_VIA34_1_2_58_52 ;
      VIA 20.628 39.15 Element_VIA23_1_3_36_36 ;
      VIA 20.628 38.61 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 38.593 20.673 38.627 ;
      VIA 20.628 38.61 Element_VIA34_1_2_58_52 ;
      VIA 20.628 38.61 Element_VIA23_1_3_36_36 ;
      VIA 20.628 38.07 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 38.053 20.673 38.087 ;
      VIA 20.628 38.07 Element_VIA34_1_2_58_52 ;
      VIA 20.628 38.07 Element_VIA23_1_3_36_36 ;
      VIA 20.628 37.53 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 37.513 20.673 37.547 ;
      VIA 20.628 37.53 Element_VIA34_1_2_58_52 ;
      VIA 20.628 37.53 Element_VIA23_1_3_36_36 ;
      VIA 20.628 36.99 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 36.973 20.673 37.007 ;
      VIA 20.628 36.99 Element_VIA34_1_2_58_52 ;
      VIA 20.628 36.99 Element_VIA23_1_3_36_36 ;
      VIA 20.628 36.45 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 36.433 20.673 36.467 ;
      VIA 20.628 36.45 Element_VIA34_1_2_58_52 ;
      VIA 20.628 36.45 Element_VIA23_1_3_36_36 ;
      VIA 20.628 35.91 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 35.893 20.673 35.927 ;
      VIA 20.628 35.91 Element_VIA34_1_2_58_52 ;
      VIA 20.628 35.91 Element_VIA23_1_3_36_36 ;
      VIA 20.628 35.37 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 35.353 20.673 35.387 ;
      VIA 20.628 35.37 Element_VIA34_1_2_58_52 ;
      VIA 20.628 35.37 Element_VIA23_1_3_36_36 ;
      VIA 20.628 34.83 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 34.813 20.673 34.847 ;
      VIA 20.628 34.83 Element_VIA34_1_2_58_52 ;
      VIA 20.628 34.83 Element_VIA23_1_3_36_36 ;
      VIA 20.628 34.29 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 34.273 20.673 34.307 ;
      VIA 20.628 34.29 Element_VIA34_1_2_58_52 ;
      VIA 20.628 34.29 Element_VIA23_1_3_36_36 ;
      VIA 20.628 33.75 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 33.733 20.673 33.767 ;
      VIA 20.628 33.75 Element_VIA34_1_2_58_52 ;
      VIA 20.628 33.75 Element_VIA23_1_3_36_36 ;
      VIA 20.628 33.21 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 33.193 20.673 33.227 ;
      VIA 20.628 33.21 Element_VIA34_1_2_58_52 ;
      VIA 20.628 33.21 Element_VIA23_1_3_36_36 ;
      VIA 20.628 32.67 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 32.653 20.673 32.687 ;
      VIA 20.628 32.67 Element_VIA34_1_2_58_52 ;
      VIA 20.628 32.67 Element_VIA23_1_3_36_36 ;
      VIA 20.628 32.13 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 32.113 20.673 32.147 ;
      VIA 20.628 32.13 Element_VIA34_1_2_58_52 ;
      VIA 20.628 32.13 Element_VIA23_1_3_36_36 ;
      VIA 20.628 31.59 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 31.573 20.673 31.607 ;
      VIA 20.628 31.59 Element_VIA34_1_2_58_52 ;
      VIA 20.628 31.59 Element_VIA23_1_3_36_36 ;
      VIA 20.628 31.05 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 31.033 20.673 31.067 ;
      VIA 20.628 31.05 Element_VIA34_1_2_58_52 ;
      VIA 20.628 31.05 Element_VIA23_1_3_36_36 ;
      VIA 20.628 30.51 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 30.493 20.673 30.527 ;
      VIA 20.628 30.51 Element_VIA34_1_2_58_52 ;
      VIA 20.628 30.51 Element_VIA23_1_3_36_36 ;
      VIA 20.628 29.97 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 29.953 20.673 29.987 ;
      VIA 20.628 29.97 Element_VIA34_1_2_58_52 ;
      VIA 20.628 29.97 Element_VIA23_1_3_36_36 ;
      VIA 20.628 29.43 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 29.413 20.673 29.447 ;
      VIA 20.628 29.43 Element_VIA34_1_2_58_52 ;
      VIA 20.628 29.43 Element_VIA23_1_3_36_36 ;
      VIA 20.628 28.89 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 28.873 20.673 28.907 ;
      VIA 20.628 28.89 Element_VIA34_1_2_58_52 ;
      VIA 20.628 28.89 Element_VIA23_1_3_36_36 ;
      VIA 20.628 28.35 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 28.333 20.673 28.367 ;
      VIA 20.628 28.35 Element_VIA34_1_2_58_52 ;
      VIA 20.628 28.35 Element_VIA23_1_3_36_36 ;
      VIA 20.628 27.81 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 27.793 20.673 27.827 ;
      VIA 20.628 27.81 Element_VIA34_1_2_58_52 ;
      VIA 20.628 27.81 Element_VIA23_1_3_36_36 ;
      VIA 20.628 27.27 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 27.253 20.673 27.287 ;
      VIA 20.628 27.27 Element_VIA34_1_2_58_52 ;
      VIA 20.628 27.27 Element_VIA23_1_3_36_36 ;
      VIA 20.628 26.73 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 26.713 20.673 26.747 ;
      VIA 20.628 26.73 Element_VIA34_1_2_58_52 ;
      VIA 20.628 26.73 Element_VIA23_1_3_36_36 ;
      VIA 20.628 26.19 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 26.173 20.673 26.207 ;
      VIA 20.628 26.19 Element_VIA34_1_2_58_52 ;
      VIA 20.628 26.19 Element_VIA23_1_3_36_36 ;
      VIA 20.628 25.65 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 25.633 20.673 25.667 ;
      VIA 20.628 25.65 Element_VIA34_1_2_58_52 ;
      VIA 20.628 25.65 Element_VIA23_1_3_36_36 ;
      VIA 20.628 25.11 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 25.093 20.673 25.127 ;
      VIA 20.628 25.11 Element_VIA34_1_2_58_52 ;
      VIA 20.628 25.11 Element_VIA23_1_3_36_36 ;
      VIA 20.628 24.57 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 24.553 20.673 24.587 ;
      VIA 20.628 24.57 Element_VIA34_1_2_58_52 ;
      VIA 20.628 24.57 Element_VIA23_1_3_36_36 ;
      VIA 20.628 24.03 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 24.013 20.673 24.047 ;
      VIA 20.628 24.03 Element_VIA34_1_2_58_52 ;
      VIA 20.628 24.03 Element_VIA23_1_3_36_36 ;
      VIA 20.628 23.49 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 23.473 20.673 23.507 ;
      VIA 20.628 23.49 Element_VIA34_1_2_58_52 ;
      VIA 20.628 23.49 Element_VIA23_1_3_36_36 ;
      VIA 20.628 22.95 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 22.933 20.673 22.967 ;
      VIA 20.628 22.95 Element_VIA34_1_2_58_52 ;
      VIA 20.628 22.95 Element_VIA23_1_3_36_36 ;
      VIA 20.628 22.41 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 22.393 20.673 22.427 ;
      VIA 20.628 22.41 Element_VIA34_1_2_58_52 ;
      VIA 20.628 22.41 Element_VIA23_1_3_36_36 ;
      VIA 20.628 21.87 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 21.853 20.673 21.887 ;
      VIA 20.628 21.87 Element_VIA34_1_2_58_52 ;
      VIA 20.628 21.87 Element_VIA23_1_3_36_36 ;
      VIA 20.628 21.33 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 21.313 20.673 21.347 ;
      VIA 20.628 21.33 Element_VIA34_1_2_58_52 ;
      VIA 20.628 21.33 Element_VIA23_1_3_36_36 ;
      VIA 20.628 20.79 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 20.773 20.673 20.807 ;
      VIA 20.628 20.79 Element_VIA34_1_2_58_52 ;
      VIA 20.628 20.79 Element_VIA23_1_3_36_36 ;
      VIA 20.628 20.25 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 20.233 20.673 20.267 ;
      VIA 20.628 20.25 Element_VIA34_1_2_58_52 ;
      VIA 20.628 20.25 Element_VIA23_1_3_36_36 ;
      VIA 20.628 19.71 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 19.693 20.673 19.727 ;
      VIA 20.628 19.71 Element_VIA34_1_2_58_52 ;
      VIA 20.628 19.71 Element_VIA23_1_3_36_36 ;
      VIA 20.628 19.17 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 19.153 20.673 19.187 ;
      VIA 20.628 19.17 Element_VIA34_1_2_58_52 ;
      VIA 20.628 19.17 Element_VIA23_1_3_36_36 ;
      VIA 20.628 18.63 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 18.613 20.673 18.647 ;
      VIA 20.628 18.63 Element_VIA34_1_2_58_52 ;
      VIA 20.628 18.63 Element_VIA23_1_3_36_36 ;
      VIA 20.628 18.09 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 18.073 20.673 18.107 ;
      VIA 20.628 18.09 Element_VIA34_1_2_58_52 ;
      VIA 20.628 18.09 Element_VIA23_1_3_36_36 ;
      VIA 20.628 17.55 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 17.533 20.673 17.567 ;
      VIA 20.628 17.55 Element_VIA34_1_2_58_52 ;
      VIA 20.628 17.55 Element_VIA23_1_3_36_36 ;
      VIA 20.628 17.01 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 16.993 20.673 17.027 ;
      VIA 20.628 17.01 Element_VIA34_1_2_58_52 ;
      VIA 20.628 17.01 Element_VIA23_1_3_36_36 ;
      VIA 20.628 16.47 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 16.453 20.673 16.487 ;
      VIA 20.628 16.47 Element_VIA34_1_2_58_52 ;
      VIA 20.628 16.47 Element_VIA23_1_3_36_36 ;
      VIA 20.628 15.93 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 15.913 20.673 15.947 ;
      VIA 20.628 15.93 Element_VIA34_1_2_58_52 ;
      VIA 20.628 15.93 Element_VIA23_1_3_36_36 ;
      VIA 20.628 15.39 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 15.373 20.673 15.407 ;
      VIA 20.628 15.39 Element_VIA34_1_2_58_52 ;
      VIA 20.628 15.39 Element_VIA23_1_3_36_36 ;
      VIA 20.628 14.85 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 14.833 20.673 14.867 ;
      VIA 20.628 14.85 Element_VIA34_1_2_58_52 ;
      VIA 20.628 14.85 Element_VIA23_1_3_36_36 ;
      VIA 20.628 14.31 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 14.293 20.673 14.327 ;
      VIA 20.628 14.31 Element_VIA34_1_2_58_52 ;
      VIA 20.628 14.31 Element_VIA23_1_3_36_36 ;
      VIA 20.628 13.77 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 13.753 20.673 13.787 ;
      VIA 20.628 13.77 Element_VIA34_1_2_58_52 ;
      VIA 20.628 13.77 Element_VIA23_1_3_36_36 ;
      VIA 20.628 13.23 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 13.213 20.673 13.247 ;
      VIA 20.628 13.23 Element_VIA34_1_2_58_52 ;
      VIA 20.628 13.23 Element_VIA23_1_3_36_36 ;
      VIA 20.628 12.69 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 12.673 20.673 12.707 ;
      VIA 20.628 12.69 Element_VIA34_1_2_58_52 ;
      VIA 20.628 12.69 Element_VIA23_1_3_36_36 ;
      VIA 20.628 12.15 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 12.133 20.673 12.167 ;
      VIA 20.628 12.15 Element_VIA34_1_2_58_52 ;
      VIA 20.628 12.15 Element_VIA23_1_3_36_36 ;
      VIA 20.628 11.61 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 11.593 20.673 11.627 ;
      VIA 20.628 11.61 Element_VIA34_1_2_58_52 ;
      VIA 20.628 11.61 Element_VIA23_1_3_36_36 ;
      VIA 20.628 11.07 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 11.053 20.673 11.087 ;
      VIA 20.628 11.07 Element_VIA34_1_2_58_52 ;
      VIA 20.628 11.07 Element_VIA23_1_3_36_36 ;
      VIA 20.628 10.53 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 10.513 20.673 10.547 ;
      VIA 20.628 10.53 Element_VIA34_1_2_58_52 ;
      VIA 20.628 10.53 Element_VIA23_1_3_36_36 ;
      VIA 20.628 9.99 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 9.973 20.673 10.007 ;
      VIA 20.628 9.99 Element_VIA34_1_2_58_52 ;
      VIA 20.628 9.99 Element_VIA23_1_3_36_36 ;
      VIA 20.628 9.45 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 9.433 20.673 9.467 ;
      VIA 20.628 9.45 Element_VIA34_1_2_58_52 ;
      VIA 20.628 9.45 Element_VIA23_1_3_36_36 ;
      VIA 20.628 8.91 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 8.893 20.673 8.927 ;
      VIA 20.628 8.91 Element_VIA34_1_2_58_52 ;
      VIA 20.628 8.91 Element_VIA23_1_3_36_36 ;
      VIA 20.628 8.37 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 8.353 20.673 8.387 ;
      VIA 20.628 8.37 Element_VIA34_1_2_58_52 ;
      VIA 20.628 8.37 Element_VIA23_1_3_36_36 ;
      VIA 20.628 7.83 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 7.813 20.673 7.847 ;
      VIA 20.628 7.83 Element_VIA34_1_2_58_52 ;
      VIA 20.628 7.83 Element_VIA23_1_3_36_36 ;
      VIA 20.628 7.29 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 7.273 20.673 7.307 ;
      VIA 20.628 7.29 Element_VIA34_1_2_58_52 ;
      VIA 20.628 7.29 Element_VIA23_1_3_36_36 ;
      VIA 20.628 6.75 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 6.733 20.673 6.767 ;
      VIA 20.628 6.75 Element_VIA34_1_2_58_52 ;
      VIA 20.628 6.75 Element_VIA23_1_3_36_36 ;
      VIA 20.628 6.21 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 6.193 20.673 6.227 ;
      VIA 20.628 6.21 Element_VIA34_1_2_58_52 ;
      VIA 20.628 6.21 Element_VIA23_1_3_36_36 ;
      VIA 20.628 5.67 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 5.653 20.673 5.687 ;
      VIA 20.628 5.67 Element_VIA34_1_2_58_52 ;
      VIA 20.628 5.67 Element_VIA23_1_3_36_36 ;
      VIA 20.628 5.13 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 5.113 20.673 5.147 ;
      VIA 20.628 5.13 Element_VIA34_1_2_58_52 ;
      VIA 20.628 5.13 Element_VIA23_1_3_36_36 ;
      VIA 20.628 4.59 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 4.573 20.673 4.607 ;
      VIA 20.628 4.59 Element_VIA34_1_2_58_52 ;
      VIA 20.628 4.59 Element_VIA23_1_3_36_36 ;
      VIA 20.628 4.05 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 4.033 20.673 4.067 ;
      VIA 20.628 4.05 Element_VIA34_1_2_58_52 ;
      VIA 20.628 4.05 Element_VIA23_1_3_36_36 ;
      VIA 20.628 3.51 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 3.493 20.673 3.527 ;
      VIA 20.628 3.51 Element_VIA34_1_2_58_52 ;
      VIA 20.628 3.51 Element_VIA23_1_3_36_36 ;
      VIA 20.628 2.97 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 2.953 20.673 2.987 ;
      VIA 20.628 2.97 Element_VIA34_1_2_58_52 ;
      VIA 20.628 2.97 Element_VIA23_1_3_36_36 ;
      VIA 20.628 2.43 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 2.413 20.673 2.447 ;
      VIA 20.628 2.43 Element_VIA34_1_2_58_52 ;
      VIA 20.628 2.43 Element_VIA23_1_3_36_36 ;
      VIA 20.628 1.89 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 1.873 20.673 1.907 ;
      VIA 20.628 1.89 Element_VIA34_1_2_58_52 ;
      VIA 20.628 1.89 Element_VIA23_1_3_36_36 ;
      VIA 20.628 1.35 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.583 1.333 20.673 1.367 ;
      VIA 20.628 1.35 Element_VIA34_1_2_58_52 ;
      VIA 20.628 1.35 Element_VIA23_1_3_36_36 ;
      VIA 17.652 41.85 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 41.833 17.697 41.867 ;
      VIA 17.652 41.85 Element_VIA34_1_2_58_52 ;
      VIA 17.652 41.85 Element_VIA23_1_3_36_36 ;
      VIA 17.652 41.31 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 41.293 17.697 41.327 ;
      VIA 17.652 41.31 Element_VIA34_1_2_58_52 ;
      VIA 17.652 41.31 Element_VIA23_1_3_36_36 ;
      VIA 17.652 40.77 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 40.753 17.697 40.787 ;
      VIA 17.652 40.77 Element_VIA34_1_2_58_52 ;
      VIA 17.652 40.77 Element_VIA23_1_3_36_36 ;
      VIA 17.652 40.23 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 40.213 17.697 40.247 ;
      VIA 17.652 40.23 Element_VIA34_1_2_58_52 ;
      VIA 17.652 40.23 Element_VIA23_1_3_36_36 ;
      VIA 17.652 39.69 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 39.673 17.697 39.707 ;
      VIA 17.652 39.69 Element_VIA34_1_2_58_52 ;
      VIA 17.652 39.69 Element_VIA23_1_3_36_36 ;
      VIA 17.652 39.15 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 39.133 17.697 39.167 ;
      VIA 17.652 39.15 Element_VIA34_1_2_58_52 ;
      VIA 17.652 39.15 Element_VIA23_1_3_36_36 ;
      VIA 17.652 38.61 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 38.593 17.697 38.627 ;
      VIA 17.652 38.61 Element_VIA34_1_2_58_52 ;
      VIA 17.652 38.61 Element_VIA23_1_3_36_36 ;
      VIA 17.652 38.07 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 38.053 17.697 38.087 ;
      VIA 17.652 38.07 Element_VIA34_1_2_58_52 ;
      VIA 17.652 38.07 Element_VIA23_1_3_36_36 ;
      VIA 17.652 37.53 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 37.513 17.697 37.547 ;
      VIA 17.652 37.53 Element_VIA34_1_2_58_52 ;
      VIA 17.652 37.53 Element_VIA23_1_3_36_36 ;
      VIA 17.652 36.99 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 36.973 17.697 37.007 ;
      VIA 17.652 36.99 Element_VIA34_1_2_58_52 ;
      VIA 17.652 36.99 Element_VIA23_1_3_36_36 ;
      VIA 17.652 36.45 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 36.433 17.697 36.467 ;
      VIA 17.652 36.45 Element_VIA34_1_2_58_52 ;
      VIA 17.652 36.45 Element_VIA23_1_3_36_36 ;
      VIA 17.652 35.91 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 35.893 17.697 35.927 ;
      VIA 17.652 35.91 Element_VIA34_1_2_58_52 ;
      VIA 17.652 35.91 Element_VIA23_1_3_36_36 ;
      VIA 17.652 35.37 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 35.353 17.697 35.387 ;
      VIA 17.652 35.37 Element_VIA34_1_2_58_52 ;
      VIA 17.652 35.37 Element_VIA23_1_3_36_36 ;
      VIA 17.652 34.83 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 34.813 17.697 34.847 ;
      VIA 17.652 34.83 Element_VIA34_1_2_58_52 ;
      VIA 17.652 34.83 Element_VIA23_1_3_36_36 ;
      VIA 17.652 34.29 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 34.273 17.697 34.307 ;
      VIA 17.652 34.29 Element_VIA34_1_2_58_52 ;
      VIA 17.652 34.29 Element_VIA23_1_3_36_36 ;
      VIA 17.652 33.75 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 33.733 17.697 33.767 ;
      VIA 17.652 33.75 Element_VIA34_1_2_58_52 ;
      VIA 17.652 33.75 Element_VIA23_1_3_36_36 ;
      VIA 17.652 33.21 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 33.193 17.697 33.227 ;
      VIA 17.652 33.21 Element_VIA34_1_2_58_52 ;
      VIA 17.652 33.21 Element_VIA23_1_3_36_36 ;
      VIA 17.652 32.67 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 32.653 17.697 32.687 ;
      VIA 17.652 32.67 Element_VIA34_1_2_58_52 ;
      VIA 17.652 32.67 Element_VIA23_1_3_36_36 ;
      VIA 17.652 32.13 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 32.113 17.697 32.147 ;
      VIA 17.652 32.13 Element_VIA34_1_2_58_52 ;
      VIA 17.652 32.13 Element_VIA23_1_3_36_36 ;
      VIA 17.652 31.59 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 31.573 17.697 31.607 ;
      VIA 17.652 31.59 Element_VIA34_1_2_58_52 ;
      VIA 17.652 31.59 Element_VIA23_1_3_36_36 ;
      VIA 17.652 31.05 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 31.033 17.697 31.067 ;
      VIA 17.652 31.05 Element_VIA34_1_2_58_52 ;
      VIA 17.652 31.05 Element_VIA23_1_3_36_36 ;
      VIA 17.652 30.51 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 30.493 17.697 30.527 ;
      VIA 17.652 30.51 Element_VIA34_1_2_58_52 ;
      VIA 17.652 30.51 Element_VIA23_1_3_36_36 ;
      VIA 17.652 29.97 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 29.953 17.697 29.987 ;
      VIA 17.652 29.97 Element_VIA34_1_2_58_52 ;
      VIA 17.652 29.97 Element_VIA23_1_3_36_36 ;
      VIA 17.652 29.43 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 29.413 17.697 29.447 ;
      VIA 17.652 29.43 Element_VIA34_1_2_58_52 ;
      VIA 17.652 29.43 Element_VIA23_1_3_36_36 ;
      VIA 17.652 28.89 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 28.873 17.697 28.907 ;
      VIA 17.652 28.89 Element_VIA34_1_2_58_52 ;
      VIA 17.652 28.89 Element_VIA23_1_3_36_36 ;
      VIA 17.652 28.35 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 28.333 17.697 28.367 ;
      VIA 17.652 28.35 Element_VIA34_1_2_58_52 ;
      VIA 17.652 28.35 Element_VIA23_1_3_36_36 ;
      VIA 17.652 27.81 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 27.793 17.697 27.827 ;
      VIA 17.652 27.81 Element_VIA34_1_2_58_52 ;
      VIA 17.652 27.81 Element_VIA23_1_3_36_36 ;
      VIA 17.652 27.27 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 27.253 17.697 27.287 ;
      VIA 17.652 27.27 Element_VIA34_1_2_58_52 ;
      VIA 17.652 27.27 Element_VIA23_1_3_36_36 ;
      VIA 17.652 26.73 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 26.713 17.697 26.747 ;
      VIA 17.652 26.73 Element_VIA34_1_2_58_52 ;
      VIA 17.652 26.73 Element_VIA23_1_3_36_36 ;
      VIA 17.652 26.19 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 26.173 17.697 26.207 ;
      VIA 17.652 26.19 Element_VIA34_1_2_58_52 ;
      VIA 17.652 26.19 Element_VIA23_1_3_36_36 ;
      VIA 17.652 25.65 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 25.633 17.697 25.667 ;
      VIA 17.652 25.65 Element_VIA34_1_2_58_52 ;
      VIA 17.652 25.65 Element_VIA23_1_3_36_36 ;
      VIA 17.652 25.11 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 25.093 17.697 25.127 ;
      VIA 17.652 25.11 Element_VIA34_1_2_58_52 ;
      VIA 17.652 25.11 Element_VIA23_1_3_36_36 ;
      VIA 17.652 24.57 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 24.553 17.697 24.587 ;
      VIA 17.652 24.57 Element_VIA34_1_2_58_52 ;
      VIA 17.652 24.57 Element_VIA23_1_3_36_36 ;
      VIA 17.652 24.03 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 24.013 17.697 24.047 ;
      VIA 17.652 24.03 Element_VIA34_1_2_58_52 ;
      VIA 17.652 24.03 Element_VIA23_1_3_36_36 ;
      VIA 17.652 23.49 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 23.473 17.697 23.507 ;
      VIA 17.652 23.49 Element_VIA34_1_2_58_52 ;
      VIA 17.652 23.49 Element_VIA23_1_3_36_36 ;
      VIA 17.652 22.95 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 22.933 17.697 22.967 ;
      VIA 17.652 22.95 Element_VIA34_1_2_58_52 ;
      VIA 17.652 22.95 Element_VIA23_1_3_36_36 ;
      VIA 17.652 22.41 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 22.393 17.697 22.427 ;
      VIA 17.652 22.41 Element_VIA34_1_2_58_52 ;
      VIA 17.652 22.41 Element_VIA23_1_3_36_36 ;
      VIA 17.652 21.87 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 21.853 17.697 21.887 ;
      VIA 17.652 21.87 Element_VIA34_1_2_58_52 ;
      VIA 17.652 21.87 Element_VIA23_1_3_36_36 ;
      VIA 17.652 21.33 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 21.313 17.697 21.347 ;
      VIA 17.652 21.33 Element_VIA34_1_2_58_52 ;
      VIA 17.652 21.33 Element_VIA23_1_3_36_36 ;
      VIA 17.652 20.79 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 20.773 17.697 20.807 ;
      VIA 17.652 20.79 Element_VIA34_1_2_58_52 ;
      VIA 17.652 20.79 Element_VIA23_1_3_36_36 ;
      VIA 17.652 20.25 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 20.233 17.697 20.267 ;
      VIA 17.652 20.25 Element_VIA34_1_2_58_52 ;
      VIA 17.652 20.25 Element_VIA23_1_3_36_36 ;
      VIA 17.652 19.71 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 19.693 17.697 19.727 ;
      VIA 17.652 19.71 Element_VIA34_1_2_58_52 ;
      VIA 17.652 19.71 Element_VIA23_1_3_36_36 ;
      VIA 17.652 19.17 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 19.153 17.697 19.187 ;
      VIA 17.652 19.17 Element_VIA34_1_2_58_52 ;
      VIA 17.652 19.17 Element_VIA23_1_3_36_36 ;
      VIA 17.652 18.63 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 18.613 17.697 18.647 ;
      VIA 17.652 18.63 Element_VIA34_1_2_58_52 ;
      VIA 17.652 18.63 Element_VIA23_1_3_36_36 ;
      VIA 17.652 18.09 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 18.073 17.697 18.107 ;
      VIA 17.652 18.09 Element_VIA34_1_2_58_52 ;
      VIA 17.652 18.09 Element_VIA23_1_3_36_36 ;
      VIA 17.652 17.55 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 17.533 17.697 17.567 ;
      VIA 17.652 17.55 Element_VIA34_1_2_58_52 ;
      VIA 17.652 17.55 Element_VIA23_1_3_36_36 ;
      VIA 17.652 17.01 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 16.993 17.697 17.027 ;
      VIA 17.652 17.01 Element_VIA34_1_2_58_52 ;
      VIA 17.652 17.01 Element_VIA23_1_3_36_36 ;
      VIA 17.652 16.47 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 16.453 17.697 16.487 ;
      VIA 17.652 16.47 Element_VIA34_1_2_58_52 ;
      VIA 17.652 16.47 Element_VIA23_1_3_36_36 ;
      VIA 17.652 15.93 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 15.913 17.697 15.947 ;
      VIA 17.652 15.93 Element_VIA34_1_2_58_52 ;
      VIA 17.652 15.93 Element_VIA23_1_3_36_36 ;
      VIA 17.652 15.39 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 15.373 17.697 15.407 ;
      VIA 17.652 15.39 Element_VIA34_1_2_58_52 ;
      VIA 17.652 15.39 Element_VIA23_1_3_36_36 ;
      VIA 17.652 14.85 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 14.833 17.697 14.867 ;
      VIA 17.652 14.85 Element_VIA34_1_2_58_52 ;
      VIA 17.652 14.85 Element_VIA23_1_3_36_36 ;
      VIA 17.652 14.31 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 14.293 17.697 14.327 ;
      VIA 17.652 14.31 Element_VIA34_1_2_58_52 ;
      VIA 17.652 14.31 Element_VIA23_1_3_36_36 ;
      VIA 17.652 13.77 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 13.753 17.697 13.787 ;
      VIA 17.652 13.77 Element_VIA34_1_2_58_52 ;
      VIA 17.652 13.77 Element_VIA23_1_3_36_36 ;
      VIA 17.652 13.23 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 13.213 17.697 13.247 ;
      VIA 17.652 13.23 Element_VIA34_1_2_58_52 ;
      VIA 17.652 13.23 Element_VIA23_1_3_36_36 ;
      VIA 17.652 12.69 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 12.673 17.697 12.707 ;
      VIA 17.652 12.69 Element_VIA34_1_2_58_52 ;
      VIA 17.652 12.69 Element_VIA23_1_3_36_36 ;
      VIA 17.652 12.15 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 12.133 17.697 12.167 ;
      VIA 17.652 12.15 Element_VIA34_1_2_58_52 ;
      VIA 17.652 12.15 Element_VIA23_1_3_36_36 ;
      VIA 17.652 11.61 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 11.593 17.697 11.627 ;
      VIA 17.652 11.61 Element_VIA34_1_2_58_52 ;
      VIA 17.652 11.61 Element_VIA23_1_3_36_36 ;
      VIA 17.652 11.07 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 11.053 17.697 11.087 ;
      VIA 17.652 11.07 Element_VIA34_1_2_58_52 ;
      VIA 17.652 11.07 Element_VIA23_1_3_36_36 ;
      VIA 17.652 10.53 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 10.513 17.697 10.547 ;
      VIA 17.652 10.53 Element_VIA34_1_2_58_52 ;
      VIA 17.652 10.53 Element_VIA23_1_3_36_36 ;
      VIA 17.652 9.99 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 9.973 17.697 10.007 ;
      VIA 17.652 9.99 Element_VIA34_1_2_58_52 ;
      VIA 17.652 9.99 Element_VIA23_1_3_36_36 ;
      VIA 17.652 9.45 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 9.433 17.697 9.467 ;
      VIA 17.652 9.45 Element_VIA34_1_2_58_52 ;
      VIA 17.652 9.45 Element_VIA23_1_3_36_36 ;
      VIA 17.652 8.91 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 8.893 17.697 8.927 ;
      VIA 17.652 8.91 Element_VIA34_1_2_58_52 ;
      VIA 17.652 8.91 Element_VIA23_1_3_36_36 ;
      VIA 17.652 8.37 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 8.353 17.697 8.387 ;
      VIA 17.652 8.37 Element_VIA34_1_2_58_52 ;
      VIA 17.652 8.37 Element_VIA23_1_3_36_36 ;
      VIA 17.652 7.83 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 7.813 17.697 7.847 ;
      VIA 17.652 7.83 Element_VIA34_1_2_58_52 ;
      VIA 17.652 7.83 Element_VIA23_1_3_36_36 ;
      VIA 17.652 7.29 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 7.273 17.697 7.307 ;
      VIA 17.652 7.29 Element_VIA34_1_2_58_52 ;
      VIA 17.652 7.29 Element_VIA23_1_3_36_36 ;
      VIA 17.652 6.75 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 6.733 17.697 6.767 ;
      VIA 17.652 6.75 Element_VIA34_1_2_58_52 ;
      VIA 17.652 6.75 Element_VIA23_1_3_36_36 ;
      VIA 17.652 6.21 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 6.193 17.697 6.227 ;
      VIA 17.652 6.21 Element_VIA34_1_2_58_52 ;
      VIA 17.652 6.21 Element_VIA23_1_3_36_36 ;
      VIA 17.652 5.67 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 5.653 17.697 5.687 ;
      VIA 17.652 5.67 Element_VIA34_1_2_58_52 ;
      VIA 17.652 5.67 Element_VIA23_1_3_36_36 ;
      VIA 17.652 5.13 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 5.113 17.697 5.147 ;
      VIA 17.652 5.13 Element_VIA34_1_2_58_52 ;
      VIA 17.652 5.13 Element_VIA23_1_3_36_36 ;
      VIA 17.652 4.59 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 4.573 17.697 4.607 ;
      VIA 17.652 4.59 Element_VIA34_1_2_58_52 ;
      VIA 17.652 4.59 Element_VIA23_1_3_36_36 ;
      VIA 17.652 4.05 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 4.033 17.697 4.067 ;
      VIA 17.652 4.05 Element_VIA34_1_2_58_52 ;
      VIA 17.652 4.05 Element_VIA23_1_3_36_36 ;
      VIA 17.652 3.51 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 3.493 17.697 3.527 ;
      VIA 17.652 3.51 Element_VIA34_1_2_58_52 ;
      VIA 17.652 3.51 Element_VIA23_1_3_36_36 ;
      VIA 17.652 2.97 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 2.953 17.697 2.987 ;
      VIA 17.652 2.97 Element_VIA34_1_2_58_52 ;
      VIA 17.652 2.97 Element_VIA23_1_3_36_36 ;
      VIA 17.652 2.43 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 2.413 17.697 2.447 ;
      VIA 17.652 2.43 Element_VIA34_1_2_58_52 ;
      VIA 17.652 2.43 Element_VIA23_1_3_36_36 ;
      VIA 17.652 1.89 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 1.873 17.697 1.907 ;
      VIA 17.652 1.89 Element_VIA34_1_2_58_52 ;
      VIA 17.652 1.89 Element_VIA23_1_3_36_36 ;
      VIA 17.652 1.35 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.607 1.333 17.697 1.367 ;
      VIA 17.652 1.35 Element_VIA34_1_2_58_52 ;
      VIA 17.652 1.35 Element_VIA23_1_3_36_36 ;
      VIA 14.676 41.85 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 41.833 14.721 41.867 ;
      VIA 14.676 41.85 Element_VIA34_1_2_58_52 ;
      VIA 14.676 41.85 Element_VIA23_1_3_36_36 ;
      VIA 14.676 41.31 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 41.293 14.721 41.327 ;
      VIA 14.676 41.31 Element_VIA34_1_2_58_52 ;
      VIA 14.676 41.31 Element_VIA23_1_3_36_36 ;
      VIA 14.676 40.77 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 40.753 14.721 40.787 ;
      VIA 14.676 40.77 Element_VIA34_1_2_58_52 ;
      VIA 14.676 40.77 Element_VIA23_1_3_36_36 ;
      VIA 14.676 40.23 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 40.213 14.721 40.247 ;
      VIA 14.676 40.23 Element_VIA34_1_2_58_52 ;
      VIA 14.676 40.23 Element_VIA23_1_3_36_36 ;
      VIA 14.676 39.69 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 39.673 14.721 39.707 ;
      VIA 14.676 39.69 Element_VIA34_1_2_58_52 ;
      VIA 14.676 39.69 Element_VIA23_1_3_36_36 ;
      VIA 14.676 39.15 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 39.133 14.721 39.167 ;
      VIA 14.676 39.15 Element_VIA34_1_2_58_52 ;
      VIA 14.676 39.15 Element_VIA23_1_3_36_36 ;
      VIA 14.676 38.61 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 38.593 14.721 38.627 ;
      VIA 14.676 38.61 Element_VIA34_1_2_58_52 ;
      VIA 14.676 38.61 Element_VIA23_1_3_36_36 ;
      VIA 14.676 38.07 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 38.053 14.721 38.087 ;
      VIA 14.676 38.07 Element_VIA34_1_2_58_52 ;
      VIA 14.676 38.07 Element_VIA23_1_3_36_36 ;
      VIA 14.676 37.53 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 37.513 14.721 37.547 ;
      VIA 14.676 37.53 Element_VIA34_1_2_58_52 ;
      VIA 14.676 37.53 Element_VIA23_1_3_36_36 ;
      VIA 14.676 36.99 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 36.973 14.721 37.007 ;
      VIA 14.676 36.99 Element_VIA34_1_2_58_52 ;
      VIA 14.676 36.99 Element_VIA23_1_3_36_36 ;
      VIA 14.676 36.45 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 36.433 14.721 36.467 ;
      VIA 14.676 36.45 Element_VIA34_1_2_58_52 ;
      VIA 14.676 36.45 Element_VIA23_1_3_36_36 ;
      VIA 14.676 35.91 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 35.893 14.721 35.927 ;
      VIA 14.676 35.91 Element_VIA34_1_2_58_52 ;
      VIA 14.676 35.91 Element_VIA23_1_3_36_36 ;
      VIA 14.676 35.37 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 35.353 14.721 35.387 ;
      VIA 14.676 35.37 Element_VIA34_1_2_58_52 ;
      VIA 14.676 35.37 Element_VIA23_1_3_36_36 ;
      VIA 14.676 34.83 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 34.813 14.721 34.847 ;
      VIA 14.676 34.83 Element_VIA34_1_2_58_52 ;
      VIA 14.676 34.83 Element_VIA23_1_3_36_36 ;
      VIA 14.676 34.29 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 34.273 14.721 34.307 ;
      VIA 14.676 34.29 Element_VIA34_1_2_58_52 ;
      VIA 14.676 34.29 Element_VIA23_1_3_36_36 ;
      VIA 14.676 33.75 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 33.733 14.721 33.767 ;
      VIA 14.676 33.75 Element_VIA34_1_2_58_52 ;
      VIA 14.676 33.75 Element_VIA23_1_3_36_36 ;
      VIA 14.676 33.21 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 33.193 14.721 33.227 ;
      VIA 14.676 33.21 Element_VIA34_1_2_58_52 ;
      VIA 14.676 33.21 Element_VIA23_1_3_36_36 ;
      VIA 14.676 32.67 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 32.653 14.721 32.687 ;
      VIA 14.676 32.67 Element_VIA34_1_2_58_52 ;
      VIA 14.676 32.67 Element_VIA23_1_3_36_36 ;
      VIA 14.676 32.13 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 32.113 14.721 32.147 ;
      VIA 14.676 32.13 Element_VIA34_1_2_58_52 ;
      VIA 14.676 32.13 Element_VIA23_1_3_36_36 ;
      VIA 14.676 31.59 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 31.573 14.721 31.607 ;
      VIA 14.676 31.59 Element_VIA34_1_2_58_52 ;
      VIA 14.676 31.59 Element_VIA23_1_3_36_36 ;
      VIA 14.676 31.05 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 31.033 14.721 31.067 ;
      VIA 14.676 31.05 Element_VIA34_1_2_58_52 ;
      VIA 14.676 31.05 Element_VIA23_1_3_36_36 ;
      VIA 14.676 30.51 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 30.493 14.721 30.527 ;
      VIA 14.676 30.51 Element_VIA34_1_2_58_52 ;
      VIA 14.676 30.51 Element_VIA23_1_3_36_36 ;
      VIA 14.676 29.97 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 29.953 14.721 29.987 ;
      VIA 14.676 29.97 Element_VIA34_1_2_58_52 ;
      VIA 14.676 29.97 Element_VIA23_1_3_36_36 ;
      VIA 14.676 29.43 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 29.413 14.721 29.447 ;
      VIA 14.676 29.43 Element_VIA34_1_2_58_52 ;
      VIA 14.676 29.43 Element_VIA23_1_3_36_36 ;
      VIA 14.676 28.89 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 28.873 14.721 28.907 ;
      VIA 14.676 28.89 Element_VIA34_1_2_58_52 ;
      VIA 14.676 28.89 Element_VIA23_1_3_36_36 ;
      VIA 14.676 28.35 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 28.333 14.721 28.367 ;
      VIA 14.676 28.35 Element_VIA34_1_2_58_52 ;
      VIA 14.676 28.35 Element_VIA23_1_3_36_36 ;
      VIA 14.676 27.81 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 27.793 14.721 27.827 ;
      VIA 14.676 27.81 Element_VIA34_1_2_58_52 ;
      VIA 14.676 27.81 Element_VIA23_1_3_36_36 ;
      VIA 14.676 27.27 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 27.253 14.721 27.287 ;
      VIA 14.676 27.27 Element_VIA34_1_2_58_52 ;
      VIA 14.676 27.27 Element_VIA23_1_3_36_36 ;
      VIA 14.676 26.73 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 26.713 14.721 26.747 ;
      VIA 14.676 26.73 Element_VIA34_1_2_58_52 ;
      VIA 14.676 26.73 Element_VIA23_1_3_36_36 ;
      VIA 14.676 26.19 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 26.173 14.721 26.207 ;
      VIA 14.676 26.19 Element_VIA34_1_2_58_52 ;
      VIA 14.676 26.19 Element_VIA23_1_3_36_36 ;
      VIA 14.676 25.65 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 25.633 14.721 25.667 ;
      VIA 14.676 25.65 Element_VIA34_1_2_58_52 ;
      VIA 14.676 25.65 Element_VIA23_1_3_36_36 ;
      VIA 14.676 25.11 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 25.093 14.721 25.127 ;
      VIA 14.676 25.11 Element_VIA34_1_2_58_52 ;
      VIA 14.676 25.11 Element_VIA23_1_3_36_36 ;
      VIA 14.676 24.57 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 24.553 14.721 24.587 ;
      VIA 14.676 24.57 Element_VIA34_1_2_58_52 ;
      VIA 14.676 24.57 Element_VIA23_1_3_36_36 ;
      VIA 14.676 24.03 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 24.013 14.721 24.047 ;
      VIA 14.676 24.03 Element_VIA34_1_2_58_52 ;
      VIA 14.676 24.03 Element_VIA23_1_3_36_36 ;
      VIA 14.676 23.49 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 23.473 14.721 23.507 ;
      VIA 14.676 23.49 Element_VIA34_1_2_58_52 ;
      VIA 14.676 23.49 Element_VIA23_1_3_36_36 ;
      VIA 14.676 22.95 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 22.933 14.721 22.967 ;
      VIA 14.676 22.95 Element_VIA34_1_2_58_52 ;
      VIA 14.676 22.95 Element_VIA23_1_3_36_36 ;
      VIA 14.676 22.41 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 22.393 14.721 22.427 ;
      VIA 14.676 22.41 Element_VIA34_1_2_58_52 ;
      VIA 14.676 22.41 Element_VIA23_1_3_36_36 ;
      VIA 14.676 21.87 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 21.853 14.721 21.887 ;
      VIA 14.676 21.87 Element_VIA34_1_2_58_52 ;
      VIA 14.676 21.87 Element_VIA23_1_3_36_36 ;
      VIA 14.676 21.33 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 21.313 14.721 21.347 ;
      VIA 14.676 21.33 Element_VIA34_1_2_58_52 ;
      VIA 14.676 21.33 Element_VIA23_1_3_36_36 ;
      VIA 14.676 20.79 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 20.773 14.721 20.807 ;
      VIA 14.676 20.79 Element_VIA34_1_2_58_52 ;
      VIA 14.676 20.79 Element_VIA23_1_3_36_36 ;
      VIA 14.676 20.25 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 20.233 14.721 20.267 ;
      VIA 14.676 20.25 Element_VIA34_1_2_58_52 ;
      VIA 14.676 20.25 Element_VIA23_1_3_36_36 ;
      VIA 14.676 19.71 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 19.693 14.721 19.727 ;
      VIA 14.676 19.71 Element_VIA34_1_2_58_52 ;
      VIA 14.676 19.71 Element_VIA23_1_3_36_36 ;
      VIA 14.676 19.17 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 19.153 14.721 19.187 ;
      VIA 14.676 19.17 Element_VIA34_1_2_58_52 ;
      VIA 14.676 19.17 Element_VIA23_1_3_36_36 ;
      VIA 14.676 18.63 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 18.613 14.721 18.647 ;
      VIA 14.676 18.63 Element_VIA34_1_2_58_52 ;
      VIA 14.676 18.63 Element_VIA23_1_3_36_36 ;
      VIA 14.676 18.09 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 18.073 14.721 18.107 ;
      VIA 14.676 18.09 Element_VIA34_1_2_58_52 ;
      VIA 14.676 18.09 Element_VIA23_1_3_36_36 ;
      VIA 14.676 17.55 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 17.533 14.721 17.567 ;
      VIA 14.676 17.55 Element_VIA34_1_2_58_52 ;
      VIA 14.676 17.55 Element_VIA23_1_3_36_36 ;
      VIA 14.676 17.01 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 16.993 14.721 17.027 ;
      VIA 14.676 17.01 Element_VIA34_1_2_58_52 ;
      VIA 14.676 17.01 Element_VIA23_1_3_36_36 ;
      VIA 14.676 16.47 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 16.453 14.721 16.487 ;
      VIA 14.676 16.47 Element_VIA34_1_2_58_52 ;
      VIA 14.676 16.47 Element_VIA23_1_3_36_36 ;
      VIA 14.676 15.93 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 15.913 14.721 15.947 ;
      VIA 14.676 15.93 Element_VIA34_1_2_58_52 ;
      VIA 14.676 15.93 Element_VIA23_1_3_36_36 ;
      VIA 14.676 15.39 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 15.373 14.721 15.407 ;
      VIA 14.676 15.39 Element_VIA34_1_2_58_52 ;
      VIA 14.676 15.39 Element_VIA23_1_3_36_36 ;
      VIA 14.676 14.85 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 14.833 14.721 14.867 ;
      VIA 14.676 14.85 Element_VIA34_1_2_58_52 ;
      VIA 14.676 14.85 Element_VIA23_1_3_36_36 ;
      VIA 14.676 14.31 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 14.293 14.721 14.327 ;
      VIA 14.676 14.31 Element_VIA34_1_2_58_52 ;
      VIA 14.676 14.31 Element_VIA23_1_3_36_36 ;
      VIA 14.676 13.77 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 13.753 14.721 13.787 ;
      VIA 14.676 13.77 Element_VIA34_1_2_58_52 ;
      VIA 14.676 13.77 Element_VIA23_1_3_36_36 ;
      VIA 14.676 13.23 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 13.213 14.721 13.247 ;
      VIA 14.676 13.23 Element_VIA34_1_2_58_52 ;
      VIA 14.676 13.23 Element_VIA23_1_3_36_36 ;
      VIA 14.676 12.69 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 12.673 14.721 12.707 ;
      VIA 14.676 12.69 Element_VIA34_1_2_58_52 ;
      VIA 14.676 12.69 Element_VIA23_1_3_36_36 ;
      VIA 14.676 12.15 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 12.133 14.721 12.167 ;
      VIA 14.676 12.15 Element_VIA34_1_2_58_52 ;
      VIA 14.676 12.15 Element_VIA23_1_3_36_36 ;
      VIA 14.676 11.61 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 11.593 14.721 11.627 ;
      VIA 14.676 11.61 Element_VIA34_1_2_58_52 ;
      VIA 14.676 11.61 Element_VIA23_1_3_36_36 ;
      VIA 14.676 11.07 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 11.053 14.721 11.087 ;
      VIA 14.676 11.07 Element_VIA34_1_2_58_52 ;
      VIA 14.676 11.07 Element_VIA23_1_3_36_36 ;
      VIA 14.676 10.53 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 10.513 14.721 10.547 ;
      VIA 14.676 10.53 Element_VIA34_1_2_58_52 ;
      VIA 14.676 10.53 Element_VIA23_1_3_36_36 ;
      VIA 14.676 9.99 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 9.973 14.721 10.007 ;
      VIA 14.676 9.99 Element_VIA34_1_2_58_52 ;
      VIA 14.676 9.99 Element_VIA23_1_3_36_36 ;
      VIA 14.676 9.45 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 9.433 14.721 9.467 ;
      VIA 14.676 9.45 Element_VIA34_1_2_58_52 ;
      VIA 14.676 9.45 Element_VIA23_1_3_36_36 ;
      VIA 14.676 8.91 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 8.893 14.721 8.927 ;
      VIA 14.676 8.91 Element_VIA34_1_2_58_52 ;
      VIA 14.676 8.91 Element_VIA23_1_3_36_36 ;
      VIA 14.676 8.37 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 8.353 14.721 8.387 ;
      VIA 14.676 8.37 Element_VIA34_1_2_58_52 ;
      VIA 14.676 8.37 Element_VIA23_1_3_36_36 ;
      VIA 14.676 7.83 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 7.813 14.721 7.847 ;
      VIA 14.676 7.83 Element_VIA34_1_2_58_52 ;
      VIA 14.676 7.83 Element_VIA23_1_3_36_36 ;
      VIA 14.676 7.29 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 7.273 14.721 7.307 ;
      VIA 14.676 7.29 Element_VIA34_1_2_58_52 ;
      VIA 14.676 7.29 Element_VIA23_1_3_36_36 ;
      VIA 14.676 6.75 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 6.733 14.721 6.767 ;
      VIA 14.676 6.75 Element_VIA34_1_2_58_52 ;
      VIA 14.676 6.75 Element_VIA23_1_3_36_36 ;
      VIA 14.676 6.21 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 6.193 14.721 6.227 ;
      VIA 14.676 6.21 Element_VIA34_1_2_58_52 ;
      VIA 14.676 6.21 Element_VIA23_1_3_36_36 ;
      VIA 14.676 5.67 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 5.653 14.721 5.687 ;
      VIA 14.676 5.67 Element_VIA34_1_2_58_52 ;
      VIA 14.676 5.67 Element_VIA23_1_3_36_36 ;
      VIA 14.676 5.13 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 5.113 14.721 5.147 ;
      VIA 14.676 5.13 Element_VIA34_1_2_58_52 ;
      VIA 14.676 5.13 Element_VIA23_1_3_36_36 ;
      VIA 14.676 4.59 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 4.573 14.721 4.607 ;
      VIA 14.676 4.59 Element_VIA34_1_2_58_52 ;
      VIA 14.676 4.59 Element_VIA23_1_3_36_36 ;
      VIA 14.676 4.05 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 4.033 14.721 4.067 ;
      VIA 14.676 4.05 Element_VIA34_1_2_58_52 ;
      VIA 14.676 4.05 Element_VIA23_1_3_36_36 ;
      VIA 14.676 3.51 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 3.493 14.721 3.527 ;
      VIA 14.676 3.51 Element_VIA34_1_2_58_52 ;
      VIA 14.676 3.51 Element_VIA23_1_3_36_36 ;
      VIA 14.676 2.97 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 2.953 14.721 2.987 ;
      VIA 14.676 2.97 Element_VIA34_1_2_58_52 ;
      VIA 14.676 2.97 Element_VIA23_1_3_36_36 ;
      VIA 14.676 2.43 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 2.413 14.721 2.447 ;
      VIA 14.676 2.43 Element_VIA34_1_2_58_52 ;
      VIA 14.676 2.43 Element_VIA23_1_3_36_36 ;
      VIA 14.676 1.89 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 1.873 14.721 1.907 ;
      VIA 14.676 1.89 Element_VIA34_1_2_58_52 ;
      VIA 14.676 1.89 Element_VIA23_1_3_36_36 ;
      VIA 14.676 1.35 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.631 1.333 14.721 1.367 ;
      VIA 14.676 1.35 Element_VIA34_1_2_58_52 ;
      VIA 14.676 1.35 Element_VIA23_1_3_36_36 ;
      VIA 11.7 41.85 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 41.833 11.745 41.867 ;
      VIA 11.7 41.85 Element_VIA34_1_2_58_52 ;
      VIA 11.7 41.85 Element_VIA23_1_3_36_36 ;
      VIA 11.7 41.31 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 41.293 11.745 41.327 ;
      VIA 11.7 41.31 Element_VIA34_1_2_58_52 ;
      VIA 11.7 41.31 Element_VIA23_1_3_36_36 ;
      VIA 11.7 40.77 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 40.753 11.745 40.787 ;
      VIA 11.7 40.77 Element_VIA34_1_2_58_52 ;
      VIA 11.7 40.77 Element_VIA23_1_3_36_36 ;
      VIA 11.7 40.23 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 40.213 11.745 40.247 ;
      VIA 11.7 40.23 Element_VIA34_1_2_58_52 ;
      VIA 11.7 40.23 Element_VIA23_1_3_36_36 ;
      VIA 11.7 39.69 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 39.673 11.745 39.707 ;
      VIA 11.7 39.69 Element_VIA34_1_2_58_52 ;
      VIA 11.7 39.69 Element_VIA23_1_3_36_36 ;
      VIA 11.7 39.15 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 39.133 11.745 39.167 ;
      VIA 11.7 39.15 Element_VIA34_1_2_58_52 ;
      VIA 11.7 39.15 Element_VIA23_1_3_36_36 ;
      VIA 11.7 38.61 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 38.593 11.745 38.627 ;
      VIA 11.7 38.61 Element_VIA34_1_2_58_52 ;
      VIA 11.7 38.61 Element_VIA23_1_3_36_36 ;
      VIA 11.7 38.07 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 38.053 11.745 38.087 ;
      VIA 11.7 38.07 Element_VIA34_1_2_58_52 ;
      VIA 11.7 38.07 Element_VIA23_1_3_36_36 ;
      VIA 11.7 37.53 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 37.513 11.745 37.547 ;
      VIA 11.7 37.53 Element_VIA34_1_2_58_52 ;
      VIA 11.7 37.53 Element_VIA23_1_3_36_36 ;
      VIA 11.7 36.99 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 36.973 11.745 37.007 ;
      VIA 11.7 36.99 Element_VIA34_1_2_58_52 ;
      VIA 11.7 36.99 Element_VIA23_1_3_36_36 ;
      VIA 11.7 36.45 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 36.433 11.745 36.467 ;
      VIA 11.7 36.45 Element_VIA34_1_2_58_52 ;
      VIA 11.7 36.45 Element_VIA23_1_3_36_36 ;
      VIA 11.7 35.91 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 35.893 11.745 35.927 ;
      VIA 11.7 35.91 Element_VIA34_1_2_58_52 ;
      VIA 11.7 35.91 Element_VIA23_1_3_36_36 ;
      VIA 11.7 35.37 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 35.353 11.745 35.387 ;
      VIA 11.7 35.37 Element_VIA34_1_2_58_52 ;
      VIA 11.7 35.37 Element_VIA23_1_3_36_36 ;
      VIA 11.7 34.83 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 34.813 11.745 34.847 ;
      VIA 11.7 34.83 Element_VIA34_1_2_58_52 ;
      VIA 11.7 34.83 Element_VIA23_1_3_36_36 ;
      VIA 11.7 34.29 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 34.273 11.745 34.307 ;
      VIA 11.7 34.29 Element_VIA34_1_2_58_52 ;
      VIA 11.7 34.29 Element_VIA23_1_3_36_36 ;
      VIA 11.7 33.75 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 33.733 11.745 33.767 ;
      VIA 11.7 33.75 Element_VIA34_1_2_58_52 ;
      VIA 11.7 33.75 Element_VIA23_1_3_36_36 ;
      VIA 11.7 33.21 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 33.193 11.745 33.227 ;
      VIA 11.7 33.21 Element_VIA34_1_2_58_52 ;
      VIA 11.7 33.21 Element_VIA23_1_3_36_36 ;
      VIA 11.7 32.67 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 32.653 11.745 32.687 ;
      VIA 11.7 32.67 Element_VIA34_1_2_58_52 ;
      VIA 11.7 32.67 Element_VIA23_1_3_36_36 ;
      VIA 11.7 32.13 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 32.113 11.745 32.147 ;
      VIA 11.7 32.13 Element_VIA34_1_2_58_52 ;
      VIA 11.7 32.13 Element_VIA23_1_3_36_36 ;
      VIA 11.7 31.59 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 31.573 11.745 31.607 ;
      VIA 11.7 31.59 Element_VIA34_1_2_58_52 ;
      VIA 11.7 31.59 Element_VIA23_1_3_36_36 ;
      VIA 11.7 31.05 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 31.033 11.745 31.067 ;
      VIA 11.7 31.05 Element_VIA34_1_2_58_52 ;
      VIA 11.7 31.05 Element_VIA23_1_3_36_36 ;
      VIA 11.7 30.51 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 30.493 11.745 30.527 ;
      VIA 11.7 30.51 Element_VIA34_1_2_58_52 ;
      VIA 11.7 30.51 Element_VIA23_1_3_36_36 ;
      VIA 11.7 29.97 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 29.953 11.745 29.987 ;
      VIA 11.7 29.97 Element_VIA34_1_2_58_52 ;
      VIA 11.7 29.97 Element_VIA23_1_3_36_36 ;
      VIA 11.7 29.43 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 29.413 11.745 29.447 ;
      VIA 11.7 29.43 Element_VIA34_1_2_58_52 ;
      VIA 11.7 29.43 Element_VIA23_1_3_36_36 ;
      VIA 11.7 28.89 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 28.873 11.745 28.907 ;
      VIA 11.7 28.89 Element_VIA34_1_2_58_52 ;
      VIA 11.7 28.89 Element_VIA23_1_3_36_36 ;
      VIA 11.7 28.35 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 28.333 11.745 28.367 ;
      VIA 11.7 28.35 Element_VIA34_1_2_58_52 ;
      VIA 11.7 28.35 Element_VIA23_1_3_36_36 ;
      VIA 11.7 27.81 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 27.793 11.745 27.827 ;
      VIA 11.7 27.81 Element_VIA34_1_2_58_52 ;
      VIA 11.7 27.81 Element_VIA23_1_3_36_36 ;
      VIA 11.7 27.27 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 27.253 11.745 27.287 ;
      VIA 11.7 27.27 Element_VIA34_1_2_58_52 ;
      VIA 11.7 27.27 Element_VIA23_1_3_36_36 ;
      VIA 11.7 26.73 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 26.713 11.745 26.747 ;
      VIA 11.7 26.73 Element_VIA34_1_2_58_52 ;
      VIA 11.7 26.73 Element_VIA23_1_3_36_36 ;
      VIA 11.7 26.19 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 26.173 11.745 26.207 ;
      VIA 11.7 26.19 Element_VIA34_1_2_58_52 ;
      VIA 11.7 26.19 Element_VIA23_1_3_36_36 ;
      VIA 11.7 25.65 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 25.633 11.745 25.667 ;
      VIA 11.7 25.65 Element_VIA34_1_2_58_52 ;
      VIA 11.7 25.65 Element_VIA23_1_3_36_36 ;
      VIA 11.7 25.11 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 25.093 11.745 25.127 ;
      VIA 11.7 25.11 Element_VIA34_1_2_58_52 ;
      VIA 11.7 25.11 Element_VIA23_1_3_36_36 ;
      VIA 11.7 24.57 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 24.553 11.745 24.587 ;
      VIA 11.7 24.57 Element_VIA34_1_2_58_52 ;
      VIA 11.7 24.57 Element_VIA23_1_3_36_36 ;
      VIA 11.7 24.03 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 24.013 11.745 24.047 ;
      VIA 11.7 24.03 Element_VIA34_1_2_58_52 ;
      VIA 11.7 24.03 Element_VIA23_1_3_36_36 ;
      VIA 11.7 23.49 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 23.473 11.745 23.507 ;
      VIA 11.7 23.49 Element_VIA34_1_2_58_52 ;
      VIA 11.7 23.49 Element_VIA23_1_3_36_36 ;
      VIA 11.7 22.95 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 22.933 11.745 22.967 ;
      VIA 11.7 22.95 Element_VIA34_1_2_58_52 ;
      VIA 11.7 22.95 Element_VIA23_1_3_36_36 ;
      VIA 11.7 22.41 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 22.393 11.745 22.427 ;
      VIA 11.7 22.41 Element_VIA34_1_2_58_52 ;
      VIA 11.7 22.41 Element_VIA23_1_3_36_36 ;
      VIA 11.7 21.87 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 21.853 11.745 21.887 ;
      VIA 11.7 21.87 Element_VIA34_1_2_58_52 ;
      VIA 11.7 21.87 Element_VIA23_1_3_36_36 ;
      VIA 11.7 21.33 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 21.313 11.745 21.347 ;
      VIA 11.7 21.33 Element_VIA34_1_2_58_52 ;
      VIA 11.7 21.33 Element_VIA23_1_3_36_36 ;
      VIA 11.7 20.79 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 20.773 11.745 20.807 ;
      VIA 11.7 20.79 Element_VIA34_1_2_58_52 ;
      VIA 11.7 20.79 Element_VIA23_1_3_36_36 ;
      VIA 11.7 20.25 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 20.233 11.745 20.267 ;
      VIA 11.7 20.25 Element_VIA34_1_2_58_52 ;
      VIA 11.7 20.25 Element_VIA23_1_3_36_36 ;
      VIA 11.7 19.71 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 19.693 11.745 19.727 ;
      VIA 11.7 19.71 Element_VIA34_1_2_58_52 ;
      VIA 11.7 19.71 Element_VIA23_1_3_36_36 ;
      VIA 11.7 19.17 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 19.153 11.745 19.187 ;
      VIA 11.7 19.17 Element_VIA34_1_2_58_52 ;
      VIA 11.7 19.17 Element_VIA23_1_3_36_36 ;
      VIA 11.7 18.63 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 18.613 11.745 18.647 ;
      VIA 11.7 18.63 Element_VIA34_1_2_58_52 ;
      VIA 11.7 18.63 Element_VIA23_1_3_36_36 ;
      VIA 11.7 18.09 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 18.073 11.745 18.107 ;
      VIA 11.7 18.09 Element_VIA34_1_2_58_52 ;
      VIA 11.7 18.09 Element_VIA23_1_3_36_36 ;
      VIA 11.7 17.55 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 17.533 11.745 17.567 ;
      VIA 11.7 17.55 Element_VIA34_1_2_58_52 ;
      VIA 11.7 17.55 Element_VIA23_1_3_36_36 ;
      VIA 11.7 17.01 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 16.993 11.745 17.027 ;
      VIA 11.7 17.01 Element_VIA34_1_2_58_52 ;
      VIA 11.7 17.01 Element_VIA23_1_3_36_36 ;
      VIA 11.7 16.47 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 16.453 11.745 16.487 ;
      VIA 11.7 16.47 Element_VIA34_1_2_58_52 ;
      VIA 11.7 16.47 Element_VIA23_1_3_36_36 ;
      VIA 11.7 15.93 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 15.913 11.745 15.947 ;
      VIA 11.7 15.93 Element_VIA34_1_2_58_52 ;
      VIA 11.7 15.93 Element_VIA23_1_3_36_36 ;
      VIA 11.7 15.39 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 15.373 11.745 15.407 ;
      VIA 11.7 15.39 Element_VIA34_1_2_58_52 ;
      VIA 11.7 15.39 Element_VIA23_1_3_36_36 ;
      VIA 11.7 14.85 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 14.833 11.745 14.867 ;
      VIA 11.7 14.85 Element_VIA34_1_2_58_52 ;
      VIA 11.7 14.85 Element_VIA23_1_3_36_36 ;
      VIA 11.7 14.31 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 14.293 11.745 14.327 ;
      VIA 11.7 14.31 Element_VIA34_1_2_58_52 ;
      VIA 11.7 14.31 Element_VIA23_1_3_36_36 ;
      VIA 11.7 13.77 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 13.753 11.745 13.787 ;
      VIA 11.7 13.77 Element_VIA34_1_2_58_52 ;
      VIA 11.7 13.77 Element_VIA23_1_3_36_36 ;
      VIA 11.7 13.23 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 13.213 11.745 13.247 ;
      VIA 11.7 13.23 Element_VIA34_1_2_58_52 ;
      VIA 11.7 13.23 Element_VIA23_1_3_36_36 ;
      VIA 11.7 12.69 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 12.673 11.745 12.707 ;
      VIA 11.7 12.69 Element_VIA34_1_2_58_52 ;
      VIA 11.7 12.69 Element_VIA23_1_3_36_36 ;
      VIA 11.7 12.15 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 12.133 11.745 12.167 ;
      VIA 11.7 12.15 Element_VIA34_1_2_58_52 ;
      VIA 11.7 12.15 Element_VIA23_1_3_36_36 ;
      VIA 11.7 11.61 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 11.593 11.745 11.627 ;
      VIA 11.7 11.61 Element_VIA34_1_2_58_52 ;
      VIA 11.7 11.61 Element_VIA23_1_3_36_36 ;
      VIA 11.7 11.07 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 11.053 11.745 11.087 ;
      VIA 11.7 11.07 Element_VIA34_1_2_58_52 ;
      VIA 11.7 11.07 Element_VIA23_1_3_36_36 ;
      VIA 11.7 10.53 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 10.513 11.745 10.547 ;
      VIA 11.7 10.53 Element_VIA34_1_2_58_52 ;
      VIA 11.7 10.53 Element_VIA23_1_3_36_36 ;
      VIA 11.7 9.99 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 9.973 11.745 10.007 ;
      VIA 11.7 9.99 Element_VIA34_1_2_58_52 ;
      VIA 11.7 9.99 Element_VIA23_1_3_36_36 ;
      VIA 11.7 9.45 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 9.433 11.745 9.467 ;
      VIA 11.7 9.45 Element_VIA34_1_2_58_52 ;
      VIA 11.7 9.45 Element_VIA23_1_3_36_36 ;
      VIA 11.7 8.91 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 8.893 11.745 8.927 ;
      VIA 11.7 8.91 Element_VIA34_1_2_58_52 ;
      VIA 11.7 8.91 Element_VIA23_1_3_36_36 ;
      VIA 11.7 8.37 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 8.353 11.745 8.387 ;
      VIA 11.7 8.37 Element_VIA34_1_2_58_52 ;
      VIA 11.7 8.37 Element_VIA23_1_3_36_36 ;
      VIA 11.7 7.83 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 7.813 11.745 7.847 ;
      VIA 11.7 7.83 Element_VIA34_1_2_58_52 ;
      VIA 11.7 7.83 Element_VIA23_1_3_36_36 ;
      VIA 11.7 7.29 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 7.273 11.745 7.307 ;
      VIA 11.7 7.29 Element_VIA34_1_2_58_52 ;
      VIA 11.7 7.29 Element_VIA23_1_3_36_36 ;
      VIA 11.7 6.75 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 6.733 11.745 6.767 ;
      VIA 11.7 6.75 Element_VIA34_1_2_58_52 ;
      VIA 11.7 6.75 Element_VIA23_1_3_36_36 ;
      VIA 11.7 6.21 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 6.193 11.745 6.227 ;
      VIA 11.7 6.21 Element_VIA34_1_2_58_52 ;
      VIA 11.7 6.21 Element_VIA23_1_3_36_36 ;
      VIA 11.7 5.67 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 5.653 11.745 5.687 ;
      VIA 11.7 5.67 Element_VIA34_1_2_58_52 ;
      VIA 11.7 5.67 Element_VIA23_1_3_36_36 ;
      VIA 11.7 5.13 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 5.113 11.745 5.147 ;
      VIA 11.7 5.13 Element_VIA34_1_2_58_52 ;
      VIA 11.7 5.13 Element_VIA23_1_3_36_36 ;
      VIA 11.7 4.59 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 4.573 11.745 4.607 ;
      VIA 11.7 4.59 Element_VIA34_1_2_58_52 ;
      VIA 11.7 4.59 Element_VIA23_1_3_36_36 ;
      VIA 11.7 4.05 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 4.033 11.745 4.067 ;
      VIA 11.7 4.05 Element_VIA34_1_2_58_52 ;
      VIA 11.7 4.05 Element_VIA23_1_3_36_36 ;
      VIA 11.7 3.51 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 3.493 11.745 3.527 ;
      VIA 11.7 3.51 Element_VIA34_1_2_58_52 ;
      VIA 11.7 3.51 Element_VIA23_1_3_36_36 ;
      VIA 11.7 2.97 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 2.953 11.745 2.987 ;
      VIA 11.7 2.97 Element_VIA34_1_2_58_52 ;
      VIA 11.7 2.97 Element_VIA23_1_3_36_36 ;
      VIA 11.7 2.43 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 2.413 11.745 2.447 ;
      VIA 11.7 2.43 Element_VIA34_1_2_58_52 ;
      VIA 11.7 2.43 Element_VIA23_1_3_36_36 ;
      VIA 11.7 1.89 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 1.873 11.745 1.907 ;
      VIA 11.7 1.89 Element_VIA34_1_2_58_52 ;
      VIA 11.7 1.89 Element_VIA23_1_3_36_36 ;
      VIA 11.7 1.35 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.655 1.333 11.745 1.367 ;
      VIA 11.7 1.35 Element_VIA34_1_2_58_52 ;
      VIA 11.7 1.35 Element_VIA23_1_3_36_36 ;
      VIA 8.724 41.85 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 41.833 8.769 41.867 ;
      VIA 8.724 41.85 Element_VIA34_1_2_58_52 ;
      VIA 8.724 41.85 Element_VIA23_1_3_36_36 ;
      VIA 8.724 41.31 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 41.293 8.769 41.327 ;
      VIA 8.724 41.31 Element_VIA34_1_2_58_52 ;
      VIA 8.724 41.31 Element_VIA23_1_3_36_36 ;
      VIA 8.724 40.77 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 40.753 8.769 40.787 ;
      VIA 8.724 40.77 Element_VIA34_1_2_58_52 ;
      VIA 8.724 40.77 Element_VIA23_1_3_36_36 ;
      VIA 8.724 40.23 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 40.213 8.769 40.247 ;
      VIA 8.724 40.23 Element_VIA34_1_2_58_52 ;
      VIA 8.724 40.23 Element_VIA23_1_3_36_36 ;
      VIA 8.724 39.69 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 39.673 8.769 39.707 ;
      VIA 8.724 39.69 Element_VIA34_1_2_58_52 ;
      VIA 8.724 39.69 Element_VIA23_1_3_36_36 ;
      VIA 8.724 39.15 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 39.133 8.769 39.167 ;
      VIA 8.724 39.15 Element_VIA34_1_2_58_52 ;
      VIA 8.724 39.15 Element_VIA23_1_3_36_36 ;
      VIA 8.724 38.61 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 38.593 8.769 38.627 ;
      VIA 8.724 38.61 Element_VIA34_1_2_58_52 ;
      VIA 8.724 38.61 Element_VIA23_1_3_36_36 ;
      VIA 8.724 38.07 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 38.053 8.769 38.087 ;
      VIA 8.724 38.07 Element_VIA34_1_2_58_52 ;
      VIA 8.724 38.07 Element_VIA23_1_3_36_36 ;
      VIA 8.724 37.53 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 37.513 8.769 37.547 ;
      VIA 8.724 37.53 Element_VIA34_1_2_58_52 ;
      VIA 8.724 37.53 Element_VIA23_1_3_36_36 ;
      VIA 8.724 36.99 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 36.973 8.769 37.007 ;
      VIA 8.724 36.99 Element_VIA34_1_2_58_52 ;
      VIA 8.724 36.99 Element_VIA23_1_3_36_36 ;
      VIA 8.724 36.45 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 36.433 8.769 36.467 ;
      VIA 8.724 36.45 Element_VIA34_1_2_58_52 ;
      VIA 8.724 36.45 Element_VIA23_1_3_36_36 ;
      VIA 8.724 35.91 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 35.893 8.769 35.927 ;
      VIA 8.724 35.91 Element_VIA34_1_2_58_52 ;
      VIA 8.724 35.91 Element_VIA23_1_3_36_36 ;
      VIA 8.724 35.37 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 35.353 8.769 35.387 ;
      VIA 8.724 35.37 Element_VIA34_1_2_58_52 ;
      VIA 8.724 35.37 Element_VIA23_1_3_36_36 ;
      VIA 8.724 34.83 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 34.813 8.769 34.847 ;
      VIA 8.724 34.83 Element_VIA34_1_2_58_52 ;
      VIA 8.724 34.83 Element_VIA23_1_3_36_36 ;
      VIA 8.724 34.29 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 34.273 8.769 34.307 ;
      VIA 8.724 34.29 Element_VIA34_1_2_58_52 ;
      VIA 8.724 34.29 Element_VIA23_1_3_36_36 ;
      VIA 8.724 33.75 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 33.733 8.769 33.767 ;
      VIA 8.724 33.75 Element_VIA34_1_2_58_52 ;
      VIA 8.724 33.75 Element_VIA23_1_3_36_36 ;
      VIA 8.724 33.21 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 33.193 8.769 33.227 ;
      VIA 8.724 33.21 Element_VIA34_1_2_58_52 ;
      VIA 8.724 33.21 Element_VIA23_1_3_36_36 ;
      VIA 8.724 32.67 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 32.653 8.769 32.687 ;
      VIA 8.724 32.67 Element_VIA34_1_2_58_52 ;
      VIA 8.724 32.67 Element_VIA23_1_3_36_36 ;
      VIA 8.724 32.13 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 32.113 8.769 32.147 ;
      VIA 8.724 32.13 Element_VIA34_1_2_58_52 ;
      VIA 8.724 32.13 Element_VIA23_1_3_36_36 ;
      VIA 8.724 31.59 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 31.573 8.769 31.607 ;
      VIA 8.724 31.59 Element_VIA34_1_2_58_52 ;
      VIA 8.724 31.59 Element_VIA23_1_3_36_36 ;
      VIA 8.724 31.05 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 31.033 8.769 31.067 ;
      VIA 8.724 31.05 Element_VIA34_1_2_58_52 ;
      VIA 8.724 31.05 Element_VIA23_1_3_36_36 ;
      VIA 8.724 30.51 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 30.493 8.769 30.527 ;
      VIA 8.724 30.51 Element_VIA34_1_2_58_52 ;
      VIA 8.724 30.51 Element_VIA23_1_3_36_36 ;
      VIA 8.724 29.97 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 29.953 8.769 29.987 ;
      VIA 8.724 29.97 Element_VIA34_1_2_58_52 ;
      VIA 8.724 29.97 Element_VIA23_1_3_36_36 ;
      VIA 8.724 29.43 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 29.413 8.769 29.447 ;
      VIA 8.724 29.43 Element_VIA34_1_2_58_52 ;
      VIA 8.724 29.43 Element_VIA23_1_3_36_36 ;
      VIA 8.724 28.89 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 28.873 8.769 28.907 ;
      VIA 8.724 28.89 Element_VIA34_1_2_58_52 ;
      VIA 8.724 28.89 Element_VIA23_1_3_36_36 ;
      VIA 8.724 28.35 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 28.333 8.769 28.367 ;
      VIA 8.724 28.35 Element_VIA34_1_2_58_52 ;
      VIA 8.724 28.35 Element_VIA23_1_3_36_36 ;
      VIA 8.724 27.81 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 27.793 8.769 27.827 ;
      VIA 8.724 27.81 Element_VIA34_1_2_58_52 ;
      VIA 8.724 27.81 Element_VIA23_1_3_36_36 ;
      VIA 8.724 27.27 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 27.253 8.769 27.287 ;
      VIA 8.724 27.27 Element_VIA34_1_2_58_52 ;
      VIA 8.724 27.27 Element_VIA23_1_3_36_36 ;
      VIA 8.724 26.73 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 26.713 8.769 26.747 ;
      VIA 8.724 26.73 Element_VIA34_1_2_58_52 ;
      VIA 8.724 26.73 Element_VIA23_1_3_36_36 ;
      VIA 8.724 26.19 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 26.173 8.769 26.207 ;
      VIA 8.724 26.19 Element_VIA34_1_2_58_52 ;
      VIA 8.724 26.19 Element_VIA23_1_3_36_36 ;
      VIA 8.724 25.65 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 25.633 8.769 25.667 ;
      VIA 8.724 25.65 Element_VIA34_1_2_58_52 ;
      VIA 8.724 25.65 Element_VIA23_1_3_36_36 ;
      VIA 8.724 25.11 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 25.093 8.769 25.127 ;
      VIA 8.724 25.11 Element_VIA34_1_2_58_52 ;
      VIA 8.724 25.11 Element_VIA23_1_3_36_36 ;
      VIA 8.724 24.57 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 24.553 8.769 24.587 ;
      VIA 8.724 24.57 Element_VIA34_1_2_58_52 ;
      VIA 8.724 24.57 Element_VIA23_1_3_36_36 ;
      VIA 8.724 24.03 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 24.013 8.769 24.047 ;
      VIA 8.724 24.03 Element_VIA34_1_2_58_52 ;
      VIA 8.724 24.03 Element_VIA23_1_3_36_36 ;
      VIA 8.724 23.49 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 23.473 8.769 23.507 ;
      VIA 8.724 23.49 Element_VIA34_1_2_58_52 ;
      VIA 8.724 23.49 Element_VIA23_1_3_36_36 ;
      VIA 8.724 22.95 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 22.933 8.769 22.967 ;
      VIA 8.724 22.95 Element_VIA34_1_2_58_52 ;
      VIA 8.724 22.95 Element_VIA23_1_3_36_36 ;
      VIA 8.724 22.41 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 22.393 8.769 22.427 ;
      VIA 8.724 22.41 Element_VIA34_1_2_58_52 ;
      VIA 8.724 22.41 Element_VIA23_1_3_36_36 ;
      VIA 8.724 21.87 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 21.853 8.769 21.887 ;
      VIA 8.724 21.87 Element_VIA34_1_2_58_52 ;
      VIA 8.724 21.87 Element_VIA23_1_3_36_36 ;
      VIA 8.724 21.33 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 21.313 8.769 21.347 ;
      VIA 8.724 21.33 Element_VIA34_1_2_58_52 ;
      VIA 8.724 21.33 Element_VIA23_1_3_36_36 ;
      VIA 8.724 20.79 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 20.773 8.769 20.807 ;
      VIA 8.724 20.79 Element_VIA34_1_2_58_52 ;
      VIA 8.724 20.79 Element_VIA23_1_3_36_36 ;
      VIA 8.724 20.25 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 20.233 8.769 20.267 ;
      VIA 8.724 20.25 Element_VIA34_1_2_58_52 ;
      VIA 8.724 20.25 Element_VIA23_1_3_36_36 ;
      VIA 8.724 19.71 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 19.693 8.769 19.727 ;
      VIA 8.724 19.71 Element_VIA34_1_2_58_52 ;
      VIA 8.724 19.71 Element_VIA23_1_3_36_36 ;
      VIA 8.724 19.17 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 19.153 8.769 19.187 ;
      VIA 8.724 19.17 Element_VIA34_1_2_58_52 ;
      VIA 8.724 19.17 Element_VIA23_1_3_36_36 ;
      VIA 8.724 18.63 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 18.613 8.769 18.647 ;
      VIA 8.724 18.63 Element_VIA34_1_2_58_52 ;
      VIA 8.724 18.63 Element_VIA23_1_3_36_36 ;
      VIA 8.724 18.09 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 18.073 8.769 18.107 ;
      VIA 8.724 18.09 Element_VIA34_1_2_58_52 ;
      VIA 8.724 18.09 Element_VIA23_1_3_36_36 ;
      VIA 8.724 17.55 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 17.533 8.769 17.567 ;
      VIA 8.724 17.55 Element_VIA34_1_2_58_52 ;
      VIA 8.724 17.55 Element_VIA23_1_3_36_36 ;
      VIA 8.724 17.01 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 16.993 8.769 17.027 ;
      VIA 8.724 17.01 Element_VIA34_1_2_58_52 ;
      VIA 8.724 17.01 Element_VIA23_1_3_36_36 ;
      VIA 8.724 16.47 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 16.453 8.769 16.487 ;
      VIA 8.724 16.47 Element_VIA34_1_2_58_52 ;
      VIA 8.724 16.47 Element_VIA23_1_3_36_36 ;
      VIA 8.724 15.93 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 15.913 8.769 15.947 ;
      VIA 8.724 15.93 Element_VIA34_1_2_58_52 ;
      VIA 8.724 15.93 Element_VIA23_1_3_36_36 ;
      VIA 8.724 15.39 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 15.373 8.769 15.407 ;
      VIA 8.724 15.39 Element_VIA34_1_2_58_52 ;
      VIA 8.724 15.39 Element_VIA23_1_3_36_36 ;
      VIA 8.724 14.85 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 14.833 8.769 14.867 ;
      VIA 8.724 14.85 Element_VIA34_1_2_58_52 ;
      VIA 8.724 14.85 Element_VIA23_1_3_36_36 ;
      VIA 8.724 14.31 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 14.293 8.769 14.327 ;
      VIA 8.724 14.31 Element_VIA34_1_2_58_52 ;
      VIA 8.724 14.31 Element_VIA23_1_3_36_36 ;
      VIA 8.724 13.77 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 13.753 8.769 13.787 ;
      VIA 8.724 13.77 Element_VIA34_1_2_58_52 ;
      VIA 8.724 13.77 Element_VIA23_1_3_36_36 ;
      VIA 8.724 13.23 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 13.213 8.769 13.247 ;
      VIA 8.724 13.23 Element_VIA34_1_2_58_52 ;
      VIA 8.724 13.23 Element_VIA23_1_3_36_36 ;
      VIA 8.724 12.69 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 12.673 8.769 12.707 ;
      VIA 8.724 12.69 Element_VIA34_1_2_58_52 ;
      VIA 8.724 12.69 Element_VIA23_1_3_36_36 ;
      VIA 8.724 12.15 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 12.133 8.769 12.167 ;
      VIA 8.724 12.15 Element_VIA34_1_2_58_52 ;
      VIA 8.724 12.15 Element_VIA23_1_3_36_36 ;
      VIA 8.724 11.61 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 11.593 8.769 11.627 ;
      VIA 8.724 11.61 Element_VIA34_1_2_58_52 ;
      VIA 8.724 11.61 Element_VIA23_1_3_36_36 ;
      VIA 8.724 11.07 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 11.053 8.769 11.087 ;
      VIA 8.724 11.07 Element_VIA34_1_2_58_52 ;
      VIA 8.724 11.07 Element_VIA23_1_3_36_36 ;
      VIA 8.724 10.53 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 10.513 8.769 10.547 ;
      VIA 8.724 10.53 Element_VIA34_1_2_58_52 ;
      VIA 8.724 10.53 Element_VIA23_1_3_36_36 ;
      VIA 8.724 9.99 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 9.973 8.769 10.007 ;
      VIA 8.724 9.99 Element_VIA34_1_2_58_52 ;
      VIA 8.724 9.99 Element_VIA23_1_3_36_36 ;
      VIA 8.724 9.45 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 9.433 8.769 9.467 ;
      VIA 8.724 9.45 Element_VIA34_1_2_58_52 ;
      VIA 8.724 9.45 Element_VIA23_1_3_36_36 ;
      VIA 8.724 8.91 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 8.893 8.769 8.927 ;
      VIA 8.724 8.91 Element_VIA34_1_2_58_52 ;
      VIA 8.724 8.91 Element_VIA23_1_3_36_36 ;
      VIA 8.724 8.37 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 8.353 8.769 8.387 ;
      VIA 8.724 8.37 Element_VIA34_1_2_58_52 ;
      VIA 8.724 8.37 Element_VIA23_1_3_36_36 ;
      VIA 8.724 7.83 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 7.813 8.769 7.847 ;
      VIA 8.724 7.83 Element_VIA34_1_2_58_52 ;
      VIA 8.724 7.83 Element_VIA23_1_3_36_36 ;
      VIA 8.724 7.29 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 7.273 8.769 7.307 ;
      VIA 8.724 7.29 Element_VIA34_1_2_58_52 ;
      VIA 8.724 7.29 Element_VIA23_1_3_36_36 ;
      VIA 8.724 6.75 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 6.733 8.769 6.767 ;
      VIA 8.724 6.75 Element_VIA34_1_2_58_52 ;
      VIA 8.724 6.75 Element_VIA23_1_3_36_36 ;
      VIA 8.724 6.21 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 6.193 8.769 6.227 ;
      VIA 8.724 6.21 Element_VIA34_1_2_58_52 ;
      VIA 8.724 6.21 Element_VIA23_1_3_36_36 ;
      VIA 8.724 5.67 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 5.653 8.769 5.687 ;
      VIA 8.724 5.67 Element_VIA34_1_2_58_52 ;
      VIA 8.724 5.67 Element_VIA23_1_3_36_36 ;
      VIA 8.724 5.13 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 5.113 8.769 5.147 ;
      VIA 8.724 5.13 Element_VIA34_1_2_58_52 ;
      VIA 8.724 5.13 Element_VIA23_1_3_36_36 ;
      VIA 8.724 4.59 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 4.573 8.769 4.607 ;
      VIA 8.724 4.59 Element_VIA34_1_2_58_52 ;
      VIA 8.724 4.59 Element_VIA23_1_3_36_36 ;
      VIA 8.724 4.05 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 4.033 8.769 4.067 ;
      VIA 8.724 4.05 Element_VIA34_1_2_58_52 ;
      VIA 8.724 4.05 Element_VIA23_1_3_36_36 ;
      VIA 8.724 3.51 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 3.493 8.769 3.527 ;
      VIA 8.724 3.51 Element_VIA34_1_2_58_52 ;
      VIA 8.724 3.51 Element_VIA23_1_3_36_36 ;
      VIA 8.724 2.97 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 2.953 8.769 2.987 ;
      VIA 8.724 2.97 Element_VIA34_1_2_58_52 ;
      VIA 8.724 2.97 Element_VIA23_1_3_36_36 ;
      VIA 8.724 2.43 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 2.413 8.769 2.447 ;
      VIA 8.724 2.43 Element_VIA34_1_2_58_52 ;
      VIA 8.724 2.43 Element_VIA23_1_3_36_36 ;
      VIA 8.724 1.89 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 1.873 8.769 1.907 ;
      VIA 8.724 1.89 Element_VIA34_1_2_58_52 ;
      VIA 8.724 1.89 Element_VIA23_1_3_36_36 ;
      VIA 8.724 1.35 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.679 1.333 8.769 1.367 ;
      VIA 8.724 1.35 Element_VIA34_1_2_58_52 ;
      VIA 8.724 1.35 Element_VIA23_1_3_36_36 ;
      VIA 5.748 41.85 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 41.833 5.793 41.867 ;
      VIA 5.748 41.85 Element_VIA34_1_2_58_52 ;
      VIA 5.748 41.85 Element_VIA23_1_3_36_36 ;
      VIA 5.748 41.31 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 41.293 5.793 41.327 ;
      VIA 5.748 41.31 Element_VIA34_1_2_58_52 ;
      VIA 5.748 41.31 Element_VIA23_1_3_36_36 ;
      VIA 5.748 40.77 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 40.753 5.793 40.787 ;
      VIA 5.748 40.77 Element_VIA34_1_2_58_52 ;
      VIA 5.748 40.77 Element_VIA23_1_3_36_36 ;
      VIA 5.748 40.23 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 40.213 5.793 40.247 ;
      VIA 5.748 40.23 Element_VIA34_1_2_58_52 ;
      VIA 5.748 40.23 Element_VIA23_1_3_36_36 ;
      VIA 5.748 39.69 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 39.673 5.793 39.707 ;
      VIA 5.748 39.69 Element_VIA34_1_2_58_52 ;
      VIA 5.748 39.69 Element_VIA23_1_3_36_36 ;
      VIA 5.748 39.15 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 39.133 5.793 39.167 ;
      VIA 5.748 39.15 Element_VIA34_1_2_58_52 ;
      VIA 5.748 39.15 Element_VIA23_1_3_36_36 ;
      VIA 5.748 38.61 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 38.593 5.793 38.627 ;
      VIA 5.748 38.61 Element_VIA34_1_2_58_52 ;
      VIA 5.748 38.61 Element_VIA23_1_3_36_36 ;
      VIA 5.748 38.07 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 38.053 5.793 38.087 ;
      VIA 5.748 38.07 Element_VIA34_1_2_58_52 ;
      VIA 5.748 38.07 Element_VIA23_1_3_36_36 ;
      VIA 5.748 37.53 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 37.513 5.793 37.547 ;
      VIA 5.748 37.53 Element_VIA34_1_2_58_52 ;
      VIA 5.748 37.53 Element_VIA23_1_3_36_36 ;
      VIA 5.748 36.99 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 36.973 5.793 37.007 ;
      VIA 5.748 36.99 Element_VIA34_1_2_58_52 ;
      VIA 5.748 36.99 Element_VIA23_1_3_36_36 ;
      VIA 5.748 36.45 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 36.433 5.793 36.467 ;
      VIA 5.748 36.45 Element_VIA34_1_2_58_52 ;
      VIA 5.748 36.45 Element_VIA23_1_3_36_36 ;
      VIA 5.748 35.91 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 35.893 5.793 35.927 ;
      VIA 5.748 35.91 Element_VIA34_1_2_58_52 ;
      VIA 5.748 35.91 Element_VIA23_1_3_36_36 ;
      VIA 5.748 35.37 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 35.353 5.793 35.387 ;
      VIA 5.748 35.37 Element_VIA34_1_2_58_52 ;
      VIA 5.748 35.37 Element_VIA23_1_3_36_36 ;
      VIA 5.748 34.83 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 34.813 5.793 34.847 ;
      VIA 5.748 34.83 Element_VIA34_1_2_58_52 ;
      VIA 5.748 34.83 Element_VIA23_1_3_36_36 ;
      VIA 5.748 34.29 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 34.273 5.793 34.307 ;
      VIA 5.748 34.29 Element_VIA34_1_2_58_52 ;
      VIA 5.748 34.29 Element_VIA23_1_3_36_36 ;
      VIA 5.748 33.75 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 33.733 5.793 33.767 ;
      VIA 5.748 33.75 Element_VIA34_1_2_58_52 ;
      VIA 5.748 33.75 Element_VIA23_1_3_36_36 ;
      VIA 5.748 33.21 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 33.193 5.793 33.227 ;
      VIA 5.748 33.21 Element_VIA34_1_2_58_52 ;
      VIA 5.748 33.21 Element_VIA23_1_3_36_36 ;
      VIA 5.748 32.67 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 32.653 5.793 32.687 ;
      VIA 5.748 32.67 Element_VIA34_1_2_58_52 ;
      VIA 5.748 32.67 Element_VIA23_1_3_36_36 ;
      VIA 5.748 32.13 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 32.113 5.793 32.147 ;
      VIA 5.748 32.13 Element_VIA34_1_2_58_52 ;
      VIA 5.748 32.13 Element_VIA23_1_3_36_36 ;
      VIA 5.748 31.59 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 31.573 5.793 31.607 ;
      VIA 5.748 31.59 Element_VIA34_1_2_58_52 ;
      VIA 5.748 31.59 Element_VIA23_1_3_36_36 ;
      VIA 5.748 31.05 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 31.033 5.793 31.067 ;
      VIA 5.748 31.05 Element_VIA34_1_2_58_52 ;
      VIA 5.748 31.05 Element_VIA23_1_3_36_36 ;
      VIA 5.748 30.51 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 30.493 5.793 30.527 ;
      VIA 5.748 30.51 Element_VIA34_1_2_58_52 ;
      VIA 5.748 30.51 Element_VIA23_1_3_36_36 ;
      VIA 5.748 29.97 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 29.953 5.793 29.987 ;
      VIA 5.748 29.97 Element_VIA34_1_2_58_52 ;
      VIA 5.748 29.97 Element_VIA23_1_3_36_36 ;
      VIA 5.748 29.43 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 29.413 5.793 29.447 ;
      VIA 5.748 29.43 Element_VIA34_1_2_58_52 ;
      VIA 5.748 29.43 Element_VIA23_1_3_36_36 ;
      VIA 5.748 28.89 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 28.873 5.793 28.907 ;
      VIA 5.748 28.89 Element_VIA34_1_2_58_52 ;
      VIA 5.748 28.89 Element_VIA23_1_3_36_36 ;
      VIA 5.748 28.35 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 28.333 5.793 28.367 ;
      VIA 5.748 28.35 Element_VIA34_1_2_58_52 ;
      VIA 5.748 28.35 Element_VIA23_1_3_36_36 ;
      VIA 5.748 27.81 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 27.793 5.793 27.827 ;
      VIA 5.748 27.81 Element_VIA34_1_2_58_52 ;
      VIA 5.748 27.81 Element_VIA23_1_3_36_36 ;
      VIA 5.748 27.27 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 27.253 5.793 27.287 ;
      VIA 5.748 27.27 Element_VIA34_1_2_58_52 ;
      VIA 5.748 27.27 Element_VIA23_1_3_36_36 ;
      VIA 5.748 26.73 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 26.713 5.793 26.747 ;
      VIA 5.748 26.73 Element_VIA34_1_2_58_52 ;
      VIA 5.748 26.73 Element_VIA23_1_3_36_36 ;
      VIA 5.748 26.19 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 26.173 5.793 26.207 ;
      VIA 5.748 26.19 Element_VIA34_1_2_58_52 ;
      VIA 5.748 26.19 Element_VIA23_1_3_36_36 ;
      VIA 5.748 25.65 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 25.633 5.793 25.667 ;
      VIA 5.748 25.65 Element_VIA34_1_2_58_52 ;
      VIA 5.748 25.65 Element_VIA23_1_3_36_36 ;
      VIA 5.748 25.11 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 25.093 5.793 25.127 ;
      VIA 5.748 25.11 Element_VIA34_1_2_58_52 ;
      VIA 5.748 25.11 Element_VIA23_1_3_36_36 ;
      VIA 5.748 24.57 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 24.553 5.793 24.587 ;
      VIA 5.748 24.57 Element_VIA34_1_2_58_52 ;
      VIA 5.748 24.57 Element_VIA23_1_3_36_36 ;
      VIA 5.748 24.03 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 24.013 5.793 24.047 ;
      VIA 5.748 24.03 Element_VIA34_1_2_58_52 ;
      VIA 5.748 24.03 Element_VIA23_1_3_36_36 ;
      VIA 5.748 23.49 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 23.473 5.793 23.507 ;
      VIA 5.748 23.49 Element_VIA34_1_2_58_52 ;
      VIA 5.748 23.49 Element_VIA23_1_3_36_36 ;
      VIA 5.748 22.95 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 22.933 5.793 22.967 ;
      VIA 5.748 22.95 Element_VIA34_1_2_58_52 ;
      VIA 5.748 22.95 Element_VIA23_1_3_36_36 ;
      VIA 5.748 22.41 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 22.393 5.793 22.427 ;
      VIA 5.748 22.41 Element_VIA34_1_2_58_52 ;
      VIA 5.748 22.41 Element_VIA23_1_3_36_36 ;
      VIA 5.748 21.87 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 21.853 5.793 21.887 ;
      VIA 5.748 21.87 Element_VIA34_1_2_58_52 ;
      VIA 5.748 21.87 Element_VIA23_1_3_36_36 ;
      VIA 5.748 21.33 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 21.313 5.793 21.347 ;
      VIA 5.748 21.33 Element_VIA34_1_2_58_52 ;
      VIA 5.748 21.33 Element_VIA23_1_3_36_36 ;
      VIA 5.748 20.79 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 20.773 5.793 20.807 ;
      VIA 5.748 20.79 Element_VIA34_1_2_58_52 ;
      VIA 5.748 20.79 Element_VIA23_1_3_36_36 ;
      VIA 5.748 20.25 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 20.233 5.793 20.267 ;
      VIA 5.748 20.25 Element_VIA34_1_2_58_52 ;
      VIA 5.748 20.25 Element_VIA23_1_3_36_36 ;
      VIA 5.748 19.71 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 19.693 5.793 19.727 ;
      VIA 5.748 19.71 Element_VIA34_1_2_58_52 ;
      VIA 5.748 19.71 Element_VIA23_1_3_36_36 ;
      VIA 5.748 19.17 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 19.153 5.793 19.187 ;
      VIA 5.748 19.17 Element_VIA34_1_2_58_52 ;
      VIA 5.748 19.17 Element_VIA23_1_3_36_36 ;
      VIA 5.748 18.63 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 18.613 5.793 18.647 ;
      VIA 5.748 18.63 Element_VIA34_1_2_58_52 ;
      VIA 5.748 18.63 Element_VIA23_1_3_36_36 ;
      VIA 5.748 18.09 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 18.073 5.793 18.107 ;
      VIA 5.748 18.09 Element_VIA34_1_2_58_52 ;
      VIA 5.748 18.09 Element_VIA23_1_3_36_36 ;
      VIA 5.748 17.55 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 17.533 5.793 17.567 ;
      VIA 5.748 17.55 Element_VIA34_1_2_58_52 ;
      VIA 5.748 17.55 Element_VIA23_1_3_36_36 ;
      VIA 5.748 17.01 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 16.993 5.793 17.027 ;
      VIA 5.748 17.01 Element_VIA34_1_2_58_52 ;
      VIA 5.748 17.01 Element_VIA23_1_3_36_36 ;
      VIA 5.748 16.47 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 16.453 5.793 16.487 ;
      VIA 5.748 16.47 Element_VIA34_1_2_58_52 ;
      VIA 5.748 16.47 Element_VIA23_1_3_36_36 ;
      VIA 5.748 15.93 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 15.913 5.793 15.947 ;
      VIA 5.748 15.93 Element_VIA34_1_2_58_52 ;
      VIA 5.748 15.93 Element_VIA23_1_3_36_36 ;
      VIA 5.748 15.39 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 15.373 5.793 15.407 ;
      VIA 5.748 15.39 Element_VIA34_1_2_58_52 ;
      VIA 5.748 15.39 Element_VIA23_1_3_36_36 ;
      VIA 5.748 14.85 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 14.833 5.793 14.867 ;
      VIA 5.748 14.85 Element_VIA34_1_2_58_52 ;
      VIA 5.748 14.85 Element_VIA23_1_3_36_36 ;
      VIA 5.748 14.31 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 14.293 5.793 14.327 ;
      VIA 5.748 14.31 Element_VIA34_1_2_58_52 ;
      VIA 5.748 14.31 Element_VIA23_1_3_36_36 ;
      VIA 5.748 13.77 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 13.753 5.793 13.787 ;
      VIA 5.748 13.77 Element_VIA34_1_2_58_52 ;
      VIA 5.748 13.77 Element_VIA23_1_3_36_36 ;
      VIA 5.748 13.23 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 13.213 5.793 13.247 ;
      VIA 5.748 13.23 Element_VIA34_1_2_58_52 ;
      VIA 5.748 13.23 Element_VIA23_1_3_36_36 ;
      VIA 5.748 12.69 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 12.673 5.793 12.707 ;
      VIA 5.748 12.69 Element_VIA34_1_2_58_52 ;
      VIA 5.748 12.69 Element_VIA23_1_3_36_36 ;
      VIA 5.748 12.15 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 12.133 5.793 12.167 ;
      VIA 5.748 12.15 Element_VIA34_1_2_58_52 ;
      VIA 5.748 12.15 Element_VIA23_1_3_36_36 ;
      VIA 5.748 11.61 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 11.593 5.793 11.627 ;
      VIA 5.748 11.61 Element_VIA34_1_2_58_52 ;
      VIA 5.748 11.61 Element_VIA23_1_3_36_36 ;
      VIA 5.748 11.07 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 11.053 5.793 11.087 ;
      VIA 5.748 11.07 Element_VIA34_1_2_58_52 ;
      VIA 5.748 11.07 Element_VIA23_1_3_36_36 ;
      VIA 5.748 10.53 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 10.513 5.793 10.547 ;
      VIA 5.748 10.53 Element_VIA34_1_2_58_52 ;
      VIA 5.748 10.53 Element_VIA23_1_3_36_36 ;
      VIA 5.748 9.99 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 9.973 5.793 10.007 ;
      VIA 5.748 9.99 Element_VIA34_1_2_58_52 ;
      VIA 5.748 9.99 Element_VIA23_1_3_36_36 ;
      VIA 5.748 9.45 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 9.433 5.793 9.467 ;
      VIA 5.748 9.45 Element_VIA34_1_2_58_52 ;
      VIA 5.748 9.45 Element_VIA23_1_3_36_36 ;
      VIA 5.748 8.91 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 8.893 5.793 8.927 ;
      VIA 5.748 8.91 Element_VIA34_1_2_58_52 ;
      VIA 5.748 8.91 Element_VIA23_1_3_36_36 ;
      VIA 5.748 8.37 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 8.353 5.793 8.387 ;
      VIA 5.748 8.37 Element_VIA34_1_2_58_52 ;
      VIA 5.748 8.37 Element_VIA23_1_3_36_36 ;
      VIA 5.748 7.83 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 7.813 5.793 7.847 ;
      VIA 5.748 7.83 Element_VIA34_1_2_58_52 ;
      VIA 5.748 7.83 Element_VIA23_1_3_36_36 ;
      VIA 5.748 7.29 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 7.273 5.793 7.307 ;
      VIA 5.748 7.29 Element_VIA34_1_2_58_52 ;
      VIA 5.748 7.29 Element_VIA23_1_3_36_36 ;
      VIA 5.748 6.75 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 6.733 5.793 6.767 ;
      VIA 5.748 6.75 Element_VIA34_1_2_58_52 ;
      VIA 5.748 6.75 Element_VIA23_1_3_36_36 ;
      VIA 5.748 6.21 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 6.193 5.793 6.227 ;
      VIA 5.748 6.21 Element_VIA34_1_2_58_52 ;
      VIA 5.748 6.21 Element_VIA23_1_3_36_36 ;
      VIA 5.748 5.67 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 5.653 5.793 5.687 ;
      VIA 5.748 5.67 Element_VIA34_1_2_58_52 ;
      VIA 5.748 5.67 Element_VIA23_1_3_36_36 ;
      VIA 5.748 5.13 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 5.113 5.793 5.147 ;
      VIA 5.748 5.13 Element_VIA34_1_2_58_52 ;
      VIA 5.748 5.13 Element_VIA23_1_3_36_36 ;
      VIA 5.748 4.59 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 4.573 5.793 4.607 ;
      VIA 5.748 4.59 Element_VIA34_1_2_58_52 ;
      VIA 5.748 4.59 Element_VIA23_1_3_36_36 ;
      VIA 5.748 4.05 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 4.033 5.793 4.067 ;
      VIA 5.748 4.05 Element_VIA34_1_2_58_52 ;
      VIA 5.748 4.05 Element_VIA23_1_3_36_36 ;
      VIA 5.748 3.51 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 3.493 5.793 3.527 ;
      VIA 5.748 3.51 Element_VIA34_1_2_58_52 ;
      VIA 5.748 3.51 Element_VIA23_1_3_36_36 ;
      VIA 5.748 2.97 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 2.953 5.793 2.987 ;
      VIA 5.748 2.97 Element_VIA34_1_2_58_52 ;
      VIA 5.748 2.97 Element_VIA23_1_3_36_36 ;
      VIA 5.748 2.43 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 2.413 5.793 2.447 ;
      VIA 5.748 2.43 Element_VIA34_1_2_58_52 ;
      VIA 5.748 2.43 Element_VIA23_1_3_36_36 ;
      VIA 5.748 1.89 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 1.873 5.793 1.907 ;
      VIA 5.748 1.89 Element_VIA34_1_2_58_52 ;
      VIA 5.748 1.89 Element_VIA23_1_3_36_36 ;
      VIA 5.748 1.35 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.703 1.333 5.793 1.367 ;
      VIA 5.748 1.35 Element_VIA34_1_2_58_52 ;
      VIA 5.748 1.35 Element_VIA23_1_3_36_36 ;
      VIA 2.772 41.85 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 41.833 2.817 41.867 ;
      VIA 2.772 41.85 Element_VIA34_1_2_58_52 ;
      VIA 2.772 41.85 Element_VIA23_1_3_36_36 ;
      VIA 2.772 41.31 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 41.293 2.817 41.327 ;
      VIA 2.772 41.31 Element_VIA34_1_2_58_52 ;
      VIA 2.772 41.31 Element_VIA23_1_3_36_36 ;
      VIA 2.772 40.77 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 40.753 2.817 40.787 ;
      VIA 2.772 40.77 Element_VIA34_1_2_58_52 ;
      VIA 2.772 40.77 Element_VIA23_1_3_36_36 ;
      VIA 2.772 40.23 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 40.213 2.817 40.247 ;
      VIA 2.772 40.23 Element_VIA34_1_2_58_52 ;
      VIA 2.772 40.23 Element_VIA23_1_3_36_36 ;
      VIA 2.772 39.69 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 39.673 2.817 39.707 ;
      VIA 2.772 39.69 Element_VIA34_1_2_58_52 ;
      VIA 2.772 39.69 Element_VIA23_1_3_36_36 ;
      VIA 2.772 39.15 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 39.133 2.817 39.167 ;
      VIA 2.772 39.15 Element_VIA34_1_2_58_52 ;
      VIA 2.772 39.15 Element_VIA23_1_3_36_36 ;
      VIA 2.772 38.61 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 38.593 2.817 38.627 ;
      VIA 2.772 38.61 Element_VIA34_1_2_58_52 ;
      VIA 2.772 38.61 Element_VIA23_1_3_36_36 ;
      VIA 2.772 38.07 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 38.053 2.817 38.087 ;
      VIA 2.772 38.07 Element_VIA34_1_2_58_52 ;
      VIA 2.772 38.07 Element_VIA23_1_3_36_36 ;
      VIA 2.772 37.53 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 37.513 2.817 37.547 ;
      VIA 2.772 37.53 Element_VIA34_1_2_58_52 ;
      VIA 2.772 37.53 Element_VIA23_1_3_36_36 ;
      VIA 2.772 36.99 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 36.973 2.817 37.007 ;
      VIA 2.772 36.99 Element_VIA34_1_2_58_52 ;
      VIA 2.772 36.99 Element_VIA23_1_3_36_36 ;
      VIA 2.772 36.45 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 36.433 2.817 36.467 ;
      VIA 2.772 36.45 Element_VIA34_1_2_58_52 ;
      VIA 2.772 36.45 Element_VIA23_1_3_36_36 ;
      VIA 2.772 35.91 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 35.893 2.817 35.927 ;
      VIA 2.772 35.91 Element_VIA34_1_2_58_52 ;
      VIA 2.772 35.91 Element_VIA23_1_3_36_36 ;
      VIA 2.772 35.37 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 35.353 2.817 35.387 ;
      VIA 2.772 35.37 Element_VIA34_1_2_58_52 ;
      VIA 2.772 35.37 Element_VIA23_1_3_36_36 ;
      VIA 2.772 34.83 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 34.813 2.817 34.847 ;
      VIA 2.772 34.83 Element_VIA34_1_2_58_52 ;
      VIA 2.772 34.83 Element_VIA23_1_3_36_36 ;
      VIA 2.772 34.29 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 34.273 2.817 34.307 ;
      VIA 2.772 34.29 Element_VIA34_1_2_58_52 ;
      VIA 2.772 34.29 Element_VIA23_1_3_36_36 ;
      VIA 2.772 33.75 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 33.733 2.817 33.767 ;
      VIA 2.772 33.75 Element_VIA34_1_2_58_52 ;
      VIA 2.772 33.75 Element_VIA23_1_3_36_36 ;
      VIA 2.772 33.21 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 33.193 2.817 33.227 ;
      VIA 2.772 33.21 Element_VIA34_1_2_58_52 ;
      VIA 2.772 33.21 Element_VIA23_1_3_36_36 ;
      VIA 2.772 32.67 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 32.653 2.817 32.687 ;
      VIA 2.772 32.67 Element_VIA34_1_2_58_52 ;
      VIA 2.772 32.67 Element_VIA23_1_3_36_36 ;
      VIA 2.772 32.13 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 32.113 2.817 32.147 ;
      VIA 2.772 32.13 Element_VIA34_1_2_58_52 ;
      VIA 2.772 32.13 Element_VIA23_1_3_36_36 ;
      VIA 2.772 31.59 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 31.573 2.817 31.607 ;
      VIA 2.772 31.59 Element_VIA34_1_2_58_52 ;
      VIA 2.772 31.59 Element_VIA23_1_3_36_36 ;
      VIA 2.772 31.05 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 31.033 2.817 31.067 ;
      VIA 2.772 31.05 Element_VIA34_1_2_58_52 ;
      VIA 2.772 31.05 Element_VIA23_1_3_36_36 ;
      VIA 2.772 30.51 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 30.493 2.817 30.527 ;
      VIA 2.772 30.51 Element_VIA34_1_2_58_52 ;
      VIA 2.772 30.51 Element_VIA23_1_3_36_36 ;
      VIA 2.772 29.97 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 29.953 2.817 29.987 ;
      VIA 2.772 29.97 Element_VIA34_1_2_58_52 ;
      VIA 2.772 29.97 Element_VIA23_1_3_36_36 ;
      VIA 2.772 29.43 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 29.413 2.817 29.447 ;
      VIA 2.772 29.43 Element_VIA34_1_2_58_52 ;
      VIA 2.772 29.43 Element_VIA23_1_3_36_36 ;
      VIA 2.772 28.89 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 28.873 2.817 28.907 ;
      VIA 2.772 28.89 Element_VIA34_1_2_58_52 ;
      VIA 2.772 28.89 Element_VIA23_1_3_36_36 ;
      VIA 2.772 28.35 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 28.333 2.817 28.367 ;
      VIA 2.772 28.35 Element_VIA34_1_2_58_52 ;
      VIA 2.772 28.35 Element_VIA23_1_3_36_36 ;
      VIA 2.772 27.81 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 27.793 2.817 27.827 ;
      VIA 2.772 27.81 Element_VIA34_1_2_58_52 ;
      VIA 2.772 27.81 Element_VIA23_1_3_36_36 ;
      VIA 2.772 27.27 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 27.253 2.817 27.287 ;
      VIA 2.772 27.27 Element_VIA34_1_2_58_52 ;
      VIA 2.772 27.27 Element_VIA23_1_3_36_36 ;
      VIA 2.772 26.73 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 26.713 2.817 26.747 ;
      VIA 2.772 26.73 Element_VIA34_1_2_58_52 ;
      VIA 2.772 26.73 Element_VIA23_1_3_36_36 ;
      VIA 2.772 26.19 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 26.173 2.817 26.207 ;
      VIA 2.772 26.19 Element_VIA34_1_2_58_52 ;
      VIA 2.772 26.19 Element_VIA23_1_3_36_36 ;
      VIA 2.772 25.65 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 25.633 2.817 25.667 ;
      VIA 2.772 25.65 Element_VIA34_1_2_58_52 ;
      VIA 2.772 25.65 Element_VIA23_1_3_36_36 ;
      VIA 2.772 25.11 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 25.093 2.817 25.127 ;
      VIA 2.772 25.11 Element_VIA34_1_2_58_52 ;
      VIA 2.772 25.11 Element_VIA23_1_3_36_36 ;
      VIA 2.772 24.57 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 24.553 2.817 24.587 ;
      VIA 2.772 24.57 Element_VIA34_1_2_58_52 ;
      VIA 2.772 24.57 Element_VIA23_1_3_36_36 ;
      VIA 2.772 24.03 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 24.013 2.817 24.047 ;
      VIA 2.772 24.03 Element_VIA34_1_2_58_52 ;
      VIA 2.772 24.03 Element_VIA23_1_3_36_36 ;
      VIA 2.772 23.49 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 23.473 2.817 23.507 ;
      VIA 2.772 23.49 Element_VIA34_1_2_58_52 ;
      VIA 2.772 23.49 Element_VIA23_1_3_36_36 ;
      VIA 2.772 22.95 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 22.933 2.817 22.967 ;
      VIA 2.772 22.95 Element_VIA34_1_2_58_52 ;
      VIA 2.772 22.95 Element_VIA23_1_3_36_36 ;
      VIA 2.772 22.41 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 22.393 2.817 22.427 ;
      VIA 2.772 22.41 Element_VIA34_1_2_58_52 ;
      VIA 2.772 22.41 Element_VIA23_1_3_36_36 ;
      VIA 2.772 21.87 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 21.853 2.817 21.887 ;
      VIA 2.772 21.87 Element_VIA34_1_2_58_52 ;
      VIA 2.772 21.87 Element_VIA23_1_3_36_36 ;
      VIA 2.772 21.33 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 21.313 2.817 21.347 ;
      VIA 2.772 21.33 Element_VIA34_1_2_58_52 ;
      VIA 2.772 21.33 Element_VIA23_1_3_36_36 ;
      VIA 2.772 20.79 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 20.773 2.817 20.807 ;
      VIA 2.772 20.79 Element_VIA34_1_2_58_52 ;
      VIA 2.772 20.79 Element_VIA23_1_3_36_36 ;
      VIA 2.772 20.25 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 20.233 2.817 20.267 ;
      VIA 2.772 20.25 Element_VIA34_1_2_58_52 ;
      VIA 2.772 20.25 Element_VIA23_1_3_36_36 ;
      VIA 2.772 19.71 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 19.693 2.817 19.727 ;
      VIA 2.772 19.71 Element_VIA34_1_2_58_52 ;
      VIA 2.772 19.71 Element_VIA23_1_3_36_36 ;
      VIA 2.772 19.17 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 19.153 2.817 19.187 ;
      VIA 2.772 19.17 Element_VIA34_1_2_58_52 ;
      VIA 2.772 19.17 Element_VIA23_1_3_36_36 ;
      VIA 2.772 18.63 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 18.613 2.817 18.647 ;
      VIA 2.772 18.63 Element_VIA34_1_2_58_52 ;
      VIA 2.772 18.63 Element_VIA23_1_3_36_36 ;
      VIA 2.772 18.09 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 18.073 2.817 18.107 ;
      VIA 2.772 18.09 Element_VIA34_1_2_58_52 ;
      VIA 2.772 18.09 Element_VIA23_1_3_36_36 ;
      VIA 2.772 17.55 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 17.533 2.817 17.567 ;
      VIA 2.772 17.55 Element_VIA34_1_2_58_52 ;
      VIA 2.772 17.55 Element_VIA23_1_3_36_36 ;
      VIA 2.772 17.01 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 16.993 2.817 17.027 ;
      VIA 2.772 17.01 Element_VIA34_1_2_58_52 ;
      VIA 2.772 17.01 Element_VIA23_1_3_36_36 ;
      VIA 2.772 16.47 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 16.453 2.817 16.487 ;
      VIA 2.772 16.47 Element_VIA34_1_2_58_52 ;
      VIA 2.772 16.47 Element_VIA23_1_3_36_36 ;
      VIA 2.772 15.93 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 15.913 2.817 15.947 ;
      VIA 2.772 15.93 Element_VIA34_1_2_58_52 ;
      VIA 2.772 15.93 Element_VIA23_1_3_36_36 ;
      VIA 2.772 15.39 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 15.373 2.817 15.407 ;
      VIA 2.772 15.39 Element_VIA34_1_2_58_52 ;
      VIA 2.772 15.39 Element_VIA23_1_3_36_36 ;
      VIA 2.772 14.85 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 14.833 2.817 14.867 ;
      VIA 2.772 14.85 Element_VIA34_1_2_58_52 ;
      VIA 2.772 14.85 Element_VIA23_1_3_36_36 ;
      VIA 2.772 14.31 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 14.293 2.817 14.327 ;
      VIA 2.772 14.31 Element_VIA34_1_2_58_52 ;
      VIA 2.772 14.31 Element_VIA23_1_3_36_36 ;
      VIA 2.772 13.77 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 13.753 2.817 13.787 ;
      VIA 2.772 13.77 Element_VIA34_1_2_58_52 ;
      VIA 2.772 13.77 Element_VIA23_1_3_36_36 ;
      VIA 2.772 13.23 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 13.213 2.817 13.247 ;
      VIA 2.772 13.23 Element_VIA34_1_2_58_52 ;
      VIA 2.772 13.23 Element_VIA23_1_3_36_36 ;
      VIA 2.772 12.69 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 12.673 2.817 12.707 ;
      VIA 2.772 12.69 Element_VIA34_1_2_58_52 ;
      VIA 2.772 12.69 Element_VIA23_1_3_36_36 ;
      VIA 2.772 12.15 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 12.133 2.817 12.167 ;
      VIA 2.772 12.15 Element_VIA34_1_2_58_52 ;
      VIA 2.772 12.15 Element_VIA23_1_3_36_36 ;
      VIA 2.772 11.61 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 11.593 2.817 11.627 ;
      VIA 2.772 11.61 Element_VIA34_1_2_58_52 ;
      VIA 2.772 11.61 Element_VIA23_1_3_36_36 ;
      VIA 2.772 11.07 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 11.053 2.817 11.087 ;
      VIA 2.772 11.07 Element_VIA34_1_2_58_52 ;
      VIA 2.772 11.07 Element_VIA23_1_3_36_36 ;
      VIA 2.772 10.53 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 10.513 2.817 10.547 ;
      VIA 2.772 10.53 Element_VIA34_1_2_58_52 ;
      VIA 2.772 10.53 Element_VIA23_1_3_36_36 ;
      VIA 2.772 9.99 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 9.973 2.817 10.007 ;
      VIA 2.772 9.99 Element_VIA34_1_2_58_52 ;
      VIA 2.772 9.99 Element_VIA23_1_3_36_36 ;
      VIA 2.772 9.45 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 9.433 2.817 9.467 ;
      VIA 2.772 9.45 Element_VIA34_1_2_58_52 ;
      VIA 2.772 9.45 Element_VIA23_1_3_36_36 ;
      VIA 2.772 8.91 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 8.893 2.817 8.927 ;
      VIA 2.772 8.91 Element_VIA34_1_2_58_52 ;
      VIA 2.772 8.91 Element_VIA23_1_3_36_36 ;
      VIA 2.772 8.37 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 8.353 2.817 8.387 ;
      VIA 2.772 8.37 Element_VIA34_1_2_58_52 ;
      VIA 2.772 8.37 Element_VIA23_1_3_36_36 ;
      VIA 2.772 7.83 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 7.813 2.817 7.847 ;
      VIA 2.772 7.83 Element_VIA34_1_2_58_52 ;
      VIA 2.772 7.83 Element_VIA23_1_3_36_36 ;
      VIA 2.772 7.29 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 7.273 2.817 7.307 ;
      VIA 2.772 7.29 Element_VIA34_1_2_58_52 ;
      VIA 2.772 7.29 Element_VIA23_1_3_36_36 ;
      VIA 2.772 6.75 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 6.733 2.817 6.767 ;
      VIA 2.772 6.75 Element_VIA34_1_2_58_52 ;
      VIA 2.772 6.75 Element_VIA23_1_3_36_36 ;
      VIA 2.772 6.21 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 6.193 2.817 6.227 ;
      VIA 2.772 6.21 Element_VIA34_1_2_58_52 ;
      VIA 2.772 6.21 Element_VIA23_1_3_36_36 ;
      VIA 2.772 5.67 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 5.653 2.817 5.687 ;
      VIA 2.772 5.67 Element_VIA34_1_2_58_52 ;
      VIA 2.772 5.67 Element_VIA23_1_3_36_36 ;
      VIA 2.772 5.13 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 5.113 2.817 5.147 ;
      VIA 2.772 5.13 Element_VIA34_1_2_58_52 ;
      VIA 2.772 5.13 Element_VIA23_1_3_36_36 ;
      VIA 2.772 4.59 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 4.573 2.817 4.607 ;
      VIA 2.772 4.59 Element_VIA34_1_2_58_52 ;
      VIA 2.772 4.59 Element_VIA23_1_3_36_36 ;
      VIA 2.772 4.05 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 4.033 2.817 4.067 ;
      VIA 2.772 4.05 Element_VIA34_1_2_58_52 ;
      VIA 2.772 4.05 Element_VIA23_1_3_36_36 ;
      VIA 2.772 3.51 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 3.493 2.817 3.527 ;
      VIA 2.772 3.51 Element_VIA34_1_2_58_52 ;
      VIA 2.772 3.51 Element_VIA23_1_3_36_36 ;
      VIA 2.772 2.97 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 2.953 2.817 2.987 ;
      VIA 2.772 2.97 Element_VIA34_1_2_58_52 ;
      VIA 2.772 2.97 Element_VIA23_1_3_36_36 ;
      VIA 2.772 2.43 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 2.413 2.817 2.447 ;
      VIA 2.772 2.43 Element_VIA34_1_2_58_52 ;
      VIA 2.772 2.43 Element_VIA23_1_3_36_36 ;
      VIA 2.772 1.89 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 1.873 2.817 1.907 ;
      VIA 2.772 1.89 Element_VIA34_1_2_58_52 ;
      VIA 2.772 1.89 Element_VIA23_1_3_36_36 ;
      VIA 2.772 1.35 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.727 1.333 2.817 1.367 ;
      VIA 2.772 1.35 Element_VIA34_1_2_58_52 ;
      VIA 2.772 1.35 Element_VIA23_1_3_36_36 ;
      VIA 21.6 41.85 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 41.31 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 40.77 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 40.23 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 39.69 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 39.15 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 38.61 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 38.07 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 37.53 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 36.99 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 36.45 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 35.91 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 35.37 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 34.83 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 34.29 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 33.75 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 33.21 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 32.67 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 32.13 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 31.59 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 31.05 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 30.51 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 29.97 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 29.43 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 28.89 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 28.35 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 27.81 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 27.27 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 26.73 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 26.19 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 25.65 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 25.11 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 24.57 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 24.03 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 23.49 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 22.95 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 22.41 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 21.87 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 21.33 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 20.79 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 20.25 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 19.71 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 19.17 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 18.63 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 18.09 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 17.55 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 17.01 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 16.47 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 15.93 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 15.39 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 14.85 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 14.31 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 13.77 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 13.23 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 12.69 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 12.15 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 11.61 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 11.07 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 10.53 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 9.99 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 9.45 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 8.91 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 8.37 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 7.83 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 7.29 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 6.75 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 6.21 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 5.67 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 5.13 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 4.59 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 4.05 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 3.51 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 2.97 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 2.43 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 1.89 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 1.35 Element_via1_2_41040_18_1_1140_36_36 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER M5 ;
        RECT  41.208 0.876 41.328 42.324 ;
        RECT  38.232 0.876 38.352 42.324 ;
        RECT  35.256 0.876 35.376 42.324 ;
        RECT  32.28 0.876 32.4 42.324 ;
        RECT  29.304 0.876 29.424 42.324 ;
        RECT  26.328 0.876 26.448 42.324 ;
        RECT  23.352 0.876 23.472 42.324 ;
        RECT  20.376 0.876 20.496 42.324 ;
        RECT  17.4 0.876 17.52 42.324 ;
        RECT  14.424 0.876 14.544 42.324 ;
        RECT  11.448 0.876 11.568 42.324 ;
        RECT  8.472 0.876 8.592 42.324 ;
        RECT  5.496 0.876 5.616 42.324 ;
        RECT  2.52 0.876 2.64 42.324 ;
      LAYER M2 ;
        RECT  1.08 42.111 42.12 42.129 ;
        RECT  1.08 41.571 42.12 41.589 ;
        RECT  1.08 41.031 42.12 41.049 ;
        RECT  1.08 40.491 42.12 40.509 ;
        RECT  1.08 39.951 42.12 39.969 ;
        RECT  1.08 39.411 42.12 39.429 ;
        RECT  1.08 38.871 42.12 38.889 ;
        RECT  1.08 38.331 42.12 38.349 ;
        RECT  1.08 37.791 42.12 37.809 ;
        RECT  1.08 37.251 42.12 37.269 ;
        RECT  1.08 36.711 42.12 36.729 ;
        RECT  1.08 36.171 42.12 36.189 ;
        RECT  1.08 35.631 42.12 35.649 ;
        RECT  1.08 35.091 42.12 35.109 ;
        RECT  1.08 34.551 42.12 34.569 ;
        RECT  1.08 34.011 42.12 34.029 ;
        RECT  1.08 33.471 42.12 33.489 ;
        RECT  1.08 32.931 42.12 32.949 ;
        RECT  1.08 32.391 42.12 32.409 ;
        RECT  1.08 31.851 42.12 31.869 ;
        RECT  1.08 31.311 42.12 31.329 ;
        RECT  1.08 30.771 42.12 30.789 ;
        RECT  1.08 30.231 42.12 30.249 ;
        RECT  1.08 29.691 42.12 29.709 ;
        RECT  1.08 29.151 42.12 29.169 ;
        RECT  1.08 28.611 42.12 28.629 ;
        RECT  1.08 28.071 42.12 28.089 ;
        RECT  1.08 27.531 42.12 27.549 ;
        RECT  1.08 26.991 42.12 27.009 ;
        RECT  1.08 26.451 42.12 26.469 ;
        RECT  1.08 25.911 42.12 25.929 ;
        RECT  1.08 25.371 42.12 25.389 ;
        RECT  1.08 24.831 42.12 24.849 ;
        RECT  1.08 24.291 42.12 24.309 ;
        RECT  1.08 23.751 42.12 23.769 ;
        RECT  1.08 23.211 42.12 23.229 ;
        RECT  1.08 22.671 42.12 22.689 ;
        RECT  1.08 22.131 42.12 22.149 ;
        RECT  1.08 21.591 42.12 21.609 ;
        RECT  1.08 21.051 42.12 21.069 ;
        RECT  1.08 20.511 42.12 20.529 ;
        RECT  1.08 19.971 42.12 19.989 ;
        RECT  1.08 19.431 42.12 19.449 ;
        RECT  1.08 18.891 42.12 18.909 ;
        RECT  1.08 18.351 42.12 18.369 ;
        RECT  1.08 17.811 42.12 17.829 ;
        RECT  1.08 17.271 42.12 17.289 ;
        RECT  1.08 16.731 42.12 16.749 ;
        RECT  1.08 16.191 42.12 16.209 ;
        RECT  1.08 15.651 42.12 15.669 ;
        RECT  1.08 15.111 42.12 15.129 ;
        RECT  1.08 14.571 42.12 14.589 ;
        RECT  1.08 14.031 42.12 14.049 ;
        RECT  1.08 13.491 42.12 13.509 ;
        RECT  1.08 12.951 42.12 12.969 ;
        RECT  1.08 12.411 42.12 12.429 ;
        RECT  1.08 11.871 42.12 11.889 ;
        RECT  1.08 11.331 42.12 11.349 ;
        RECT  1.08 10.791 42.12 10.809 ;
        RECT  1.08 10.251 42.12 10.269 ;
        RECT  1.08 9.711 42.12 9.729 ;
        RECT  1.08 9.171 42.12 9.189 ;
        RECT  1.08 8.631 42.12 8.649 ;
        RECT  1.08 8.091 42.12 8.109 ;
        RECT  1.08 7.551 42.12 7.569 ;
        RECT  1.08 7.011 42.12 7.029 ;
        RECT  1.08 6.471 42.12 6.489 ;
        RECT  1.08 5.931 42.12 5.949 ;
        RECT  1.08 5.391 42.12 5.409 ;
        RECT  1.08 4.851 42.12 4.869 ;
        RECT  1.08 4.311 42.12 4.329 ;
        RECT  1.08 3.771 42.12 3.789 ;
        RECT  1.08 3.231 42.12 3.249 ;
        RECT  1.08 2.691 42.12 2.709 ;
        RECT  1.08 2.151 42.12 2.169 ;
        RECT  1.08 1.611 42.12 1.629 ;
        RECT  1.08 1.071 42.12 1.089 ;
      LAYER M1 ;
        RECT  1.08 42.111 42.12 42.129 ;
        RECT  1.08 41.571 42.12 41.589 ;
        RECT  1.08 41.031 42.12 41.049 ;
        RECT  1.08 40.491 42.12 40.509 ;
        RECT  1.08 39.951 42.12 39.969 ;
        RECT  1.08 39.411 42.12 39.429 ;
        RECT  1.08 38.871 42.12 38.889 ;
        RECT  1.08 38.331 42.12 38.349 ;
        RECT  1.08 37.791 42.12 37.809 ;
        RECT  1.08 37.251 42.12 37.269 ;
        RECT  1.08 36.711 42.12 36.729 ;
        RECT  1.08 36.171 42.12 36.189 ;
        RECT  1.08 35.631 42.12 35.649 ;
        RECT  1.08 35.091 42.12 35.109 ;
        RECT  1.08 34.551 42.12 34.569 ;
        RECT  1.08 34.011 42.12 34.029 ;
        RECT  1.08 33.471 42.12 33.489 ;
        RECT  1.08 32.931 42.12 32.949 ;
        RECT  1.08 32.391 42.12 32.409 ;
        RECT  1.08 31.851 42.12 31.869 ;
        RECT  1.08 31.311 42.12 31.329 ;
        RECT  1.08 30.771 42.12 30.789 ;
        RECT  1.08 30.231 42.12 30.249 ;
        RECT  1.08 29.691 42.12 29.709 ;
        RECT  1.08 29.151 42.12 29.169 ;
        RECT  1.08 28.611 42.12 28.629 ;
        RECT  1.08 28.071 42.12 28.089 ;
        RECT  1.08 27.531 42.12 27.549 ;
        RECT  1.08 26.991 42.12 27.009 ;
        RECT  1.08 26.451 42.12 26.469 ;
        RECT  1.08 25.911 42.12 25.929 ;
        RECT  1.08 25.371 42.12 25.389 ;
        RECT  1.08 24.831 42.12 24.849 ;
        RECT  1.08 24.291 42.12 24.309 ;
        RECT  1.08 23.751 42.12 23.769 ;
        RECT  1.08 23.211 42.12 23.229 ;
        RECT  1.08 22.671 42.12 22.689 ;
        RECT  1.08 22.131 42.12 22.149 ;
        RECT  1.08 21.591 42.12 21.609 ;
        RECT  1.08 21.051 42.12 21.069 ;
        RECT  1.08 20.511 42.12 20.529 ;
        RECT  1.08 19.971 42.12 19.989 ;
        RECT  1.08 19.431 42.12 19.449 ;
        RECT  1.08 18.891 42.12 18.909 ;
        RECT  1.08 18.351 42.12 18.369 ;
        RECT  1.08 17.811 42.12 17.829 ;
        RECT  1.08 17.271 42.12 17.289 ;
        RECT  1.08 16.731 42.12 16.749 ;
        RECT  1.08 16.191 42.12 16.209 ;
        RECT  1.08 15.651 42.12 15.669 ;
        RECT  1.08 15.111 42.12 15.129 ;
        RECT  1.08 14.571 42.12 14.589 ;
        RECT  1.08 14.031 42.12 14.049 ;
        RECT  1.08 13.491 42.12 13.509 ;
        RECT  1.08 12.951 42.12 12.969 ;
        RECT  1.08 12.411 42.12 12.429 ;
        RECT  1.08 11.871 42.12 11.889 ;
        RECT  1.08 11.331 42.12 11.349 ;
        RECT  1.08 10.791 42.12 10.809 ;
        RECT  1.08 10.251 42.12 10.269 ;
        RECT  1.08 9.711 42.12 9.729 ;
        RECT  1.08 9.171 42.12 9.189 ;
        RECT  1.08 8.631 42.12 8.649 ;
        RECT  1.08 8.091 42.12 8.109 ;
        RECT  1.08 7.551 42.12 7.569 ;
        RECT  1.08 7.011 42.12 7.029 ;
        RECT  1.08 6.471 42.12 6.489 ;
        RECT  1.08 5.931 42.12 5.949 ;
        RECT  1.08 5.391 42.12 5.409 ;
        RECT  1.08 4.851 42.12 4.869 ;
        RECT  1.08 4.311 42.12 4.329 ;
        RECT  1.08 3.771 42.12 3.789 ;
        RECT  1.08 3.231 42.12 3.249 ;
        RECT  1.08 2.691 42.12 2.709 ;
        RECT  1.08 2.151 42.12 2.169 ;
        RECT  1.08 1.611 42.12 1.629 ;
        RECT  1.08 1.071 42.12 1.089 ;
      LAYER M5 ;
        RECT  42.204 0.876 42.324 42.324 ;
      LAYER M4 ;
        RECT  0.876 42.204 42.324 42.324 ;
        RECT  0.876 0.876 42.324 0.996 ;
      LAYER M5 ;
        RECT  0.876 0.876 0.996 42.324 ;
      VIA 42.264 42.264 Element_VIA45_2_2_58_58 ;
      VIA 42.264 0.936 Element_VIA45_2_2_58_58 ;
      VIA 41.268 42.264 Element_VIA45_2_2_58_58 ;
      VIA 41.268 0.936 Element_VIA45_2_2_58_58 ;
      VIA 38.292 42.264 Element_VIA45_2_2_58_58 ;
      VIA 38.292 0.936 Element_VIA45_2_2_58_58 ;
      VIA 35.316 42.264 Element_VIA45_2_2_58_58 ;
      VIA 35.316 0.936 Element_VIA45_2_2_58_58 ;
      VIA 32.34 42.264 Element_VIA45_2_2_58_58 ;
      VIA 32.34 0.936 Element_VIA45_2_2_58_58 ;
      VIA 29.364 42.264 Element_VIA45_2_2_58_58 ;
      VIA 29.364 0.936 Element_VIA45_2_2_58_58 ;
      VIA 26.388 42.264 Element_VIA45_2_2_58_58 ;
      VIA 26.388 0.936 Element_VIA45_2_2_58_58 ;
      VIA 23.412 42.264 Element_VIA45_2_2_58_58 ;
      VIA 23.412 0.936 Element_VIA45_2_2_58_58 ;
      VIA 20.436 42.264 Element_VIA45_2_2_58_58 ;
      VIA 20.436 0.936 Element_VIA45_2_2_58_58 ;
      VIA 17.46 42.264 Element_VIA45_2_2_58_58 ;
      VIA 17.46 0.936 Element_VIA45_2_2_58_58 ;
      VIA 14.484 42.264 Element_VIA45_2_2_58_58 ;
      VIA 14.484 0.936 Element_VIA45_2_2_58_58 ;
      VIA 11.508 42.264 Element_VIA45_2_2_58_58 ;
      VIA 11.508 0.936 Element_VIA45_2_2_58_58 ;
      VIA 8.532 42.264 Element_VIA45_2_2_58_58 ;
      VIA 8.532 0.936 Element_VIA45_2_2_58_58 ;
      VIA 5.556 42.264 Element_VIA45_2_2_58_58 ;
      VIA 5.556 0.936 Element_VIA45_2_2_58_58 ;
      VIA 2.58 42.264 Element_VIA45_2_2_58_58 ;
      VIA 2.58 0.936 Element_VIA45_2_2_58_58 ;
      VIA 0.936 42.264 Element_VIA45_2_2_58_58 ;
      VIA 0.936 0.936 Element_VIA45_2_2_58_58 ;
      VIA 41.268 42.12 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 42.103 41.313 42.137 ;
      VIA 41.268 42.12 Element_VIA34_1_2_58_52 ;
      VIA 41.268 42.12 Element_VIA23_1_3_36_36 ;
      VIA 41.268 41.58 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 41.563 41.313 41.597 ;
      VIA 41.268 41.58 Element_VIA34_1_2_58_52 ;
      VIA 41.268 41.58 Element_VIA23_1_3_36_36 ;
      VIA 41.268 41.04 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 41.023 41.313 41.057 ;
      VIA 41.268 41.04 Element_VIA34_1_2_58_52 ;
      VIA 41.268 41.04 Element_VIA23_1_3_36_36 ;
      VIA 41.268 40.5 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 40.483 41.313 40.517 ;
      VIA 41.268 40.5 Element_VIA34_1_2_58_52 ;
      VIA 41.268 40.5 Element_VIA23_1_3_36_36 ;
      VIA 41.268 39.96 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 39.943 41.313 39.977 ;
      VIA 41.268 39.96 Element_VIA34_1_2_58_52 ;
      VIA 41.268 39.96 Element_VIA23_1_3_36_36 ;
      VIA 41.268 39.42 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 39.403 41.313 39.437 ;
      VIA 41.268 39.42 Element_VIA34_1_2_58_52 ;
      VIA 41.268 39.42 Element_VIA23_1_3_36_36 ;
      VIA 41.268 38.88 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 38.863 41.313 38.897 ;
      VIA 41.268 38.88 Element_VIA34_1_2_58_52 ;
      VIA 41.268 38.88 Element_VIA23_1_3_36_36 ;
      VIA 41.268 38.34 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 38.323 41.313 38.357 ;
      VIA 41.268 38.34 Element_VIA34_1_2_58_52 ;
      VIA 41.268 38.34 Element_VIA23_1_3_36_36 ;
      VIA 41.268 37.8 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 37.783 41.313 37.817 ;
      VIA 41.268 37.8 Element_VIA34_1_2_58_52 ;
      VIA 41.268 37.8 Element_VIA23_1_3_36_36 ;
      VIA 41.268 37.26 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 37.243 41.313 37.277 ;
      VIA 41.268 37.26 Element_VIA34_1_2_58_52 ;
      VIA 41.268 37.26 Element_VIA23_1_3_36_36 ;
      VIA 41.268 36.72 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 36.703 41.313 36.737 ;
      VIA 41.268 36.72 Element_VIA34_1_2_58_52 ;
      VIA 41.268 36.72 Element_VIA23_1_3_36_36 ;
      VIA 41.268 36.18 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 36.163 41.313 36.197 ;
      VIA 41.268 36.18 Element_VIA34_1_2_58_52 ;
      VIA 41.268 36.18 Element_VIA23_1_3_36_36 ;
      VIA 41.268 35.64 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 35.623 41.313 35.657 ;
      VIA 41.268 35.64 Element_VIA34_1_2_58_52 ;
      VIA 41.268 35.64 Element_VIA23_1_3_36_36 ;
      VIA 41.268 35.1 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 35.083 41.313 35.117 ;
      VIA 41.268 35.1 Element_VIA34_1_2_58_52 ;
      VIA 41.268 35.1 Element_VIA23_1_3_36_36 ;
      VIA 41.268 34.56 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 34.543 41.313 34.577 ;
      VIA 41.268 34.56 Element_VIA34_1_2_58_52 ;
      VIA 41.268 34.56 Element_VIA23_1_3_36_36 ;
      VIA 41.268 34.02 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 34.003 41.313 34.037 ;
      VIA 41.268 34.02 Element_VIA34_1_2_58_52 ;
      VIA 41.268 34.02 Element_VIA23_1_3_36_36 ;
      VIA 41.268 33.48 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 33.463 41.313 33.497 ;
      VIA 41.268 33.48 Element_VIA34_1_2_58_52 ;
      VIA 41.268 33.48 Element_VIA23_1_3_36_36 ;
      VIA 41.268 32.94 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 32.923 41.313 32.957 ;
      VIA 41.268 32.94 Element_VIA34_1_2_58_52 ;
      VIA 41.268 32.94 Element_VIA23_1_3_36_36 ;
      VIA 41.268 32.4 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 32.383 41.313 32.417 ;
      VIA 41.268 32.4 Element_VIA34_1_2_58_52 ;
      VIA 41.268 32.4 Element_VIA23_1_3_36_36 ;
      VIA 41.268 31.86 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 31.843 41.313 31.877 ;
      VIA 41.268 31.86 Element_VIA34_1_2_58_52 ;
      VIA 41.268 31.86 Element_VIA23_1_3_36_36 ;
      VIA 41.268 31.32 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 31.303 41.313 31.337 ;
      VIA 41.268 31.32 Element_VIA34_1_2_58_52 ;
      VIA 41.268 31.32 Element_VIA23_1_3_36_36 ;
      VIA 41.268 30.78 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 30.763 41.313 30.797 ;
      VIA 41.268 30.78 Element_VIA34_1_2_58_52 ;
      VIA 41.268 30.78 Element_VIA23_1_3_36_36 ;
      VIA 41.268 30.24 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 30.223 41.313 30.257 ;
      VIA 41.268 30.24 Element_VIA34_1_2_58_52 ;
      VIA 41.268 30.24 Element_VIA23_1_3_36_36 ;
      VIA 41.268 29.7 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 29.683 41.313 29.717 ;
      VIA 41.268 29.7 Element_VIA34_1_2_58_52 ;
      VIA 41.268 29.7 Element_VIA23_1_3_36_36 ;
      VIA 41.268 29.16 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 29.143 41.313 29.177 ;
      VIA 41.268 29.16 Element_VIA34_1_2_58_52 ;
      VIA 41.268 29.16 Element_VIA23_1_3_36_36 ;
      VIA 41.268 28.62 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 28.603 41.313 28.637 ;
      VIA 41.268 28.62 Element_VIA34_1_2_58_52 ;
      VIA 41.268 28.62 Element_VIA23_1_3_36_36 ;
      VIA 41.268 28.08 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 28.063 41.313 28.097 ;
      VIA 41.268 28.08 Element_VIA34_1_2_58_52 ;
      VIA 41.268 28.08 Element_VIA23_1_3_36_36 ;
      VIA 41.268 27.54 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 27.523 41.313 27.557 ;
      VIA 41.268 27.54 Element_VIA34_1_2_58_52 ;
      VIA 41.268 27.54 Element_VIA23_1_3_36_36 ;
      VIA 41.268 27 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 26.983 41.313 27.017 ;
      VIA 41.268 27 Element_VIA34_1_2_58_52 ;
      VIA 41.268 27 Element_VIA23_1_3_36_36 ;
      VIA 41.268 26.46 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 26.443 41.313 26.477 ;
      VIA 41.268 26.46 Element_VIA34_1_2_58_52 ;
      VIA 41.268 26.46 Element_VIA23_1_3_36_36 ;
      VIA 41.268 25.92 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 25.903 41.313 25.937 ;
      VIA 41.268 25.92 Element_VIA34_1_2_58_52 ;
      VIA 41.268 25.92 Element_VIA23_1_3_36_36 ;
      VIA 41.268 25.38 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 25.363 41.313 25.397 ;
      VIA 41.268 25.38 Element_VIA34_1_2_58_52 ;
      VIA 41.268 25.38 Element_VIA23_1_3_36_36 ;
      VIA 41.268 24.84 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 24.823 41.313 24.857 ;
      VIA 41.268 24.84 Element_VIA34_1_2_58_52 ;
      VIA 41.268 24.84 Element_VIA23_1_3_36_36 ;
      VIA 41.268 24.3 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 24.283 41.313 24.317 ;
      VIA 41.268 24.3 Element_VIA34_1_2_58_52 ;
      VIA 41.268 24.3 Element_VIA23_1_3_36_36 ;
      VIA 41.268 23.76 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 23.743 41.313 23.777 ;
      VIA 41.268 23.76 Element_VIA34_1_2_58_52 ;
      VIA 41.268 23.76 Element_VIA23_1_3_36_36 ;
      VIA 41.268 23.22 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 23.203 41.313 23.237 ;
      VIA 41.268 23.22 Element_VIA34_1_2_58_52 ;
      VIA 41.268 23.22 Element_VIA23_1_3_36_36 ;
      VIA 41.268 22.68 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 22.663 41.313 22.697 ;
      VIA 41.268 22.68 Element_VIA34_1_2_58_52 ;
      VIA 41.268 22.68 Element_VIA23_1_3_36_36 ;
      VIA 41.268 22.14 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 22.123 41.313 22.157 ;
      VIA 41.268 22.14 Element_VIA34_1_2_58_52 ;
      VIA 41.268 22.14 Element_VIA23_1_3_36_36 ;
      VIA 41.268 21.6 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 21.583 41.313 21.617 ;
      VIA 41.268 21.6 Element_VIA34_1_2_58_52 ;
      VIA 41.268 21.6 Element_VIA23_1_3_36_36 ;
      VIA 41.268 21.06 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 21.043 41.313 21.077 ;
      VIA 41.268 21.06 Element_VIA34_1_2_58_52 ;
      VIA 41.268 21.06 Element_VIA23_1_3_36_36 ;
      VIA 41.268 20.52 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 20.503 41.313 20.537 ;
      VIA 41.268 20.52 Element_VIA34_1_2_58_52 ;
      VIA 41.268 20.52 Element_VIA23_1_3_36_36 ;
      VIA 41.268 19.98 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 19.963 41.313 19.997 ;
      VIA 41.268 19.98 Element_VIA34_1_2_58_52 ;
      VIA 41.268 19.98 Element_VIA23_1_3_36_36 ;
      VIA 41.268 19.44 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 19.423 41.313 19.457 ;
      VIA 41.268 19.44 Element_VIA34_1_2_58_52 ;
      VIA 41.268 19.44 Element_VIA23_1_3_36_36 ;
      VIA 41.268 18.9 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 18.883 41.313 18.917 ;
      VIA 41.268 18.9 Element_VIA34_1_2_58_52 ;
      VIA 41.268 18.9 Element_VIA23_1_3_36_36 ;
      VIA 41.268 18.36 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 18.343 41.313 18.377 ;
      VIA 41.268 18.36 Element_VIA34_1_2_58_52 ;
      VIA 41.268 18.36 Element_VIA23_1_3_36_36 ;
      VIA 41.268 17.82 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 17.803 41.313 17.837 ;
      VIA 41.268 17.82 Element_VIA34_1_2_58_52 ;
      VIA 41.268 17.82 Element_VIA23_1_3_36_36 ;
      VIA 41.268 17.28 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 17.263 41.313 17.297 ;
      VIA 41.268 17.28 Element_VIA34_1_2_58_52 ;
      VIA 41.268 17.28 Element_VIA23_1_3_36_36 ;
      VIA 41.268 16.74 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 16.723 41.313 16.757 ;
      VIA 41.268 16.74 Element_VIA34_1_2_58_52 ;
      VIA 41.268 16.74 Element_VIA23_1_3_36_36 ;
      VIA 41.268 16.2 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 16.183 41.313 16.217 ;
      VIA 41.268 16.2 Element_VIA34_1_2_58_52 ;
      VIA 41.268 16.2 Element_VIA23_1_3_36_36 ;
      VIA 41.268 15.66 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 15.643 41.313 15.677 ;
      VIA 41.268 15.66 Element_VIA34_1_2_58_52 ;
      VIA 41.268 15.66 Element_VIA23_1_3_36_36 ;
      VIA 41.268 15.12 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 15.103 41.313 15.137 ;
      VIA 41.268 15.12 Element_VIA34_1_2_58_52 ;
      VIA 41.268 15.12 Element_VIA23_1_3_36_36 ;
      VIA 41.268 14.58 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 14.563 41.313 14.597 ;
      VIA 41.268 14.58 Element_VIA34_1_2_58_52 ;
      VIA 41.268 14.58 Element_VIA23_1_3_36_36 ;
      VIA 41.268 14.04 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 14.023 41.313 14.057 ;
      VIA 41.268 14.04 Element_VIA34_1_2_58_52 ;
      VIA 41.268 14.04 Element_VIA23_1_3_36_36 ;
      VIA 41.268 13.5 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 13.483 41.313 13.517 ;
      VIA 41.268 13.5 Element_VIA34_1_2_58_52 ;
      VIA 41.268 13.5 Element_VIA23_1_3_36_36 ;
      VIA 41.268 12.96 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 12.943 41.313 12.977 ;
      VIA 41.268 12.96 Element_VIA34_1_2_58_52 ;
      VIA 41.268 12.96 Element_VIA23_1_3_36_36 ;
      VIA 41.268 12.42 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 12.403 41.313 12.437 ;
      VIA 41.268 12.42 Element_VIA34_1_2_58_52 ;
      VIA 41.268 12.42 Element_VIA23_1_3_36_36 ;
      VIA 41.268 11.88 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 11.863 41.313 11.897 ;
      VIA 41.268 11.88 Element_VIA34_1_2_58_52 ;
      VIA 41.268 11.88 Element_VIA23_1_3_36_36 ;
      VIA 41.268 11.34 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 11.323 41.313 11.357 ;
      VIA 41.268 11.34 Element_VIA34_1_2_58_52 ;
      VIA 41.268 11.34 Element_VIA23_1_3_36_36 ;
      VIA 41.268 10.8 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 10.783 41.313 10.817 ;
      VIA 41.268 10.8 Element_VIA34_1_2_58_52 ;
      VIA 41.268 10.8 Element_VIA23_1_3_36_36 ;
      VIA 41.268 10.26 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 10.243 41.313 10.277 ;
      VIA 41.268 10.26 Element_VIA34_1_2_58_52 ;
      VIA 41.268 10.26 Element_VIA23_1_3_36_36 ;
      VIA 41.268 9.72 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 9.703 41.313 9.737 ;
      VIA 41.268 9.72 Element_VIA34_1_2_58_52 ;
      VIA 41.268 9.72 Element_VIA23_1_3_36_36 ;
      VIA 41.268 9.18 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 9.163 41.313 9.197 ;
      VIA 41.268 9.18 Element_VIA34_1_2_58_52 ;
      VIA 41.268 9.18 Element_VIA23_1_3_36_36 ;
      VIA 41.268 8.64 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 8.623 41.313 8.657 ;
      VIA 41.268 8.64 Element_VIA34_1_2_58_52 ;
      VIA 41.268 8.64 Element_VIA23_1_3_36_36 ;
      VIA 41.268 8.1 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 8.083 41.313 8.117 ;
      VIA 41.268 8.1 Element_VIA34_1_2_58_52 ;
      VIA 41.268 8.1 Element_VIA23_1_3_36_36 ;
      VIA 41.268 7.56 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 7.543 41.313 7.577 ;
      VIA 41.268 7.56 Element_VIA34_1_2_58_52 ;
      VIA 41.268 7.56 Element_VIA23_1_3_36_36 ;
      VIA 41.268 7.02 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 7.003 41.313 7.037 ;
      VIA 41.268 7.02 Element_VIA34_1_2_58_52 ;
      VIA 41.268 7.02 Element_VIA23_1_3_36_36 ;
      VIA 41.268 6.48 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 6.463 41.313 6.497 ;
      VIA 41.268 6.48 Element_VIA34_1_2_58_52 ;
      VIA 41.268 6.48 Element_VIA23_1_3_36_36 ;
      VIA 41.268 5.94 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 5.923 41.313 5.957 ;
      VIA 41.268 5.94 Element_VIA34_1_2_58_52 ;
      VIA 41.268 5.94 Element_VIA23_1_3_36_36 ;
      VIA 41.268 5.4 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 5.383 41.313 5.417 ;
      VIA 41.268 5.4 Element_VIA34_1_2_58_52 ;
      VIA 41.268 5.4 Element_VIA23_1_3_36_36 ;
      VIA 41.268 4.86 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 4.843 41.313 4.877 ;
      VIA 41.268 4.86 Element_VIA34_1_2_58_52 ;
      VIA 41.268 4.86 Element_VIA23_1_3_36_36 ;
      VIA 41.268 4.32 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 4.303 41.313 4.337 ;
      VIA 41.268 4.32 Element_VIA34_1_2_58_52 ;
      VIA 41.268 4.32 Element_VIA23_1_3_36_36 ;
      VIA 41.268 3.78 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 3.763 41.313 3.797 ;
      VIA 41.268 3.78 Element_VIA34_1_2_58_52 ;
      VIA 41.268 3.78 Element_VIA23_1_3_36_36 ;
      VIA 41.268 3.24 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 3.223 41.313 3.257 ;
      VIA 41.268 3.24 Element_VIA34_1_2_58_52 ;
      VIA 41.268 3.24 Element_VIA23_1_3_36_36 ;
      VIA 41.268 2.7 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 2.683 41.313 2.717 ;
      VIA 41.268 2.7 Element_VIA34_1_2_58_52 ;
      VIA 41.268 2.7 Element_VIA23_1_3_36_36 ;
      VIA 41.268 2.16 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 2.143 41.313 2.177 ;
      VIA 41.268 2.16 Element_VIA34_1_2_58_52 ;
      VIA 41.268 2.16 Element_VIA23_1_3_36_36 ;
      VIA 41.268 1.62 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 1.603 41.313 1.637 ;
      VIA 41.268 1.62 Element_VIA34_1_2_58_52 ;
      VIA 41.268 1.62 Element_VIA23_1_3_36_36 ;
      VIA 41.268 1.08 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  41.223 1.063 41.313 1.097 ;
      VIA 41.268 1.08 Element_VIA34_1_2_58_52 ;
      VIA 41.268 1.08 Element_VIA23_1_3_36_36 ;
      VIA 38.292 42.12 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 42.103 38.337 42.137 ;
      VIA 38.292 42.12 Element_VIA34_1_2_58_52 ;
      VIA 38.292 42.12 Element_VIA23_1_3_36_36 ;
      VIA 38.292 41.58 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 41.563 38.337 41.597 ;
      VIA 38.292 41.58 Element_VIA34_1_2_58_52 ;
      VIA 38.292 41.58 Element_VIA23_1_3_36_36 ;
      VIA 38.292 41.04 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 41.023 38.337 41.057 ;
      VIA 38.292 41.04 Element_VIA34_1_2_58_52 ;
      VIA 38.292 41.04 Element_VIA23_1_3_36_36 ;
      VIA 38.292 40.5 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 40.483 38.337 40.517 ;
      VIA 38.292 40.5 Element_VIA34_1_2_58_52 ;
      VIA 38.292 40.5 Element_VIA23_1_3_36_36 ;
      VIA 38.292 39.96 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 39.943 38.337 39.977 ;
      VIA 38.292 39.96 Element_VIA34_1_2_58_52 ;
      VIA 38.292 39.96 Element_VIA23_1_3_36_36 ;
      VIA 38.292 39.42 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 39.403 38.337 39.437 ;
      VIA 38.292 39.42 Element_VIA34_1_2_58_52 ;
      VIA 38.292 39.42 Element_VIA23_1_3_36_36 ;
      VIA 38.292 38.88 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 38.863 38.337 38.897 ;
      VIA 38.292 38.88 Element_VIA34_1_2_58_52 ;
      VIA 38.292 38.88 Element_VIA23_1_3_36_36 ;
      VIA 38.292 38.34 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 38.323 38.337 38.357 ;
      VIA 38.292 38.34 Element_VIA34_1_2_58_52 ;
      VIA 38.292 38.34 Element_VIA23_1_3_36_36 ;
      VIA 38.292 37.8 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 37.783 38.337 37.817 ;
      VIA 38.292 37.8 Element_VIA34_1_2_58_52 ;
      VIA 38.292 37.8 Element_VIA23_1_3_36_36 ;
      VIA 38.292 37.26 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 37.243 38.337 37.277 ;
      VIA 38.292 37.26 Element_VIA34_1_2_58_52 ;
      VIA 38.292 37.26 Element_VIA23_1_3_36_36 ;
      VIA 38.292 36.72 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 36.703 38.337 36.737 ;
      VIA 38.292 36.72 Element_VIA34_1_2_58_52 ;
      VIA 38.292 36.72 Element_VIA23_1_3_36_36 ;
      VIA 38.292 36.18 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 36.163 38.337 36.197 ;
      VIA 38.292 36.18 Element_VIA34_1_2_58_52 ;
      VIA 38.292 36.18 Element_VIA23_1_3_36_36 ;
      VIA 38.292 35.64 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 35.623 38.337 35.657 ;
      VIA 38.292 35.64 Element_VIA34_1_2_58_52 ;
      VIA 38.292 35.64 Element_VIA23_1_3_36_36 ;
      VIA 38.292 35.1 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 35.083 38.337 35.117 ;
      VIA 38.292 35.1 Element_VIA34_1_2_58_52 ;
      VIA 38.292 35.1 Element_VIA23_1_3_36_36 ;
      VIA 38.292 34.56 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 34.543 38.337 34.577 ;
      VIA 38.292 34.56 Element_VIA34_1_2_58_52 ;
      VIA 38.292 34.56 Element_VIA23_1_3_36_36 ;
      VIA 38.292 34.02 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 34.003 38.337 34.037 ;
      VIA 38.292 34.02 Element_VIA34_1_2_58_52 ;
      VIA 38.292 34.02 Element_VIA23_1_3_36_36 ;
      VIA 38.292 33.48 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 33.463 38.337 33.497 ;
      VIA 38.292 33.48 Element_VIA34_1_2_58_52 ;
      VIA 38.292 33.48 Element_VIA23_1_3_36_36 ;
      VIA 38.292 32.94 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 32.923 38.337 32.957 ;
      VIA 38.292 32.94 Element_VIA34_1_2_58_52 ;
      VIA 38.292 32.94 Element_VIA23_1_3_36_36 ;
      VIA 38.292 32.4 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 32.383 38.337 32.417 ;
      VIA 38.292 32.4 Element_VIA34_1_2_58_52 ;
      VIA 38.292 32.4 Element_VIA23_1_3_36_36 ;
      VIA 38.292 31.86 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 31.843 38.337 31.877 ;
      VIA 38.292 31.86 Element_VIA34_1_2_58_52 ;
      VIA 38.292 31.86 Element_VIA23_1_3_36_36 ;
      VIA 38.292 31.32 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 31.303 38.337 31.337 ;
      VIA 38.292 31.32 Element_VIA34_1_2_58_52 ;
      VIA 38.292 31.32 Element_VIA23_1_3_36_36 ;
      VIA 38.292 30.78 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 30.763 38.337 30.797 ;
      VIA 38.292 30.78 Element_VIA34_1_2_58_52 ;
      VIA 38.292 30.78 Element_VIA23_1_3_36_36 ;
      VIA 38.292 30.24 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 30.223 38.337 30.257 ;
      VIA 38.292 30.24 Element_VIA34_1_2_58_52 ;
      VIA 38.292 30.24 Element_VIA23_1_3_36_36 ;
      VIA 38.292 29.7 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 29.683 38.337 29.717 ;
      VIA 38.292 29.7 Element_VIA34_1_2_58_52 ;
      VIA 38.292 29.7 Element_VIA23_1_3_36_36 ;
      VIA 38.292 29.16 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 29.143 38.337 29.177 ;
      VIA 38.292 29.16 Element_VIA34_1_2_58_52 ;
      VIA 38.292 29.16 Element_VIA23_1_3_36_36 ;
      VIA 38.292 28.62 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 28.603 38.337 28.637 ;
      VIA 38.292 28.62 Element_VIA34_1_2_58_52 ;
      VIA 38.292 28.62 Element_VIA23_1_3_36_36 ;
      VIA 38.292 28.08 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 28.063 38.337 28.097 ;
      VIA 38.292 28.08 Element_VIA34_1_2_58_52 ;
      VIA 38.292 28.08 Element_VIA23_1_3_36_36 ;
      VIA 38.292 27.54 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 27.523 38.337 27.557 ;
      VIA 38.292 27.54 Element_VIA34_1_2_58_52 ;
      VIA 38.292 27.54 Element_VIA23_1_3_36_36 ;
      VIA 38.292 27 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 26.983 38.337 27.017 ;
      VIA 38.292 27 Element_VIA34_1_2_58_52 ;
      VIA 38.292 27 Element_VIA23_1_3_36_36 ;
      VIA 38.292 26.46 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 26.443 38.337 26.477 ;
      VIA 38.292 26.46 Element_VIA34_1_2_58_52 ;
      VIA 38.292 26.46 Element_VIA23_1_3_36_36 ;
      VIA 38.292 25.92 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 25.903 38.337 25.937 ;
      VIA 38.292 25.92 Element_VIA34_1_2_58_52 ;
      VIA 38.292 25.92 Element_VIA23_1_3_36_36 ;
      VIA 38.292 25.38 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 25.363 38.337 25.397 ;
      VIA 38.292 25.38 Element_VIA34_1_2_58_52 ;
      VIA 38.292 25.38 Element_VIA23_1_3_36_36 ;
      VIA 38.292 24.84 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 24.823 38.337 24.857 ;
      VIA 38.292 24.84 Element_VIA34_1_2_58_52 ;
      VIA 38.292 24.84 Element_VIA23_1_3_36_36 ;
      VIA 38.292 24.3 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 24.283 38.337 24.317 ;
      VIA 38.292 24.3 Element_VIA34_1_2_58_52 ;
      VIA 38.292 24.3 Element_VIA23_1_3_36_36 ;
      VIA 38.292 23.76 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 23.743 38.337 23.777 ;
      VIA 38.292 23.76 Element_VIA34_1_2_58_52 ;
      VIA 38.292 23.76 Element_VIA23_1_3_36_36 ;
      VIA 38.292 23.22 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 23.203 38.337 23.237 ;
      VIA 38.292 23.22 Element_VIA34_1_2_58_52 ;
      VIA 38.292 23.22 Element_VIA23_1_3_36_36 ;
      VIA 38.292 22.68 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 22.663 38.337 22.697 ;
      VIA 38.292 22.68 Element_VIA34_1_2_58_52 ;
      VIA 38.292 22.68 Element_VIA23_1_3_36_36 ;
      VIA 38.292 22.14 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 22.123 38.337 22.157 ;
      VIA 38.292 22.14 Element_VIA34_1_2_58_52 ;
      VIA 38.292 22.14 Element_VIA23_1_3_36_36 ;
      VIA 38.292 21.6 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 21.583 38.337 21.617 ;
      VIA 38.292 21.6 Element_VIA34_1_2_58_52 ;
      VIA 38.292 21.6 Element_VIA23_1_3_36_36 ;
      VIA 38.292 21.06 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 21.043 38.337 21.077 ;
      VIA 38.292 21.06 Element_VIA34_1_2_58_52 ;
      VIA 38.292 21.06 Element_VIA23_1_3_36_36 ;
      VIA 38.292 20.52 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 20.503 38.337 20.537 ;
      VIA 38.292 20.52 Element_VIA34_1_2_58_52 ;
      VIA 38.292 20.52 Element_VIA23_1_3_36_36 ;
      VIA 38.292 19.98 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 19.963 38.337 19.997 ;
      VIA 38.292 19.98 Element_VIA34_1_2_58_52 ;
      VIA 38.292 19.98 Element_VIA23_1_3_36_36 ;
      VIA 38.292 19.44 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 19.423 38.337 19.457 ;
      VIA 38.292 19.44 Element_VIA34_1_2_58_52 ;
      VIA 38.292 19.44 Element_VIA23_1_3_36_36 ;
      VIA 38.292 18.9 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 18.883 38.337 18.917 ;
      VIA 38.292 18.9 Element_VIA34_1_2_58_52 ;
      VIA 38.292 18.9 Element_VIA23_1_3_36_36 ;
      VIA 38.292 18.36 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 18.343 38.337 18.377 ;
      VIA 38.292 18.36 Element_VIA34_1_2_58_52 ;
      VIA 38.292 18.36 Element_VIA23_1_3_36_36 ;
      VIA 38.292 17.82 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 17.803 38.337 17.837 ;
      VIA 38.292 17.82 Element_VIA34_1_2_58_52 ;
      VIA 38.292 17.82 Element_VIA23_1_3_36_36 ;
      VIA 38.292 17.28 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 17.263 38.337 17.297 ;
      VIA 38.292 17.28 Element_VIA34_1_2_58_52 ;
      VIA 38.292 17.28 Element_VIA23_1_3_36_36 ;
      VIA 38.292 16.74 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 16.723 38.337 16.757 ;
      VIA 38.292 16.74 Element_VIA34_1_2_58_52 ;
      VIA 38.292 16.74 Element_VIA23_1_3_36_36 ;
      VIA 38.292 16.2 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 16.183 38.337 16.217 ;
      VIA 38.292 16.2 Element_VIA34_1_2_58_52 ;
      VIA 38.292 16.2 Element_VIA23_1_3_36_36 ;
      VIA 38.292 15.66 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 15.643 38.337 15.677 ;
      VIA 38.292 15.66 Element_VIA34_1_2_58_52 ;
      VIA 38.292 15.66 Element_VIA23_1_3_36_36 ;
      VIA 38.292 15.12 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 15.103 38.337 15.137 ;
      VIA 38.292 15.12 Element_VIA34_1_2_58_52 ;
      VIA 38.292 15.12 Element_VIA23_1_3_36_36 ;
      VIA 38.292 14.58 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 14.563 38.337 14.597 ;
      VIA 38.292 14.58 Element_VIA34_1_2_58_52 ;
      VIA 38.292 14.58 Element_VIA23_1_3_36_36 ;
      VIA 38.292 14.04 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 14.023 38.337 14.057 ;
      VIA 38.292 14.04 Element_VIA34_1_2_58_52 ;
      VIA 38.292 14.04 Element_VIA23_1_3_36_36 ;
      VIA 38.292 13.5 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 13.483 38.337 13.517 ;
      VIA 38.292 13.5 Element_VIA34_1_2_58_52 ;
      VIA 38.292 13.5 Element_VIA23_1_3_36_36 ;
      VIA 38.292 12.96 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 12.943 38.337 12.977 ;
      VIA 38.292 12.96 Element_VIA34_1_2_58_52 ;
      VIA 38.292 12.96 Element_VIA23_1_3_36_36 ;
      VIA 38.292 12.42 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 12.403 38.337 12.437 ;
      VIA 38.292 12.42 Element_VIA34_1_2_58_52 ;
      VIA 38.292 12.42 Element_VIA23_1_3_36_36 ;
      VIA 38.292 11.88 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 11.863 38.337 11.897 ;
      VIA 38.292 11.88 Element_VIA34_1_2_58_52 ;
      VIA 38.292 11.88 Element_VIA23_1_3_36_36 ;
      VIA 38.292 11.34 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 11.323 38.337 11.357 ;
      VIA 38.292 11.34 Element_VIA34_1_2_58_52 ;
      VIA 38.292 11.34 Element_VIA23_1_3_36_36 ;
      VIA 38.292 10.8 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 10.783 38.337 10.817 ;
      VIA 38.292 10.8 Element_VIA34_1_2_58_52 ;
      VIA 38.292 10.8 Element_VIA23_1_3_36_36 ;
      VIA 38.292 10.26 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 10.243 38.337 10.277 ;
      VIA 38.292 10.26 Element_VIA34_1_2_58_52 ;
      VIA 38.292 10.26 Element_VIA23_1_3_36_36 ;
      VIA 38.292 9.72 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 9.703 38.337 9.737 ;
      VIA 38.292 9.72 Element_VIA34_1_2_58_52 ;
      VIA 38.292 9.72 Element_VIA23_1_3_36_36 ;
      VIA 38.292 9.18 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 9.163 38.337 9.197 ;
      VIA 38.292 9.18 Element_VIA34_1_2_58_52 ;
      VIA 38.292 9.18 Element_VIA23_1_3_36_36 ;
      VIA 38.292 8.64 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 8.623 38.337 8.657 ;
      VIA 38.292 8.64 Element_VIA34_1_2_58_52 ;
      VIA 38.292 8.64 Element_VIA23_1_3_36_36 ;
      VIA 38.292 8.1 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 8.083 38.337 8.117 ;
      VIA 38.292 8.1 Element_VIA34_1_2_58_52 ;
      VIA 38.292 8.1 Element_VIA23_1_3_36_36 ;
      VIA 38.292 7.56 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 7.543 38.337 7.577 ;
      VIA 38.292 7.56 Element_VIA34_1_2_58_52 ;
      VIA 38.292 7.56 Element_VIA23_1_3_36_36 ;
      VIA 38.292 7.02 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 7.003 38.337 7.037 ;
      VIA 38.292 7.02 Element_VIA34_1_2_58_52 ;
      VIA 38.292 7.02 Element_VIA23_1_3_36_36 ;
      VIA 38.292 6.48 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 6.463 38.337 6.497 ;
      VIA 38.292 6.48 Element_VIA34_1_2_58_52 ;
      VIA 38.292 6.48 Element_VIA23_1_3_36_36 ;
      VIA 38.292 5.94 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 5.923 38.337 5.957 ;
      VIA 38.292 5.94 Element_VIA34_1_2_58_52 ;
      VIA 38.292 5.94 Element_VIA23_1_3_36_36 ;
      VIA 38.292 5.4 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 5.383 38.337 5.417 ;
      VIA 38.292 5.4 Element_VIA34_1_2_58_52 ;
      VIA 38.292 5.4 Element_VIA23_1_3_36_36 ;
      VIA 38.292 4.86 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 4.843 38.337 4.877 ;
      VIA 38.292 4.86 Element_VIA34_1_2_58_52 ;
      VIA 38.292 4.86 Element_VIA23_1_3_36_36 ;
      VIA 38.292 4.32 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 4.303 38.337 4.337 ;
      VIA 38.292 4.32 Element_VIA34_1_2_58_52 ;
      VIA 38.292 4.32 Element_VIA23_1_3_36_36 ;
      VIA 38.292 3.78 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 3.763 38.337 3.797 ;
      VIA 38.292 3.78 Element_VIA34_1_2_58_52 ;
      VIA 38.292 3.78 Element_VIA23_1_3_36_36 ;
      VIA 38.292 3.24 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 3.223 38.337 3.257 ;
      VIA 38.292 3.24 Element_VIA34_1_2_58_52 ;
      VIA 38.292 3.24 Element_VIA23_1_3_36_36 ;
      VIA 38.292 2.7 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 2.683 38.337 2.717 ;
      VIA 38.292 2.7 Element_VIA34_1_2_58_52 ;
      VIA 38.292 2.7 Element_VIA23_1_3_36_36 ;
      VIA 38.292 2.16 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 2.143 38.337 2.177 ;
      VIA 38.292 2.16 Element_VIA34_1_2_58_52 ;
      VIA 38.292 2.16 Element_VIA23_1_3_36_36 ;
      VIA 38.292 1.62 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 1.603 38.337 1.637 ;
      VIA 38.292 1.62 Element_VIA34_1_2_58_52 ;
      VIA 38.292 1.62 Element_VIA23_1_3_36_36 ;
      VIA 38.292 1.08 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  38.247 1.063 38.337 1.097 ;
      VIA 38.292 1.08 Element_VIA34_1_2_58_52 ;
      VIA 38.292 1.08 Element_VIA23_1_3_36_36 ;
      VIA 35.316 42.12 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 42.103 35.361 42.137 ;
      VIA 35.316 42.12 Element_VIA34_1_2_58_52 ;
      VIA 35.316 42.12 Element_VIA23_1_3_36_36 ;
      VIA 35.316 41.58 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 41.563 35.361 41.597 ;
      VIA 35.316 41.58 Element_VIA34_1_2_58_52 ;
      VIA 35.316 41.58 Element_VIA23_1_3_36_36 ;
      VIA 35.316 41.04 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 41.023 35.361 41.057 ;
      VIA 35.316 41.04 Element_VIA34_1_2_58_52 ;
      VIA 35.316 41.04 Element_VIA23_1_3_36_36 ;
      VIA 35.316 40.5 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 40.483 35.361 40.517 ;
      VIA 35.316 40.5 Element_VIA34_1_2_58_52 ;
      VIA 35.316 40.5 Element_VIA23_1_3_36_36 ;
      VIA 35.316 39.96 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 39.943 35.361 39.977 ;
      VIA 35.316 39.96 Element_VIA34_1_2_58_52 ;
      VIA 35.316 39.96 Element_VIA23_1_3_36_36 ;
      VIA 35.316 39.42 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 39.403 35.361 39.437 ;
      VIA 35.316 39.42 Element_VIA34_1_2_58_52 ;
      VIA 35.316 39.42 Element_VIA23_1_3_36_36 ;
      VIA 35.316 38.88 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 38.863 35.361 38.897 ;
      VIA 35.316 38.88 Element_VIA34_1_2_58_52 ;
      VIA 35.316 38.88 Element_VIA23_1_3_36_36 ;
      VIA 35.316 38.34 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 38.323 35.361 38.357 ;
      VIA 35.316 38.34 Element_VIA34_1_2_58_52 ;
      VIA 35.316 38.34 Element_VIA23_1_3_36_36 ;
      VIA 35.316 37.8 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 37.783 35.361 37.817 ;
      VIA 35.316 37.8 Element_VIA34_1_2_58_52 ;
      VIA 35.316 37.8 Element_VIA23_1_3_36_36 ;
      VIA 35.316 37.26 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 37.243 35.361 37.277 ;
      VIA 35.316 37.26 Element_VIA34_1_2_58_52 ;
      VIA 35.316 37.26 Element_VIA23_1_3_36_36 ;
      VIA 35.316 36.72 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 36.703 35.361 36.737 ;
      VIA 35.316 36.72 Element_VIA34_1_2_58_52 ;
      VIA 35.316 36.72 Element_VIA23_1_3_36_36 ;
      VIA 35.316 36.18 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 36.163 35.361 36.197 ;
      VIA 35.316 36.18 Element_VIA34_1_2_58_52 ;
      VIA 35.316 36.18 Element_VIA23_1_3_36_36 ;
      VIA 35.316 35.64 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 35.623 35.361 35.657 ;
      VIA 35.316 35.64 Element_VIA34_1_2_58_52 ;
      VIA 35.316 35.64 Element_VIA23_1_3_36_36 ;
      VIA 35.316 35.1 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 35.083 35.361 35.117 ;
      VIA 35.316 35.1 Element_VIA34_1_2_58_52 ;
      VIA 35.316 35.1 Element_VIA23_1_3_36_36 ;
      VIA 35.316 34.56 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 34.543 35.361 34.577 ;
      VIA 35.316 34.56 Element_VIA34_1_2_58_52 ;
      VIA 35.316 34.56 Element_VIA23_1_3_36_36 ;
      VIA 35.316 34.02 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 34.003 35.361 34.037 ;
      VIA 35.316 34.02 Element_VIA34_1_2_58_52 ;
      VIA 35.316 34.02 Element_VIA23_1_3_36_36 ;
      VIA 35.316 33.48 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 33.463 35.361 33.497 ;
      VIA 35.316 33.48 Element_VIA34_1_2_58_52 ;
      VIA 35.316 33.48 Element_VIA23_1_3_36_36 ;
      VIA 35.316 32.94 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 32.923 35.361 32.957 ;
      VIA 35.316 32.94 Element_VIA34_1_2_58_52 ;
      VIA 35.316 32.94 Element_VIA23_1_3_36_36 ;
      VIA 35.316 32.4 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 32.383 35.361 32.417 ;
      VIA 35.316 32.4 Element_VIA34_1_2_58_52 ;
      VIA 35.316 32.4 Element_VIA23_1_3_36_36 ;
      VIA 35.316 31.86 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 31.843 35.361 31.877 ;
      VIA 35.316 31.86 Element_VIA34_1_2_58_52 ;
      VIA 35.316 31.86 Element_VIA23_1_3_36_36 ;
      VIA 35.316 31.32 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 31.303 35.361 31.337 ;
      VIA 35.316 31.32 Element_VIA34_1_2_58_52 ;
      VIA 35.316 31.32 Element_VIA23_1_3_36_36 ;
      VIA 35.316 30.78 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 30.763 35.361 30.797 ;
      VIA 35.316 30.78 Element_VIA34_1_2_58_52 ;
      VIA 35.316 30.78 Element_VIA23_1_3_36_36 ;
      VIA 35.316 30.24 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 30.223 35.361 30.257 ;
      VIA 35.316 30.24 Element_VIA34_1_2_58_52 ;
      VIA 35.316 30.24 Element_VIA23_1_3_36_36 ;
      VIA 35.316 29.7 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 29.683 35.361 29.717 ;
      VIA 35.316 29.7 Element_VIA34_1_2_58_52 ;
      VIA 35.316 29.7 Element_VIA23_1_3_36_36 ;
      VIA 35.316 29.16 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 29.143 35.361 29.177 ;
      VIA 35.316 29.16 Element_VIA34_1_2_58_52 ;
      VIA 35.316 29.16 Element_VIA23_1_3_36_36 ;
      VIA 35.316 28.62 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 28.603 35.361 28.637 ;
      VIA 35.316 28.62 Element_VIA34_1_2_58_52 ;
      VIA 35.316 28.62 Element_VIA23_1_3_36_36 ;
      VIA 35.316 28.08 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 28.063 35.361 28.097 ;
      VIA 35.316 28.08 Element_VIA34_1_2_58_52 ;
      VIA 35.316 28.08 Element_VIA23_1_3_36_36 ;
      VIA 35.316 27.54 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 27.523 35.361 27.557 ;
      VIA 35.316 27.54 Element_VIA34_1_2_58_52 ;
      VIA 35.316 27.54 Element_VIA23_1_3_36_36 ;
      VIA 35.316 27 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 26.983 35.361 27.017 ;
      VIA 35.316 27 Element_VIA34_1_2_58_52 ;
      VIA 35.316 27 Element_VIA23_1_3_36_36 ;
      VIA 35.316 26.46 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 26.443 35.361 26.477 ;
      VIA 35.316 26.46 Element_VIA34_1_2_58_52 ;
      VIA 35.316 26.46 Element_VIA23_1_3_36_36 ;
      VIA 35.316 25.92 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 25.903 35.361 25.937 ;
      VIA 35.316 25.92 Element_VIA34_1_2_58_52 ;
      VIA 35.316 25.92 Element_VIA23_1_3_36_36 ;
      VIA 35.316 25.38 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 25.363 35.361 25.397 ;
      VIA 35.316 25.38 Element_VIA34_1_2_58_52 ;
      VIA 35.316 25.38 Element_VIA23_1_3_36_36 ;
      VIA 35.316 24.84 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 24.823 35.361 24.857 ;
      VIA 35.316 24.84 Element_VIA34_1_2_58_52 ;
      VIA 35.316 24.84 Element_VIA23_1_3_36_36 ;
      VIA 35.316 24.3 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 24.283 35.361 24.317 ;
      VIA 35.316 24.3 Element_VIA34_1_2_58_52 ;
      VIA 35.316 24.3 Element_VIA23_1_3_36_36 ;
      VIA 35.316 23.76 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 23.743 35.361 23.777 ;
      VIA 35.316 23.76 Element_VIA34_1_2_58_52 ;
      VIA 35.316 23.76 Element_VIA23_1_3_36_36 ;
      VIA 35.316 23.22 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 23.203 35.361 23.237 ;
      VIA 35.316 23.22 Element_VIA34_1_2_58_52 ;
      VIA 35.316 23.22 Element_VIA23_1_3_36_36 ;
      VIA 35.316 22.68 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 22.663 35.361 22.697 ;
      VIA 35.316 22.68 Element_VIA34_1_2_58_52 ;
      VIA 35.316 22.68 Element_VIA23_1_3_36_36 ;
      VIA 35.316 22.14 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 22.123 35.361 22.157 ;
      VIA 35.316 22.14 Element_VIA34_1_2_58_52 ;
      VIA 35.316 22.14 Element_VIA23_1_3_36_36 ;
      VIA 35.316 21.6 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 21.583 35.361 21.617 ;
      VIA 35.316 21.6 Element_VIA34_1_2_58_52 ;
      VIA 35.316 21.6 Element_VIA23_1_3_36_36 ;
      VIA 35.316 21.06 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 21.043 35.361 21.077 ;
      VIA 35.316 21.06 Element_VIA34_1_2_58_52 ;
      VIA 35.316 21.06 Element_VIA23_1_3_36_36 ;
      VIA 35.316 20.52 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 20.503 35.361 20.537 ;
      VIA 35.316 20.52 Element_VIA34_1_2_58_52 ;
      VIA 35.316 20.52 Element_VIA23_1_3_36_36 ;
      VIA 35.316 19.98 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 19.963 35.361 19.997 ;
      VIA 35.316 19.98 Element_VIA34_1_2_58_52 ;
      VIA 35.316 19.98 Element_VIA23_1_3_36_36 ;
      VIA 35.316 19.44 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 19.423 35.361 19.457 ;
      VIA 35.316 19.44 Element_VIA34_1_2_58_52 ;
      VIA 35.316 19.44 Element_VIA23_1_3_36_36 ;
      VIA 35.316 18.9 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 18.883 35.361 18.917 ;
      VIA 35.316 18.9 Element_VIA34_1_2_58_52 ;
      VIA 35.316 18.9 Element_VIA23_1_3_36_36 ;
      VIA 35.316 18.36 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 18.343 35.361 18.377 ;
      VIA 35.316 18.36 Element_VIA34_1_2_58_52 ;
      VIA 35.316 18.36 Element_VIA23_1_3_36_36 ;
      VIA 35.316 17.82 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 17.803 35.361 17.837 ;
      VIA 35.316 17.82 Element_VIA34_1_2_58_52 ;
      VIA 35.316 17.82 Element_VIA23_1_3_36_36 ;
      VIA 35.316 17.28 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 17.263 35.361 17.297 ;
      VIA 35.316 17.28 Element_VIA34_1_2_58_52 ;
      VIA 35.316 17.28 Element_VIA23_1_3_36_36 ;
      VIA 35.316 16.74 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 16.723 35.361 16.757 ;
      VIA 35.316 16.74 Element_VIA34_1_2_58_52 ;
      VIA 35.316 16.74 Element_VIA23_1_3_36_36 ;
      VIA 35.316 16.2 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 16.183 35.361 16.217 ;
      VIA 35.316 16.2 Element_VIA34_1_2_58_52 ;
      VIA 35.316 16.2 Element_VIA23_1_3_36_36 ;
      VIA 35.316 15.66 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 15.643 35.361 15.677 ;
      VIA 35.316 15.66 Element_VIA34_1_2_58_52 ;
      VIA 35.316 15.66 Element_VIA23_1_3_36_36 ;
      VIA 35.316 15.12 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 15.103 35.361 15.137 ;
      VIA 35.316 15.12 Element_VIA34_1_2_58_52 ;
      VIA 35.316 15.12 Element_VIA23_1_3_36_36 ;
      VIA 35.316 14.58 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 14.563 35.361 14.597 ;
      VIA 35.316 14.58 Element_VIA34_1_2_58_52 ;
      VIA 35.316 14.58 Element_VIA23_1_3_36_36 ;
      VIA 35.316 14.04 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 14.023 35.361 14.057 ;
      VIA 35.316 14.04 Element_VIA34_1_2_58_52 ;
      VIA 35.316 14.04 Element_VIA23_1_3_36_36 ;
      VIA 35.316 13.5 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 13.483 35.361 13.517 ;
      VIA 35.316 13.5 Element_VIA34_1_2_58_52 ;
      VIA 35.316 13.5 Element_VIA23_1_3_36_36 ;
      VIA 35.316 12.96 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 12.943 35.361 12.977 ;
      VIA 35.316 12.96 Element_VIA34_1_2_58_52 ;
      VIA 35.316 12.96 Element_VIA23_1_3_36_36 ;
      VIA 35.316 12.42 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 12.403 35.361 12.437 ;
      VIA 35.316 12.42 Element_VIA34_1_2_58_52 ;
      VIA 35.316 12.42 Element_VIA23_1_3_36_36 ;
      VIA 35.316 11.88 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 11.863 35.361 11.897 ;
      VIA 35.316 11.88 Element_VIA34_1_2_58_52 ;
      VIA 35.316 11.88 Element_VIA23_1_3_36_36 ;
      VIA 35.316 11.34 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 11.323 35.361 11.357 ;
      VIA 35.316 11.34 Element_VIA34_1_2_58_52 ;
      VIA 35.316 11.34 Element_VIA23_1_3_36_36 ;
      VIA 35.316 10.8 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 10.783 35.361 10.817 ;
      VIA 35.316 10.8 Element_VIA34_1_2_58_52 ;
      VIA 35.316 10.8 Element_VIA23_1_3_36_36 ;
      VIA 35.316 10.26 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 10.243 35.361 10.277 ;
      VIA 35.316 10.26 Element_VIA34_1_2_58_52 ;
      VIA 35.316 10.26 Element_VIA23_1_3_36_36 ;
      VIA 35.316 9.72 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 9.703 35.361 9.737 ;
      VIA 35.316 9.72 Element_VIA34_1_2_58_52 ;
      VIA 35.316 9.72 Element_VIA23_1_3_36_36 ;
      VIA 35.316 9.18 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 9.163 35.361 9.197 ;
      VIA 35.316 9.18 Element_VIA34_1_2_58_52 ;
      VIA 35.316 9.18 Element_VIA23_1_3_36_36 ;
      VIA 35.316 8.64 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 8.623 35.361 8.657 ;
      VIA 35.316 8.64 Element_VIA34_1_2_58_52 ;
      VIA 35.316 8.64 Element_VIA23_1_3_36_36 ;
      VIA 35.316 8.1 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 8.083 35.361 8.117 ;
      VIA 35.316 8.1 Element_VIA34_1_2_58_52 ;
      VIA 35.316 8.1 Element_VIA23_1_3_36_36 ;
      VIA 35.316 7.56 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 7.543 35.361 7.577 ;
      VIA 35.316 7.56 Element_VIA34_1_2_58_52 ;
      VIA 35.316 7.56 Element_VIA23_1_3_36_36 ;
      VIA 35.316 7.02 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 7.003 35.361 7.037 ;
      VIA 35.316 7.02 Element_VIA34_1_2_58_52 ;
      VIA 35.316 7.02 Element_VIA23_1_3_36_36 ;
      VIA 35.316 6.48 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 6.463 35.361 6.497 ;
      VIA 35.316 6.48 Element_VIA34_1_2_58_52 ;
      VIA 35.316 6.48 Element_VIA23_1_3_36_36 ;
      VIA 35.316 5.94 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 5.923 35.361 5.957 ;
      VIA 35.316 5.94 Element_VIA34_1_2_58_52 ;
      VIA 35.316 5.94 Element_VIA23_1_3_36_36 ;
      VIA 35.316 5.4 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 5.383 35.361 5.417 ;
      VIA 35.316 5.4 Element_VIA34_1_2_58_52 ;
      VIA 35.316 5.4 Element_VIA23_1_3_36_36 ;
      VIA 35.316 4.86 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 4.843 35.361 4.877 ;
      VIA 35.316 4.86 Element_VIA34_1_2_58_52 ;
      VIA 35.316 4.86 Element_VIA23_1_3_36_36 ;
      VIA 35.316 4.32 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 4.303 35.361 4.337 ;
      VIA 35.316 4.32 Element_VIA34_1_2_58_52 ;
      VIA 35.316 4.32 Element_VIA23_1_3_36_36 ;
      VIA 35.316 3.78 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 3.763 35.361 3.797 ;
      VIA 35.316 3.78 Element_VIA34_1_2_58_52 ;
      VIA 35.316 3.78 Element_VIA23_1_3_36_36 ;
      VIA 35.316 3.24 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 3.223 35.361 3.257 ;
      VIA 35.316 3.24 Element_VIA34_1_2_58_52 ;
      VIA 35.316 3.24 Element_VIA23_1_3_36_36 ;
      VIA 35.316 2.7 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 2.683 35.361 2.717 ;
      VIA 35.316 2.7 Element_VIA34_1_2_58_52 ;
      VIA 35.316 2.7 Element_VIA23_1_3_36_36 ;
      VIA 35.316 2.16 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 2.143 35.361 2.177 ;
      VIA 35.316 2.16 Element_VIA34_1_2_58_52 ;
      VIA 35.316 2.16 Element_VIA23_1_3_36_36 ;
      VIA 35.316 1.62 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 1.603 35.361 1.637 ;
      VIA 35.316 1.62 Element_VIA34_1_2_58_52 ;
      VIA 35.316 1.62 Element_VIA23_1_3_36_36 ;
      VIA 35.316 1.08 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  35.271 1.063 35.361 1.097 ;
      VIA 35.316 1.08 Element_VIA34_1_2_58_52 ;
      VIA 35.316 1.08 Element_VIA23_1_3_36_36 ;
      VIA 32.34 42.12 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 42.103 32.385 42.137 ;
      VIA 32.34 42.12 Element_VIA34_1_2_58_52 ;
      VIA 32.34 42.12 Element_VIA23_1_3_36_36 ;
      VIA 32.34 41.58 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 41.563 32.385 41.597 ;
      VIA 32.34 41.58 Element_VIA34_1_2_58_52 ;
      VIA 32.34 41.58 Element_VIA23_1_3_36_36 ;
      VIA 32.34 41.04 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 41.023 32.385 41.057 ;
      VIA 32.34 41.04 Element_VIA34_1_2_58_52 ;
      VIA 32.34 41.04 Element_VIA23_1_3_36_36 ;
      VIA 32.34 40.5 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 40.483 32.385 40.517 ;
      VIA 32.34 40.5 Element_VIA34_1_2_58_52 ;
      VIA 32.34 40.5 Element_VIA23_1_3_36_36 ;
      VIA 32.34 39.96 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 39.943 32.385 39.977 ;
      VIA 32.34 39.96 Element_VIA34_1_2_58_52 ;
      VIA 32.34 39.96 Element_VIA23_1_3_36_36 ;
      VIA 32.34 39.42 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 39.403 32.385 39.437 ;
      VIA 32.34 39.42 Element_VIA34_1_2_58_52 ;
      VIA 32.34 39.42 Element_VIA23_1_3_36_36 ;
      VIA 32.34 38.88 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 38.863 32.385 38.897 ;
      VIA 32.34 38.88 Element_VIA34_1_2_58_52 ;
      VIA 32.34 38.88 Element_VIA23_1_3_36_36 ;
      VIA 32.34 38.34 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 38.323 32.385 38.357 ;
      VIA 32.34 38.34 Element_VIA34_1_2_58_52 ;
      VIA 32.34 38.34 Element_VIA23_1_3_36_36 ;
      VIA 32.34 37.8 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 37.783 32.385 37.817 ;
      VIA 32.34 37.8 Element_VIA34_1_2_58_52 ;
      VIA 32.34 37.8 Element_VIA23_1_3_36_36 ;
      VIA 32.34 37.26 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 37.243 32.385 37.277 ;
      VIA 32.34 37.26 Element_VIA34_1_2_58_52 ;
      VIA 32.34 37.26 Element_VIA23_1_3_36_36 ;
      VIA 32.34 36.72 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 36.703 32.385 36.737 ;
      VIA 32.34 36.72 Element_VIA34_1_2_58_52 ;
      VIA 32.34 36.72 Element_VIA23_1_3_36_36 ;
      VIA 32.34 36.18 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 36.163 32.385 36.197 ;
      VIA 32.34 36.18 Element_VIA34_1_2_58_52 ;
      VIA 32.34 36.18 Element_VIA23_1_3_36_36 ;
      VIA 32.34 35.64 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 35.623 32.385 35.657 ;
      VIA 32.34 35.64 Element_VIA34_1_2_58_52 ;
      VIA 32.34 35.64 Element_VIA23_1_3_36_36 ;
      VIA 32.34 35.1 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 35.083 32.385 35.117 ;
      VIA 32.34 35.1 Element_VIA34_1_2_58_52 ;
      VIA 32.34 35.1 Element_VIA23_1_3_36_36 ;
      VIA 32.34 34.56 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 34.543 32.385 34.577 ;
      VIA 32.34 34.56 Element_VIA34_1_2_58_52 ;
      VIA 32.34 34.56 Element_VIA23_1_3_36_36 ;
      VIA 32.34 34.02 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 34.003 32.385 34.037 ;
      VIA 32.34 34.02 Element_VIA34_1_2_58_52 ;
      VIA 32.34 34.02 Element_VIA23_1_3_36_36 ;
      VIA 32.34 33.48 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 33.463 32.385 33.497 ;
      VIA 32.34 33.48 Element_VIA34_1_2_58_52 ;
      VIA 32.34 33.48 Element_VIA23_1_3_36_36 ;
      VIA 32.34 32.94 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 32.923 32.385 32.957 ;
      VIA 32.34 32.94 Element_VIA34_1_2_58_52 ;
      VIA 32.34 32.94 Element_VIA23_1_3_36_36 ;
      VIA 32.34 32.4 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 32.383 32.385 32.417 ;
      VIA 32.34 32.4 Element_VIA34_1_2_58_52 ;
      VIA 32.34 32.4 Element_VIA23_1_3_36_36 ;
      VIA 32.34 31.86 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 31.843 32.385 31.877 ;
      VIA 32.34 31.86 Element_VIA34_1_2_58_52 ;
      VIA 32.34 31.86 Element_VIA23_1_3_36_36 ;
      VIA 32.34 31.32 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 31.303 32.385 31.337 ;
      VIA 32.34 31.32 Element_VIA34_1_2_58_52 ;
      VIA 32.34 31.32 Element_VIA23_1_3_36_36 ;
      VIA 32.34 30.78 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 30.763 32.385 30.797 ;
      VIA 32.34 30.78 Element_VIA34_1_2_58_52 ;
      VIA 32.34 30.78 Element_VIA23_1_3_36_36 ;
      VIA 32.34 30.24 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 30.223 32.385 30.257 ;
      VIA 32.34 30.24 Element_VIA34_1_2_58_52 ;
      VIA 32.34 30.24 Element_VIA23_1_3_36_36 ;
      VIA 32.34 29.7 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 29.683 32.385 29.717 ;
      VIA 32.34 29.7 Element_VIA34_1_2_58_52 ;
      VIA 32.34 29.7 Element_VIA23_1_3_36_36 ;
      VIA 32.34 29.16 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 29.143 32.385 29.177 ;
      VIA 32.34 29.16 Element_VIA34_1_2_58_52 ;
      VIA 32.34 29.16 Element_VIA23_1_3_36_36 ;
      VIA 32.34 28.62 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 28.603 32.385 28.637 ;
      VIA 32.34 28.62 Element_VIA34_1_2_58_52 ;
      VIA 32.34 28.62 Element_VIA23_1_3_36_36 ;
      VIA 32.34 28.08 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 28.063 32.385 28.097 ;
      VIA 32.34 28.08 Element_VIA34_1_2_58_52 ;
      VIA 32.34 28.08 Element_VIA23_1_3_36_36 ;
      VIA 32.34 27.54 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 27.523 32.385 27.557 ;
      VIA 32.34 27.54 Element_VIA34_1_2_58_52 ;
      VIA 32.34 27.54 Element_VIA23_1_3_36_36 ;
      VIA 32.34 27 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 26.983 32.385 27.017 ;
      VIA 32.34 27 Element_VIA34_1_2_58_52 ;
      VIA 32.34 27 Element_VIA23_1_3_36_36 ;
      VIA 32.34 26.46 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 26.443 32.385 26.477 ;
      VIA 32.34 26.46 Element_VIA34_1_2_58_52 ;
      VIA 32.34 26.46 Element_VIA23_1_3_36_36 ;
      VIA 32.34 25.92 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 25.903 32.385 25.937 ;
      VIA 32.34 25.92 Element_VIA34_1_2_58_52 ;
      VIA 32.34 25.92 Element_VIA23_1_3_36_36 ;
      VIA 32.34 25.38 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 25.363 32.385 25.397 ;
      VIA 32.34 25.38 Element_VIA34_1_2_58_52 ;
      VIA 32.34 25.38 Element_VIA23_1_3_36_36 ;
      VIA 32.34 24.84 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 24.823 32.385 24.857 ;
      VIA 32.34 24.84 Element_VIA34_1_2_58_52 ;
      VIA 32.34 24.84 Element_VIA23_1_3_36_36 ;
      VIA 32.34 24.3 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 24.283 32.385 24.317 ;
      VIA 32.34 24.3 Element_VIA34_1_2_58_52 ;
      VIA 32.34 24.3 Element_VIA23_1_3_36_36 ;
      VIA 32.34 23.76 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 23.743 32.385 23.777 ;
      VIA 32.34 23.76 Element_VIA34_1_2_58_52 ;
      VIA 32.34 23.76 Element_VIA23_1_3_36_36 ;
      VIA 32.34 23.22 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 23.203 32.385 23.237 ;
      VIA 32.34 23.22 Element_VIA34_1_2_58_52 ;
      VIA 32.34 23.22 Element_VIA23_1_3_36_36 ;
      VIA 32.34 22.68 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 22.663 32.385 22.697 ;
      VIA 32.34 22.68 Element_VIA34_1_2_58_52 ;
      VIA 32.34 22.68 Element_VIA23_1_3_36_36 ;
      VIA 32.34 22.14 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 22.123 32.385 22.157 ;
      VIA 32.34 22.14 Element_VIA34_1_2_58_52 ;
      VIA 32.34 22.14 Element_VIA23_1_3_36_36 ;
      VIA 32.34 21.6 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 21.583 32.385 21.617 ;
      VIA 32.34 21.6 Element_VIA34_1_2_58_52 ;
      VIA 32.34 21.6 Element_VIA23_1_3_36_36 ;
      VIA 32.34 21.06 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 21.043 32.385 21.077 ;
      VIA 32.34 21.06 Element_VIA34_1_2_58_52 ;
      VIA 32.34 21.06 Element_VIA23_1_3_36_36 ;
      VIA 32.34 20.52 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 20.503 32.385 20.537 ;
      VIA 32.34 20.52 Element_VIA34_1_2_58_52 ;
      VIA 32.34 20.52 Element_VIA23_1_3_36_36 ;
      VIA 32.34 19.98 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 19.963 32.385 19.997 ;
      VIA 32.34 19.98 Element_VIA34_1_2_58_52 ;
      VIA 32.34 19.98 Element_VIA23_1_3_36_36 ;
      VIA 32.34 19.44 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 19.423 32.385 19.457 ;
      VIA 32.34 19.44 Element_VIA34_1_2_58_52 ;
      VIA 32.34 19.44 Element_VIA23_1_3_36_36 ;
      VIA 32.34 18.9 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 18.883 32.385 18.917 ;
      VIA 32.34 18.9 Element_VIA34_1_2_58_52 ;
      VIA 32.34 18.9 Element_VIA23_1_3_36_36 ;
      VIA 32.34 18.36 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 18.343 32.385 18.377 ;
      VIA 32.34 18.36 Element_VIA34_1_2_58_52 ;
      VIA 32.34 18.36 Element_VIA23_1_3_36_36 ;
      VIA 32.34 17.82 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 17.803 32.385 17.837 ;
      VIA 32.34 17.82 Element_VIA34_1_2_58_52 ;
      VIA 32.34 17.82 Element_VIA23_1_3_36_36 ;
      VIA 32.34 17.28 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 17.263 32.385 17.297 ;
      VIA 32.34 17.28 Element_VIA34_1_2_58_52 ;
      VIA 32.34 17.28 Element_VIA23_1_3_36_36 ;
      VIA 32.34 16.74 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 16.723 32.385 16.757 ;
      VIA 32.34 16.74 Element_VIA34_1_2_58_52 ;
      VIA 32.34 16.74 Element_VIA23_1_3_36_36 ;
      VIA 32.34 16.2 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 16.183 32.385 16.217 ;
      VIA 32.34 16.2 Element_VIA34_1_2_58_52 ;
      VIA 32.34 16.2 Element_VIA23_1_3_36_36 ;
      VIA 32.34 15.66 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 15.643 32.385 15.677 ;
      VIA 32.34 15.66 Element_VIA34_1_2_58_52 ;
      VIA 32.34 15.66 Element_VIA23_1_3_36_36 ;
      VIA 32.34 15.12 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 15.103 32.385 15.137 ;
      VIA 32.34 15.12 Element_VIA34_1_2_58_52 ;
      VIA 32.34 15.12 Element_VIA23_1_3_36_36 ;
      VIA 32.34 14.58 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 14.563 32.385 14.597 ;
      VIA 32.34 14.58 Element_VIA34_1_2_58_52 ;
      VIA 32.34 14.58 Element_VIA23_1_3_36_36 ;
      VIA 32.34 14.04 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 14.023 32.385 14.057 ;
      VIA 32.34 14.04 Element_VIA34_1_2_58_52 ;
      VIA 32.34 14.04 Element_VIA23_1_3_36_36 ;
      VIA 32.34 13.5 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 13.483 32.385 13.517 ;
      VIA 32.34 13.5 Element_VIA34_1_2_58_52 ;
      VIA 32.34 13.5 Element_VIA23_1_3_36_36 ;
      VIA 32.34 12.96 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 12.943 32.385 12.977 ;
      VIA 32.34 12.96 Element_VIA34_1_2_58_52 ;
      VIA 32.34 12.96 Element_VIA23_1_3_36_36 ;
      VIA 32.34 12.42 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 12.403 32.385 12.437 ;
      VIA 32.34 12.42 Element_VIA34_1_2_58_52 ;
      VIA 32.34 12.42 Element_VIA23_1_3_36_36 ;
      VIA 32.34 11.88 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 11.863 32.385 11.897 ;
      VIA 32.34 11.88 Element_VIA34_1_2_58_52 ;
      VIA 32.34 11.88 Element_VIA23_1_3_36_36 ;
      VIA 32.34 11.34 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 11.323 32.385 11.357 ;
      VIA 32.34 11.34 Element_VIA34_1_2_58_52 ;
      VIA 32.34 11.34 Element_VIA23_1_3_36_36 ;
      VIA 32.34 10.8 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 10.783 32.385 10.817 ;
      VIA 32.34 10.8 Element_VIA34_1_2_58_52 ;
      VIA 32.34 10.8 Element_VIA23_1_3_36_36 ;
      VIA 32.34 10.26 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 10.243 32.385 10.277 ;
      VIA 32.34 10.26 Element_VIA34_1_2_58_52 ;
      VIA 32.34 10.26 Element_VIA23_1_3_36_36 ;
      VIA 32.34 9.72 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 9.703 32.385 9.737 ;
      VIA 32.34 9.72 Element_VIA34_1_2_58_52 ;
      VIA 32.34 9.72 Element_VIA23_1_3_36_36 ;
      VIA 32.34 9.18 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 9.163 32.385 9.197 ;
      VIA 32.34 9.18 Element_VIA34_1_2_58_52 ;
      VIA 32.34 9.18 Element_VIA23_1_3_36_36 ;
      VIA 32.34 8.64 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 8.623 32.385 8.657 ;
      VIA 32.34 8.64 Element_VIA34_1_2_58_52 ;
      VIA 32.34 8.64 Element_VIA23_1_3_36_36 ;
      VIA 32.34 8.1 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 8.083 32.385 8.117 ;
      VIA 32.34 8.1 Element_VIA34_1_2_58_52 ;
      VIA 32.34 8.1 Element_VIA23_1_3_36_36 ;
      VIA 32.34 7.56 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 7.543 32.385 7.577 ;
      VIA 32.34 7.56 Element_VIA34_1_2_58_52 ;
      VIA 32.34 7.56 Element_VIA23_1_3_36_36 ;
      VIA 32.34 7.02 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 7.003 32.385 7.037 ;
      VIA 32.34 7.02 Element_VIA34_1_2_58_52 ;
      VIA 32.34 7.02 Element_VIA23_1_3_36_36 ;
      VIA 32.34 6.48 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 6.463 32.385 6.497 ;
      VIA 32.34 6.48 Element_VIA34_1_2_58_52 ;
      VIA 32.34 6.48 Element_VIA23_1_3_36_36 ;
      VIA 32.34 5.94 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 5.923 32.385 5.957 ;
      VIA 32.34 5.94 Element_VIA34_1_2_58_52 ;
      VIA 32.34 5.94 Element_VIA23_1_3_36_36 ;
      VIA 32.34 5.4 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 5.383 32.385 5.417 ;
      VIA 32.34 5.4 Element_VIA34_1_2_58_52 ;
      VIA 32.34 5.4 Element_VIA23_1_3_36_36 ;
      VIA 32.34 4.86 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 4.843 32.385 4.877 ;
      VIA 32.34 4.86 Element_VIA34_1_2_58_52 ;
      VIA 32.34 4.86 Element_VIA23_1_3_36_36 ;
      VIA 32.34 4.32 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 4.303 32.385 4.337 ;
      VIA 32.34 4.32 Element_VIA34_1_2_58_52 ;
      VIA 32.34 4.32 Element_VIA23_1_3_36_36 ;
      VIA 32.34 3.78 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 3.763 32.385 3.797 ;
      VIA 32.34 3.78 Element_VIA34_1_2_58_52 ;
      VIA 32.34 3.78 Element_VIA23_1_3_36_36 ;
      VIA 32.34 3.24 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 3.223 32.385 3.257 ;
      VIA 32.34 3.24 Element_VIA34_1_2_58_52 ;
      VIA 32.34 3.24 Element_VIA23_1_3_36_36 ;
      VIA 32.34 2.7 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 2.683 32.385 2.717 ;
      VIA 32.34 2.7 Element_VIA34_1_2_58_52 ;
      VIA 32.34 2.7 Element_VIA23_1_3_36_36 ;
      VIA 32.34 2.16 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 2.143 32.385 2.177 ;
      VIA 32.34 2.16 Element_VIA34_1_2_58_52 ;
      VIA 32.34 2.16 Element_VIA23_1_3_36_36 ;
      VIA 32.34 1.62 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 1.603 32.385 1.637 ;
      VIA 32.34 1.62 Element_VIA34_1_2_58_52 ;
      VIA 32.34 1.62 Element_VIA23_1_3_36_36 ;
      VIA 32.34 1.08 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  32.295 1.063 32.385 1.097 ;
      VIA 32.34 1.08 Element_VIA34_1_2_58_52 ;
      VIA 32.34 1.08 Element_VIA23_1_3_36_36 ;
      VIA 29.364 42.12 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 42.103 29.409 42.137 ;
      VIA 29.364 42.12 Element_VIA34_1_2_58_52 ;
      VIA 29.364 42.12 Element_VIA23_1_3_36_36 ;
      VIA 29.364 41.58 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 41.563 29.409 41.597 ;
      VIA 29.364 41.58 Element_VIA34_1_2_58_52 ;
      VIA 29.364 41.58 Element_VIA23_1_3_36_36 ;
      VIA 29.364 41.04 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 41.023 29.409 41.057 ;
      VIA 29.364 41.04 Element_VIA34_1_2_58_52 ;
      VIA 29.364 41.04 Element_VIA23_1_3_36_36 ;
      VIA 29.364 40.5 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 40.483 29.409 40.517 ;
      VIA 29.364 40.5 Element_VIA34_1_2_58_52 ;
      VIA 29.364 40.5 Element_VIA23_1_3_36_36 ;
      VIA 29.364 39.96 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 39.943 29.409 39.977 ;
      VIA 29.364 39.96 Element_VIA34_1_2_58_52 ;
      VIA 29.364 39.96 Element_VIA23_1_3_36_36 ;
      VIA 29.364 39.42 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 39.403 29.409 39.437 ;
      VIA 29.364 39.42 Element_VIA34_1_2_58_52 ;
      VIA 29.364 39.42 Element_VIA23_1_3_36_36 ;
      VIA 29.364 38.88 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 38.863 29.409 38.897 ;
      VIA 29.364 38.88 Element_VIA34_1_2_58_52 ;
      VIA 29.364 38.88 Element_VIA23_1_3_36_36 ;
      VIA 29.364 38.34 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 38.323 29.409 38.357 ;
      VIA 29.364 38.34 Element_VIA34_1_2_58_52 ;
      VIA 29.364 38.34 Element_VIA23_1_3_36_36 ;
      VIA 29.364 37.8 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 37.783 29.409 37.817 ;
      VIA 29.364 37.8 Element_VIA34_1_2_58_52 ;
      VIA 29.364 37.8 Element_VIA23_1_3_36_36 ;
      VIA 29.364 37.26 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 37.243 29.409 37.277 ;
      VIA 29.364 37.26 Element_VIA34_1_2_58_52 ;
      VIA 29.364 37.26 Element_VIA23_1_3_36_36 ;
      VIA 29.364 36.72 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 36.703 29.409 36.737 ;
      VIA 29.364 36.72 Element_VIA34_1_2_58_52 ;
      VIA 29.364 36.72 Element_VIA23_1_3_36_36 ;
      VIA 29.364 36.18 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 36.163 29.409 36.197 ;
      VIA 29.364 36.18 Element_VIA34_1_2_58_52 ;
      VIA 29.364 36.18 Element_VIA23_1_3_36_36 ;
      VIA 29.364 35.64 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 35.623 29.409 35.657 ;
      VIA 29.364 35.64 Element_VIA34_1_2_58_52 ;
      VIA 29.364 35.64 Element_VIA23_1_3_36_36 ;
      VIA 29.364 35.1 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 35.083 29.409 35.117 ;
      VIA 29.364 35.1 Element_VIA34_1_2_58_52 ;
      VIA 29.364 35.1 Element_VIA23_1_3_36_36 ;
      VIA 29.364 34.56 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 34.543 29.409 34.577 ;
      VIA 29.364 34.56 Element_VIA34_1_2_58_52 ;
      VIA 29.364 34.56 Element_VIA23_1_3_36_36 ;
      VIA 29.364 34.02 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 34.003 29.409 34.037 ;
      VIA 29.364 34.02 Element_VIA34_1_2_58_52 ;
      VIA 29.364 34.02 Element_VIA23_1_3_36_36 ;
      VIA 29.364 33.48 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 33.463 29.409 33.497 ;
      VIA 29.364 33.48 Element_VIA34_1_2_58_52 ;
      VIA 29.364 33.48 Element_VIA23_1_3_36_36 ;
      VIA 29.364 32.94 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 32.923 29.409 32.957 ;
      VIA 29.364 32.94 Element_VIA34_1_2_58_52 ;
      VIA 29.364 32.94 Element_VIA23_1_3_36_36 ;
      VIA 29.364 32.4 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 32.383 29.409 32.417 ;
      VIA 29.364 32.4 Element_VIA34_1_2_58_52 ;
      VIA 29.364 32.4 Element_VIA23_1_3_36_36 ;
      VIA 29.364 31.86 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 31.843 29.409 31.877 ;
      VIA 29.364 31.86 Element_VIA34_1_2_58_52 ;
      VIA 29.364 31.86 Element_VIA23_1_3_36_36 ;
      VIA 29.364 31.32 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 31.303 29.409 31.337 ;
      VIA 29.364 31.32 Element_VIA34_1_2_58_52 ;
      VIA 29.364 31.32 Element_VIA23_1_3_36_36 ;
      VIA 29.364 30.78 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 30.763 29.409 30.797 ;
      VIA 29.364 30.78 Element_VIA34_1_2_58_52 ;
      VIA 29.364 30.78 Element_VIA23_1_3_36_36 ;
      VIA 29.364 30.24 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 30.223 29.409 30.257 ;
      VIA 29.364 30.24 Element_VIA34_1_2_58_52 ;
      VIA 29.364 30.24 Element_VIA23_1_3_36_36 ;
      VIA 29.364 29.7 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 29.683 29.409 29.717 ;
      VIA 29.364 29.7 Element_VIA34_1_2_58_52 ;
      VIA 29.364 29.7 Element_VIA23_1_3_36_36 ;
      VIA 29.364 29.16 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 29.143 29.409 29.177 ;
      VIA 29.364 29.16 Element_VIA34_1_2_58_52 ;
      VIA 29.364 29.16 Element_VIA23_1_3_36_36 ;
      VIA 29.364 28.62 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 28.603 29.409 28.637 ;
      VIA 29.364 28.62 Element_VIA34_1_2_58_52 ;
      VIA 29.364 28.62 Element_VIA23_1_3_36_36 ;
      VIA 29.364 28.08 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 28.063 29.409 28.097 ;
      VIA 29.364 28.08 Element_VIA34_1_2_58_52 ;
      VIA 29.364 28.08 Element_VIA23_1_3_36_36 ;
      VIA 29.364 27.54 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 27.523 29.409 27.557 ;
      VIA 29.364 27.54 Element_VIA34_1_2_58_52 ;
      VIA 29.364 27.54 Element_VIA23_1_3_36_36 ;
      VIA 29.364 27 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 26.983 29.409 27.017 ;
      VIA 29.364 27 Element_VIA34_1_2_58_52 ;
      VIA 29.364 27 Element_VIA23_1_3_36_36 ;
      VIA 29.364 26.46 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 26.443 29.409 26.477 ;
      VIA 29.364 26.46 Element_VIA34_1_2_58_52 ;
      VIA 29.364 26.46 Element_VIA23_1_3_36_36 ;
      VIA 29.364 25.92 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 25.903 29.409 25.937 ;
      VIA 29.364 25.92 Element_VIA34_1_2_58_52 ;
      VIA 29.364 25.92 Element_VIA23_1_3_36_36 ;
      VIA 29.364 25.38 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 25.363 29.409 25.397 ;
      VIA 29.364 25.38 Element_VIA34_1_2_58_52 ;
      VIA 29.364 25.38 Element_VIA23_1_3_36_36 ;
      VIA 29.364 24.84 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 24.823 29.409 24.857 ;
      VIA 29.364 24.84 Element_VIA34_1_2_58_52 ;
      VIA 29.364 24.84 Element_VIA23_1_3_36_36 ;
      VIA 29.364 24.3 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 24.283 29.409 24.317 ;
      VIA 29.364 24.3 Element_VIA34_1_2_58_52 ;
      VIA 29.364 24.3 Element_VIA23_1_3_36_36 ;
      VIA 29.364 23.76 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 23.743 29.409 23.777 ;
      VIA 29.364 23.76 Element_VIA34_1_2_58_52 ;
      VIA 29.364 23.76 Element_VIA23_1_3_36_36 ;
      VIA 29.364 23.22 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 23.203 29.409 23.237 ;
      VIA 29.364 23.22 Element_VIA34_1_2_58_52 ;
      VIA 29.364 23.22 Element_VIA23_1_3_36_36 ;
      VIA 29.364 22.68 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 22.663 29.409 22.697 ;
      VIA 29.364 22.68 Element_VIA34_1_2_58_52 ;
      VIA 29.364 22.68 Element_VIA23_1_3_36_36 ;
      VIA 29.364 22.14 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 22.123 29.409 22.157 ;
      VIA 29.364 22.14 Element_VIA34_1_2_58_52 ;
      VIA 29.364 22.14 Element_VIA23_1_3_36_36 ;
      VIA 29.364 21.6 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 21.583 29.409 21.617 ;
      VIA 29.364 21.6 Element_VIA34_1_2_58_52 ;
      VIA 29.364 21.6 Element_VIA23_1_3_36_36 ;
      VIA 29.364 21.06 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 21.043 29.409 21.077 ;
      VIA 29.364 21.06 Element_VIA34_1_2_58_52 ;
      VIA 29.364 21.06 Element_VIA23_1_3_36_36 ;
      VIA 29.364 20.52 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 20.503 29.409 20.537 ;
      VIA 29.364 20.52 Element_VIA34_1_2_58_52 ;
      VIA 29.364 20.52 Element_VIA23_1_3_36_36 ;
      VIA 29.364 19.98 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 19.963 29.409 19.997 ;
      VIA 29.364 19.98 Element_VIA34_1_2_58_52 ;
      VIA 29.364 19.98 Element_VIA23_1_3_36_36 ;
      VIA 29.364 19.44 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 19.423 29.409 19.457 ;
      VIA 29.364 19.44 Element_VIA34_1_2_58_52 ;
      VIA 29.364 19.44 Element_VIA23_1_3_36_36 ;
      VIA 29.364 18.9 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 18.883 29.409 18.917 ;
      VIA 29.364 18.9 Element_VIA34_1_2_58_52 ;
      VIA 29.364 18.9 Element_VIA23_1_3_36_36 ;
      VIA 29.364 18.36 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 18.343 29.409 18.377 ;
      VIA 29.364 18.36 Element_VIA34_1_2_58_52 ;
      VIA 29.364 18.36 Element_VIA23_1_3_36_36 ;
      VIA 29.364 17.82 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 17.803 29.409 17.837 ;
      VIA 29.364 17.82 Element_VIA34_1_2_58_52 ;
      VIA 29.364 17.82 Element_VIA23_1_3_36_36 ;
      VIA 29.364 17.28 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 17.263 29.409 17.297 ;
      VIA 29.364 17.28 Element_VIA34_1_2_58_52 ;
      VIA 29.364 17.28 Element_VIA23_1_3_36_36 ;
      VIA 29.364 16.74 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 16.723 29.409 16.757 ;
      VIA 29.364 16.74 Element_VIA34_1_2_58_52 ;
      VIA 29.364 16.74 Element_VIA23_1_3_36_36 ;
      VIA 29.364 16.2 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 16.183 29.409 16.217 ;
      VIA 29.364 16.2 Element_VIA34_1_2_58_52 ;
      VIA 29.364 16.2 Element_VIA23_1_3_36_36 ;
      VIA 29.364 15.66 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 15.643 29.409 15.677 ;
      VIA 29.364 15.66 Element_VIA34_1_2_58_52 ;
      VIA 29.364 15.66 Element_VIA23_1_3_36_36 ;
      VIA 29.364 15.12 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 15.103 29.409 15.137 ;
      VIA 29.364 15.12 Element_VIA34_1_2_58_52 ;
      VIA 29.364 15.12 Element_VIA23_1_3_36_36 ;
      VIA 29.364 14.58 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 14.563 29.409 14.597 ;
      VIA 29.364 14.58 Element_VIA34_1_2_58_52 ;
      VIA 29.364 14.58 Element_VIA23_1_3_36_36 ;
      VIA 29.364 14.04 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 14.023 29.409 14.057 ;
      VIA 29.364 14.04 Element_VIA34_1_2_58_52 ;
      VIA 29.364 14.04 Element_VIA23_1_3_36_36 ;
      VIA 29.364 13.5 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 13.483 29.409 13.517 ;
      VIA 29.364 13.5 Element_VIA34_1_2_58_52 ;
      VIA 29.364 13.5 Element_VIA23_1_3_36_36 ;
      VIA 29.364 12.96 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 12.943 29.409 12.977 ;
      VIA 29.364 12.96 Element_VIA34_1_2_58_52 ;
      VIA 29.364 12.96 Element_VIA23_1_3_36_36 ;
      VIA 29.364 12.42 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 12.403 29.409 12.437 ;
      VIA 29.364 12.42 Element_VIA34_1_2_58_52 ;
      VIA 29.364 12.42 Element_VIA23_1_3_36_36 ;
      VIA 29.364 11.88 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 11.863 29.409 11.897 ;
      VIA 29.364 11.88 Element_VIA34_1_2_58_52 ;
      VIA 29.364 11.88 Element_VIA23_1_3_36_36 ;
      VIA 29.364 11.34 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 11.323 29.409 11.357 ;
      VIA 29.364 11.34 Element_VIA34_1_2_58_52 ;
      VIA 29.364 11.34 Element_VIA23_1_3_36_36 ;
      VIA 29.364 10.8 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 10.783 29.409 10.817 ;
      VIA 29.364 10.8 Element_VIA34_1_2_58_52 ;
      VIA 29.364 10.8 Element_VIA23_1_3_36_36 ;
      VIA 29.364 10.26 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 10.243 29.409 10.277 ;
      VIA 29.364 10.26 Element_VIA34_1_2_58_52 ;
      VIA 29.364 10.26 Element_VIA23_1_3_36_36 ;
      VIA 29.364 9.72 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 9.703 29.409 9.737 ;
      VIA 29.364 9.72 Element_VIA34_1_2_58_52 ;
      VIA 29.364 9.72 Element_VIA23_1_3_36_36 ;
      VIA 29.364 9.18 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 9.163 29.409 9.197 ;
      VIA 29.364 9.18 Element_VIA34_1_2_58_52 ;
      VIA 29.364 9.18 Element_VIA23_1_3_36_36 ;
      VIA 29.364 8.64 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 8.623 29.409 8.657 ;
      VIA 29.364 8.64 Element_VIA34_1_2_58_52 ;
      VIA 29.364 8.64 Element_VIA23_1_3_36_36 ;
      VIA 29.364 8.1 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 8.083 29.409 8.117 ;
      VIA 29.364 8.1 Element_VIA34_1_2_58_52 ;
      VIA 29.364 8.1 Element_VIA23_1_3_36_36 ;
      VIA 29.364 7.56 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 7.543 29.409 7.577 ;
      VIA 29.364 7.56 Element_VIA34_1_2_58_52 ;
      VIA 29.364 7.56 Element_VIA23_1_3_36_36 ;
      VIA 29.364 7.02 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 7.003 29.409 7.037 ;
      VIA 29.364 7.02 Element_VIA34_1_2_58_52 ;
      VIA 29.364 7.02 Element_VIA23_1_3_36_36 ;
      VIA 29.364 6.48 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 6.463 29.409 6.497 ;
      VIA 29.364 6.48 Element_VIA34_1_2_58_52 ;
      VIA 29.364 6.48 Element_VIA23_1_3_36_36 ;
      VIA 29.364 5.94 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 5.923 29.409 5.957 ;
      VIA 29.364 5.94 Element_VIA34_1_2_58_52 ;
      VIA 29.364 5.94 Element_VIA23_1_3_36_36 ;
      VIA 29.364 5.4 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 5.383 29.409 5.417 ;
      VIA 29.364 5.4 Element_VIA34_1_2_58_52 ;
      VIA 29.364 5.4 Element_VIA23_1_3_36_36 ;
      VIA 29.364 4.86 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 4.843 29.409 4.877 ;
      VIA 29.364 4.86 Element_VIA34_1_2_58_52 ;
      VIA 29.364 4.86 Element_VIA23_1_3_36_36 ;
      VIA 29.364 4.32 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 4.303 29.409 4.337 ;
      VIA 29.364 4.32 Element_VIA34_1_2_58_52 ;
      VIA 29.364 4.32 Element_VIA23_1_3_36_36 ;
      VIA 29.364 3.78 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 3.763 29.409 3.797 ;
      VIA 29.364 3.78 Element_VIA34_1_2_58_52 ;
      VIA 29.364 3.78 Element_VIA23_1_3_36_36 ;
      VIA 29.364 3.24 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 3.223 29.409 3.257 ;
      VIA 29.364 3.24 Element_VIA34_1_2_58_52 ;
      VIA 29.364 3.24 Element_VIA23_1_3_36_36 ;
      VIA 29.364 2.7 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 2.683 29.409 2.717 ;
      VIA 29.364 2.7 Element_VIA34_1_2_58_52 ;
      VIA 29.364 2.7 Element_VIA23_1_3_36_36 ;
      VIA 29.364 2.16 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 2.143 29.409 2.177 ;
      VIA 29.364 2.16 Element_VIA34_1_2_58_52 ;
      VIA 29.364 2.16 Element_VIA23_1_3_36_36 ;
      VIA 29.364 1.62 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 1.603 29.409 1.637 ;
      VIA 29.364 1.62 Element_VIA34_1_2_58_52 ;
      VIA 29.364 1.62 Element_VIA23_1_3_36_36 ;
      VIA 29.364 1.08 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  29.319 1.063 29.409 1.097 ;
      VIA 29.364 1.08 Element_VIA34_1_2_58_52 ;
      VIA 29.364 1.08 Element_VIA23_1_3_36_36 ;
      VIA 26.388 42.12 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 42.103 26.433 42.137 ;
      VIA 26.388 42.12 Element_VIA34_1_2_58_52 ;
      VIA 26.388 42.12 Element_VIA23_1_3_36_36 ;
      VIA 26.388 41.58 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 41.563 26.433 41.597 ;
      VIA 26.388 41.58 Element_VIA34_1_2_58_52 ;
      VIA 26.388 41.58 Element_VIA23_1_3_36_36 ;
      VIA 26.388 41.04 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 41.023 26.433 41.057 ;
      VIA 26.388 41.04 Element_VIA34_1_2_58_52 ;
      VIA 26.388 41.04 Element_VIA23_1_3_36_36 ;
      VIA 26.388 40.5 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 40.483 26.433 40.517 ;
      VIA 26.388 40.5 Element_VIA34_1_2_58_52 ;
      VIA 26.388 40.5 Element_VIA23_1_3_36_36 ;
      VIA 26.388 39.96 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 39.943 26.433 39.977 ;
      VIA 26.388 39.96 Element_VIA34_1_2_58_52 ;
      VIA 26.388 39.96 Element_VIA23_1_3_36_36 ;
      VIA 26.388 39.42 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 39.403 26.433 39.437 ;
      VIA 26.388 39.42 Element_VIA34_1_2_58_52 ;
      VIA 26.388 39.42 Element_VIA23_1_3_36_36 ;
      VIA 26.388 38.88 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 38.863 26.433 38.897 ;
      VIA 26.388 38.88 Element_VIA34_1_2_58_52 ;
      VIA 26.388 38.88 Element_VIA23_1_3_36_36 ;
      VIA 26.388 38.34 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 38.323 26.433 38.357 ;
      VIA 26.388 38.34 Element_VIA34_1_2_58_52 ;
      VIA 26.388 38.34 Element_VIA23_1_3_36_36 ;
      VIA 26.388 37.8 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 37.783 26.433 37.817 ;
      VIA 26.388 37.8 Element_VIA34_1_2_58_52 ;
      VIA 26.388 37.8 Element_VIA23_1_3_36_36 ;
      VIA 26.388 37.26 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 37.243 26.433 37.277 ;
      VIA 26.388 37.26 Element_VIA34_1_2_58_52 ;
      VIA 26.388 37.26 Element_VIA23_1_3_36_36 ;
      VIA 26.388 36.72 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 36.703 26.433 36.737 ;
      VIA 26.388 36.72 Element_VIA34_1_2_58_52 ;
      VIA 26.388 36.72 Element_VIA23_1_3_36_36 ;
      VIA 26.388 36.18 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 36.163 26.433 36.197 ;
      VIA 26.388 36.18 Element_VIA34_1_2_58_52 ;
      VIA 26.388 36.18 Element_VIA23_1_3_36_36 ;
      VIA 26.388 35.64 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 35.623 26.433 35.657 ;
      VIA 26.388 35.64 Element_VIA34_1_2_58_52 ;
      VIA 26.388 35.64 Element_VIA23_1_3_36_36 ;
      VIA 26.388 35.1 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 35.083 26.433 35.117 ;
      VIA 26.388 35.1 Element_VIA34_1_2_58_52 ;
      VIA 26.388 35.1 Element_VIA23_1_3_36_36 ;
      VIA 26.388 34.56 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 34.543 26.433 34.577 ;
      VIA 26.388 34.56 Element_VIA34_1_2_58_52 ;
      VIA 26.388 34.56 Element_VIA23_1_3_36_36 ;
      VIA 26.388 34.02 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 34.003 26.433 34.037 ;
      VIA 26.388 34.02 Element_VIA34_1_2_58_52 ;
      VIA 26.388 34.02 Element_VIA23_1_3_36_36 ;
      VIA 26.388 33.48 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 33.463 26.433 33.497 ;
      VIA 26.388 33.48 Element_VIA34_1_2_58_52 ;
      VIA 26.388 33.48 Element_VIA23_1_3_36_36 ;
      VIA 26.388 32.94 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 32.923 26.433 32.957 ;
      VIA 26.388 32.94 Element_VIA34_1_2_58_52 ;
      VIA 26.388 32.94 Element_VIA23_1_3_36_36 ;
      VIA 26.388 32.4 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 32.383 26.433 32.417 ;
      VIA 26.388 32.4 Element_VIA34_1_2_58_52 ;
      VIA 26.388 32.4 Element_VIA23_1_3_36_36 ;
      VIA 26.388 31.86 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 31.843 26.433 31.877 ;
      VIA 26.388 31.86 Element_VIA34_1_2_58_52 ;
      VIA 26.388 31.86 Element_VIA23_1_3_36_36 ;
      VIA 26.388 31.32 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 31.303 26.433 31.337 ;
      VIA 26.388 31.32 Element_VIA34_1_2_58_52 ;
      VIA 26.388 31.32 Element_VIA23_1_3_36_36 ;
      VIA 26.388 30.78 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 30.763 26.433 30.797 ;
      VIA 26.388 30.78 Element_VIA34_1_2_58_52 ;
      VIA 26.388 30.78 Element_VIA23_1_3_36_36 ;
      VIA 26.388 30.24 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 30.223 26.433 30.257 ;
      VIA 26.388 30.24 Element_VIA34_1_2_58_52 ;
      VIA 26.388 30.24 Element_VIA23_1_3_36_36 ;
      VIA 26.388 29.7 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 29.683 26.433 29.717 ;
      VIA 26.388 29.7 Element_VIA34_1_2_58_52 ;
      VIA 26.388 29.7 Element_VIA23_1_3_36_36 ;
      VIA 26.388 29.16 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 29.143 26.433 29.177 ;
      VIA 26.388 29.16 Element_VIA34_1_2_58_52 ;
      VIA 26.388 29.16 Element_VIA23_1_3_36_36 ;
      VIA 26.388 28.62 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 28.603 26.433 28.637 ;
      VIA 26.388 28.62 Element_VIA34_1_2_58_52 ;
      VIA 26.388 28.62 Element_VIA23_1_3_36_36 ;
      VIA 26.388 28.08 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 28.063 26.433 28.097 ;
      VIA 26.388 28.08 Element_VIA34_1_2_58_52 ;
      VIA 26.388 28.08 Element_VIA23_1_3_36_36 ;
      VIA 26.388 27.54 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 27.523 26.433 27.557 ;
      VIA 26.388 27.54 Element_VIA34_1_2_58_52 ;
      VIA 26.388 27.54 Element_VIA23_1_3_36_36 ;
      VIA 26.388 27 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 26.983 26.433 27.017 ;
      VIA 26.388 27 Element_VIA34_1_2_58_52 ;
      VIA 26.388 27 Element_VIA23_1_3_36_36 ;
      VIA 26.388 26.46 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 26.443 26.433 26.477 ;
      VIA 26.388 26.46 Element_VIA34_1_2_58_52 ;
      VIA 26.388 26.46 Element_VIA23_1_3_36_36 ;
      VIA 26.388 25.92 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 25.903 26.433 25.937 ;
      VIA 26.388 25.92 Element_VIA34_1_2_58_52 ;
      VIA 26.388 25.92 Element_VIA23_1_3_36_36 ;
      VIA 26.388 25.38 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 25.363 26.433 25.397 ;
      VIA 26.388 25.38 Element_VIA34_1_2_58_52 ;
      VIA 26.388 25.38 Element_VIA23_1_3_36_36 ;
      VIA 26.388 24.84 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 24.823 26.433 24.857 ;
      VIA 26.388 24.84 Element_VIA34_1_2_58_52 ;
      VIA 26.388 24.84 Element_VIA23_1_3_36_36 ;
      VIA 26.388 24.3 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 24.283 26.433 24.317 ;
      VIA 26.388 24.3 Element_VIA34_1_2_58_52 ;
      VIA 26.388 24.3 Element_VIA23_1_3_36_36 ;
      VIA 26.388 23.76 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 23.743 26.433 23.777 ;
      VIA 26.388 23.76 Element_VIA34_1_2_58_52 ;
      VIA 26.388 23.76 Element_VIA23_1_3_36_36 ;
      VIA 26.388 23.22 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 23.203 26.433 23.237 ;
      VIA 26.388 23.22 Element_VIA34_1_2_58_52 ;
      VIA 26.388 23.22 Element_VIA23_1_3_36_36 ;
      VIA 26.388 22.68 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 22.663 26.433 22.697 ;
      VIA 26.388 22.68 Element_VIA34_1_2_58_52 ;
      VIA 26.388 22.68 Element_VIA23_1_3_36_36 ;
      VIA 26.388 22.14 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 22.123 26.433 22.157 ;
      VIA 26.388 22.14 Element_VIA34_1_2_58_52 ;
      VIA 26.388 22.14 Element_VIA23_1_3_36_36 ;
      VIA 26.388 21.6 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 21.583 26.433 21.617 ;
      VIA 26.388 21.6 Element_VIA34_1_2_58_52 ;
      VIA 26.388 21.6 Element_VIA23_1_3_36_36 ;
      VIA 26.388 21.06 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 21.043 26.433 21.077 ;
      VIA 26.388 21.06 Element_VIA34_1_2_58_52 ;
      VIA 26.388 21.06 Element_VIA23_1_3_36_36 ;
      VIA 26.388 20.52 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 20.503 26.433 20.537 ;
      VIA 26.388 20.52 Element_VIA34_1_2_58_52 ;
      VIA 26.388 20.52 Element_VIA23_1_3_36_36 ;
      VIA 26.388 19.98 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 19.963 26.433 19.997 ;
      VIA 26.388 19.98 Element_VIA34_1_2_58_52 ;
      VIA 26.388 19.98 Element_VIA23_1_3_36_36 ;
      VIA 26.388 19.44 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 19.423 26.433 19.457 ;
      VIA 26.388 19.44 Element_VIA34_1_2_58_52 ;
      VIA 26.388 19.44 Element_VIA23_1_3_36_36 ;
      VIA 26.388 18.9 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 18.883 26.433 18.917 ;
      VIA 26.388 18.9 Element_VIA34_1_2_58_52 ;
      VIA 26.388 18.9 Element_VIA23_1_3_36_36 ;
      VIA 26.388 18.36 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 18.343 26.433 18.377 ;
      VIA 26.388 18.36 Element_VIA34_1_2_58_52 ;
      VIA 26.388 18.36 Element_VIA23_1_3_36_36 ;
      VIA 26.388 17.82 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 17.803 26.433 17.837 ;
      VIA 26.388 17.82 Element_VIA34_1_2_58_52 ;
      VIA 26.388 17.82 Element_VIA23_1_3_36_36 ;
      VIA 26.388 17.28 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 17.263 26.433 17.297 ;
      VIA 26.388 17.28 Element_VIA34_1_2_58_52 ;
      VIA 26.388 17.28 Element_VIA23_1_3_36_36 ;
      VIA 26.388 16.74 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 16.723 26.433 16.757 ;
      VIA 26.388 16.74 Element_VIA34_1_2_58_52 ;
      VIA 26.388 16.74 Element_VIA23_1_3_36_36 ;
      VIA 26.388 16.2 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 16.183 26.433 16.217 ;
      VIA 26.388 16.2 Element_VIA34_1_2_58_52 ;
      VIA 26.388 16.2 Element_VIA23_1_3_36_36 ;
      VIA 26.388 15.66 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 15.643 26.433 15.677 ;
      VIA 26.388 15.66 Element_VIA34_1_2_58_52 ;
      VIA 26.388 15.66 Element_VIA23_1_3_36_36 ;
      VIA 26.388 15.12 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 15.103 26.433 15.137 ;
      VIA 26.388 15.12 Element_VIA34_1_2_58_52 ;
      VIA 26.388 15.12 Element_VIA23_1_3_36_36 ;
      VIA 26.388 14.58 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 14.563 26.433 14.597 ;
      VIA 26.388 14.58 Element_VIA34_1_2_58_52 ;
      VIA 26.388 14.58 Element_VIA23_1_3_36_36 ;
      VIA 26.388 14.04 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 14.023 26.433 14.057 ;
      VIA 26.388 14.04 Element_VIA34_1_2_58_52 ;
      VIA 26.388 14.04 Element_VIA23_1_3_36_36 ;
      VIA 26.388 13.5 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 13.483 26.433 13.517 ;
      VIA 26.388 13.5 Element_VIA34_1_2_58_52 ;
      VIA 26.388 13.5 Element_VIA23_1_3_36_36 ;
      VIA 26.388 12.96 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 12.943 26.433 12.977 ;
      VIA 26.388 12.96 Element_VIA34_1_2_58_52 ;
      VIA 26.388 12.96 Element_VIA23_1_3_36_36 ;
      VIA 26.388 12.42 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 12.403 26.433 12.437 ;
      VIA 26.388 12.42 Element_VIA34_1_2_58_52 ;
      VIA 26.388 12.42 Element_VIA23_1_3_36_36 ;
      VIA 26.388 11.88 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 11.863 26.433 11.897 ;
      VIA 26.388 11.88 Element_VIA34_1_2_58_52 ;
      VIA 26.388 11.88 Element_VIA23_1_3_36_36 ;
      VIA 26.388 11.34 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 11.323 26.433 11.357 ;
      VIA 26.388 11.34 Element_VIA34_1_2_58_52 ;
      VIA 26.388 11.34 Element_VIA23_1_3_36_36 ;
      VIA 26.388 10.8 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 10.783 26.433 10.817 ;
      VIA 26.388 10.8 Element_VIA34_1_2_58_52 ;
      VIA 26.388 10.8 Element_VIA23_1_3_36_36 ;
      VIA 26.388 10.26 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 10.243 26.433 10.277 ;
      VIA 26.388 10.26 Element_VIA34_1_2_58_52 ;
      VIA 26.388 10.26 Element_VIA23_1_3_36_36 ;
      VIA 26.388 9.72 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 9.703 26.433 9.737 ;
      VIA 26.388 9.72 Element_VIA34_1_2_58_52 ;
      VIA 26.388 9.72 Element_VIA23_1_3_36_36 ;
      VIA 26.388 9.18 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 9.163 26.433 9.197 ;
      VIA 26.388 9.18 Element_VIA34_1_2_58_52 ;
      VIA 26.388 9.18 Element_VIA23_1_3_36_36 ;
      VIA 26.388 8.64 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 8.623 26.433 8.657 ;
      VIA 26.388 8.64 Element_VIA34_1_2_58_52 ;
      VIA 26.388 8.64 Element_VIA23_1_3_36_36 ;
      VIA 26.388 8.1 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 8.083 26.433 8.117 ;
      VIA 26.388 8.1 Element_VIA34_1_2_58_52 ;
      VIA 26.388 8.1 Element_VIA23_1_3_36_36 ;
      VIA 26.388 7.56 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 7.543 26.433 7.577 ;
      VIA 26.388 7.56 Element_VIA34_1_2_58_52 ;
      VIA 26.388 7.56 Element_VIA23_1_3_36_36 ;
      VIA 26.388 7.02 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 7.003 26.433 7.037 ;
      VIA 26.388 7.02 Element_VIA34_1_2_58_52 ;
      VIA 26.388 7.02 Element_VIA23_1_3_36_36 ;
      VIA 26.388 6.48 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 6.463 26.433 6.497 ;
      VIA 26.388 6.48 Element_VIA34_1_2_58_52 ;
      VIA 26.388 6.48 Element_VIA23_1_3_36_36 ;
      VIA 26.388 5.94 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 5.923 26.433 5.957 ;
      VIA 26.388 5.94 Element_VIA34_1_2_58_52 ;
      VIA 26.388 5.94 Element_VIA23_1_3_36_36 ;
      VIA 26.388 5.4 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 5.383 26.433 5.417 ;
      VIA 26.388 5.4 Element_VIA34_1_2_58_52 ;
      VIA 26.388 5.4 Element_VIA23_1_3_36_36 ;
      VIA 26.388 4.86 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 4.843 26.433 4.877 ;
      VIA 26.388 4.86 Element_VIA34_1_2_58_52 ;
      VIA 26.388 4.86 Element_VIA23_1_3_36_36 ;
      VIA 26.388 4.32 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 4.303 26.433 4.337 ;
      VIA 26.388 4.32 Element_VIA34_1_2_58_52 ;
      VIA 26.388 4.32 Element_VIA23_1_3_36_36 ;
      VIA 26.388 3.78 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 3.763 26.433 3.797 ;
      VIA 26.388 3.78 Element_VIA34_1_2_58_52 ;
      VIA 26.388 3.78 Element_VIA23_1_3_36_36 ;
      VIA 26.388 3.24 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 3.223 26.433 3.257 ;
      VIA 26.388 3.24 Element_VIA34_1_2_58_52 ;
      VIA 26.388 3.24 Element_VIA23_1_3_36_36 ;
      VIA 26.388 2.7 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 2.683 26.433 2.717 ;
      VIA 26.388 2.7 Element_VIA34_1_2_58_52 ;
      VIA 26.388 2.7 Element_VIA23_1_3_36_36 ;
      VIA 26.388 2.16 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 2.143 26.433 2.177 ;
      VIA 26.388 2.16 Element_VIA34_1_2_58_52 ;
      VIA 26.388 2.16 Element_VIA23_1_3_36_36 ;
      VIA 26.388 1.62 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 1.603 26.433 1.637 ;
      VIA 26.388 1.62 Element_VIA34_1_2_58_52 ;
      VIA 26.388 1.62 Element_VIA23_1_3_36_36 ;
      VIA 26.388 1.08 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  26.343 1.063 26.433 1.097 ;
      VIA 26.388 1.08 Element_VIA34_1_2_58_52 ;
      VIA 26.388 1.08 Element_VIA23_1_3_36_36 ;
      VIA 23.412 42.12 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 42.103 23.457 42.137 ;
      VIA 23.412 42.12 Element_VIA34_1_2_58_52 ;
      VIA 23.412 42.12 Element_VIA23_1_3_36_36 ;
      VIA 23.412 41.58 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 41.563 23.457 41.597 ;
      VIA 23.412 41.58 Element_VIA34_1_2_58_52 ;
      VIA 23.412 41.58 Element_VIA23_1_3_36_36 ;
      VIA 23.412 41.04 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 41.023 23.457 41.057 ;
      VIA 23.412 41.04 Element_VIA34_1_2_58_52 ;
      VIA 23.412 41.04 Element_VIA23_1_3_36_36 ;
      VIA 23.412 40.5 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 40.483 23.457 40.517 ;
      VIA 23.412 40.5 Element_VIA34_1_2_58_52 ;
      VIA 23.412 40.5 Element_VIA23_1_3_36_36 ;
      VIA 23.412 39.96 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 39.943 23.457 39.977 ;
      VIA 23.412 39.96 Element_VIA34_1_2_58_52 ;
      VIA 23.412 39.96 Element_VIA23_1_3_36_36 ;
      VIA 23.412 39.42 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 39.403 23.457 39.437 ;
      VIA 23.412 39.42 Element_VIA34_1_2_58_52 ;
      VIA 23.412 39.42 Element_VIA23_1_3_36_36 ;
      VIA 23.412 38.88 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 38.863 23.457 38.897 ;
      VIA 23.412 38.88 Element_VIA34_1_2_58_52 ;
      VIA 23.412 38.88 Element_VIA23_1_3_36_36 ;
      VIA 23.412 38.34 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 38.323 23.457 38.357 ;
      VIA 23.412 38.34 Element_VIA34_1_2_58_52 ;
      VIA 23.412 38.34 Element_VIA23_1_3_36_36 ;
      VIA 23.412 37.8 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 37.783 23.457 37.817 ;
      VIA 23.412 37.8 Element_VIA34_1_2_58_52 ;
      VIA 23.412 37.8 Element_VIA23_1_3_36_36 ;
      VIA 23.412 37.26 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 37.243 23.457 37.277 ;
      VIA 23.412 37.26 Element_VIA34_1_2_58_52 ;
      VIA 23.412 37.26 Element_VIA23_1_3_36_36 ;
      VIA 23.412 36.72 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 36.703 23.457 36.737 ;
      VIA 23.412 36.72 Element_VIA34_1_2_58_52 ;
      VIA 23.412 36.72 Element_VIA23_1_3_36_36 ;
      VIA 23.412 36.18 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 36.163 23.457 36.197 ;
      VIA 23.412 36.18 Element_VIA34_1_2_58_52 ;
      VIA 23.412 36.18 Element_VIA23_1_3_36_36 ;
      VIA 23.412 35.64 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 35.623 23.457 35.657 ;
      VIA 23.412 35.64 Element_VIA34_1_2_58_52 ;
      VIA 23.412 35.64 Element_VIA23_1_3_36_36 ;
      VIA 23.412 35.1 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 35.083 23.457 35.117 ;
      VIA 23.412 35.1 Element_VIA34_1_2_58_52 ;
      VIA 23.412 35.1 Element_VIA23_1_3_36_36 ;
      VIA 23.412 34.56 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 34.543 23.457 34.577 ;
      VIA 23.412 34.56 Element_VIA34_1_2_58_52 ;
      VIA 23.412 34.56 Element_VIA23_1_3_36_36 ;
      VIA 23.412 34.02 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 34.003 23.457 34.037 ;
      VIA 23.412 34.02 Element_VIA34_1_2_58_52 ;
      VIA 23.412 34.02 Element_VIA23_1_3_36_36 ;
      VIA 23.412 33.48 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 33.463 23.457 33.497 ;
      VIA 23.412 33.48 Element_VIA34_1_2_58_52 ;
      VIA 23.412 33.48 Element_VIA23_1_3_36_36 ;
      VIA 23.412 32.94 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 32.923 23.457 32.957 ;
      VIA 23.412 32.94 Element_VIA34_1_2_58_52 ;
      VIA 23.412 32.94 Element_VIA23_1_3_36_36 ;
      VIA 23.412 32.4 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 32.383 23.457 32.417 ;
      VIA 23.412 32.4 Element_VIA34_1_2_58_52 ;
      VIA 23.412 32.4 Element_VIA23_1_3_36_36 ;
      VIA 23.412 31.86 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 31.843 23.457 31.877 ;
      VIA 23.412 31.86 Element_VIA34_1_2_58_52 ;
      VIA 23.412 31.86 Element_VIA23_1_3_36_36 ;
      VIA 23.412 31.32 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 31.303 23.457 31.337 ;
      VIA 23.412 31.32 Element_VIA34_1_2_58_52 ;
      VIA 23.412 31.32 Element_VIA23_1_3_36_36 ;
      VIA 23.412 30.78 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 30.763 23.457 30.797 ;
      VIA 23.412 30.78 Element_VIA34_1_2_58_52 ;
      VIA 23.412 30.78 Element_VIA23_1_3_36_36 ;
      VIA 23.412 30.24 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 30.223 23.457 30.257 ;
      VIA 23.412 30.24 Element_VIA34_1_2_58_52 ;
      VIA 23.412 30.24 Element_VIA23_1_3_36_36 ;
      VIA 23.412 29.7 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 29.683 23.457 29.717 ;
      VIA 23.412 29.7 Element_VIA34_1_2_58_52 ;
      VIA 23.412 29.7 Element_VIA23_1_3_36_36 ;
      VIA 23.412 29.16 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 29.143 23.457 29.177 ;
      VIA 23.412 29.16 Element_VIA34_1_2_58_52 ;
      VIA 23.412 29.16 Element_VIA23_1_3_36_36 ;
      VIA 23.412 28.62 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 28.603 23.457 28.637 ;
      VIA 23.412 28.62 Element_VIA34_1_2_58_52 ;
      VIA 23.412 28.62 Element_VIA23_1_3_36_36 ;
      VIA 23.412 28.08 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 28.063 23.457 28.097 ;
      VIA 23.412 28.08 Element_VIA34_1_2_58_52 ;
      VIA 23.412 28.08 Element_VIA23_1_3_36_36 ;
      VIA 23.412 27.54 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 27.523 23.457 27.557 ;
      VIA 23.412 27.54 Element_VIA34_1_2_58_52 ;
      VIA 23.412 27.54 Element_VIA23_1_3_36_36 ;
      VIA 23.412 27 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 26.983 23.457 27.017 ;
      VIA 23.412 27 Element_VIA34_1_2_58_52 ;
      VIA 23.412 27 Element_VIA23_1_3_36_36 ;
      VIA 23.412 26.46 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 26.443 23.457 26.477 ;
      VIA 23.412 26.46 Element_VIA34_1_2_58_52 ;
      VIA 23.412 26.46 Element_VIA23_1_3_36_36 ;
      VIA 23.412 25.92 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 25.903 23.457 25.937 ;
      VIA 23.412 25.92 Element_VIA34_1_2_58_52 ;
      VIA 23.412 25.92 Element_VIA23_1_3_36_36 ;
      VIA 23.412 25.38 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 25.363 23.457 25.397 ;
      VIA 23.412 25.38 Element_VIA34_1_2_58_52 ;
      VIA 23.412 25.38 Element_VIA23_1_3_36_36 ;
      VIA 23.412 24.84 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 24.823 23.457 24.857 ;
      VIA 23.412 24.84 Element_VIA34_1_2_58_52 ;
      VIA 23.412 24.84 Element_VIA23_1_3_36_36 ;
      VIA 23.412 24.3 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 24.283 23.457 24.317 ;
      VIA 23.412 24.3 Element_VIA34_1_2_58_52 ;
      VIA 23.412 24.3 Element_VIA23_1_3_36_36 ;
      VIA 23.412 23.76 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 23.743 23.457 23.777 ;
      VIA 23.412 23.76 Element_VIA34_1_2_58_52 ;
      VIA 23.412 23.76 Element_VIA23_1_3_36_36 ;
      VIA 23.412 23.22 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 23.203 23.457 23.237 ;
      VIA 23.412 23.22 Element_VIA34_1_2_58_52 ;
      VIA 23.412 23.22 Element_VIA23_1_3_36_36 ;
      VIA 23.412 22.68 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 22.663 23.457 22.697 ;
      VIA 23.412 22.68 Element_VIA34_1_2_58_52 ;
      VIA 23.412 22.68 Element_VIA23_1_3_36_36 ;
      VIA 23.412 22.14 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 22.123 23.457 22.157 ;
      VIA 23.412 22.14 Element_VIA34_1_2_58_52 ;
      VIA 23.412 22.14 Element_VIA23_1_3_36_36 ;
      VIA 23.412 21.6 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 21.583 23.457 21.617 ;
      VIA 23.412 21.6 Element_VIA34_1_2_58_52 ;
      VIA 23.412 21.6 Element_VIA23_1_3_36_36 ;
      VIA 23.412 21.06 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 21.043 23.457 21.077 ;
      VIA 23.412 21.06 Element_VIA34_1_2_58_52 ;
      VIA 23.412 21.06 Element_VIA23_1_3_36_36 ;
      VIA 23.412 20.52 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 20.503 23.457 20.537 ;
      VIA 23.412 20.52 Element_VIA34_1_2_58_52 ;
      VIA 23.412 20.52 Element_VIA23_1_3_36_36 ;
      VIA 23.412 19.98 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 19.963 23.457 19.997 ;
      VIA 23.412 19.98 Element_VIA34_1_2_58_52 ;
      VIA 23.412 19.98 Element_VIA23_1_3_36_36 ;
      VIA 23.412 19.44 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 19.423 23.457 19.457 ;
      VIA 23.412 19.44 Element_VIA34_1_2_58_52 ;
      VIA 23.412 19.44 Element_VIA23_1_3_36_36 ;
      VIA 23.412 18.9 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 18.883 23.457 18.917 ;
      VIA 23.412 18.9 Element_VIA34_1_2_58_52 ;
      VIA 23.412 18.9 Element_VIA23_1_3_36_36 ;
      VIA 23.412 18.36 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 18.343 23.457 18.377 ;
      VIA 23.412 18.36 Element_VIA34_1_2_58_52 ;
      VIA 23.412 18.36 Element_VIA23_1_3_36_36 ;
      VIA 23.412 17.82 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 17.803 23.457 17.837 ;
      VIA 23.412 17.82 Element_VIA34_1_2_58_52 ;
      VIA 23.412 17.82 Element_VIA23_1_3_36_36 ;
      VIA 23.412 17.28 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 17.263 23.457 17.297 ;
      VIA 23.412 17.28 Element_VIA34_1_2_58_52 ;
      VIA 23.412 17.28 Element_VIA23_1_3_36_36 ;
      VIA 23.412 16.74 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 16.723 23.457 16.757 ;
      VIA 23.412 16.74 Element_VIA34_1_2_58_52 ;
      VIA 23.412 16.74 Element_VIA23_1_3_36_36 ;
      VIA 23.412 16.2 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 16.183 23.457 16.217 ;
      VIA 23.412 16.2 Element_VIA34_1_2_58_52 ;
      VIA 23.412 16.2 Element_VIA23_1_3_36_36 ;
      VIA 23.412 15.66 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 15.643 23.457 15.677 ;
      VIA 23.412 15.66 Element_VIA34_1_2_58_52 ;
      VIA 23.412 15.66 Element_VIA23_1_3_36_36 ;
      VIA 23.412 15.12 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 15.103 23.457 15.137 ;
      VIA 23.412 15.12 Element_VIA34_1_2_58_52 ;
      VIA 23.412 15.12 Element_VIA23_1_3_36_36 ;
      VIA 23.412 14.58 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 14.563 23.457 14.597 ;
      VIA 23.412 14.58 Element_VIA34_1_2_58_52 ;
      VIA 23.412 14.58 Element_VIA23_1_3_36_36 ;
      VIA 23.412 14.04 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 14.023 23.457 14.057 ;
      VIA 23.412 14.04 Element_VIA34_1_2_58_52 ;
      VIA 23.412 14.04 Element_VIA23_1_3_36_36 ;
      VIA 23.412 13.5 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 13.483 23.457 13.517 ;
      VIA 23.412 13.5 Element_VIA34_1_2_58_52 ;
      VIA 23.412 13.5 Element_VIA23_1_3_36_36 ;
      VIA 23.412 12.96 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 12.943 23.457 12.977 ;
      VIA 23.412 12.96 Element_VIA34_1_2_58_52 ;
      VIA 23.412 12.96 Element_VIA23_1_3_36_36 ;
      VIA 23.412 12.42 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 12.403 23.457 12.437 ;
      VIA 23.412 12.42 Element_VIA34_1_2_58_52 ;
      VIA 23.412 12.42 Element_VIA23_1_3_36_36 ;
      VIA 23.412 11.88 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 11.863 23.457 11.897 ;
      VIA 23.412 11.88 Element_VIA34_1_2_58_52 ;
      VIA 23.412 11.88 Element_VIA23_1_3_36_36 ;
      VIA 23.412 11.34 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 11.323 23.457 11.357 ;
      VIA 23.412 11.34 Element_VIA34_1_2_58_52 ;
      VIA 23.412 11.34 Element_VIA23_1_3_36_36 ;
      VIA 23.412 10.8 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 10.783 23.457 10.817 ;
      VIA 23.412 10.8 Element_VIA34_1_2_58_52 ;
      VIA 23.412 10.8 Element_VIA23_1_3_36_36 ;
      VIA 23.412 10.26 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 10.243 23.457 10.277 ;
      VIA 23.412 10.26 Element_VIA34_1_2_58_52 ;
      VIA 23.412 10.26 Element_VIA23_1_3_36_36 ;
      VIA 23.412 9.72 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 9.703 23.457 9.737 ;
      VIA 23.412 9.72 Element_VIA34_1_2_58_52 ;
      VIA 23.412 9.72 Element_VIA23_1_3_36_36 ;
      VIA 23.412 9.18 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 9.163 23.457 9.197 ;
      VIA 23.412 9.18 Element_VIA34_1_2_58_52 ;
      VIA 23.412 9.18 Element_VIA23_1_3_36_36 ;
      VIA 23.412 8.64 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 8.623 23.457 8.657 ;
      VIA 23.412 8.64 Element_VIA34_1_2_58_52 ;
      VIA 23.412 8.64 Element_VIA23_1_3_36_36 ;
      VIA 23.412 8.1 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 8.083 23.457 8.117 ;
      VIA 23.412 8.1 Element_VIA34_1_2_58_52 ;
      VIA 23.412 8.1 Element_VIA23_1_3_36_36 ;
      VIA 23.412 7.56 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 7.543 23.457 7.577 ;
      VIA 23.412 7.56 Element_VIA34_1_2_58_52 ;
      VIA 23.412 7.56 Element_VIA23_1_3_36_36 ;
      VIA 23.412 7.02 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 7.003 23.457 7.037 ;
      VIA 23.412 7.02 Element_VIA34_1_2_58_52 ;
      VIA 23.412 7.02 Element_VIA23_1_3_36_36 ;
      VIA 23.412 6.48 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 6.463 23.457 6.497 ;
      VIA 23.412 6.48 Element_VIA34_1_2_58_52 ;
      VIA 23.412 6.48 Element_VIA23_1_3_36_36 ;
      VIA 23.412 5.94 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 5.923 23.457 5.957 ;
      VIA 23.412 5.94 Element_VIA34_1_2_58_52 ;
      VIA 23.412 5.94 Element_VIA23_1_3_36_36 ;
      VIA 23.412 5.4 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 5.383 23.457 5.417 ;
      VIA 23.412 5.4 Element_VIA34_1_2_58_52 ;
      VIA 23.412 5.4 Element_VIA23_1_3_36_36 ;
      VIA 23.412 4.86 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 4.843 23.457 4.877 ;
      VIA 23.412 4.86 Element_VIA34_1_2_58_52 ;
      VIA 23.412 4.86 Element_VIA23_1_3_36_36 ;
      VIA 23.412 4.32 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 4.303 23.457 4.337 ;
      VIA 23.412 4.32 Element_VIA34_1_2_58_52 ;
      VIA 23.412 4.32 Element_VIA23_1_3_36_36 ;
      VIA 23.412 3.78 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 3.763 23.457 3.797 ;
      VIA 23.412 3.78 Element_VIA34_1_2_58_52 ;
      VIA 23.412 3.78 Element_VIA23_1_3_36_36 ;
      VIA 23.412 3.24 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 3.223 23.457 3.257 ;
      VIA 23.412 3.24 Element_VIA34_1_2_58_52 ;
      VIA 23.412 3.24 Element_VIA23_1_3_36_36 ;
      VIA 23.412 2.7 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 2.683 23.457 2.717 ;
      VIA 23.412 2.7 Element_VIA34_1_2_58_52 ;
      VIA 23.412 2.7 Element_VIA23_1_3_36_36 ;
      VIA 23.412 2.16 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 2.143 23.457 2.177 ;
      VIA 23.412 2.16 Element_VIA34_1_2_58_52 ;
      VIA 23.412 2.16 Element_VIA23_1_3_36_36 ;
      VIA 23.412 1.62 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 1.603 23.457 1.637 ;
      VIA 23.412 1.62 Element_VIA34_1_2_58_52 ;
      VIA 23.412 1.62 Element_VIA23_1_3_36_36 ;
      VIA 23.412 1.08 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  23.367 1.063 23.457 1.097 ;
      VIA 23.412 1.08 Element_VIA34_1_2_58_52 ;
      VIA 23.412 1.08 Element_VIA23_1_3_36_36 ;
      VIA 20.436 42.12 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 42.103 20.481 42.137 ;
      VIA 20.436 42.12 Element_VIA34_1_2_58_52 ;
      VIA 20.436 42.12 Element_VIA23_1_3_36_36 ;
      VIA 20.436 41.58 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 41.563 20.481 41.597 ;
      VIA 20.436 41.58 Element_VIA34_1_2_58_52 ;
      VIA 20.436 41.58 Element_VIA23_1_3_36_36 ;
      VIA 20.436 41.04 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 41.023 20.481 41.057 ;
      VIA 20.436 41.04 Element_VIA34_1_2_58_52 ;
      VIA 20.436 41.04 Element_VIA23_1_3_36_36 ;
      VIA 20.436 40.5 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 40.483 20.481 40.517 ;
      VIA 20.436 40.5 Element_VIA34_1_2_58_52 ;
      VIA 20.436 40.5 Element_VIA23_1_3_36_36 ;
      VIA 20.436 39.96 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 39.943 20.481 39.977 ;
      VIA 20.436 39.96 Element_VIA34_1_2_58_52 ;
      VIA 20.436 39.96 Element_VIA23_1_3_36_36 ;
      VIA 20.436 39.42 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 39.403 20.481 39.437 ;
      VIA 20.436 39.42 Element_VIA34_1_2_58_52 ;
      VIA 20.436 39.42 Element_VIA23_1_3_36_36 ;
      VIA 20.436 38.88 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 38.863 20.481 38.897 ;
      VIA 20.436 38.88 Element_VIA34_1_2_58_52 ;
      VIA 20.436 38.88 Element_VIA23_1_3_36_36 ;
      VIA 20.436 38.34 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 38.323 20.481 38.357 ;
      VIA 20.436 38.34 Element_VIA34_1_2_58_52 ;
      VIA 20.436 38.34 Element_VIA23_1_3_36_36 ;
      VIA 20.436 37.8 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 37.783 20.481 37.817 ;
      VIA 20.436 37.8 Element_VIA34_1_2_58_52 ;
      VIA 20.436 37.8 Element_VIA23_1_3_36_36 ;
      VIA 20.436 37.26 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 37.243 20.481 37.277 ;
      VIA 20.436 37.26 Element_VIA34_1_2_58_52 ;
      VIA 20.436 37.26 Element_VIA23_1_3_36_36 ;
      VIA 20.436 36.72 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 36.703 20.481 36.737 ;
      VIA 20.436 36.72 Element_VIA34_1_2_58_52 ;
      VIA 20.436 36.72 Element_VIA23_1_3_36_36 ;
      VIA 20.436 36.18 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 36.163 20.481 36.197 ;
      VIA 20.436 36.18 Element_VIA34_1_2_58_52 ;
      VIA 20.436 36.18 Element_VIA23_1_3_36_36 ;
      VIA 20.436 35.64 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 35.623 20.481 35.657 ;
      VIA 20.436 35.64 Element_VIA34_1_2_58_52 ;
      VIA 20.436 35.64 Element_VIA23_1_3_36_36 ;
      VIA 20.436 35.1 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 35.083 20.481 35.117 ;
      VIA 20.436 35.1 Element_VIA34_1_2_58_52 ;
      VIA 20.436 35.1 Element_VIA23_1_3_36_36 ;
      VIA 20.436 34.56 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 34.543 20.481 34.577 ;
      VIA 20.436 34.56 Element_VIA34_1_2_58_52 ;
      VIA 20.436 34.56 Element_VIA23_1_3_36_36 ;
      VIA 20.436 34.02 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 34.003 20.481 34.037 ;
      VIA 20.436 34.02 Element_VIA34_1_2_58_52 ;
      VIA 20.436 34.02 Element_VIA23_1_3_36_36 ;
      VIA 20.436 33.48 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 33.463 20.481 33.497 ;
      VIA 20.436 33.48 Element_VIA34_1_2_58_52 ;
      VIA 20.436 33.48 Element_VIA23_1_3_36_36 ;
      VIA 20.436 32.94 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 32.923 20.481 32.957 ;
      VIA 20.436 32.94 Element_VIA34_1_2_58_52 ;
      VIA 20.436 32.94 Element_VIA23_1_3_36_36 ;
      VIA 20.436 32.4 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 32.383 20.481 32.417 ;
      VIA 20.436 32.4 Element_VIA34_1_2_58_52 ;
      VIA 20.436 32.4 Element_VIA23_1_3_36_36 ;
      VIA 20.436 31.86 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 31.843 20.481 31.877 ;
      VIA 20.436 31.86 Element_VIA34_1_2_58_52 ;
      VIA 20.436 31.86 Element_VIA23_1_3_36_36 ;
      VIA 20.436 31.32 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 31.303 20.481 31.337 ;
      VIA 20.436 31.32 Element_VIA34_1_2_58_52 ;
      VIA 20.436 31.32 Element_VIA23_1_3_36_36 ;
      VIA 20.436 30.78 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 30.763 20.481 30.797 ;
      VIA 20.436 30.78 Element_VIA34_1_2_58_52 ;
      VIA 20.436 30.78 Element_VIA23_1_3_36_36 ;
      VIA 20.436 30.24 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 30.223 20.481 30.257 ;
      VIA 20.436 30.24 Element_VIA34_1_2_58_52 ;
      VIA 20.436 30.24 Element_VIA23_1_3_36_36 ;
      VIA 20.436 29.7 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 29.683 20.481 29.717 ;
      VIA 20.436 29.7 Element_VIA34_1_2_58_52 ;
      VIA 20.436 29.7 Element_VIA23_1_3_36_36 ;
      VIA 20.436 29.16 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 29.143 20.481 29.177 ;
      VIA 20.436 29.16 Element_VIA34_1_2_58_52 ;
      VIA 20.436 29.16 Element_VIA23_1_3_36_36 ;
      VIA 20.436 28.62 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 28.603 20.481 28.637 ;
      VIA 20.436 28.62 Element_VIA34_1_2_58_52 ;
      VIA 20.436 28.62 Element_VIA23_1_3_36_36 ;
      VIA 20.436 28.08 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 28.063 20.481 28.097 ;
      VIA 20.436 28.08 Element_VIA34_1_2_58_52 ;
      VIA 20.436 28.08 Element_VIA23_1_3_36_36 ;
      VIA 20.436 27.54 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 27.523 20.481 27.557 ;
      VIA 20.436 27.54 Element_VIA34_1_2_58_52 ;
      VIA 20.436 27.54 Element_VIA23_1_3_36_36 ;
      VIA 20.436 27 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 26.983 20.481 27.017 ;
      VIA 20.436 27 Element_VIA34_1_2_58_52 ;
      VIA 20.436 27 Element_VIA23_1_3_36_36 ;
      VIA 20.436 26.46 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 26.443 20.481 26.477 ;
      VIA 20.436 26.46 Element_VIA34_1_2_58_52 ;
      VIA 20.436 26.46 Element_VIA23_1_3_36_36 ;
      VIA 20.436 25.92 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 25.903 20.481 25.937 ;
      VIA 20.436 25.92 Element_VIA34_1_2_58_52 ;
      VIA 20.436 25.92 Element_VIA23_1_3_36_36 ;
      VIA 20.436 25.38 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 25.363 20.481 25.397 ;
      VIA 20.436 25.38 Element_VIA34_1_2_58_52 ;
      VIA 20.436 25.38 Element_VIA23_1_3_36_36 ;
      VIA 20.436 24.84 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 24.823 20.481 24.857 ;
      VIA 20.436 24.84 Element_VIA34_1_2_58_52 ;
      VIA 20.436 24.84 Element_VIA23_1_3_36_36 ;
      VIA 20.436 24.3 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 24.283 20.481 24.317 ;
      VIA 20.436 24.3 Element_VIA34_1_2_58_52 ;
      VIA 20.436 24.3 Element_VIA23_1_3_36_36 ;
      VIA 20.436 23.76 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 23.743 20.481 23.777 ;
      VIA 20.436 23.76 Element_VIA34_1_2_58_52 ;
      VIA 20.436 23.76 Element_VIA23_1_3_36_36 ;
      VIA 20.436 23.22 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 23.203 20.481 23.237 ;
      VIA 20.436 23.22 Element_VIA34_1_2_58_52 ;
      VIA 20.436 23.22 Element_VIA23_1_3_36_36 ;
      VIA 20.436 22.68 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 22.663 20.481 22.697 ;
      VIA 20.436 22.68 Element_VIA34_1_2_58_52 ;
      VIA 20.436 22.68 Element_VIA23_1_3_36_36 ;
      VIA 20.436 22.14 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 22.123 20.481 22.157 ;
      VIA 20.436 22.14 Element_VIA34_1_2_58_52 ;
      VIA 20.436 22.14 Element_VIA23_1_3_36_36 ;
      VIA 20.436 21.6 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 21.583 20.481 21.617 ;
      VIA 20.436 21.6 Element_VIA34_1_2_58_52 ;
      VIA 20.436 21.6 Element_VIA23_1_3_36_36 ;
      VIA 20.436 21.06 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 21.043 20.481 21.077 ;
      VIA 20.436 21.06 Element_VIA34_1_2_58_52 ;
      VIA 20.436 21.06 Element_VIA23_1_3_36_36 ;
      VIA 20.436 20.52 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 20.503 20.481 20.537 ;
      VIA 20.436 20.52 Element_VIA34_1_2_58_52 ;
      VIA 20.436 20.52 Element_VIA23_1_3_36_36 ;
      VIA 20.436 19.98 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 19.963 20.481 19.997 ;
      VIA 20.436 19.98 Element_VIA34_1_2_58_52 ;
      VIA 20.436 19.98 Element_VIA23_1_3_36_36 ;
      VIA 20.436 19.44 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 19.423 20.481 19.457 ;
      VIA 20.436 19.44 Element_VIA34_1_2_58_52 ;
      VIA 20.436 19.44 Element_VIA23_1_3_36_36 ;
      VIA 20.436 18.9 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 18.883 20.481 18.917 ;
      VIA 20.436 18.9 Element_VIA34_1_2_58_52 ;
      VIA 20.436 18.9 Element_VIA23_1_3_36_36 ;
      VIA 20.436 18.36 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 18.343 20.481 18.377 ;
      VIA 20.436 18.36 Element_VIA34_1_2_58_52 ;
      VIA 20.436 18.36 Element_VIA23_1_3_36_36 ;
      VIA 20.436 17.82 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 17.803 20.481 17.837 ;
      VIA 20.436 17.82 Element_VIA34_1_2_58_52 ;
      VIA 20.436 17.82 Element_VIA23_1_3_36_36 ;
      VIA 20.436 17.28 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 17.263 20.481 17.297 ;
      VIA 20.436 17.28 Element_VIA34_1_2_58_52 ;
      VIA 20.436 17.28 Element_VIA23_1_3_36_36 ;
      VIA 20.436 16.74 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 16.723 20.481 16.757 ;
      VIA 20.436 16.74 Element_VIA34_1_2_58_52 ;
      VIA 20.436 16.74 Element_VIA23_1_3_36_36 ;
      VIA 20.436 16.2 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 16.183 20.481 16.217 ;
      VIA 20.436 16.2 Element_VIA34_1_2_58_52 ;
      VIA 20.436 16.2 Element_VIA23_1_3_36_36 ;
      VIA 20.436 15.66 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 15.643 20.481 15.677 ;
      VIA 20.436 15.66 Element_VIA34_1_2_58_52 ;
      VIA 20.436 15.66 Element_VIA23_1_3_36_36 ;
      VIA 20.436 15.12 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 15.103 20.481 15.137 ;
      VIA 20.436 15.12 Element_VIA34_1_2_58_52 ;
      VIA 20.436 15.12 Element_VIA23_1_3_36_36 ;
      VIA 20.436 14.58 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 14.563 20.481 14.597 ;
      VIA 20.436 14.58 Element_VIA34_1_2_58_52 ;
      VIA 20.436 14.58 Element_VIA23_1_3_36_36 ;
      VIA 20.436 14.04 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 14.023 20.481 14.057 ;
      VIA 20.436 14.04 Element_VIA34_1_2_58_52 ;
      VIA 20.436 14.04 Element_VIA23_1_3_36_36 ;
      VIA 20.436 13.5 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 13.483 20.481 13.517 ;
      VIA 20.436 13.5 Element_VIA34_1_2_58_52 ;
      VIA 20.436 13.5 Element_VIA23_1_3_36_36 ;
      VIA 20.436 12.96 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 12.943 20.481 12.977 ;
      VIA 20.436 12.96 Element_VIA34_1_2_58_52 ;
      VIA 20.436 12.96 Element_VIA23_1_3_36_36 ;
      VIA 20.436 12.42 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 12.403 20.481 12.437 ;
      VIA 20.436 12.42 Element_VIA34_1_2_58_52 ;
      VIA 20.436 12.42 Element_VIA23_1_3_36_36 ;
      VIA 20.436 11.88 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 11.863 20.481 11.897 ;
      VIA 20.436 11.88 Element_VIA34_1_2_58_52 ;
      VIA 20.436 11.88 Element_VIA23_1_3_36_36 ;
      VIA 20.436 11.34 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 11.323 20.481 11.357 ;
      VIA 20.436 11.34 Element_VIA34_1_2_58_52 ;
      VIA 20.436 11.34 Element_VIA23_1_3_36_36 ;
      VIA 20.436 10.8 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 10.783 20.481 10.817 ;
      VIA 20.436 10.8 Element_VIA34_1_2_58_52 ;
      VIA 20.436 10.8 Element_VIA23_1_3_36_36 ;
      VIA 20.436 10.26 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 10.243 20.481 10.277 ;
      VIA 20.436 10.26 Element_VIA34_1_2_58_52 ;
      VIA 20.436 10.26 Element_VIA23_1_3_36_36 ;
      VIA 20.436 9.72 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 9.703 20.481 9.737 ;
      VIA 20.436 9.72 Element_VIA34_1_2_58_52 ;
      VIA 20.436 9.72 Element_VIA23_1_3_36_36 ;
      VIA 20.436 9.18 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 9.163 20.481 9.197 ;
      VIA 20.436 9.18 Element_VIA34_1_2_58_52 ;
      VIA 20.436 9.18 Element_VIA23_1_3_36_36 ;
      VIA 20.436 8.64 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 8.623 20.481 8.657 ;
      VIA 20.436 8.64 Element_VIA34_1_2_58_52 ;
      VIA 20.436 8.64 Element_VIA23_1_3_36_36 ;
      VIA 20.436 8.1 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 8.083 20.481 8.117 ;
      VIA 20.436 8.1 Element_VIA34_1_2_58_52 ;
      VIA 20.436 8.1 Element_VIA23_1_3_36_36 ;
      VIA 20.436 7.56 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 7.543 20.481 7.577 ;
      VIA 20.436 7.56 Element_VIA34_1_2_58_52 ;
      VIA 20.436 7.56 Element_VIA23_1_3_36_36 ;
      VIA 20.436 7.02 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 7.003 20.481 7.037 ;
      VIA 20.436 7.02 Element_VIA34_1_2_58_52 ;
      VIA 20.436 7.02 Element_VIA23_1_3_36_36 ;
      VIA 20.436 6.48 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 6.463 20.481 6.497 ;
      VIA 20.436 6.48 Element_VIA34_1_2_58_52 ;
      VIA 20.436 6.48 Element_VIA23_1_3_36_36 ;
      VIA 20.436 5.94 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 5.923 20.481 5.957 ;
      VIA 20.436 5.94 Element_VIA34_1_2_58_52 ;
      VIA 20.436 5.94 Element_VIA23_1_3_36_36 ;
      VIA 20.436 5.4 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 5.383 20.481 5.417 ;
      VIA 20.436 5.4 Element_VIA34_1_2_58_52 ;
      VIA 20.436 5.4 Element_VIA23_1_3_36_36 ;
      VIA 20.436 4.86 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 4.843 20.481 4.877 ;
      VIA 20.436 4.86 Element_VIA34_1_2_58_52 ;
      VIA 20.436 4.86 Element_VIA23_1_3_36_36 ;
      VIA 20.436 4.32 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 4.303 20.481 4.337 ;
      VIA 20.436 4.32 Element_VIA34_1_2_58_52 ;
      VIA 20.436 4.32 Element_VIA23_1_3_36_36 ;
      VIA 20.436 3.78 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 3.763 20.481 3.797 ;
      VIA 20.436 3.78 Element_VIA34_1_2_58_52 ;
      VIA 20.436 3.78 Element_VIA23_1_3_36_36 ;
      VIA 20.436 3.24 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 3.223 20.481 3.257 ;
      VIA 20.436 3.24 Element_VIA34_1_2_58_52 ;
      VIA 20.436 3.24 Element_VIA23_1_3_36_36 ;
      VIA 20.436 2.7 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 2.683 20.481 2.717 ;
      VIA 20.436 2.7 Element_VIA34_1_2_58_52 ;
      VIA 20.436 2.7 Element_VIA23_1_3_36_36 ;
      VIA 20.436 2.16 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 2.143 20.481 2.177 ;
      VIA 20.436 2.16 Element_VIA34_1_2_58_52 ;
      VIA 20.436 2.16 Element_VIA23_1_3_36_36 ;
      VIA 20.436 1.62 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 1.603 20.481 1.637 ;
      VIA 20.436 1.62 Element_VIA34_1_2_58_52 ;
      VIA 20.436 1.62 Element_VIA23_1_3_36_36 ;
      VIA 20.436 1.08 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  20.391 1.063 20.481 1.097 ;
      VIA 20.436 1.08 Element_VIA34_1_2_58_52 ;
      VIA 20.436 1.08 Element_VIA23_1_3_36_36 ;
      VIA 17.46 42.12 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 42.103 17.505 42.137 ;
      VIA 17.46 42.12 Element_VIA34_1_2_58_52 ;
      VIA 17.46 42.12 Element_VIA23_1_3_36_36 ;
      VIA 17.46 41.58 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 41.563 17.505 41.597 ;
      VIA 17.46 41.58 Element_VIA34_1_2_58_52 ;
      VIA 17.46 41.58 Element_VIA23_1_3_36_36 ;
      VIA 17.46 41.04 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 41.023 17.505 41.057 ;
      VIA 17.46 41.04 Element_VIA34_1_2_58_52 ;
      VIA 17.46 41.04 Element_VIA23_1_3_36_36 ;
      VIA 17.46 40.5 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 40.483 17.505 40.517 ;
      VIA 17.46 40.5 Element_VIA34_1_2_58_52 ;
      VIA 17.46 40.5 Element_VIA23_1_3_36_36 ;
      VIA 17.46 39.96 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 39.943 17.505 39.977 ;
      VIA 17.46 39.96 Element_VIA34_1_2_58_52 ;
      VIA 17.46 39.96 Element_VIA23_1_3_36_36 ;
      VIA 17.46 39.42 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 39.403 17.505 39.437 ;
      VIA 17.46 39.42 Element_VIA34_1_2_58_52 ;
      VIA 17.46 39.42 Element_VIA23_1_3_36_36 ;
      VIA 17.46 38.88 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 38.863 17.505 38.897 ;
      VIA 17.46 38.88 Element_VIA34_1_2_58_52 ;
      VIA 17.46 38.88 Element_VIA23_1_3_36_36 ;
      VIA 17.46 38.34 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 38.323 17.505 38.357 ;
      VIA 17.46 38.34 Element_VIA34_1_2_58_52 ;
      VIA 17.46 38.34 Element_VIA23_1_3_36_36 ;
      VIA 17.46 37.8 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 37.783 17.505 37.817 ;
      VIA 17.46 37.8 Element_VIA34_1_2_58_52 ;
      VIA 17.46 37.8 Element_VIA23_1_3_36_36 ;
      VIA 17.46 37.26 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 37.243 17.505 37.277 ;
      VIA 17.46 37.26 Element_VIA34_1_2_58_52 ;
      VIA 17.46 37.26 Element_VIA23_1_3_36_36 ;
      VIA 17.46 36.72 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 36.703 17.505 36.737 ;
      VIA 17.46 36.72 Element_VIA34_1_2_58_52 ;
      VIA 17.46 36.72 Element_VIA23_1_3_36_36 ;
      VIA 17.46 36.18 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 36.163 17.505 36.197 ;
      VIA 17.46 36.18 Element_VIA34_1_2_58_52 ;
      VIA 17.46 36.18 Element_VIA23_1_3_36_36 ;
      VIA 17.46 35.64 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 35.623 17.505 35.657 ;
      VIA 17.46 35.64 Element_VIA34_1_2_58_52 ;
      VIA 17.46 35.64 Element_VIA23_1_3_36_36 ;
      VIA 17.46 35.1 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 35.083 17.505 35.117 ;
      VIA 17.46 35.1 Element_VIA34_1_2_58_52 ;
      VIA 17.46 35.1 Element_VIA23_1_3_36_36 ;
      VIA 17.46 34.56 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 34.543 17.505 34.577 ;
      VIA 17.46 34.56 Element_VIA34_1_2_58_52 ;
      VIA 17.46 34.56 Element_VIA23_1_3_36_36 ;
      VIA 17.46 34.02 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 34.003 17.505 34.037 ;
      VIA 17.46 34.02 Element_VIA34_1_2_58_52 ;
      VIA 17.46 34.02 Element_VIA23_1_3_36_36 ;
      VIA 17.46 33.48 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 33.463 17.505 33.497 ;
      VIA 17.46 33.48 Element_VIA34_1_2_58_52 ;
      VIA 17.46 33.48 Element_VIA23_1_3_36_36 ;
      VIA 17.46 32.94 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 32.923 17.505 32.957 ;
      VIA 17.46 32.94 Element_VIA34_1_2_58_52 ;
      VIA 17.46 32.94 Element_VIA23_1_3_36_36 ;
      VIA 17.46 32.4 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 32.383 17.505 32.417 ;
      VIA 17.46 32.4 Element_VIA34_1_2_58_52 ;
      VIA 17.46 32.4 Element_VIA23_1_3_36_36 ;
      VIA 17.46 31.86 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 31.843 17.505 31.877 ;
      VIA 17.46 31.86 Element_VIA34_1_2_58_52 ;
      VIA 17.46 31.86 Element_VIA23_1_3_36_36 ;
      VIA 17.46 31.32 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 31.303 17.505 31.337 ;
      VIA 17.46 31.32 Element_VIA34_1_2_58_52 ;
      VIA 17.46 31.32 Element_VIA23_1_3_36_36 ;
      VIA 17.46 30.78 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 30.763 17.505 30.797 ;
      VIA 17.46 30.78 Element_VIA34_1_2_58_52 ;
      VIA 17.46 30.78 Element_VIA23_1_3_36_36 ;
      VIA 17.46 30.24 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 30.223 17.505 30.257 ;
      VIA 17.46 30.24 Element_VIA34_1_2_58_52 ;
      VIA 17.46 30.24 Element_VIA23_1_3_36_36 ;
      VIA 17.46 29.7 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 29.683 17.505 29.717 ;
      VIA 17.46 29.7 Element_VIA34_1_2_58_52 ;
      VIA 17.46 29.7 Element_VIA23_1_3_36_36 ;
      VIA 17.46 29.16 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 29.143 17.505 29.177 ;
      VIA 17.46 29.16 Element_VIA34_1_2_58_52 ;
      VIA 17.46 29.16 Element_VIA23_1_3_36_36 ;
      VIA 17.46 28.62 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 28.603 17.505 28.637 ;
      VIA 17.46 28.62 Element_VIA34_1_2_58_52 ;
      VIA 17.46 28.62 Element_VIA23_1_3_36_36 ;
      VIA 17.46 28.08 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 28.063 17.505 28.097 ;
      VIA 17.46 28.08 Element_VIA34_1_2_58_52 ;
      VIA 17.46 28.08 Element_VIA23_1_3_36_36 ;
      VIA 17.46 27.54 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 27.523 17.505 27.557 ;
      VIA 17.46 27.54 Element_VIA34_1_2_58_52 ;
      VIA 17.46 27.54 Element_VIA23_1_3_36_36 ;
      VIA 17.46 27 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 26.983 17.505 27.017 ;
      VIA 17.46 27 Element_VIA34_1_2_58_52 ;
      VIA 17.46 27 Element_VIA23_1_3_36_36 ;
      VIA 17.46 26.46 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 26.443 17.505 26.477 ;
      VIA 17.46 26.46 Element_VIA34_1_2_58_52 ;
      VIA 17.46 26.46 Element_VIA23_1_3_36_36 ;
      VIA 17.46 25.92 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 25.903 17.505 25.937 ;
      VIA 17.46 25.92 Element_VIA34_1_2_58_52 ;
      VIA 17.46 25.92 Element_VIA23_1_3_36_36 ;
      VIA 17.46 25.38 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 25.363 17.505 25.397 ;
      VIA 17.46 25.38 Element_VIA34_1_2_58_52 ;
      VIA 17.46 25.38 Element_VIA23_1_3_36_36 ;
      VIA 17.46 24.84 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 24.823 17.505 24.857 ;
      VIA 17.46 24.84 Element_VIA34_1_2_58_52 ;
      VIA 17.46 24.84 Element_VIA23_1_3_36_36 ;
      VIA 17.46 24.3 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 24.283 17.505 24.317 ;
      VIA 17.46 24.3 Element_VIA34_1_2_58_52 ;
      VIA 17.46 24.3 Element_VIA23_1_3_36_36 ;
      VIA 17.46 23.76 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 23.743 17.505 23.777 ;
      VIA 17.46 23.76 Element_VIA34_1_2_58_52 ;
      VIA 17.46 23.76 Element_VIA23_1_3_36_36 ;
      VIA 17.46 23.22 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 23.203 17.505 23.237 ;
      VIA 17.46 23.22 Element_VIA34_1_2_58_52 ;
      VIA 17.46 23.22 Element_VIA23_1_3_36_36 ;
      VIA 17.46 22.68 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 22.663 17.505 22.697 ;
      VIA 17.46 22.68 Element_VIA34_1_2_58_52 ;
      VIA 17.46 22.68 Element_VIA23_1_3_36_36 ;
      VIA 17.46 22.14 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 22.123 17.505 22.157 ;
      VIA 17.46 22.14 Element_VIA34_1_2_58_52 ;
      VIA 17.46 22.14 Element_VIA23_1_3_36_36 ;
      VIA 17.46 21.6 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 21.583 17.505 21.617 ;
      VIA 17.46 21.6 Element_VIA34_1_2_58_52 ;
      VIA 17.46 21.6 Element_VIA23_1_3_36_36 ;
      VIA 17.46 21.06 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 21.043 17.505 21.077 ;
      VIA 17.46 21.06 Element_VIA34_1_2_58_52 ;
      VIA 17.46 21.06 Element_VIA23_1_3_36_36 ;
      VIA 17.46 20.52 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 20.503 17.505 20.537 ;
      VIA 17.46 20.52 Element_VIA34_1_2_58_52 ;
      VIA 17.46 20.52 Element_VIA23_1_3_36_36 ;
      VIA 17.46 19.98 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 19.963 17.505 19.997 ;
      VIA 17.46 19.98 Element_VIA34_1_2_58_52 ;
      VIA 17.46 19.98 Element_VIA23_1_3_36_36 ;
      VIA 17.46 19.44 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 19.423 17.505 19.457 ;
      VIA 17.46 19.44 Element_VIA34_1_2_58_52 ;
      VIA 17.46 19.44 Element_VIA23_1_3_36_36 ;
      VIA 17.46 18.9 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 18.883 17.505 18.917 ;
      VIA 17.46 18.9 Element_VIA34_1_2_58_52 ;
      VIA 17.46 18.9 Element_VIA23_1_3_36_36 ;
      VIA 17.46 18.36 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 18.343 17.505 18.377 ;
      VIA 17.46 18.36 Element_VIA34_1_2_58_52 ;
      VIA 17.46 18.36 Element_VIA23_1_3_36_36 ;
      VIA 17.46 17.82 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 17.803 17.505 17.837 ;
      VIA 17.46 17.82 Element_VIA34_1_2_58_52 ;
      VIA 17.46 17.82 Element_VIA23_1_3_36_36 ;
      VIA 17.46 17.28 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 17.263 17.505 17.297 ;
      VIA 17.46 17.28 Element_VIA34_1_2_58_52 ;
      VIA 17.46 17.28 Element_VIA23_1_3_36_36 ;
      VIA 17.46 16.74 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 16.723 17.505 16.757 ;
      VIA 17.46 16.74 Element_VIA34_1_2_58_52 ;
      VIA 17.46 16.74 Element_VIA23_1_3_36_36 ;
      VIA 17.46 16.2 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 16.183 17.505 16.217 ;
      VIA 17.46 16.2 Element_VIA34_1_2_58_52 ;
      VIA 17.46 16.2 Element_VIA23_1_3_36_36 ;
      VIA 17.46 15.66 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 15.643 17.505 15.677 ;
      VIA 17.46 15.66 Element_VIA34_1_2_58_52 ;
      VIA 17.46 15.66 Element_VIA23_1_3_36_36 ;
      VIA 17.46 15.12 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 15.103 17.505 15.137 ;
      VIA 17.46 15.12 Element_VIA34_1_2_58_52 ;
      VIA 17.46 15.12 Element_VIA23_1_3_36_36 ;
      VIA 17.46 14.58 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 14.563 17.505 14.597 ;
      VIA 17.46 14.58 Element_VIA34_1_2_58_52 ;
      VIA 17.46 14.58 Element_VIA23_1_3_36_36 ;
      VIA 17.46 14.04 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 14.023 17.505 14.057 ;
      VIA 17.46 14.04 Element_VIA34_1_2_58_52 ;
      VIA 17.46 14.04 Element_VIA23_1_3_36_36 ;
      VIA 17.46 13.5 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 13.483 17.505 13.517 ;
      VIA 17.46 13.5 Element_VIA34_1_2_58_52 ;
      VIA 17.46 13.5 Element_VIA23_1_3_36_36 ;
      VIA 17.46 12.96 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 12.943 17.505 12.977 ;
      VIA 17.46 12.96 Element_VIA34_1_2_58_52 ;
      VIA 17.46 12.96 Element_VIA23_1_3_36_36 ;
      VIA 17.46 12.42 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 12.403 17.505 12.437 ;
      VIA 17.46 12.42 Element_VIA34_1_2_58_52 ;
      VIA 17.46 12.42 Element_VIA23_1_3_36_36 ;
      VIA 17.46 11.88 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 11.863 17.505 11.897 ;
      VIA 17.46 11.88 Element_VIA34_1_2_58_52 ;
      VIA 17.46 11.88 Element_VIA23_1_3_36_36 ;
      VIA 17.46 11.34 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 11.323 17.505 11.357 ;
      VIA 17.46 11.34 Element_VIA34_1_2_58_52 ;
      VIA 17.46 11.34 Element_VIA23_1_3_36_36 ;
      VIA 17.46 10.8 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 10.783 17.505 10.817 ;
      VIA 17.46 10.8 Element_VIA34_1_2_58_52 ;
      VIA 17.46 10.8 Element_VIA23_1_3_36_36 ;
      VIA 17.46 10.26 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 10.243 17.505 10.277 ;
      VIA 17.46 10.26 Element_VIA34_1_2_58_52 ;
      VIA 17.46 10.26 Element_VIA23_1_3_36_36 ;
      VIA 17.46 9.72 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 9.703 17.505 9.737 ;
      VIA 17.46 9.72 Element_VIA34_1_2_58_52 ;
      VIA 17.46 9.72 Element_VIA23_1_3_36_36 ;
      VIA 17.46 9.18 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 9.163 17.505 9.197 ;
      VIA 17.46 9.18 Element_VIA34_1_2_58_52 ;
      VIA 17.46 9.18 Element_VIA23_1_3_36_36 ;
      VIA 17.46 8.64 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 8.623 17.505 8.657 ;
      VIA 17.46 8.64 Element_VIA34_1_2_58_52 ;
      VIA 17.46 8.64 Element_VIA23_1_3_36_36 ;
      VIA 17.46 8.1 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 8.083 17.505 8.117 ;
      VIA 17.46 8.1 Element_VIA34_1_2_58_52 ;
      VIA 17.46 8.1 Element_VIA23_1_3_36_36 ;
      VIA 17.46 7.56 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 7.543 17.505 7.577 ;
      VIA 17.46 7.56 Element_VIA34_1_2_58_52 ;
      VIA 17.46 7.56 Element_VIA23_1_3_36_36 ;
      VIA 17.46 7.02 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 7.003 17.505 7.037 ;
      VIA 17.46 7.02 Element_VIA34_1_2_58_52 ;
      VIA 17.46 7.02 Element_VIA23_1_3_36_36 ;
      VIA 17.46 6.48 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 6.463 17.505 6.497 ;
      VIA 17.46 6.48 Element_VIA34_1_2_58_52 ;
      VIA 17.46 6.48 Element_VIA23_1_3_36_36 ;
      VIA 17.46 5.94 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 5.923 17.505 5.957 ;
      VIA 17.46 5.94 Element_VIA34_1_2_58_52 ;
      VIA 17.46 5.94 Element_VIA23_1_3_36_36 ;
      VIA 17.46 5.4 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 5.383 17.505 5.417 ;
      VIA 17.46 5.4 Element_VIA34_1_2_58_52 ;
      VIA 17.46 5.4 Element_VIA23_1_3_36_36 ;
      VIA 17.46 4.86 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 4.843 17.505 4.877 ;
      VIA 17.46 4.86 Element_VIA34_1_2_58_52 ;
      VIA 17.46 4.86 Element_VIA23_1_3_36_36 ;
      VIA 17.46 4.32 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 4.303 17.505 4.337 ;
      VIA 17.46 4.32 Element_VIA34_1_2_58_52 ;
      VIA 17.46 4.32 Element_VIA23_1_3_36_36 ;
      VIA 17.46 3.78 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 3.763 17.505 3.797 ;
      VIA 17.46 3.78 Element_VIA34_1_2_58_52 ;
      VIA 17.46 3.78 Element_VIA23_1_3_36_36 ;
      VIA 17.46 3.24 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 3.223 17.505 3.257 ;
      VIA 17.46 3.24 Element_VIA34_1_2_58_52 ;
      VIA 17.46 3.24 Element_VIA23_1_3_36_36 ;
      VIA 17.46 2.7 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 2.683 17.505 2.717 ;
      VIA 17.46 2.7 Element_VIA34_1_2_58_52 ;
      VIA 17.46 2.7 Element_VIA23_1_3_36_36 ;
      VIA 17.46 2.16 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 2.143 17.505 2.177 ;
      VIA 17.46 2.16 Element_VIA34_1_2_58_52 ;
      VIA 17.46 2.16 Element_VIA23_1_3_36_36 ;
      VIA 17.46 1.62 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 1.603 17.505 1.637 ;
      VIA 17.46 1.62 Element_VIA34_1_2_58_52 ;
      VIA 17.46 1.62 Element_VIA23_1_3_36_36 ;
      VIA 17.46 1.08 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  17.415 1.063 17.505 1.097 ;
      VIA 17.46 1.08 Element_VIA34_1_2_58_52 ;
      VIA 17.46 1.08 Element_VIA23_1_3_36_36 ;
      VIA 14.484 42.12 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 42.103 14.529 42.137 ;
      VIA 14.484 42.12 Element_VIA34_1_2_58_52 ;
      VIA 14.484 42.12 Element_VIA23_1_3_36_36 ;
      VIA 14.484 41.58 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 41.563 14.529 41.597 ;
      VIA 14.484 41.58 Element_VIA34_1_2_58_52 ;
      VIA 14.484 41.58 Element_VIA23_1_3_36_36 ;
      VIA 14.484 41.04 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 41.023 14.529 41.057 ;
      VIA 14.484 41.04 Element_VIA34_1_2_58_52 ;
      VIA 14.484 41.04 Element_VIA23_1_3_36_36 ;
      VIA 14.484 40.5 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 40.483 14.529 40.517 ;
      VIA 14.484 40.5 Element_VIA34_1_2_58_52 ;
      VIA 14.484 40.5 Element_VIA23_1_3_36_36 ;
      VIA 14.484 39.96 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 39.943 14.529 39.977 ;
      VIA 14.484 39.96 Element_VIA34_1_2_58_52 ;
      VIA 14.484 39.96 Element_VIA23_1_3_36_36 ;
      VIA 14.484 39.42 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 39.403 14.529 39.437 ;
      VIA 14.484 39.42 Element_VIA34_1_2_58_52 ;
      VIA 14.484 39.42 Element_VIA23_1_3_36_36 ;
      VIA 14.484 38.88 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 38.863 14.529 38.897 ;
      VIA 14.484 38.88 Element_VIA34_1_2_58_52 ;
      VIA 14.484 38.88 Element_VIA23_1_3_36_36 ;
      VIA 14.484 38.34 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 38.323 14.529 38.357 ;
      VIA 14.484 38.34 Element_VIA34_1_2_58_52 ;
      VIA 14.484 38.34 Element_VIA23_1_3_36_36 ;
      VIA 14.484 37.8 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 37.783 14.529 37.817 ;
      VIA 14.484 37.8 Element_VIA34_1_2_58_52 ;
      VIA 14.484 37.8 Element_VIA23_1_3_36_36 ;
      VIA 14.484 37.26 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 37.243 14.529 37.277 ;
      VIA 14.484 37.26 Element_VIA34_1_2_58_52 ;
      VIA 14.484 37.26 Element_VIA23_1_3_36_36 ;
      VIA 14.484 36.72 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 36.703 14.529 36.737 ;
      VIA 14.484 36.72 Element_VIA34_1_2_58_52 ;
      VIA 14.484 36.72 Element_VIA23_1_3_36_36 ;
      VIA 14.484 36.18 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 36.163 14.529 36.197 ;
      VIA 14.484 36.18 Element_VIA34_1_2_58_52 ;
      VIA 14.484 36.18 Element_VIA23_1_3_36_36 ;
      VIA 14.484 35.64 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 35.623 14.529 35.657 ;
      VIA 14.484 35.64 Element_VIA34_1_2_58_52 ;
      VIA 14.484 35.64 Element_VIA23_1_3_36_36 ;
      VIA 14.484 35.1 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 35.083 14.529 35.117 ;
      VIA 14.484 35.1 Element_VIA34_1_2_58_52 ;
      VIA 14.484 35.1 Element_VIA23_1_3_36_36 ;
      VIA 14.484 34.56 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 34.543 14.529 34.577 ;
      VIA 14.484 34.56 Element_VIA34_1_2_58_52 ;
      VIA 14.484 34.56 Element_VIA23_1_3_36_36 ;
      VIA 14.484 34.02 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 34.003 14.529 34.037 ;
      VIA 14.484 34.02 Element_VIA34_1_2_58_52 ;
      VIA 14.484 34.02 Element_VIA23_1_3_36_36 ;
      VIA 14.484 33.48 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 33.463 14.529 33.497 ;
      VIA 14.484 33.48 Element_VIA34_1_2_58_52 ;
      VIA 14.484 33.48 Element_VIA23_1_3_36_36 ;
      VIA 14.484 32.94 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 32.923 14.529 32.957 ;
      VIA 14.484 32.94 Element_VIA34_1_2_58_52 ;
      VIA 14.484 32.94 Element_VIA23_1_3_36_36 ;
      VIA 14.484 32.4 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 32.383 14.529 32.417 ;
      VIA 14.484 32.4 Element_VIA34_1_2_58_52 ;
      VIA 14.484 32.4 Element_VIA23_1_3_36_36 ;
      VIA 14.484 31.86 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 31.843 14.529 31.877 ;
      VIA 14.484 31.86 Element_VIA34_1_2_58_52 ;
      VIA 14.484 31.86 Element_VIA23_1_3_36_36 ;
      VIA 14.484 31.32 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 31.303 14.529 31.337 ;
      VIA 14.484 31.32 Element_VIA34_1_2_58_52 ;
      VIA 14.484 31.32 Element_VIA23_1_3_36_36 ;
      VIA 14.484 30.78 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 30.763 14.529 30.797 ;
      VIA 14.484 30.78 Element_VIA34_1_2_58_52 ;
      VIA 14.484 30.78 Element_VIA23_1_3_36_36 ;
      VIA 14.484 30.24 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 30.223 14.529 30.257 ;
      VIA 14.484 30.24 Element_VIA34_1_2_58_52 ;
      VIA 14.484 30.24 Element_VIA23_1_3_36_36 ;
      VIA 14.484 29.7 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 29.683 14.529 29.717 ;
      VIA 14.484 29.7 Element_VIA34_1_2_58_52 ;
      VIA 14.484 29.7 Element_VIA23_1_3_36_36 ;
      VIA 14.484 29.16 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 29.143 14.529 29.177 ;
      VIA 14.484 29.16 Element_VIA34_1_2_58_52 ;
      VIA 14.484 29.16 Element_VIA23_1_3_36_36 ;
      VIA 14.484 28.62 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 28.603 14.529 28.637 ;
      VIA 14.484 28.62 Element_VIA34_1_2_58_52 ;
      VIA 14.484 28.62 Element_VIA23_1_3_36_36 ;
      VIA 14.484 28.08 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 28.063 14.529 28.097 ;
      VIA 14.484 28.08 Element_VIA34_1_2_58_52 ;
      VIA 14.484 28.08 Element_VIA23_1_3_36_36 ;
      VIA 14.484 27.54 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 27.523 14.529 27.557 ;
      VIA 14.484 27.54 Element_VIA34_1_2_58_52 ;
      VIA 14.484 27.54 Element_VIA23_1_3_36_36 ;
      VIA 14.484 27 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 26.983 14.529 27.017 ;
      VIA 14.484 27 Element_VIA34_1_2_58_52 ;
      VIA 14.484 27 Element_VIA23_1_3_36_36 ;
      VIA 14.484 26.46 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 26.443 14.529 26.477 ;
      VIA 14.484 26.46 Element_VIA34_1_2_58_52 ;
      VIA 14.484 26.46 Element_VIA23_1_3_36_36 ;
      VIA 14.484 25.92 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 25.903 14.529 25.937 ;
      VIA 14.484 25.92 Element_VIA34_1_2_58_52 ;
      VIA 14.484 25.92 Element_VIA23_1_3_36_36 ;
      VIA 14.484 25.38 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 25.363 14.529 25.397 ;
      VIA 14.484 25.38 Element_VIA34_1_2_58_52 ;
      VIA 14.484 25.38 Element_VIA23_1_3_36_36 ;
      VIA 14.484 24.84 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 24.823 14.529 24.857 ;
      VIA 14.484 24.84 Element_VIA34_1_2_58_52 ;
      VIA 14.484 24.84 Element_VIA23_1_3_36_36 ;
      VIA 14.484 24.3 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 24.283 14.529 24.317 ;
      VIA 14.484 24.3 Element_VIA34_1_2_58_52 ;
      VIA 14.484 24.3 Element_VIA23_1_3_36_36 ;
      VIA 14.484 23.76 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 23.743 14.529 23.777 ;
      VIA 14.484 23.76 Element_VIA34_1_2_58_52 ;
      VIA 14.484 23.76 Element_VIA23_1_3_36_36 ;
      VIA 14.484 23.22 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 23.203 14.529 23.237 ;
      VIA 14.484 23.22 Element_VIA34_1_2_58_52 ;
      VIA 14.484 23.22 Element_VIA23_1_3_36_36 ;
      VIA 14.484 22.68 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 22.663 14.529 22.697 ;
      VIA 14.484 22.68 Element_VIA34_1_2_58_52 ;
      VIA 14.484 22.68 Element_VIA23_1_3_36_36 ;
      VIA 14.484 22.14 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 22.123 14.529 22.157 ;
      VIA 14.484 22.14 Element_VIA34_1_2_58_52 ;
      VIA 14.484 22.14 Element_VIA23_1_3_36_36 ;
      VIA 14.484 21.6 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 21.583 14.529 21.617 ;
      VIA 14.484 21.6 Element_VIA34_1_2_58_52 ;
      VIA 14.484 21.6 Element_VIA23_1_3_36_36 ;
      VIA 14.484 21.06 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 21.043 14.529 21.077 ;
      VIA 14.484 21.06 Element_VIA34_1_2_58_52 ;
      VIA 14.484 21.06 Element_VIA23_1_3_36_36 ;
      VIA 14.484 20.52 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 20.503 14.529 20.537 ;
      VIA 14.484 20.52 Element_VIA34_1_2_58_52 ;
      VIA 14.484 20.52 Element_VIA23_1_3_36_36 ;
      VIA 14.484 19.98 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 19.963 14.529 19.997 ;
      VIA 14.484 19.98 Element_VIA34_1_2_58_52 ;
      VIA 14.484 19.98 Element_VIA23_1_3_36_36 ;
      VIA 14.484 19.44 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 19.423 14.529 19.457 ;
      VIA 14.484 19.44 Element_VIA34_1_2_58_52 ;
      VIA 14.484 19.44 Element_VIA23_1_3_36_36 ;
      VIA 14.484 18.9 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 18.883 14.529 18.917 ;
      VIA 14.484 18.9 Element_VIA34_1_2_58_52 ;
      VIA 14.484 18.9 Element_VIA23_1_3_36_36 ;
      VIA 14.484 18.36 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 18.343 14.529 18.377 ;
      VIA 14.484 18.36 Element_VIA34_1_2_58_52 ;
      VIA 14.484 18.36 Element_VIA23_1_3_36_36 ;
      VIA 14.484 17.82 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 17.803 14.529 17.837 ;
      VIA 14.484 17.82 Element_VIA34_1_2_58_52 ;
      VIA 14.484 17.82 Element_VIA23_1_3_36_36 ;
      VIA 14.484 17.28 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 17.263 14.529 17.297 ;
      VIA 14.484 17.28 Element_VIA34_1_2_58_52 ;
      VIA 14.484 17.28 Element_VIA23_1_3_36_36 ;
      VIA 14.484 16.74 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 16.723 14.529 16.757 ;
      VIA 14.484 16.74 Element_VIA34_1_2_58_52 ;
      VIA 14.484 16.74 Element_VIA23_1_3_36_36 ;
      VIA 14.484 16.2 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 16.183 14.529 16.217 ;
      VIA 14.484 16.2 Element_VIA34_1_2_58_52 ;
      VIA 14.484 16.2 Element_VIA23_1_3_36_36 ;
      VIA 14.484 15.66 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 15.643 14.529 15.677 ;
      VIA 14.484 15.66 Element_VIA34_1_2_58_52 ;
      VIA 14.484 15.66 Element_VIA23_1_3_36_36 ;
      VIA 14.484 15.12 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 15.103 14.529 15.137 ;
      VIA 14.484 15.12 Element_VIA34_1_2_58_52 ;
      VIA 14.484 15.12 Element_VIA23_1_3_36_36 ;
      VIA 14.484 14.58 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 14.563 14.529 14.597 ;
      VIA 14.484 14.58 Element_VIA34_1_2_58_52 ;
      VIA 14.484 14.58 Element_VIA23_1_3_36_36 ;
      VIA 14.484 14.04 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 14.023 14.529 14.057 ;
      VIA 14.484 14.04 Element_VIA34_1_2_58_52 ;
      VIA 14.484 14.04 Element_VIA23_1_3_36_36 ;
      VIA 14.484 13.5 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 13.483 14.529 13.517 ;
      VIA 14.484 13.5 Element_VIA34_1_2_58_52 ;
      VIA 14.484 13.5 Element_VIA23_1_3_36_36 ;
      VIA 14.484 12.96 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 12.943 14.529 12.977 ;
      VIA 14.484 12.96 Element_VIA34_1_2_58_52 ;
      VIA 14.484 12.96 Element_VIA23_1_3_36_36 ;
      VIA 14.484 12.42 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 12.403 14.529 12.437 ;
      VIA 14.484 12.42 Element_VIA34_1_2_58_52 ;
      VIA 14.484 12.42 Element_VIA23_1_3_36_36 ;
      VIA 14.484 11.88 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 11.863 14.529 11.897 ;
      VIA 14.484 11.88 Element_VIA34_1_2_58_52 ;
      VIA 14.484 11.88 Element_VIA23_1_3_36_36 ;
      VIA 14.484 11.34 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 11.323 14.529 11.357 ;
      VIA 14.484 11.34 Element_VIA34_1_2_58_52 ;
      VIA 14.484 11.34 Element_VIA23_1_3_36_36 ;
      VIA 14.484 10.8 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 10.783 14.529 10.817 ;
      VIA 14.484 10.8 Element_VIA34_1_2_58_52 ;
      VIA 14.484 10.8 Element_VIA23_1_3_36_36 ;
      VIA 14.484 10.26 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 10.243 14.529 10.277 ;
      VIA 14.484 10.26 Element_VIA34_1_2_58_52 ;
      VIA 14.484 10.26 Element_VIA23_1_3_36_36 ;
      VIA 14.484 9.72 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 9.703 14.529 9.737 ;
      VIA 14.484 9.72 Element_VIA34_1_2_58_52 ;
      VIA 14.484 9.72 Element_VIA23_1_3_36_36 ;
      VIA 14.484 9.18 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 9.163 14.529 9.197 ;
      VIA 14.484 9.18 Element_VIA34_1_2_58_52 ;
      VIA 14.484 9.18 Element_VIA23_1_3_36_36 ;
      VIA 14.484 8.64 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 8.623 14.529 8.657 ;
      VIA 14.484 8.64 Element_VIA34_1_2_58_52 ;
      VIA 14.484 8.64 Element_VIA23_1_3_36_36 ;
      VIA 14.484 8.1 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 8.083 14.529 8.117 ;
      VIA 14.484 8.1 Element_VIA34_1_2_58_52 ;
      VIA 14.484 8.1 Element_VIA23_1_3_36_36 ;
      VIA 14.484 7.56 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 7.543 14.529 7.577 ;
      VIA 14.484 7.56 Element_VIA34_1_2_58_52 ;
      VIA 14.484 7.56 Element_VIA23_1_3_36_36 ;
      VIA 14.484 7.02 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 7.003 14.529 7.037 ;
      VIA 14.484 7.02 Element_VIA34_1_2_58_52 ;
      VIA 14.484 7.02 Element_VIA23_1_3_36_36 ;
      VIA 14.484 6.48 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 6.463 14.529 6.497 ;
      VIA 14.484 6.48 Element_VIA34_1_2_58_52 ;
      VIA 14.484 6.48 Element_VIA23_1_3_36_36 ;
      VIA 14.484 5.94 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 5.923 14.529 5.957 ;
      VIA 14.484 5.94 Element_VIA34_1_2_58_52 ;
      VIA 14.484 5.94 Element_VIA23_1_3_36_36 ;
      VIA 14.484 5.4 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 5.383 14.529 5.417 ;
      VIA 14.484 5.4 Element_VIA34_1_2_58_52 ;
      VIA 14.484 5.4 Element_VIA23_1_3_36_36 ;
      VIA 14.484 4.86 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 4.843 14.529 4.877 ;
      VIA 14.484 4.86 Element_VIA34_1_2_58_52 ;
      VIA 14.484 4.86 Element_VIA23_1_3_36_36 ;
      VIA 14.484 4.32 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 4.303 14.529 4.337 ;
      VIA 14.484 4.32 Element_VIA34_1_2_58_52 ;
      VIA 14.484 4.32 Element_VIA23_1_3_36_36 ;
      VIA 14.484 3.78 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 3.763 14.529 3.797 ;
      VIA 14.484 3.78 Element_VIA34_1_2_58_52 ;
      VIA 14.484 3.78 Element_VIA23_1_3_36_36 ;
      VIA 14.484 3.24 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 3.223 14.529 3.257 ;
      VIA 14.484 3.24 Element_VIA34_1_2_58_52 ;
      VIA 14.484 3.24 Element_VIA23_1_3_36_36 ;
      VIA 14.484 2.7 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 2.683 14.529 2.717 ;
      VIA 14.484 2.7 Element_VIA34_1_2_58_52 ;
      VIA 14.484 2.7 Element_VIA23_1_3_36_36 ;
      VIA 14.484 2.16 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 2.143 14.529 2.177 ;
      VIA 14.484 2.16 Element_VIA34_1_2_58_52 ;
      VIA 14.484 2.16 Element_VIA23_1_3_36_36 ;
      VIA 14.484 1.62 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 1.603 14.529 1.637 ;
      VIA 14.484 1.62 Element_VIA34_1_2_58_52 ;
      VIA 14.484 1.62 Element_VIA23_1_3_36_36 ;
      VIA 14.484 1.08 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  14.439 1.063 14.529 1.097 ;
      VIA 14.484 1.08 Element_VIA34_1_2_58_52 ;
      VIA 14.484 1.08 Element_VIA23_1_3_36_36 ;
      VIA 11.508 42.12 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 42.103 11.553 42.137 ;
      VIA 11.508 42.12 Element_VIA34_1_2_58_52 ;
      VIA 11.508 42.12 Element_VIA23_1_3_36_36 ;
      VIA 11.508 41.58 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 41.563 11.553 41.597 ;
      VIA 11.508 41.58 Element_VIA34_1_2_58_52 ;
      VIA 11.508 41.58 Element_VIA23_1_3_36_36 ;
      VIA 11.508 41.04 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 41.023 11.553 41.057 ;
      VIA 11.508 41.04 Element_VIA34_1_2_58_52 ;
      VIA 11.508 41.04 Element_VIA23_1_3_36_36 ;
      VIA 11.508 40.5 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 40.483 11.553 40.517 ;
      VIA 11.508 40.5 Element_VIA34_1_2_58_52 ;
      VIA 11.508 40.5 Element_VIA23_1_3_36_36 ;
      VIA 11.508 39.96 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 39.943 11.553 39.977 ;
      VIA 11.508 39.96 Element_VIA34_1_2_58_52 ;
      VIA 11.508 39.96 Element_VIA23_1_3_36_36 ;
      VIA 11.508 39.42 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 39.403 11.553 39.437 ;
      VIA 11.508 39.42 Element_VIA34_1_2_58_52 ;
      VIA 11.508 39.42 Element_VIA23_1_3_36_36 ;
      VIA 11.508 38.88 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 38.863 11.553 38.897 ;
      VIA 11.508 38.88 Element_VIA34_1_2_58_52 ;
      VIA 11.508 38.88 Element_VIA23_1_3_36_36 ;
      VIA 11.508 38.34 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 38.323 11.553 38.357 ;
      VIA 11.508 38.34 Element_VIA34_1_2_58_52 ;
      VIA 11.508 38.34 Element_VIA23_1_3_36_36 ;
      VIA 11.508 37.8 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 37.783 11.553 37.817 ;
      VIA 11.508 37.8 Element_VIA34_1_2_58_52 ;
      VIA 11.508 37.8 Element_VIA23_1_3_36_36 ;
      VIA 11.508 37.26 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 37.243 11.553 37.277 ;
      VIA 11.508 37.26 Element_VIA34_1_2_58_52 ;
      VIA 11.508 37.26 Element_VIA23_1_3_36_36 ;
      VIA 11.508 36.72 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 36.703 11.553 36.737 ;
      VIA 11.508 36.72 Element_VIA34_1_2_58_52 ;
      VIA 11.508 36.72 Element_VIA23_1_3_36_36 ;
      VIA 11.508 36.18 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 36.163 11.553 36.197 ;
      VIA 11.508 36.18 Element_VIA34_1_2_58_52 ;
      VIA 11.508 36.18 Element_VIA23_1_3_36_36 ;
      VIA 11.508 35.64 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 35.623 11.553 35.657 ;
      VIA 11.508 35.64 Element_VIA34_1_2_58_52 ;
      VIA 11.508 35.64 Element_VIA23_1_3_36_36 ;
      VIA 11.508 35.1 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 35.083 11.553 35.117 ;
      VIA 11.508 35.1 Element_VIA34_1_2_58_52 ;
      VIA 11.508 35.1 Element_VIA23_1_3_36_36 ;
      VIA 11.508 34.56 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 34.543 11.553 34.577 ;
      VIA 11.508 34.56 Element_VIA34_1_2_58_52 ;
      VIA 11.508 34.56 Element_VIA23_1_3_36_36 ;
      VIA 11.508 34.02 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 34.003 11.553 34.037 ;
      VIA 11.508 34.02 Element_VIA34_1_2_58_52 ;
      VIA 11.508 34.02 Element_VIA23_1_3_36_36 ;
      VIA 11.508 33.48 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 33.463 11.553 33.497 ;
      VIA 11.508 33.48 Element_VIA34_1_2_58_52 ;
      VIA 11.508 33.48 Element_VIA23_1_3_36_36 ;
      VIA 11.508 32.94 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 32.923 11.553 32.957 ;
      VIA 11.508 32.94 Element_VIA34_1_2_58_52 ;
      VIA 11.508 32.94 Element_VIA23_1_3_36_36 ;
      VIA 11.508 32.4 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 32.383 11.553 32.417 ;
      VIA 11.508 32.4 Element_VIA34_1_2_58_52 ;
      VIA 11.508 32.4 Element_VIA23_1_3_36_36 ;
      VIA 11.508 31.86 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 31.843 11.553 31.877 ;
      VIA 11.508 31.86 Element_VIA34_1_2_58_52 ;
      VIA 11.508 31.86 Element_VIA23_1_3_36_36 ;
      VIA 11.508 31.32 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 31.303 11.553 31.337 ;
      VIA 11.508 31.32 Element_VIA34_1_2_58_52 ;
      VIA 11.508 31.32 Element_VIA23_1_3_36_36 ;
      VIA 11.508 30.78 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 30.763 11.553 30.797 ;
      VIA 11.508 30.78 Element_VIA34_1_2_58_52 ;
      VIA 11.508 30.78 Element_VIA23_1_3_36_36 ;
      VIA 11.508 30.24 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 30.223 11.553 30.257 ;
      VIA 11.508 30.24 Element_VIA34_1_2_58_52 ;
      VIA 11.508 30.24 Element_VIA23_1_3_36_36 ;
      VIA 11.508 29.7 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 29.683 11.553 29.717 ;
      VIA 11.508 29.7 Element_VIA34_1_2_58_52 ;
      VIA 11.508 29.7 Element_VIA23_1_3_36_36 ;
      VIA 11.508 29.16 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 29.143 11.553 29.177 ;
      VIA 11.508 29.16 Element_VIA34_1_2_58_52 ;
      VIA 11.508 29.16 Element_VIA23_1_3_36_36 ;
      VIA 11.508 28.62 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 28.603 11.553 28.637 ;
      VIA 11.508 28.62 Element_VIA34_1_2_58_52 ;
      VIA 11.508 28.62 Element_VIA23_1_3_36_36 ;
      VIA 11.508 28.08 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 28.063 11.553 28.097 ;
      VIA 11.508 28.08 Element_VIA34_1_2_58_52 ;
      VIA 11.508 28.08 Element_VIA23_1_3_36_36 ;
      VIA 11.508 27.54 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 27.523 11.553 27.557 ;
      VIA 11.508 27.54 Element_VIA34_1_2_58_52 ;
      VIA 11.508 27.54 Element_VIA23_1_3_36_36 ;
      VIA 11.508 27 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 26.983 11.553 27.017 ;
      VIA 11.508 27 Element_VIA34_1_2_58_52 ;
      VIA 11.508 27 Element_VIA23_1_3_36_36 ;
      VIA 11.508 26.46 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 26.443 11.553 26.477 ;
      VIA 11.508 26.46 Element_VIA34_1_2_58_52 ;
      VIA 11.508 26.46 Element_VIA23_1_3_36_36 ;
      VIA 11.508 25.92 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 25.903 11.553 25.937 ;
      VIA 11.508 25.92 Element_VIA34_1_2_58_52 ;
      VIA 11.508 25.92 Element_VIA23_1_3_36_36 ;
      VIA 11.508 25.38 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 25.363 11.553 25.397 ;
      VIA 11.508 25.38 Element_VIA34_1_2_58_52 ;
      VIA 11.508 25.38 Element_VIA23_1_3_36_36 ;
      VIA 11.508 24.84 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 24.823 11.553 24.857 ;
      VIA 11.508 24.84 Element_VIA34_1_2_58_52 ;
      VIA 11.508 24.84 Element_VIA23_1_3_36_36 ;
      VIA 11.508 24.3 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 24.283 11.553 24.317 ;
      VIA 11.508 24.3 Element_VIA34_1_2_58_52 ;
      VIA 11.508 24.3 Element_VIA23_1_3_36_36 ;
      VIA 11.508 23.76 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 23.743 11.553 23.777 ;
      VIA 11.508 23.76 Element_VIA34_1_2_58_52 ;
      VIA 11.508 23.76 Element_VIA23_1_3_36_36 ;
      VIA 11.508 23.22 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 23.203 11.553 23.237 ;
      VIA 11.508 23.22 Element_VIA34_1_2_58_52 ;
      VIA 11.508 23.22 Element_VIA23_1_3_36_36 ;
      VIA 11.508 22.68 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 22.663 11.553 22.697 ;
      VIA 11.508 22.68 Element_VIA34_1_2_58_52 ;
      VIA 11.508 22.68 Element_VIA23_1_3_36_36 ;
      VIA 11.508 22.14 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 22.123 11.553 22.157 ;
      VIA 11.508 22.14 Element_VIA34_1_2_58_52 ;
      VIA 11.508 22.14 Element_VIA23_1_3_36_36 ;
      VIA 11.508 21.6 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 21.583 11.553 21.617 ;
      VIA 11.508 21.6 Element_VIA34_1_2_58_52 ;
      VIA 11.508 21.6 Element_VIA23_1_3_36_36 ;
      VIA 11.508 21.06 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 21.043 11.553 21.077 ;
      VIA 11.508 21.06 Element_VIA34_1_2_58_52 ;
      VIA 11.508 21.06 Element_VIA23_1_3_36_36 ;
      VIA 11.508 20.52 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 20.503 11.553 20.537 ;
      VIA 11.508 20.52 Element_VIA34_1_2_58_52 ;
      VIA 11.508 20.52 Element_VIA23_1_3_36_36 ;
      VIA 11.508 19.98 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 19.963 11.553 19.997 ;
      VIA 11.508 19.98 Element_VIA34_1_2_58_52 ;
      VIA 11.508 19.98 Element_VIA23_1_3_36_36 ;
      VIA 11.508 19.44 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 19.423 11.553 19.457 ;
      VIA 11.508 19.44 Element_VIA34_1_2_58_52 ;
      VIA 11.508 19.44 Element_VIA23_1_3_36_36 ;
      VIA 11.508 18.9 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 18.883 11.553 18.917 ;
      VIA 11.508 18.9 Element_VIA34_1_2_58_52 ;
      VIA 11.508 18.9 Element_VIA23_1_3_36_36 ;
      VIA 11.508 18.36 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 18.343 11.553 18.377 ;
      VIA 11.508 18.36 Element_VIA34_1_2_58_52 ;
      VIA 11.508 18.36 Element_VIA23_1_3_36_36 ;
      VIA 11.508 17.82 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 17.803 11.553 17.837 ;
      VIA 11.508 17.82 Element_VIA34_1_2_58_52 ;
      VIA 11.508 17.82 Element_VIA23_1_3_36_36 ;
      VIA 11.508 17.28 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 17.263 11.553 17.297 ;
      VIA 11.508 17.28 Element_VIA34_1_2_58_52 ;
      VIA 11.508 17.28 Element_VIA23_1_3_36_36 ;
      VIA 11.508 16.74 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 16.723 11.553 16.757 ;
      VIA 11.508 16.74 Element_VIA34_1_2_58_52 ;
      VIA 11.508 16.74 Element_VIA23_1_3_36_36 ;
      VIA 11.508 16.2 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 16.183 11.553 16.217 ;
      VIA 11.508 16.2 Element_VIA34_1_2_58_52 ;
      VIA 11.508 16.2 Element_VIA23_1_3_36_36 ;
      VIA 11.508 15.66 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 15.643 11.553 15.677 ;
      VIA 11.508 15.66 Element_VIA34_1_2_58_52 ;
      VIA 11.508 15.66 Element_VIA23_1_3_36_36 ;
      VIA 11.508 15.12 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 15.103 11.553 15.137 ;
      VIA 11.508 15.12 Element_VIA34_1_2_58_52 ;
      VIA 11.508 15.12 Element_VIA23_1_3_36_36 ;
      VIA 11.508 14.58 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 14.563 11.553 14.597 ;
      VIA 11.508 14.58 Element_VIA34_1_2_58_52 ;
      VIA 11.508 14.58 Element_VIA23_1_3_36_36 ;
      VIA 11.508 14.04 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 14.023 11.553 14.057 ;
      VIA 11.508 14.04 Element_VIA34_1_2_58_52 ;
      VIA 11.508 14.04 Element_VIA23_1_3_36_36 ;
      VIA 11.508 13.5 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 13.483 11.553 13.517 ;
      VIA 11.508 13.5 Element_VIA34_1_2_58_52 ;
      VIA 11.508 13.5 Element_VIA23_1_3_36_36 ;
      VIA 11.508 12.96 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 12.943 11.553 12.977 ;
      VIA 11.508 12.96 Element_VIA34_1_2_58_52 ;
      VIA 11.508 12.96 Element_VIA23_1_3_36_36 ;
      VIA 11.508 12.42 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 12.403 11.553 12.437 ;
      VIA 11.508 12.42 Element_VIA34_1_2_58_52 ;
      VIA 11.508 12.42 Element_VIA23_1_3_36_36 ;
      VIA 11.508 11.88 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 11.863 11.553 11.897 ;
      VIA 11.508 11.88 Element_VIA34_1_2_58_52 ;
      VIA 11.508 11.88 Element_VIA23_1_3_36_36 ;
      VIA 11.508 11.34 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 11.323 11.553 11.357 ;
      VIA 11.508 11.34 Element_VIA34_1_2_58_52 ;
      VIA 11.508 11.34 Element_VIA23_1_3_36_36 ;
      VIA 11.508 10.8 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 10.783 11.553 10.817 ;
      VIA 11.508 10.8 Element_VIA34_1_2_58_52 ;
      VIA 11.508 10.8 Element_VIA23_1_3_36_36 ;
      VIA 11.508 10.26 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 10.243 11.553 10.277 ;
      VIA 11.508 10.26 Element_VIA34_1_2_58_52 ;
      VIA 11.508 10.26 Element_VIA23_1_3_36_36 ;
      VIA 11.508 9.72 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 9.703 11.553 9.737 ;
      VIA 11.508 9.72 Element_VIA34_1_2_58_52 ;
      VIA 11.508 9.72 Element_VIA23_1_3_36_36 ;
      VIA 11.508 9.18 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 9.163 11.553 9.197 ;
      VIA 11.508 9.18 Element_VIA34_1_2_58_52 ;
      VIA 11.508 9.18 Element_VIA23_1_3_36_36 ;
      VIA 11.508 8.64 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 8.623 11.553 8.657 ;
      VIA 11.508 8.64 Element_VIA34_1_2_58_52 ;
      VIA 11.508 8.64 Element_VIA23_1_3_36_36 ;
      VIA 11.508 8.1 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 8.083 11.553 8.117 ;
      VIA 11.508 8.1 Element_VIA34_1_2_58_52 ;
      VIA 11.508 8.1 Element_VIA23_1_3_36_36 ;
      VIA 11.508 7.56 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 7.543 11.553 7.577 ;
      VIA 11.508 7.56 Element_VIA34_1_2_58_52 ;
      VIA 11.508 7.56 Element_VIA23_1_3_36_36 ;
      VIA 11.508 7.02 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 7.003 11.553 7.037 ;
      VIA 11.508 7.02 Element_VIA34_1_2_58_52 ;
      VIA 11.508 7.02 Element_VIA23_1_3_36_36 ;
      VIA 11.508 6.48 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 6.463 11.553 6.497 ;
      VIA 11.508 6.48 Element_VIA34_1_2_58_52 ;
      VIA 11.508 6.48 Element_VIA23_1_3_36_36 ;
      VIA 11.508 5.94 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 5.923 11.553 5.957 ;
      VIA 11.508 5.94 Element_VIA34_1_2_58_52 ;
      VIA 11.508 5.94 Element_VIA23_1_3_36_36 ;
      VIA 11.508 5.4 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 5.383 11.553 5.417 ;
      VIA 11.508 5.4 Element_VIA34_1_2_58_52 ;
      VIA 11.508 5.4 Element_VIA23_1_3_36_36 ;
      VIA 11.508 4.86 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 4.843 11.553 4.877 ;
      VIA 11.508 4.86 Element_VIA34_1_2_58_52 ;
      VIA 11.508 4.86 Element_VIA23_1_3_36_36 ;
      VIA 11.508 4.32 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 4.303 11.553 4.337 ;
      VIA 11.508 4.32 Element_VIA34_1_2_58_52 ;
      VIA 11.508 4.32 Element_VIA23_1_3_36_36 ;
      VIA 11.508 3.78 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 3.763 11.553 3.797 ;
      VIA 11.508 3.78 Element_VIA34_1_2_58_52 ;
      VIA 11.508 3.78 Element_VIA23_1_3_36_36 ;
      VIA 11.508 3.24 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 3.223 11.553 3.257 ;
      VIA 11.508 3.24 Element_VIA34_1_2_58_52 ;
      VIA 11.508 3.24 Element_VIA23_1_3_36_36 ;
      VIA 11.508 2.7 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 2.683 11.553 2.717 ;
      VIA 11.508 2.7 Element_VIA34_1_2_58_52 ;
      VIA 11.508 2.7 Element_VIA23_1_3_36_36 ;
      VIA 11.508 2.16 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 2.143 11.553 2.177 ;
      VIA 11.508 2.16 Element_VIA34_1_2_58_52 ;
      VIA 11.508 2.16 Element_VIA23_1_3_36_36 ;
      VIA 11.508 1.62 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 1.603 11.553 1.637 ;
      VIA 11.508 1.62 Element_VIA34_1_2_58_52 ;
      VIA 11.508 1.62 Element_VIA23_1_3_36_36 ;
      VIA 11.508 1.08 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  11.463 1.063 11.553 1.097 ;
      VIA 11.508 1.08 Element_VIA34_1_2_58_52 ;
      VIA 11.508 1.08 Element_VIA23_1_3_36_36 ;
      VIA 8.532 42.12 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 42.103 8.577 42.137 ;
      VIA 8.532 42.12 Element_VIA34_1_2_58_52 ;
      VIA 8.532 42.12 Element_VIA23_1_3_36_36 ;
      VIA 8.532 41.58 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 41.563 8.577 41.597 ;
      VIA 8.532 41.58 Element_VIA34_1_2_58_52 ;
      VIA 8.532 41.58 Element_VIA23_1_3_36_36 ;
      VIA 8.532 41.04 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 41.023 8.577 41.057 ;
      VIA 8.532 41.04 Element_VIA34_1_2_58_52 ;
      VIA 8.532 41.04 Element_VIA23_1_3_36_36 ;
      VIA 8.532 40.5 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 40.483 8.577 40.517 ;
      VIA 8.532 40.5 Element_VIA34_1_2_58_52 ;
      VIA 8.532 40.5 Element_VIA23_1_3_36_36 ;
      VIA 8.532 39.96 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 39.943 8.577 39.977 ;
      VIA 8.532 39.96 Element_VIA34_1_2_58_52 ;
      VIA 8.532 39.96 Element_VIA23_1_3_36_36 ;
      VIA 8.532 39.42 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 39.403 8.577 39.437 ;
      VIA 8.532 39.42 Element_VIA34_1_2_58_52 ;
      VIA 8.532 39.42 Element_VIA23_1_3_36_36 ;
      VIA 8.532 38.88 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 38.863 8.577 38.897 ;
      VIA 8.532 38.88 Element_VIA34_1_2_58_52 ;
      VIA 8.532 38.88 Element_VIA23_1_3_36_36 ;
      VIA 8.532 38.34 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 38.323 8.577 38.357 ;
      VIA 8.532 38.34 Element_VIA34_1_2_58_52 ;
      VIA 8.532 38.34 Element_VIA23_1_3_36_36 ;
      VIA 8.532 37.8 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 37.783 8.577 37.817 ;
      VIA 8.532 37.8 Element_VIA34_1_2_58_52 ;
      VIA 8.532 37.8 Element_VIA23_1_3_36_36 ;
      VIA 8.532 37.26 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 37.243 8.577 37.277 ;
      VIA 8.532 37.26 Element_VIA34_1_2_58_52 ;
      VIA 8.532 37.26 Element_VIA23_1_3_36_36 ;
      VIA 8.532 36.72 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 36.703 8.577 36.737 ;
      VIA 8.532 36.72 Element_VIA34_1_2_58_52 ;
      VIA 8.532 36.72 Element_VIA23_1_3_36_36 ;
      VIA 8.532 36.18 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 36.163 8.577 36.197 ;
      VIA 8.532 36.18 Element_VIA34_1_2_58_52 ;
      VIA 8.532 36.18 Element_VIA23_1_3_36_36 ;
      VIA 8.532 35.64 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 35.623 8.577 35.657 ;
      VIA 8.532 35.64 Element_VIA34_1_2_58_52 ;
      VIA 8.532 35.64 Element_VIA23_1_3_36_36 ;
      VIA 8.532 35.1 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 35.083 8.577 35.117 ;
      VIA 8.532 35.1 Element_VIA34_1_2_58_52 ;
      VIA 8.532 35.1 Element_VIA23_1_3_36_36 ;
      VIA 8.532 34.56 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 34.543 8.577 34.577 ;
      VIA 8.532 34.56 Element_VIA34_1_2_58_52 ;
      VIA 8.532 34.56 Element_VIA23_1_3_36_36 ;
      VIA 8.532 34.02 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 34.003 8.577 34.037 ;
      VIA 8.532 34.02 Element_VIA34_1_2_58_52 ;
      VIA 8.532 34.02 Element_VIA23_1_3_36_36 ;
      VIA 8.532 33.48 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 33.463 8.577 33.497 ;
      VIA 8.532 33.48 Element_VIA34_1_2_58_52 ;
      VIA 8.532 33.48 Element_VIA23_1_3_36_36 ;
      VIA 8.532 32.94 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 32.923 8.577 32.957 ;
      VIA 8.532 32.94 Element_VIA34_1_2_58_52 ;
      VIA 8.532 32.94 Element_VIA23_1_3_36_36 ;
      VIA 8.532 32.4 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 32.383 8.577 32.417 ;
      VIA 8.532 32.4 Element_VIA34_1_2_58_52 ;
      VIA 8.532 32.4 Element_VIA23_1_3_36_36 ;
      VIA 8.532 31.86 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 31.843 8.577 31.877 ;
      VIA 8.532 31.86 Element_VIA34_1_2_58_52 ;
      VIA 8.532 31.86 Element_VIA23_1_3_36_36 ;
      VIA 8.532 31.32 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 31.303 8.577 31.337 ;
      VIA 8.532 31.32 Element_VIA34_1_2_58_52 ;
      VIA 8.532 31.32 Element_VIA23_1_3_36_36 ;
      VIA 8.532 30.78 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 30.763 8.577 30.797 ;
      VIA 8.532 30.78 Element_VIA34_1_2_58_52 ;
      VIA 8.532 30.78 Element_VIA23_1_3_36_36 ;
      VIA 8.532 30.24 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 30.223 8.577 30.257 ;
      VIA 8.532 30.24 Element_VIA34_1_2_58_52 ;
      VIA 8.532 30.24 Element_VIA23_1_3_36_36 ;
      VIA 8.532 29.7 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 29.683 8.577 29.717 ;
      VIA 8.532 29.7 Element_VIA34_1_2_58_52 ;
      VIA 8.532 29.7 Element_VIA23_1_3_36_36 ;
      VIA 8.532 29.16 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 29.143 8.577 29.177 ;
      VIA 8.532 29.16 Element_VIA34_1_2_58_52 ;
      VIA 8.532 29.16 Element_VIA23_1_3_36_36 ;
      VIA 8.532 28.62 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 28.603 8.577 28.637 ;
      VIA 8.532 28.62 Element_VIA34_1_2_58_52 ;
      VIA 8.532 28.62 Element_VIA23_1_3_36_36 ;
      VIA 8.532 28.08 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 28.063 8.577 28.097 ;
      VIA 8.532 28.08 Element_VIA34_1_2_58_52 ;
      VIA 8.532 28.08 Element_VIA23_1_3_36_36 ;
      VIA 8.532 27.54 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 27.523 8.577 27.557 ;
      VIA 8.532 27.54 Element_VIA34_1_2_58_52 ;
      VIA 8.532 27.54 Element_VIA23_1_3_36_36 ;
      VIA 8.532 27 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 26.983 8.577 27.017 ;
      VIA 8.532 27 Element_VIA34_1_2_58_52 ;
      VIA 8.532 27 Element_VIA23_1_3_36_36 ;
      VIA 8.532 26.46 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 26.443 8.577 26.477 ;
      VIA 8.532 26.46 Element_VIA34_1_2_58_52 ;
      VIA 8.532 26.46 Element_VIA23_1_3_36_36 ;
      VIA 8.532 25.92 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 25.903 8.577 25.937 ;
      VIA 8.532 25.92 Element_VIA34_1_2_58_52 ;
      VIA 8.532 25.92 Element_VIA23_1_3_36_36 ;
      VIA 8.532 25.38 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 25.363 8.577 25.397 ;
      VIA 8.532 25.38 Element_VIA34_1_2_58_52 ;
      VIA 8.532 25.38 Element_VIA23_1_3_36_36 ;
      VIA 8.532 24.84 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 24.823 8.577 24.857 ;
      VIA 8.532 24.84 Element_VIA34_1_2_58_52 ;
      VIA 8.532 24.84 Element_VIA23_1_3_36_36 ;
      VIA 8.532 24.3 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 24.283 8.577 24.317 ;
      VIA 8.532 24.3 Element_VIA34_1_2_58_52 ;
      VIA 8.532 24.3 Element_VIA23_1_3_36_36 ;
      VIA 8.532 23.76 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 23.743 8.577 23.777 ;
      VIA 8.532 23.76 Element_VIA34_1_2_58_52 ;
      VIA 8.532 23.76 Element_VIA23_1_3_36_36 ;
      VIA 8.532 23.22 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 23.203 8.577 23.237 ;
      VIA 8.532 23.22 Element_VIA34_1_2_58_52 ;
      VIA 8.532 23.22 Element_VIA23_1_3_36_36 ;
      VIA 8.532 22.68 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 22.663 8.577 22.697 ;
      VIA 8.532 22.68 Element_VIA34_1_2_58_52 ;
      VIA 8.532 22.68 Element_VIA23_1_3_36_36 ;
      VIA 8.532 22.14 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 22.123 8.577 22.157 ;
      VIA 8.532 22.14 Element_VIA34_1_2_58_52 ;
      VIA 8.532 22.14 Element_VIA23_1_3_36_36 ;
      VIA 8.532 21.6 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 21.583 8.577 21.617 ;
      VIA 8.532 21.6 Element_VIA34_1_2_58_52 ;
      VIA 8.532 21.6 Element_VIA23_1_3_36_36 ;
      VIA 8.532 21.06 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 21.043 8.577 21.077 ;
      VIA 8.532 21.06 Element_VIA34_1_2_58_52 ;
      VIA 8.532 21.06 Element_VIA23_1_3_36_36 ;
      VIA 8.532 20.52 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 20.503 8.577 20.537 ;
      VIA 8.532 20.52 Element_VIA34_1_2_58_52 ;
      VIA 8.532 20.52 Element_VIA23_1_3_36_36 ;
      VIA 8.532 19.98 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 19.963 8.577 19.997 ;
      VIA 8.532 19.98 Element_VIA34_1_2_58_52 ;
      VIA 8.532 19.98 Element_VIA23_1_3_36_36 ;
      VIA 8.532 19.44 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 19.423 8.577 19.457 ;
      VIA 8.532 19.44 Element_VIA34_1_2_58_52 ;
      VIA 8.532 19.44 Element_VIA23_1_3_36_36 ;
      VIA 8.532 18.9 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 18.883 8.577 18.917 ;
      VIA 8.532 18.9 Element_VIA34_1_2_58_52 ;
      VIA 8.532 18.9 Element_VIA23_1_3_36_36 ;
      VIA 8.532 18.36 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 18.343 8.577 18.377 ;
      VIA 8.532 18.36 Element_VIA34_1_2_58_52 ;
      VIA 8.532 18.36 Element_VIA23_1_3_36_36 ;
      VIA 8.532 17.82 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 17.803 8.577 17.837 ;
      VIA 8.532 17.82 Element_VIA34_1_2_58_52 ;
      VIA 8.532 17.82 Element_VIA23_1_3_36_36 ;
      VIA 8.532 17.28 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 17.263 8.577 17.297 ;
      VIA 8.532 17.28 Element_VIA34_1_2_58_52 ;
      VIA 8.532 17.28 Element_VIA23_1_3_36_36 ;
      VIA 8.532 16.74 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 16.723 8.577 16.757 ;
      VIA 8.532 16.74 Element_VIA34_1_2_58_52 ;
      VIA 8.532 16.74 Element_VIA23_1_3_36_36 ;
      VIA 8.532 16.2 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 16.183 8.577 16.217 ;
      VIA 8.532 16.2 Element_VIA34_1_2_58_52 ;
      VIA 8.532 16.2 Element_VIA23_1_3_36_36 ;
      VIA 8.532 15.66 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 15.643 8.577 15.677 ;
      VIA 8.532 15.66 Element_VIA34_1_2_58_52 ;
      VIA 8.532 15.66 Element_VIA23_1_3_36_36 ;
      VIA 8.532 15.12 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 15.103 8.577 15.137 ;
      VIA 8.532 15.12 Element_VIA34_1_2_58_52 ;
      VIA 8.532 15.12 Element_VIA23_1_3_36_36 ;
      VIA 8.532 14.58 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 14.563 8.577 14.597 ;
      VIA 8.532 14.58 Element_VIA34_1_2_58_52 ;
      VIA 8.532 14.58 Element_VIA23_1_3_36_36 ;
      VIA 8.532 14.04 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 14.023 8.577 14.057 ;
      VIA 8.532 14.04 Element_VIA34_1_2_58_52 ;
      VIA 8.532 14.04 Element_VIA23_1_3_36_36 ;
      VIA 8.532 13.5 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 13.483 8.577 13.517 ;
      VIA 8.532 13.5 Element_VIA34_1_2_58_52 ;
      VIA 8.532 13.5 Element_VIA23_1_3_36_36 ;
      VIA 8.532 12.96 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 12.943 8.577 12.977 ;
      VIA 8.532 12.96 Element_VIA34_1_2_58_52 ;
      VIA 8.532 12.96 Element_VIA23_1_3_36_36 ;
      VIA 8.532 12.42 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 12.403 8.577 12.437 ;
      VIA 8.532 12.42 Element_VIA34_1_2_58_52 ;
      VIA 8.532 12.42 Element_VIA23_1_3_36_36 ;
      VIA 8.532 11.88 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 11.863 8.577 11.897 ;
      VIA 8.532 11.88 Element_VIA34_1_2_58_52 ;
      VIA 8.532 11.88 Element_VIA23_1_3_36_36 ;
      VIA 8.532 11.34 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 11.323 8.577 11.357 ;
      VIA 8.532 11.34 Element_VIA34_1_2_58_52 ;
      VIA 8.532 11.34 Element_VIA23_1_3_36_36 ;
      VIA 8.532 10.8 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 10.783 8.577 10.817 ;
      VIA 8.532 10.8 Element_VIA34_1_2_58_52 ;
      VIA 8.532 10.8 Element_VIA23_1_3_36_36 ;
      VIA 8.532 10.26 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 10.243 8.577 10.277 ;
      VIA 8.532 10.26 Element_VIA34_1_2_58_52 ;
      VIA 8.532 10.26 Element_VIA23_1_3_36_36 ;
      VIA 8.532 9.72 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 9.703 8.577 9.737 ;
      VIA 8.532 9.72 Element_VIA34_1_2_58_52 ;
      VIA 8.532 9.72 Element_VIA23_1_3_36_36 ;
      VIA 8.532 9.18 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 9.163 8.577 9.197 ;
      VIA 8.532 9.18 Element_VIA34_1_2_58_52 ;
      VIA 8.532 9.18 Element_VIA23_1_3_36_36 ;
      VIA 8.532 8.64 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 8.623 8.577 8.657 ;
      VIA 8.532 8.64 Element_VIA34_1_2_58_52 ;
      VIA 8.532 8.64 Element_VIA23_1_3_36_36 ;
      VIA 8.532 8.1 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 8.083 8.577 8.117 ;
      VIA 8.532 8.1 Element_VIA34_1_2_58_52 ;
      VIA 8.532 8.1 Element_VIA23_1_3_36_36 ;
      VIA 8.532 7.56 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 7.543 8.577 7.577 ;
      VIA 8.532 7.56 Element_VIA34_1_2_58_52 ;
      VIA 8.532 7.56 Element_VIA23_1_3_36_36 ;
      VIA 8.532 7.02 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 7.003 8.577 7.037 ;
      VIA 8.532 7.02 Element_VIA34_1_2_58_52 ;
      VIA 8.532 7.02 Element_VIA23_1_3_36_36 ;
      VIA 8.532 6.48 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 6.463 8.577 6.497 ;
      VIA 8.532 6.48 Element_VIA34_1_2_58_52 ;
      VIA 8.532 6.48 Element_VIA23_1_3_36_36 ;
      VIA 8.532 5.94 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 5.923 8.577 5.957 ;
      VIA 8.532 5.94 Element_VIA34_1_2_58_52 ;
      VIA 8.532 5.94 Element_VIA23_1_3_36_36 ;
      VIA 8.532 5.4 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 5.383 8.577 5.417 ;
      VIA 8.532 5.4 Element_VIA34_1_2_58_52 ;
      VIA 8.532 5.4 Element_VIA23_1_3_36_36 ;
      VIA 8.532 4.86 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 4.843 8.577 4.877 ;
      VIA 8.532 4.86 Element_VIA34_1_2_58_52 ;
      VIA 8.532 4.86 Element_VIA23_1_3_36_36 ;
      VIA 8.532 4.32 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 4.303 8.577 4.337 ;
      VIA 8.532 4.32 Element_VIA34_1_2_58_52 ;
      VIA 8.532 4.32 Element_VIA23_1_3_36_36 ;
      VIA 8.532 3.78 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 3.763 8.577 3.797 ;
      VIA 8.532 3.78 Element_VIA34_1_2_58_52 ;
      VIA 8.532 3.78 Element_VIA23_1_3_36_36 ;
      VIA 8.532 3.24 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 3.223 8.577 3.257 ;
      VIA 8.532 3.24 Element_VIA34_1_2_58_52 ;
      VIA 8.532 3.24 Element_VIA23_1_3_36_36 ;
      VIA 8.532 2.7 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 2.683 8.577 2.717 ;
      VIA 8.532 2.7 Element_VIA34_1_2_58_52 ;
      VIA 8.532 2.7 Element_VIA23_1_3_36_36 ;
      VIA 8.532 2.16 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 2.143 8.577 2.177 ;
      VIA 8.532 2.16 Element_VIA34_1_2_58_52 ;
      VIA 8.532 2.16 Element_VIA23_1_3_36_36 ;
      VIA 8.532 1.62 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 1.603 8.577 1.637 ;
      VIA 8.532 1.62 Element_VIA34_1_2_58_52 ;
      VIA 8.532 1.62 Element_VIA23_1_3_36_36 ;
      VIA 8.532 1.08 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  8.487 1.063 8.577 1.097 ;
      VIA 8.532 1.08 Element_VIA34_1_2_58_52 ;
      VIA 8.532 1.08 Element_VIA23_1_3_36_36 ;
      VIA 5.556 42.12 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 42.103 5.601 42.137 ;
      VIA 5.556 42.12 Element_VIA34_1_2_58_52 ;
      VIA 5.556 42.12 Element_VIA23_1_3_36_36 ;
      VIA 5.556 41.58 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 41.563 5.601 41.597 ;
      VIA 5.556 41.58 Element_VIA34_1_2_58_52 ;
      VIA 5.556 41.58 Element_VIA23_1_3_36_36 ;
      VIA 5.556 41.04 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 41.023 5.601 41.057 ;
      VIA 5.556 41.04 Element_VIA34_1_2_58_52 ;
      VIA 5.556 41.04 Element_VIA23_1_3_36_36 ;
      VIA 5.556 40.5 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 40.483 5.601 40.517 ;
      VIA 5.556 40.5 Element_VIA34_1_2_58_52 ;
      VIA 5.556 40.5 Element_VIA23_1_3_36_36 ;
      VIA 5.556 39.96 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 39.943 5.601 39.977 ;
      VIA 5.556 39.96 Element_VIA34_1_2_58_52 ;
      VIA 5.556 39.96 Element_VIA23_1_3_36_36 ;
      VIA 5.556 39.42 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 39.403 5.601 39.437 ;
      VIA 5.556 39.42 Element_VIA34_1_2_58_52 ;
      VIA 5.556 39.42 Element_VIA23_1_3_36_36 ;
      VIA 5.556 38.88 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 38.863 5.601 38.897 ;
      VIA 5.556 38.88 Element_VIA34_1_2_58_52 ;
      VIA 5.556 38.88 Element_VIA23_1_3_36_36 ;
      VIA 5.556 38.34 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 38.323 5.601 38.357 ;
      VIA 5.556 38.34 Element_VIA34_1_2_58_52 ;
      VIA 5.556 38.34 Element_VIA23_1_3_36_36 ;
      VIA 5.556 37.8 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 37.783 5.601 37.817 ;
      VIA 5.556 37.8 Element_VIA34_1_2_58_52 ;
      VIA 5.556 37.8 Element_VIA23_1_3_36_36 ;
      VIA 5.556 37.26 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 37.243 5.601 37.277 ;
      VIA 5.556 37.26 Element_VIA34_1_2_58_52 ;
      VIA 5.556 37.26 Element_VIA23_1_3_36_36 ;
      VIA 5.556 36.72 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 36.703 5.601 36.737 ;
      VIA 5.556 36.72 Element_VIA34_1_2_58_52 ;
      VIA 5.556 36.72 Element_VIA23_1_3_36_36 ;
      VIA 5.556 36.18 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 36.163 5.601 36.197 ;
      VIA 5.556 36.18 Element_VIA34_1_2_58_52 ;
      VIA 5.556 36.18 Element_VIA23_1_3_36_36 ;
      VIA 5.556 35.64 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 35.623 5.601 35.657 ;
      VIA 5.556 35.64 Element_VIA34_1_2_58_52 ;
      VIA 5.556 35.64 Element_VIA23_1_3_36_36 ;
      VIA 5.556 35.1 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 35.083 5.601 35.117 ;
      VIA 5.556 35.1 Element_VIA34_1_2_58_52 ;
      VIA 5.556 35.1 Element_VIA23_1_3_36_36 ;
      VIA 5.556 34.56 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 34.543 5.601 34.577 ;
      VIA 5.556 34.56 Element_VIA34_1_2_58_52 ;
      VIA 5.556 34.56 Element_VIA23_1_3_36_36 ;
      VIA 5.556 34.02 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 34.003 5.601 34.037 ;
      VIA 5.556 34.02 Element_VIA34_1_2_58_52 ;
      VIA 5.556 34.02 Element_VIA23_1_3_36_36 ;
      VIA 5.556 33.48 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 33.463 5.601 33.497 ;
      VIA 5.556 33.48 Element_VIA34_1_2_58_52 ;
      VIA 5.556 33.48 Element_VIA23_1_3_36_36 ;
      VIA 5.556 32.94 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 32.923 5.601 32.957 ;
      VIA 5.556 32.94 Element_VIA34_1_2_58_52 ;
      VIA 5.556 32.94 Element_VIA23_1_3_36_36 ;
      VIA 5.556 32.4 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 32.383 5.601 32.417 ;
      VIA 5.556 32.4 Element_VIA34_1_2_58_52 ;
      VIA 5.556 32.4 Element_VIA23_1_3_36_36 ;
      VIA 5.556 31.86 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 31.843 5.601 31.877 ;
      VIA 5.556 31.86 Element_VIA34_1_2_58_52 ;
      VIA 5.556 31.86 Element_VIA23_1_3_36_36 ;
      VIA 5.556 31.32 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 31.303 5.601 31.337 ;
      VIA 5.556 31.32 Element_VIA34_1_2_58_52 ;
      VIA 5.556 31.32 Element_VIA23_1_3_36_36 ;
      VIA 5.556 30.78 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 30.763 5.601 30.797 ;
      VIA 5.556 30.78 Element_VIA34_1_2_58_52 ;
      VIA 5.556 30.78 Element_VIA23_1_3_36_36 ;
      VIA 5.556 30.24 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 30.223 5.601 30.257 ;
      VIA 5.556 30.24 Element_VIA34_1_2_58_52 ;
      VIA 5.556 30.24 Element_VIA23_1_3_36_36 ;
      VIA 5.556 29.7 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 29.683 5.601 29.717 ;
      VIA 5.556 29.7 Element_VIA34_1_2_58_52 ;
      VIA 5.556 29.7 Element_VIA23_1_3_36_36 ;
      VIA 5.556 29.16 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 29.143 5.601 29.177 ;
      VIA 5.556 29.16 Element_VIA34_1_2_58_52 ;
      VIA 5.556 29.16 Element_VIA23_1_3_36_36 ;
      VIA 5.556 28.62 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 28.603 5.601 28.637 ;
      VIA 5.556 28.62 Element_VIA34_1_2_58_52 ;
      VIA 5.556 28.62 Element_VIA23_1_3_36_36 ;
      VIA 5.556 28.08 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 28.063 5.601 28.097 ;
      VIA 5.556 28.08 Element_VIA34_1_2_58_52 ;
      VIA 5.556 28.08 Element_VIA23_1_3_36_36 ;
      VIA 5.556 27.54 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 27.523 5.601 27.557 ;
      VIA 5.556 27.54 Element_VIA34_1_2_58_52 ;
      VIA 5.556 27.54 Element_VIA23_1_3_36_36 ;
      VIA 5.556 27 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 26.983 5.601 27.017 ;
      VIA 5.556 27 Element_VIA34_1_2_58_52 ;
      VIA 5.556 27 Element_VIA23_1_3_36_36 ;
      VIA 5.556 26.46 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 26.443 5.601 26.477 ;
      VIA 5.556 26.46 Element_VIA34_1_2_58_52 ;
      VIA 5.556 26.46 Element_VIA23_1_3_36_36 ;
      VIA 5.556 25.92 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 25.903 5.601 25.937 ;
      VIA 5.556 25.92 Element_VIA34_1_2_58_52 ;
      VIA 5.556 25.92 Element_VIA23_1_3_36_36 ;
      VIA 5.556 25.38 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 25.363 5.601 25.397 ;
      VIA 5.556 25.38 Element_VIA34_1_2_58_52 ;
      VIA 5.556 25.38 Element_VIA23_1_3_36_36 ;
      VIA 5.556 24.84 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 24.823 5.601 24.857 ;
      VIA 5.556 24.84 Element_VIA34_1_2_58_52 ;
      VIA 5.556 24.84 Element_VIA23_1_3_36_36 ;
      VIA 5.556 24.3 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 24.283 5.601 24.317 ;
      VIA 5.556 24.3 Element_VIA34_1_2_58_52 ;
      VIA 5.556 24.3 Element_VIA23_1_3_36_36 ;
      VIA 5.556 23.76 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 23.743 5.601 23.777 ;
      VIA 5.556 23.76 Element_VIA34_1_2_58_52 ;
      VIA 5.556 23.76 Element_VIA23_1_3_36_36 ;
      VIA 5.556 23.22 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 23.203 5.601 23.237 ;
      VIA 5.556 23.22 Element_VIA34_1_2_58_52 ;
      VIA 5.556 23.22 Element_VIA23_1_3_36_36 ;
      VIA 5.556 22.68 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 22.663 5.601 22.697 ;
      VIA 5.556 22.68 Element_VIA34_1_2_58_52 ;
      VIA 5.556 22.68 Element_VIA23_1_3_36_36 ;
      VIA 5.556 22.14 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 22.123 5.601 22.157 ;
      VIA 5.556 22.14 Element_VIA34_1_2_58_52 ;
      VIA 5.556 22.14 Element_VIA23_1_3_36_36 ;
      VIA 5.556 21.6 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 21.583 5.601 21.617 ;
      VIA 5.556 21.6 Element_VIA34_1_2_58_52 ;
      VIA 5.556 21.6 Element_VIA23_1_3_36_36 ;
      VIA 5.556 21.06 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 21.043 5.601 21.077 ;
      VIA 5.556 21.06 Element_VIA34_1_2_58_52 ;
      VIA 5.556 21.06 Element_VIA23_1_3_36_36 ;
      VIA 5.556 20.52 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 20.503 5.601 20.537 ;
      VIA 5.556 20.52 Element_VIA34_1_2_58_52 ;
      VIA 5.556 20.52 Element_VIA23_1_3_36_36 ;
      VIA 5.556 19.98 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 19.963 5.601 19.997 ;
      VIA 5.556 19.98 Element_VIA34_1_2_58_52 ;
      VIA 5.556 19.98 Element_VIA23_1_3_36_36 ;
      VIA 5.556 19.44 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 19.423 5.601 19.457 ;
      VIA 5.556 19.44 Element_VIA34_1_2_58_52 ;
      VIA 5.556 19.44 Element_VIA23_1_3_36_36 ;
      VIA 5.556 18.9 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 18.883 5.601 18.917 ;
      VIA 5.556 18.9 Element_VIA34_1_2_58_52 ;
      VIA 5.556 18.9 Element_VIA23_1_3_36_36 ;
      VIA 5.556 18.36 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 18.343 5.601 18.377 ;
      VIA 5.556 18.36 Element_VIA34_1_2_58_52 ;
      VIA 5.556 18.36 Element_VIA23_1_3_36_36 ;
      VIA 5.556 17.82 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 17.803 5.601 17.837 ;
      VIA 5.556 17.82 Element_VIA34_1_2_58_52 ;
      VIA 5.556 17.82 Element_VIA23_1_3_36_36 ;
      VIA 5.556 17.28 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 17.263 5.601 17.297 ;
      VIA 5.556 17.28 Element_VIA34_1_2_58_52 ;
      VIA 5.556 17.28 Element_VIA23_1_3_36_36 ;
      VIA 5.556 16.74 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 16.723 5.601 16.757 ;
      VIA 5.556 16.74 Element_VIA34_1_2_58_52 ;
      VIA 5.556 16.74 Element_VIA23_1_3_36_36 ;
      VIA 5.556 16.2 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 16.183 5.601 16.217 ;
      VIA 5.556 16.2 Element_VIA34_1_2_58_52 ;
      VIA 5.556 16.2 Element_VIA23_1_3_36_36 ;
      VIA 5.556 15.66 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 15.643 5.601 15.677 ;
      VIA 5.556 15.66 Element_VIA34_1_2_58_52 ;
      VIA 5.556 15.66 Element_VIA23_1_3_36_36 ;
      VIA 5.556 15.12 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 15.103 5.601 15.137 ;
      VIA 5.556 15.12 Element_VIA34_1_2_58_52 ;
      VIA 5.556 15.12 Element_VIA23_1_3_36_36 ;
      VIA 5.556 14.58 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 14.563 5.601 14.597 ;
      VIA 5.556 14.58 Element_VIA34_1_2_58_52 ;
      VIA 5.556 14.58 Element_VIA23_1_3_36_36 ;
      VIA 5.556 14.04 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 14.023 5.601 14.057 ;
      VIA 5.556 14.04 Element_VIA34_1_2_58_52 ;
      VIA 5.556 14.04 Element_VIA23_1_3_36_36 ;
      VIA 5.556 13.5 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 13.483 5.601 13.517 ;
      VIA 5.556 13.5 Element_VIA34_1_2_58_52 ;
      VIA 5.556 13.5 Element_VIA23_1_3_36_36 ;
      VIA 5.556 12.96 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 12.943 5.601 12.977 ;
      VIA 5.556 12.96 Element_VIA34_1_2_58_52 ;
      VIA 5.556 12.96 Element_VIA23_1_3_36_36 ;
      VIA 5.556 12.42 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 12.403 5.601 12.437 ;
      VIA 5.556 12.42 Element_VIA34_1_2_58_52 ;
      VIA 5.556 12.42 Element_VIA23_1_3_36_36 ;
      VIA 5.556 11.88 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 11.863 5.601 11.897 ;
      VIA 5.556 11.88 Element_VIA34_1_2_58_52 ;
      VIA 5.556 11.88 Element_VIA23_1_3_36_36 ;
      VIA 5.556 11.34 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 11.323 5.601 11.357 ;
      VIA 5.556 11.34 Element_VIA34_1_2_58_52 ;
      VIA 5.556 11.34 Element_VIA23_1_3_36_36 ;
      VIA 5.556 10.8 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 10.783 5.601 10.817 ;
      VIA 5.556 10.8 Element_VIA34_1_2_58_52 ;
      VIA 5.556 10.8 Element_VIA23_1_3_36_36 ;
      VIA 5.556 10.26 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 10.243 5.601 10.277 ;
      VIA 5.556 10.26 Element_VIA34_1_2_58_52 ;
      VIA 5.556 10.26 Element_VIA23_1_3_36_36 ;
      VIA 5.556 9.72 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 9.703 5.601 9.737 ;
      VIA 5.556 9.72 Element_VIA34_1_2_58_52 ;
      VIA 5.556 9.72 Element_VIA23_1_3_36_36 ;
      VIA 5.556 9.18 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 9.163 5.601 9.197 ;
      VIA 5.556 9.18 Element_VIA34_1_2_58_52 ;
      VIA 5.556 9.18 Element_VIA23_1_3_36_36 ;
      VIA 5.556 8.64 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 8.623 5.601 8.657 ;
      VIA 5.556 8.64 Element_VIA34_1_2_58_52 ;
      VIA 5.556 8.64 Element_VIA23_1_3_36_36 ;
      VIA 5.556 8.1 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 8.083 5.601 8.117 ;
      VIA 5.556 8.1 Element_VIA34_1_2_58_52 ;
      VIA 5.556 8.1 Element_VIA23_1_3_36_36 ;
      VIA 5.556 7.56 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 7.543 5.601 7.577 ;
      VIA 5.556 7.56 Element_VIA34_1_2_58_52 ;
      VIA 5.556 7.56 Element_VIA23_1_3_36_36 ;
      VIA 5.556 7.02 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 7.003 5.601 7.037 ;
      VIA 5.556 7.02 Element_VIA34_1_2_58_52 ;
      VIA 5.556 7.02 Element_VIA23_1_3_36_36 ;
      VIA 5.556 6.48 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 6.463 5.601 6.497 ;
      VIA 5.556 6.48 Element_VIA34_1_2_58_52 ;
      VIA 5.556 6.48 Element_VIA23_1_3_36_36 ;
      VIA 5.556 5.94 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 5.923 5.601 5.957 ;
      VIA 5.556 5.94 Element_VIA34_1_2_58_52 ;
      VIA 5.556 5.94 Element_VIA23_1_3_36_36 ;
      VIA 5.556 5.4 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 5.383 5.601 5.417 ;
      VIA 5.556 5.4 Element_VIA34_1_2_58_52 ;
      VIA 5.556 5.4 Element_VIA23_1_3_36_36 ;
      VIA 5.556 4.86 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 4.843 5.601 4.877 ;
      VIA 5.556 4.86 Element_VIA34_1_2_58_52 ;
      VIA 5.556 4.86 Element_VIA23_1_3_36_36 ;
      VIA 5.556 4.32 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 4.303 5.601 4.337 ;
      VIA 5.556 4.32 Element_VIA34_1_2_58_52 ;
      VIA 5.556 4.32 Element_VIA23_1_3_36_36 ;
      VIA 5.556 3.78 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 3.763 5.601 3.797 ;
      VIA 5.556 3.78 Element_VIA34_1_2_58_52 ;
      VIA 5.556 3.78 Element_VIA23_1_3_36_36 ;
      VIA 5.556 3.24 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 3.223 5.601 3.257 ;
      VIA 5.556 3.24 Element_VIA34_1_2_58_52 ;
      VIA 5.556 3.24 Element_VIA23_1_3_36_36 ;
      VIA 5.556 2.7 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 2.683 5.601 2.717 ;
      VIA 5.556 2.7 Element_VIA34_1_2_58_52 ;
      VIA 5.556 2.7 Element_VIA23_1_3_36_36 ;
      VIA 5.556 2.16 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 2.143 5.601 2.177 ;
      VIA 5.556 2.16 Element_VIA34_1_2_58_52 ;
      VIA 5.556 2.16 Element_VIA23_1_3_36_36 ;
      VIA 5.556 1.62 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 1.603 5.601 1.637 ;
      VIA 5.556 1.62 Element_VIA34_1_2_58_52 ;
      VIA 5.556 1.62 Element_VIA23_1_3_36_36 ;
      VIA 5.556 1.08 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  5.511 1.063 5.601 1.097 ;
      VIA 5.556 1.08 Element_VIA34_1_2_58_52 ;
      VIA 5.556 1.08 Element_VIA23_1_3_36_36 ;
      VIA 2.58 42.12 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 42.103 2.625 42.137 ;
      VIA 2.58 42.12 Element_VIA34_1_2_58_52 ;
      VIA 2.58 42.12 Element_VIA23_1_3_36_36 ;
      VIA 2.58 41.58 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 41.563 2.625 41.597 ;
      VIA 2.58 41.58 Element_VIA34_1_2_58_52 ;
      VIA 2.58 41.58 Element_VIA23_1_3_36_36 ;
      VIA 2.58 41.04 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 41.023 2.625 41.057 ;
      VIA 2.58 41.04 Element_VIA34_1_2_58_52 ;
      VIA 2.58 41.04 Element_VIA23_1_3_36_36 ;
      VIA 2.58 40.5 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 40.483 2.625 40.517 ;
      VIA 2.58 40.5 Element_VIA34_1_2_58_52 ;
      VIA 2.58 40.5 Element_VIA23_1_3_36_36 ;
      VIA 2.58 39.96 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 39.943 2.625 39.977 ;
      VIA 2.58 39.96 Element_VIA34_1_2_58_52 ;
      VIA 2.58 39.96 Element_VIA23_1_3_36_36 ;
      VIA 2.58 39.42 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 39.403 2.625 39.437 ;
      VIA 2.58 39.42 Element_VIA34_1_2_58_52 ;
      VIA 2.58 39.42 Element_VIA23_1_3_36_36 ;
      VIA 2.58 38.88 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 38.863 2.625 38.897 ;
      VIA 2.58 38.88 Element_VIA34_1_2_58_52 ;
      VIA 2.58 38.88 Element_VIA23_1_3_36_36 ;
      VIA 2.58 38.34 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 38.323 2.625 38.357 ;
      VIA 2.58 38.34 Element_VIA34_1_2_58_52 ;
      VIA 2.58 38.34 Element_VIA23_1_3_36_36 ;
      VIA 2.58 37.8 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 37.783 2.625 37.817 ;
      VIA 2.58 37.8 Element_VIA34_1_2_58_52 ;
      VIA 2.58 37.8 Element_VIA23_1_3_36_36 ;
      VIA 2.58 37.26 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 37.243 2.625 37.277 ;
      VIA 2.58 37.26 Element_VIA34_1_2_58_52 ;
      VIA 2.58 37.26 Element_VIA23_1_3_36_36 ;
      VIA 2.58 36.72 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 36.703 2.625 36.737 ;
      VIA 2.58 36.72 Element_VIA34_1_2_58_52 ;
      VIA 2.58 36.72 Element_VIA23_1_3_36_36 ;
      VIA 2.58 36.18 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 36.163 2.625 36.197 ;
      VIA 2.58 36.18 Element_VIA34_1_2_58_52 ;
      VIA 2.58 36.18 Element_VIA23_1_3_36_36 ;
      VIA 2.58 35.64 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 35.623 2.625 35.657 ;
      VIA 2.58 35.64 Element_VIA34_1_2_58_52 ;
      VIA 2.58 35.64 Element_VIA23_1_3_36_36 ;
      VIA 2.58 35.1 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 35.083 2.625 35.117 ;
      VIA 2.58 35.1 Element_VIA34_1_2_58_52 ;
      VIA 2.58 35.1 Element_VIA23_1_3_36_36 ;
      VIA 2.58 34.56 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 34.543 2.625 34.577 ;
      VIA 2.58 34.56 Element_VIA34_1_2_58_52 ;
      VIA 2.58 34.56 Element_VIA23_1_3_36_36 ;
      VIA 2.58 34.02 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 34.003 2.625 34.037 ;
      VIA 2.58 34.02 Element_VIA34_1_2_58_52 ;
      VIA 2.58 34.02 Element_VIA23_1_3_36_36 ;
      VIA 2.58 33.48 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 33.463 2.625 33.497 ;
      VIA 2.58 33.48 Element_VIA34_1_2_58_52 ;
      VIA 2.58 33.48 Element_VIA23_1_3_36_36 ;
      VIA 2.58 32.94 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 32.923 2.625 32.957 ;
      VIA 2.58 32.94 Element_VIA34_1_2_58_52 ;
      VIA 2.58 32.94 Element_VIA23_1_3_36_36 ;
      VIA 2.58 32.4 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 32.383 2.625 32.417 ;
      VIA 2.58 32.4 Element_VIA34_1_2_58_52 ;
      VIA 2.58 32.4 Element_VIA23_1_3_36_36 ;
      VIA 2.58 31.86 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 31.843 2.625 31.877 ;
      VIA 2.58 31.86 Element_VIA34_1_2_58_52 ;
      VIA 2.58 31.86 Element_VIA23_1_3_36_36 ;
      VIA 2.58 31.32 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 31.303 2.625 31.337 ;
      VIA 2.58 31.32 Element_VIA34_1_2_58_52 ;
      VIA 2.58 31.32 Element_VIA23_1_3_36_36 ;
      VIA 2.58 30.78 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 30.763 2.625 30.797 ;
      VIA 2.58 30.78 Element_VIA34_1_2_58_52 ;
      VIA 2.58 30.78 Element_VIA23_1_3_36_36 ;
      VIA 2.58 30.24 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 30.223 2.625 30.257 ;
      VIA 2.58 30.24 Element_VIA34_1_2_58_52 ;
      VIA 2.58 30.24 Element_VIA23_1_3_36_36 ;
      VIA 2.58 29.7 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 29.683 2.625 29.717 ;
      VIA 2.58 29.7 Element_VIA34_1_2_58_52 ;
      VIA 2.58 29.7 Element_VIA23_1_3_36_36 ;
      VIA 2.58 29.16 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 29.143 2.625 29.177 ;
      VIA 2.58 29.16 Element_VIA34_1_2_58_52 ;
      VIA 2.58 29.16 Element_VIA23_1_3_36_36 ;
      VIA 2.58 28.62 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 28.603 2.625 28.637 ;
      VIA 2.58 28.62 Element_VIA34_1_2_58_52 ;
      VIA 2.58 28.62 Element_VIA23_1_3_36_36 ;
      VIA 2.58 28.08 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 28.063 2.625 28.097 ;
      VIA 2.58 28.08 Element_VIA34_1_2_58_52 ;
      VIA 2.58 28.08 Element_VIA23_1_3_36_36 ;
      VIA 2.58 27.54 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 27.523 2.625 27.557 ;
      VIA 2.58 27.54 Element_VIA34_1_2_58_52 ;
      VIA 2.58 27.54 Element_VIA23_1_3_36_36 ;
      VIA 2.58 27 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 26.983 2.625 27.017 ;
      VIA 2.58 27 Element_VIA34_1_2_58_52 ;
      VIA 2.58 27 Element_VIA23_1_3_36_36 ;
      VIA 2.58 26.46 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 26.443 2.625 26.477 ;
      VIA 2.58 26.46 Element_VIA34_1_2_58_52 ;
      VIA 2.58 26.46 Element_VIA23_1_3_36_36 ;
      VIA 2.58 25.92 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 25.903 2.625 25.937 ;
      VIA 2.58 25.92 Element_VIA34_1_2_58_52 ;
      VIA 2.58 25.92 Element_VIA23_1_3_36_36 ;
      VIA 2.58 25.38 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 25.363 2.625 25.397 ;
      VIA 2.58 25.38 Element_VIA34_1_2_58_52 ;
      VIA 2.58 25.38 Element_VIA23_1_3_36_36 ;
      VIA 2.58 24.84 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 24.823 2.625 24.857 ;
      VIA 2.58 24.84 Element_VIA34_1_2_58_52 ;
      VIA 2.58 24.84 Element_VIA23_1_3_36_36 ;
      VIA 2.58 24.3 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 24.283 2.625 24.317 ;
      VIA 2.58 24.3 Element_VIA34_1_2_58_52 ;
      VIA 2.58 24.3 Element_VIA23_1_3_36_36 ;
      VIA 2.58 23.76 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 23.743 2.625 23.777 ;
      VIA 2.58 23.76 Element_VIA34_1_2_58_52 ;
      VIA 2.58 23.76 Element_VIA23_1_3_36_36 ;
      VIA 2.58 23.22 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 23.203 2.625 23.237 ;
      VIA 2.58 23.22 Element_VIA34_1_2_58_52 ;
      VIA 2.58 23.22 Element_VIA23_1_3_36_36 ;
      VIA 2.58 22.68 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 22.663 2.625 22.697 ;
      VIA 2.58 22.68 Element_VIA34_1_2_58_52 ;
      VIA 2.58 22.68 Element_VIA23_1_3_36_36 ;
      VIA 2.58 22.14 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 22.123 2.625 22.157 ;
      VIA 2.58 22.14 Element_VIA34_1_2_58_52 ;
      VIA 2.58 22.14 Element_VIA23_1_3_36_36 ;
      VIA 2.58 21.6 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 21.583 2.625 21.617 ;
      VIA 2.58 21.6 Element_VIA34_1_2_58_52 ;
      VIA 2.58 21.6 Element_VIA23_1_3_36_36 ;
      VIA 2.58 21.06 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 21.043 2.625 21.077 ;
      VIA 2.58 21.06 Element_VIA34_1_2_58_52 ;
      VIA 2.58 21.06 Element_VIA23_1_3_36_36 ;
      VIA 2.58 20.52 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 20.503 2.625 20.537 ;
      VIA 2.58 20.52 Element_VIA34_1_2_58_52 ;
      VIA 2.58 20.52 Element_VIA23_1_3_36_36 ;
      VIA 2.58 19.98 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 19.963 2.625 19.997 ;
      VIA 2.58 19.98 Element_VIA34_1_2_58_52 ;
      VIA 2.58 19.98 Element_VIA23_1_3_36_36 ;
      VIA 2.58 19.44 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 19.423 2.625 19.457 ;
      VIA 2.58 19.44 Element_VIA34_1_2_58_52 ;
      VIA 2.58 19.44 Element_VIA23_1_3_36_36 ;
      VIA 2.58 18.9 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 18.883 2.625 18.917 ;
      VIA 2.58 18.9 Element_VIA34_1_2_58_52 ;
      VIA 2.58 18.9 Element_VIA23_1_3_36_36 ;
      VIA 2.58 18.36 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 18.343 2.625 18.377 ;
      VIA 2.58 18.36 Element_VIA34_1_2_58_52 ;
      VIA 2.58 18.36 Element_VIA23_1_3_36_36 ;
      VIA 2.58 17.82 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 17.803 2.625 17.837 ;
      VIA 2.58 17.82 Element_VIA34_1_2_58_52 ;
      VIA 2.58 17.82 Element_VIA23_1_3_36_36 ;
      VIA 2.58 17.28 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 17.263 2.625 17.297 ;
      VIA 2.58 17.28 Element_VIA34_1_2_58_52 ;
      VIA 2.58 17.28 Element_VIA23_1_3_36_36 ;
      VIA 2.58 16.74 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 16.723 2.625 16.757 ;
      VIA 2.58 16.74 Element_VIA34_1_2_58_52 ;
      VIA 2.58 16.74 Element_VIA23_1_3_36_36 ;
      VIA 2.58 16.2 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 16.183 2.625 16.217 ;
      VIA 2.58 16.2 Element_VIA34_1_2_58_52 ;
      VIA 2.58 16.2 Element_VIA23_1_3_36_36 ;
      VIA 2.58 15.66 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 15.643 2.625 15.677 ;
      VIA 2.58 15.66 Element_VIA34_1_2_58_52 ;
      VIA 2.58 15.66 Element_VIA23_1_3_36_36 ;
      VIA 2.58 15.12 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 15.103 2.625 15.137 ;
      VIA 2.58 15.12 Element_VIA34_1_2_58_52 ;
      VIA 2.58 15.12 Element_VIA23_1_3_36_36 ;
      VIA 2.58 14.58 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 14.563 2.625 14.597 ;
      VIA 2.58 14.58 Element_VIA34_1_2_58_52 ;
      VIA 2.58 14.58 Element_VIA23_1_3_36_36 ;
      VIA 2.58 14.04 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 14.023 2.625 14.057 ;
      VIA 2.58 14.04 Element_VIA34_1_2_58_52 ;
      VIA 2.58 14.04 Element_VIA23_1_3_36_36 ;
      VIA 2.58 13.5 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 13.483 2.625 13.517 ;
      VIA 2.58 13.5 Element_VIA34_1_2_58_52 ;
      VIA 2.58 13.5 Element_VIA23_1_3_36_36 ;
      VIA 2.58 12.96 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 12.943 2.625 12.977 ;
      VIA 2.58 12.96 Element_VIA34_1_2_58_52 ;
      VIA 2.58 12.96 Element_VIA23_1_3_36_36 ;
      VIA 2.58 12.42 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 12.403 2.625 12.437 ;
      VIA 2.58 12.42 Element_VIA34_1_2_58_52 ;
      VIA 2.58 12.42 Element_VIA23_1_3_36_36 ;
      VIA 2.58 11.88 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 11.863 2.625 11.897 ;
      VIA 2.58 11.88 Element_VIA34_1_2_58_52 ;
      VIA 2.58 11.88 Element_VIA23_1_3_36_36 ;
      VIA 2.58 11.34 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 11.323 2.625 11.357 ;
      VIA 2.58 11.34 Element_VIA34_1_2_58_52 ;
      VIA 2.58 11.34 Element_VIA23_1_3_36_36 ;
      VIA 2.58 10.8 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 10.783 2.625 10.817 ;
      VIA 2.58 10.8 Element_VIA34_1_2_58_52 ;
      VIA 2.58 10.8 Element_VIA23_1_3_36_36 ;
      VIA 2.58 10.26 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 10.243 2.625 10.277 ;
      VIA 2.58 10.26 Element_VIA34_1_2_58_52 ;
      VIA 2.58 10.26 Element_VIA23_1_3_36_36 ;
      VIA 2.58 9.72 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 9.703 2.625 9.737 ;
      VIA 2.58 9.72 Element_VIA34_1_2_58_52 ;
      VIA 2.58 9.72 Element_VIA23_1_3_36_36 ;
      VIA 2.58 9.18 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 9.163 2.625 9.197 ;
      VIA 2.58 9.18 Element_VIA34_1_2_58_52 ;
      VIA 2.58 9.18 Element_VIA23_1_3_36_36 ;
      VIA 2.58 8.64 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 8.623 2.625 8.657 ;
      VIA 2.58 8.64 Element_VIA34_1_2_58_52 ;
      VIA 2.58 8.64 Element_VIA23_1_3_36_36 ;
      VIA 2.58 8.1 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 8.083 2.625 8.117 ;
      VIA 2.58 8.1 Element_VIA34_1_2_58_52 ;
      VIA 2.58 8.1 Element_VIA23_1_3_36_36 ;
      VIA 2.58 7.56 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 7.543 2.625 7.577 ;
      VIA 2.58 7.56 Element_VIA34_1_2_58_52 ;
      VIA 2.58 7.56 Element_VIA23_1_3_36_36 ;
      VIA 2.58 7.02 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 7.003 2.625 7.037 ;
      VIA 2.58 7.02 Element_VIA34_1_2_58_52 ;
      VIA 2.58 7.02 Element_VIA23_1_3_36_36 ;
      VIA 2.58 6.48 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 6.463 2.625 6.497 ;
      VIA 2.58 6.48 Element_VIA34_1_2_58_52 ;
      VIA 2.58 6.48 Element_VIA23_1_3_36_36 ;
      VIA 2.58 5.94 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 5.923 2.625 5.957 ;
      VIA 2.58 5.94 Element_VIA34_1_2_58_52 ;
      VIA 2.58 5.94 Element_VIA23_1_3_36_36 ;
      VIA 2.58 5.4 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 5.383 2.625 5.417 ;
      VIA 2.58 5.4 Element_VIA34_1_2_58_52 ;
      VIA 2.58 5.4 Element_VIA23_1_3_36_36 ;
      VIA 2.58 4.86 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 4.843 2.625 4.877 ;
      VIA 2.58 4.86 Element_VIA34_1_2_58_52 ;
      VIA 2.58 4.86 Element_VIA23_1_3_36_36 ;
      VIA 2.58 4.32 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 4.303 2.625 4.337 ;
      VIA 2.58 4.32 Element_VIA34_1_2_58_52 ;
      VIA 2.58 4.32 Element_VIA23_1_3_36_36 ;
      VIA 2.58 3.78 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 3.763 2.625 3.797 ;
      VIA 2.58 3.78 Element_VIA34_1_2_58_52 ;
      VIA 2.58 3.78 Element_VIA23_1_3_36_36 ;
      VIA 2.58 3.24 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 3.223 2.625 3.257 ;
      VIA 2.58 3.24 Element_VIA34_1_2_58_52 ;
      VIA 2.58 3.24 Element_VIA23_1_3_36_36 ;
      VIA 2.58 2.7 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 2.683 2.625 2.717 ;
      VIA 2.58 2.7 Element_VIA34_1_2_58_52 ;
      VIA 2.58 2.7 Element_VIA23_1_3_36_36 ;
      VIA 2.58 2.16 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 2.143 2.625 2.177 ;
      VIA 2.58 2.16 Element_VIA34_1_2_58_52 ;
      VIA 2.58 2.16 Element_VIA23_1_3_36_36 ;
      VIA 2.58 1.62 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 1.603 2.625 1.637 ;
      VIA 2.58 1.62 Element_VIA34_1_2_58_52 ;
      VIA 2.58 1.62 Element_VIA23_1_3_36_36 ;
      VIA 2.58 1.08 Element_VIA45_1_2_58_58 ;
      LAYER M3 ;
        RECT  2.535 1.063 2.625 1.097 ;
      VIA 2.58 1.08 Element_VIA34_1_2_58_52 ;
      VIA 2.58 1.08 Element_VIA23_1_3_36_36 ;
      VIA 21.6 42.12 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 41.58 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 41.04 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 40.5 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 39.96 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 39.42 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 38.88 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 38.34 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 37.8 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 37.26 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 36.72 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 36.18 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 35.64 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 35.1 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 34.56 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 34.02 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 33.48 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 32.94 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 32.4 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 31.86 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 31.32 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 30.78 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 30.24 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 29.7 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 29.16 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 28.62 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 28.08 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 27.54 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 27 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 26.46 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 25.92 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 25.38 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 24.84 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 24.3 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 23.76 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 23.22 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 22.68 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 22.14 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 21.6 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 21.06 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 20.52 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 19.98 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 19.44 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 18.9 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 18.36 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 17.82 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 17.28 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 16.74 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 16.2 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 15.66 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 15.12 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 14.58 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 14.04 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 13.5 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 12.96 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 12.42 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 11.88 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 11.34 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 10.8 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 10.26 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 9.72 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 9.18 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 8.64 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 8.1 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 7.56 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 7.02 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 6.48 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 5.94 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 5.4 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 4.86 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 4.32 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 3.78 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 3.24 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 2.7 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 2.16 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 1.62 Element_via1_2_41040_18_1_1140_36_36 ;
      VIA 21.6 1.08 Element_via1_2_41040_18_1_1140_36_36 ;
    END
  END VSS
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  25.272 43.163 25.29 43.2 ;
    END
  END clock
  PIN io_ins_down[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  24.48 43.116 24.504 43.2 ;
    END
  END io_ins_down[0]
  PIN io_ins_down[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  21.672 43.163 21.69 43.2 ;
    END
  END io_ins_down[10]
  PIN io_ins_down[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  21.24 43.163 21.258 43.2 ;
    END
  END io_ins_down[11]
  PIN io_ins_down[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  20.256 43.116 20.28 43.2 ;
    END
  END io_ins_down[12]
  PIN io_ins_down[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  19.224 43.163 19.242 43.2 ;
    END
  END io_ins_down[13]
  PIN io_ins_down[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  20.088 43.163 20.106 43.2 ;
    END
  END io_ins_down[14]
  PIN io_ins_down[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  18.936 43.163 18.954 43.2 ;
    END
  END io_ins_down[15]
  PIN io_ins_down[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.12 43.116 9.144 43.2 ;
    END
  END io_ins_down[16]
  PIN io_ins_down[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  7.56 43.163 7.578 43.2 ;
    END
  END io_ins_down[17]
  PIN io_ins_down[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.064 43.116 8.088 43.2 ;
    END
  END io_ins_down[18]
  PIN io_ins_down[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  9.144 43.163 9.162 43.2 ;
    END
  END io_ins_down[19]
  PIN io_ins_down[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  21.024 43.163 21.042 43.2 ;
    END
  END io_ins_down[1]
  PIN io_ins_down[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  9.72 43.163 9.738 43.2 ;
    END
  END io_ins_down[20]
  PIN io_ins_down[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.752 43.116 10.776 43.2 ;
    END
  END io_ins_down[21]
  PIN io_ins_down[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  8.928 43.163 8.946 43.2 ;
    END
  END io_ins_down[22]
  PIN io_ins_down[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  8.352 43.163 8.37 43.2 ;
    END
  END io_ins_down[23]
  PIN io_ins_down[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  9 43.163 9.018 43.2 ;
    END
  END io_ins_down[24]
  PIN io_ins_down[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  10.296 43.163 10.314 43.2 ;
    END
  END io_ins_down[25]
  PIN io_ins_down[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.448 43.116 8.472 43.2 ;
    END
  END io_ins_down[26]
  PIN io_ins_down[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  7.776 43.163 7.794 43.2 ;
    END
  END io_ins_down[27]
  PIN io_ins_down[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.56 43.116 10.584 43.2 ;
    END
  END io_ins_down[28]
  PIN io_ins_down[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.736 43.116 8.76 43.2 ;
    END
  END io_ins_down[29]
  PIN io_ins_down[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.848 43.116 22.872 43.2 ;
    END
  END io_ins_down[2]
  PIN io_ins_down[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  10.656 43.163 10.674 43.2 ;
    END
  END io_ins_down[30]
  PIN io_ins_down[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  11.016 43.163 11.034 43.2 ;
    END
  END io_ins_down[31]
  PIN io_ins_down[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  9.36 43.163 9.378 43.2 ;
    END
  END io_ins_down[32]
  PIN io_ins_down[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  8.496 43.163 8.514 43.2 ;
    END
  END io_ins_down[33]
  PIN io_ins_down[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  10.8 43.163 10.818 43.2 ;
    END
  END io_ins_down[34]
  PIN io_ins_down[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  8.568 43.163 8.586 43.2 ;
    END
  END io_ins_down[35]
  PIN io_ins_down[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.944 43.116 10.968 43.2 ;
    END
  END io_ins_down[36]
  PIN io_ins_down[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  10.224 43.163 10.242 43.2 ;
    END
  END io_ins_down[37]
  PIN io_ins_down[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  9.216 43.163 9.234 43.2 ;
    END
  END io_ins_down[38]
  PIN io_ins_down[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  8.424 43.163 8.442 43.2 ;
    END
  END io_ins_down[39]
  PIN io_ins_down[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.696 43.116 21.72 43.2 ;
    END
  END io_ins_down[3]
  PIN io_ins_down[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  11.232 43.163 11.25 43.2 ;
    END
  END io_ins_down[40]
  PIN io_ins_down[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  9.288 43.163 9.306 43.2 ;
    END
  END io_ins_down[41]
  PIN io_ins_down[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  10.584 43.163 10.602 43.2 ;
    END
  END io_ins_down[42]
  PIN io_ins_down[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  10.152 43.163 10.17 43.2 ;
    END
  END io_ins_down[43]
  PIN io_ins_down[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  7.392 43.116 7.416 43.2 ;
    END
  END io_ins_down[44]
  PIN io_ins_down[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  9.792 43.163 9.81 43.2 ;
    END
  END io_ins_down[45]
  PIN io_ins_down[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.848 43.116 10.872 43.2 ;
    END
  END io_ins_down[46]
  PIN io_ins_down[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.176 43.116 10.2 43.2 ;
    END
  END io_ins_down[47]
  PIN io_ins_down[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  11.304 43.163 11.322 43.2 ;
    END
  END io_ins_down[48]
  PIN io_ins_down[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  9.504 43.163 9.522 43.2 ;
    END
  END io_ins_down[49]
  PIN io_ins_down[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.12 43.116 21.144 43.2 ;
    END
  END io_ins_down[4]
  PIN io_ins_down[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  10.368 43.163 10.386 43.2 ;
    END
  END io_ins_down[50]
  PIN io_ins_down[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  10.08 43.163 10.098 43.2 ;
    END
  END io_ins_down[51]
  PIN io_ins_down[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.16 43.116 8.184 43.2 ;
    END
  END io_ins_down[52]
  PIN io_ins_down[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.544 43.116 8.568 43.2 ;
    END
  END io_ins_down[53]
  PIN io_ins_down[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  8.64 43.163 8.658 43.2 ;
    END
  END io_ins_down[54]
  PIN io_ins_down[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  9.648 43.163 9.666 43.2 ;
    END
  END io_ins_down[55]
  PIN io_ins_down[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  7.416 43.163 7.434 43.2 ;
    END
  END io_ins_down[56]
  PIN io_ins_down[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.696 43.116 9.72 43.2 ;
    END
  END io_ins_down[57]
  PIN io_ins_down[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  9.072 43.163 9.09 43.2 ;
    END
  END io_ins_down[58]
  PIN io_ins_down[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  9.576 43.163 9.594 43.2 ;
    END
  END io_ins_down[59]
  PIN io_ins_down[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.52 43.116 23.544 43.2 ;
    END
  END io_ins_down[5]
  PIN io_ins_down[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  7.992 43.163 8.01 43.2 ;
    END
  END io_ins_down[60]
  PIN io_ins_down[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.6 43.116 9.624 43.2 ;
    END
  END io_ins_down[61]
  PIN io_ins_down[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.08 43.116 10.104 43.2 ;
    END
  END io_ins_down[62]
  PIN io_ins_down[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.888 43.116 9.912 43.2 ;
    END
  END io_ins_down[63]
  PIN io_ins_down[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  23.832 43.163 23.85 43.2 ;
    END
  END io_ins_down[6]
  PIN io_ins_down[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.752 43.116 22.776 43.2 ;
    END
  END io_ins_down[7]
  PIN io_ins_down[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.984 43.116 22.008 43.2 ;
    END
  END io_ins_down[8]
  PIN io_ins_down[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  21.888 43.163 21.906 43.2 ;
    END
  END io_ins_down[9]
  PIN io_ins_left[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 13.221 43.2 13.239 ;
    END
  END io_ins_left[0]
  PIN io_ins_left[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 16.308 43.2 16.326 ;
    END
  END io_ins_left[10]
  PIN io_ins_left[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 16.38 43.2 16.398 ;
    END
  END io_ins_left[11]
  PIN io_ins_left[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 18.504 43.2 18.522 ;
    END
  END io_ins_left[12]
  PIN io_ins_left[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 16.224 43.2 16.248 ;
    END
  END io_ins_left[13]
  PIN io_ins_left[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 19.776 43.2 19.8 ;
    END
  END io_ins_left[14]
  PIN io_ins_left[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 18.936 43.2 18.954 ;
    END
  END io_ins_left[15]
  PIN io_ins_left[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 11.448 43.2 11.466 ;
    END
  END io_ins_left[16]
  PIN io_ins_left[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 10.656 43.2 10.68 ;
    END
  END io_ins_left[17]
  PIN io_ins_left[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 29.844 43.2 29.862 ;
    END
  END io_ins_left[18]
  PIN io_ins_left[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 12.096 43.2 12.12 ;
    END
  END io_ins_left[19]
  PIN io_ins_left[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 12.288 43.2 12.312 ;
    END
  END io_ins_left[1]
  PIN io_ins_left[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 17.001 43.2 17.019 ;
    END
  END io_ins_left[20]
  PIN io_ins_left[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 25.056 43.2 25.08 ;
    END
  END io_ins_left[21]
  PIN io_ins_left[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 26.4 43.2 26.424 ;
    END
  END io_ins_left[22]
  PIN io_ins_left[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 20.352 43.2 20.376 ;
    END
  END io_ins_left[23]
  PIN io_ins_left[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 29.76 43.2 29.784 ;
    END
  END io_ins_left[24]
  PIN io_ins_left[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 18.54 43.2 18.558 ;
    END
  END io_ins_left[25]
  PIN io_ins_left[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 23.616 43.2 23.64 ;
    END
  END io_ins_left[26]
  PIN io_ins_left[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 11.412 43.2 11.43 ;
    END
  END io_ins_left[27]
  PIN io_ins_left[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 22.716 43.2 22.734 ;
    END
  END io_ins_left[28]
  PIN io_ins_left[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 11.424 43.2 11.448 ;
    END
  END io_ins_left[29]
  PIN io_ins_left[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 15.228 43.2 15.246 ;
    END
  END io_ins_left[2]
  PIN io_ins_left[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 29.568 43.2 29.592 ;
    END
  END io_ins_left[30]
  PIN io_ins_left[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 13.248 43.2 13.272 ;
    END
  END io_ins_left[31]
  PIN io_ins_left[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 21.321 43.2 21.339 ;
    END
  END io_ins_left[32]
  PIN io_ins_left[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 29.961 43.2 29.979 ;
    END
  END io_ins_left[33]
  PIN io_ins_left[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 13.92 43.2 13.944 ;
    END
  END io_ins_left[34]
  PIN io_ins_left[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 26.181 43.2 26.199 ;
    END
  END io_ins_left[35]
  PIN io_ins_left[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 26.304 43.2 26.328 ;
    END
  END io_ins_left[36]
  PIN io_ins_left[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 21.984 43.2 22.008 ;
    END
  END io_ins_left[37]
  PIN io_ins_left[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 18.912 43.2 18.936 ;
    END
  END io_ins_left[38]
  PIN io_ins_left[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 10.944 43.2 10.962 ;
    END
  END io_ins_left[39]
  PIN io_ins_left[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 13.608 43.2 13.626 ;
    END
  END io_ins_left[3]
  PIN io_ins_left[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 12.192 43.2 12.216 ;
    END
  END io_ins_left[40]
  PIN io_ins_left[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 22.788 43.2 22.806 ;
    END
  END io_ins_left[41]
  PIN io_ins_left[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 10.836 43.2 10.854 ;
    END
  END io_ins_left[42]
  PIN io_ins_left[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 22.752 43.2 22.77 ;
    END
  END io_ins_left[43]
  PIN io_ins_left[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 12.024 43.2 12.042 ;
    END
  END io_ins_left[44]
  PIN io_ins_left[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 26.208 43.2 26.232 ;
    END
  END io_ins_left[45]
  PIN io_ins_left[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 26.532 43.2 26.55 ;
    END
  END io_ins_left[46]
  PIN io_ins_left[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 16.032 43.2 16.056 ;
    END
  END io_ins_left[47]
  PIN io_ins_left[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 28.8 43.2 28.818 ;
    END
  END io_ins_left[48]
  PIN io_ins_left[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 18.624 43.2 18.648 ;
    END
  END io_ins_left[49]
  PIN io_ins_left[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 17.184 43.2 17.208 ;
    END
  END io_ins_left[4]
  PIN io_ins_left[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 24.021 43.2 24.039 ;
    END
  END io_ins_left[50]
  PIN io_ins_left[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 15.921 43.2 15.939 ;
    END
  END io_ins_left[51]
  PIN io_ins_left[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 14.148 43.2 14.166 ;
    END
  END io_ins_left[52]
  PIN io_ins_left[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 11.712 43.2 11.736 ;
    END
  END io_ins_left[53]
  PIN io_ins_left[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 15.456 43.2 15.48 ;
    END
  END io_ins_left[54]
  PIN io_ins_left[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 26.88 43.2 26.904 ;
    END
  END io_ins_left[55]
  PIN io_ins_left[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 26.064 43.2 26.082 ;
    END
  END io_ins_left[56]
  PIN io_ins_left[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 11.376 43.2 11.394 ;
    END
  END io_ins_left[57]
  PIN io_ins_left[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 27.84 43.2 27.864 ;
    END
  END io_ins_left[58]
  PIN io_ins_left[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 10.908 43.2 10.926 ;
    END
  END io_ins_left[59]
  PIN io_ins_left[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 14.301 43.2 14.319 ;
    END
  END io_ins_left[5]
  PIN io_ins_left[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 12.96 43.2 12.984 ;
    END
  END io_ins_left[60]
  PIN io_ins_left[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 10.752 43.2 10.776 ;
    END
  END io_ins_left[61]
  PIN io_ins_left[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 18.816 43.2 18.84 ;
    END
  END io_ins_left[62]
  PIN io_ins_left[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 11.988 43.2 12.006 ;
    END
  END io_ins_left[63]
  PIN io_ins_left[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 15.732 43.2 15.75 ;
    END
  END io_ins_left[6]
  PIN io_ins_left[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 15.156 43.2 15.174 ;
    END
  END io_ins_left[7]
  PIN io_ins_left[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 17.28 43.2 17.304 ;
    END
  END io_ins_left[8]
  PIN io_ins_left[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 15.381 43.2 15.399 ;
    END
  END io_ins_left[9]
  PIN io_ins_right[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 26.028 0.037 26.046 ;
    END
  END io_ins_right[0]
  PIN io_ins_right[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 28.296 0.037 28.314 ;
    END
  END io_ins_right[10]
  PIN io_ins_right[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 31.428 0.037 31.446 ;
    END
  END io_ins_right[11]
  PIN io_ins_right[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 28.152 0.037 28.17 ;
    END
  END io_ins_right[12]
  PIN io_ins_right[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 24.48 0.084 24.504 ;
    END
  END io_ins_right[13]
  PIN io_ins_right[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 24.672 0.084 24.696 ;
    END
  END io_ins_right[14]
  PIN io_ins_right[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 24.516 0.037 24.534 ;
    END
  END io_ins_right[15]
  PIN io_ins_right[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 12.141 0.037 12.159 ;
    END
  END io_ins_right[16]
  PIN io_ins_right[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 11.484 0.037 11.502 ;
    END
  END io_ins_right[17]
  PIN io_ins_right[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 19.296 0.084 19.32 ;
    END
  END io_ins_right[18]
  PIN io_ins_right[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 11.04 0.084 11.064 ;
    END
  END io_ins_right[19]
  PIN io_ins_right[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 22.248 0.037 22.266 ;
    END
  END io_ins_right[1]
  PIN io_ins_right[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 25.02 0.037 25.038 ;
    END
  END io_ins_right[20]
  PIN io_ins_right[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 12.636 0.037 12.654 ;
    END
  END io_ins_right[21]
  PIN io_ins_right[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 14.076 0.037 14.094 ;
    END
  END io_ins_right[22]
  PIN io_ins_right[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 14.112 0.037 14.13 ;
    END
  END io_ins_right[23]
  PIN io_ins_right[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 21.504 0.084 21.528 ;
    END
  END io_ins_right[24]
  PIN io_ins_right[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 17.664 0.084 17.688 ;
    END
  END io_ins_right[25]
  PIN io_ins_right[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 23.136 0.084 23.16 ;
    END
  END io_ins_right[26]
  PIN io_ins_right[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 24.864 0.084 24.888 ;
    END
  END io_ins_right[27]
  PIN io_ins_right[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 11.061 0.037 11.079 ;
    END
  END io_ins_right[28]
  PIN io_ins_right[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 19.968 0.084 19.992 ;
    END
  END io_ins_right[29]
  PIN io_ins_right[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 24.192 0.084 24.216 ;
    END
  END io_ins_right[2]
  PIN io_ins_right[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 10.872 0.037 10.89 ;
    END
  END io_ins_right[30]
  PIN io_ins_right[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 11.016 0.037 11.034 ;
    END
  END io_ins_right[31]
  PIN io_ins_right[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 29.952 0.084 29.976 ;
    END
  END io_ins_right[32]
  PIN io_ins_right[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 27.612 0.037 27.63 ;
    END
  END io_ins_right[33]
  PIN io_ins_right[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 10.848 0.084 10.872 ;
    END
  END io_ins_right[34]
  PIN io_ins_right[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 28.032 0.084 28.056 ;
    END
  END io_ins_right[35]
  PIN io_ins_right[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 20.016 0.037 20.034 ;
    END
  END io_ins_right[36]
  PIN io_ins_right[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 18.144 0.084 18.168 ;
    END
  END io_ins_right[37]
  PIN io_ins_right[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 13.68 0.037 13.698 ;
    END
  END io_ins_right[38]
  PIN io_ins_right[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 17.76 0.084 17.784 ;
    END
  END io_ins_right[39]
  PIN io_ins_right[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 25.488 0.037 25.506 ;
    END
  END io_ins_right[3]
  PIN io_ins_right[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 21.408 0.084 21.432 ;
    END
  END io_ins_right[40]
  PIN io_ins_right[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 23.436 0.037 23.454 ;
    END
  END io_ins_right[41]
  PIN io_ins_right[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 11.328 0.084 11.352 ;
    END
  END io_ins_right[42]
  PIN io_ins_right[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 29.664 0.084 29.688 ;
    END
  END io_ins_right[43]
  PIN io_ins_right[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 23.52 0.084 23.544 ;
    END
  END io_ins_right[44]
  PIN io_ins_right[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 27.108 0.037 27.126 ;
    END
  END io_ins_right[45]
  PIN io_ins_right[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 23.481 0.037 23.499 ;
    END
  END io_ins_right[46]
  PIN io_ins_right[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 15.936 0.084 15.96 ;
    END
  END io_ins_right[47]
  PIN io_ins_right[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 29.808 0.037 29.826 ;
    END
  END io_ins_right[48]
  PIN io_ins_right[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 15.876 0.037 15.894 ;
    END
  END io_ins_right[49]
  PIN io_ins_right[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 32.352 0.084 32.376 ;
    END
  END io_ins_right[4]
  PIN io_ins_right[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 10.944 0.084 10.968 ;
    END
  END io_ins_right[50]
  PIN io_ins_right[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 14.652 0.037 14.67 ;
    END
  END io_ins_right[51]
  PIN io_ins_right[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 15.552 0.084 15.576 ;
    END
  END io_ins_right[52]
  PIN io_ins_right[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 11.952 0.037 11.97 ;
    END
  END io_ins_right[53]
  PIN io_ins_right[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 11.136 0.084 11.16 ;
    END
  END io_ins_right[54]
  PIN io_ins_right[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 11.808 0.084 11.832 ;
    END
  END io_ins_right[55]
  PIN io_ins_right[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 18.048 0.084 18.072 ;
    END
  END io_ins_right[56]
  PIN io_ins_right[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 20.928 0.084 20.952 ;
    END
  END io_ins_right[57]
  PIN io_ins_right[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 11.232 0.084 11.256 ;
    END
  END io_ins_right[58]
  PIN io_ins_right[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 10.98 0.037 10.998 ;
    END
  END io_ins_right[59]
  PIN io_ins_right[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 25.92 0.084 25.944 ;
    END
  END io_ins_right[5]
  PIN io_ins_right[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 14.976 0.084 15 ;
    END
  END io_ins_right[60]
  PIN io_ins_right[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 30.144 0.084 30.168 ;
    END
  END io_ins_right[61]
  PIN io_ins_right[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 14.112 0.084 14.136 ;
    END
  END io_ins_right[62]
  PIN io_ins_right[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 29.916 0.037 29.934 ;
    END
  END io_ins_right[63]
  PIN io_ins_right[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 30.42 0.037 30.438 ;
    END
  END io_ins_right[6]
  PIN io_ins_right[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 30.348 0.037 30.366 ;
    END
  END io_ins_right[7]
  PIN io_ins_right[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 32.448 0.084 32.472 ;
    END
  END io_ins_right[8]
  PIN io_ins_right[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 33.084 0.037 33.102 ;
    END
  END io_ins_right[9]
  PIN io_ins_up[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  30.528 0 30.546 0.037 ;
    END
  END io_ins_up[0]
  PIN io_ins_up[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.264 0 15.288 0.084 ;
    END
  END io_ins_up[10]
  PIN io_ins_up[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  26.4 0 26.424 0.084 ;
    END
  END io_ins_up[11]
  PIN io_ins_up[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  15.768 0 15.786 0.037 ;
    END
  END io_ins_up[12]
  PIN io_ins_up[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.176 0 22.2 0.084 ;
    END
  END io_ins_up[13]
  PIN io_ins_up[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.36 0 15.384 0.084 ;
    END
  END io_ins_up[14]
  PIN io_ins_up[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  26.064 0 26.082 0.037 ;
    END
  END io_ins_up[15]
  PIN io_ins_up[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  10.872 0 10.89 0.037 ;
    END
  END io_ins_up[16]
  PIN io_ins_up[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.272 0 10.296 0.084 ;
    END
  END io_ins_up[17]
  PIN io_ins_up[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.464 0 10.488 0.084 ;
    END
  END io_ins_up[18]
  PIN io_ins_up[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  8.712 0 8.73 0.037 ;
    END
  END io_ins_up[19]
  PIN io_ins_up[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  20.352 0 20.376 0.084 ;
    END
  END io_ins_up[1]
  PIN io_ins_up[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.64 0 8.664 0.084 ;
    END
  END io_ins_up[20]
  PIN io_ins_up[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.216 0 9.24 0.084 ;
    END
  END io_ins_up[21]
  PIN io_ins_up[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  9.936 0 9.954 0.037 ;
    END
  END io_ins_up[22]
  PIN io_ins_up[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.256 0 8.28 0.084 ;
    END
  END io_ins_up[23]
  PIN io_ins_up[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.408 0 9.432 0.084 ;
    END
  END io_ins_up[24]
  PIN io_ins_up[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  7.848 0 7.866 0.037 ;
    END
  END io_ins_up[25]
  PIN io_ins_up[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  7.92 0 7.938 0.037 ;
    END
  END io_ins_up[26]
  PIN io_ins_up[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  8.208 0 8.226 0.037 ;
    END
  END io_ins_up[27]
  PIN io_ins_up[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  10.44 0 10.458 0.037 ;
    END
  END io_ins_up[28]
  PIN io_ins_up[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  7.872 0 7.896 0.084 ;
    END
  END io_ins_up[29]
  PIN io_ins_up[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  20.736 0 20.754 0.037 ;
    END
  END io_ins_up[2]
  PIN io_ins_up[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.928 0 8.952 0.084 ;
    END
  END io_ins_up[30]
  PIN io_ins_up[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.368 0 10.392 0.084 ;
    END
  END io_ins_up[31]
  PIN io_ins_up[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  11.04 0 11.064 0.084 ;
    END
  END io_ins_up[32]
  PIN io_ins_up[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.504 0 9.528 0.084 ;
    END
  END io_ins_up[33]
  PIN io_ins_up[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.312 0 9.336 0.084 ;
    END
  END io_ins_up[34]
  PIN io_ins_up[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  8.784 0 8.802 0.037 ;
    END
  END io_ins_up[35]
  PIN io_ins_up[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.024 0 9.048 0.084 ;
    END
  END io_ins_up[36]
  PIN io_ins_up[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  11.088 0 11.106 0.037 ;
    END
  END io_ins_up[37]
  PIN io_ins_up[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  9.432 0 9.45 0.037 ;
    END
  END io_ins_up[38]
  PIN io_ins_up[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  7.632 0 7.65 0.037 ;
    END
  END io_ins_up[39]
  PIN io_ins_up[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  20.808 0 20.826 0.037 ;
    END
  END io_ins_up[3]
  PIN io_ins_up[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  8.136 0 8.154 0.037 ;
    END
  END io_ins_up[40]
  PIN io_ins_up[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  7.68 0 7.704 0.084 ;
    END
  END io_ins_up[41]
  PIN io_ins_up[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.832 0 8.856 0.084 ;
    END
  END io_ins_up[42]
  PIN io_ins_up[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.352 0 8.376 0.084 ;
    END
  END io_ins_up[43]
  PIN io_ins_up[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  10.728 0 10.746 0.037 ;
    END
  END io_ins_up[44]
  PIN io_ins_up[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  9.864 0 9.882 0.037 ;
    END
  END io_ins_up[45]
  PIN io_ins_up[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  7.968 0 7.992 0.084 ;
    END
  END io_ins_up[46]
  PIN io_ins_up[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  10.512 0 10.53 0.037 ;
    END
  END io_ins_up[47]
  PIN io_ins_up[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  10.944 0 10.962 0.037 ;
    END
  END io_ins_up[48]
  PIN io_ins_up[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  10.008 0 10.026 0.037 ;
    END
  END io_ins_up[49]
  PIN io_ins_up[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  19.392 0 19.416 0.084 ;
    END
  END io_ins_up[4]
  PIN io_ins_up[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  8.856 0 8.874 0.037 ;
    END
  END io_ins_up[50]
  PIN io_ins_up[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  7.584 0 7.608 0.084 ;
    END
  END io_ins_up[51]
  PIN io_ins_up[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  8.28 0 8.298 0.037 ;
    END
  END io_ins_up[52]
  PIN io_ins_up[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.984 0 10.008 0.084 ;
    END
  END io_ins_up[53]
  PIN io_ins_up[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  7.776 0 7.8 0.084 ;
    END
  END io_ins_up[54]
  PIN io_ins_up[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  7.488 0 7.506 0.037 ;
    END
  END io_ins_up[55]
  PIN io_ins_up[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.792 0 9.816 0.084 ;
    END
  END io_ins_up[56]
  PIN io_ins_up[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  11.16 0 11.178 0.037 ;
    END
  END io_ins_up[57]
  PIN io_ins_up[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  8.064 0 8.082 0.037 ;
    END
  END io_ins_up[58]
  PIN io_ins_up[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  11.136 0 11.16 0.084 ;
    END
  END io_ins_up[59]
  PIN io_ins_up[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  24.672 0 24.696 0.084 ;
    END
  END io_ins_up[5]
  PIN io_ins_up[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  7.704 0 7.722 0.037 ;
    END
  END io_ins_up[60]
  PIN io_ins_up[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.656 0 10.68 0.084 ;
    END
  END io_ins_up[61]
  PIN io_ins_up[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  7.488 0 7.512 0.084 ;
    END
  END io_ins_up[62]
  PIN io_ins_up[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  11.232 0 11.256 0.084 ;
    END
  END io_ins_up[63]
  PIN io_ins_up[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  27.504 0 27.522 0.037 ;
    END
  END io_ins_up[6]
  PIN io_ins_up[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  19.104 0 19.128 0.084 ;
    END
  END io_ins_up[7]
  PIN io_ins_up[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  18.792 0 18.81 0.037 ;
    END
  END io_ins_up[8]
  PIN io_ins_up[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  19.2 0 19.224 0.084 ;
    END
  END io_ins_up[9]
  PIN io_lsbIns_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 18.72 0.084 18.744 ;
    END
  END io_lsbIns_1
  PIN io_lsbIns_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 1.728 0.084 1.752 ;
    END
  END io_lsbIns_2
  PIN io_lsbIns_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 4.392 0.037 4.41 ;
    END
  END io_lsbIns_3
  PIN io_lsbIns_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 7.164 0.037 7.182 ;
    END
  END io_lsbIns_4
  PIN io_lsbIns_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 1.632 0.084 1.656 ;
    END
  END io_lsbIns_5
  PIN io_lsbIns_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 37.728 0.084 37.752 ;
    END
  END io_lsbIns_6
  PIN io_lsbIns_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 25.524 0.037 25.542 ;
    END
  END io_lsbIns_7
  PIN io_lsbOuts_0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 40.32 43.2 40.344 ;
    END
  END io_lsbOuts_0
  PIN io_lsbOuts_1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 18.72 43.2 18.744 ;
    END
  END io_lsbOuts_1
  PIN io_lsbOuts_2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 1.728 43.2 1.752 ;
    END
  END io_lsbOuts_2
  PIN io_lsbOuts_3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 4.392 43.2 4.41 ;
    END
  END io_lsbOuts_3
  PIN io_lsbOuts_4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 7.164 43.2 7.182 ;
    END
  END io_lsbOuts_4
  PIN io_lsbOuts_5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 1.632 43.2 1.656 ;
    END
  END io_lsbOuts_5
  PIN io_lsbOuts_6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 37.728 43.2 37.752 ;
    END
  END io_lsbOuts_6
  PIN io_lsbOuts_7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 25.524 43.2 25.542 ;
    END
  END io_lsbOuts_7
  PIN io_outs_down[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  24.48 0 24.504 0.084 ;
    END
  END io_outs_down[0]
  PIN io_outs_down[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  21.672 0 21.69 0.037 ;
    END
  END io_outs_down[10]
  PIN io_outs_down[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  21.24 0 21.258 0.037 ;
    END
  END io_outs_down[11]
  PIN io_outs_down[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  20.256 0 20.28 0.084 ;
    END
  END io_outs_down[12]
  PIN io_outs_down[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  19.224 0 19.242 0.037 ;
    END
  END io_outs_down[13]
  PIN io_outs_down[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  20.088 0 20.106 0.037 ;
    END
  END io_outs_down[14]
  PIN io_outs_down[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  18.936 0 18.954 0.037 ;
    END
  END io_outs_down[15]
  PIN io_outs_down[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.12 0 9.144 0.084 ;
    END
  END io_outs_down[16]
  PIN io_outs_down[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  7.56 0 7.578 0.037 ;
    END
  END io_outs_down[17]
  PIN io_outs_down[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.064 0 8.088 0.084 ;
    END
  END io_outs_down[18]
  PIN io_outs_down[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  9.144 0 9.162 0.037 ;
    END
  END io_outs_down[19]
  PIN io_outs_down[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  21.024 0 21.042 0.037 ;
    END
  END io_outs_down[1]
  PIN io_outs_down[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  9.72 0 9.738 0.037 ;
    END
  END io_outs_down[20]
  PIN io_outs_down[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.752 0 10.776 0.084 ;
    END
  END io_outs_down[21]
  PIN io_outs_down[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  8.928 0 8.946 0.037 ;
    END
  END io_outs_down[22]
  PIN io_outs_down[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  8.352 0 8.37 0.037 ;
    END
  END io_outs_down[23]
  PIN io_outs_down[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  9 0 9.018 0.037 ;
    END
  END io_outs_down[24]
  PIN io_outs_down[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  10.296 0 10.314 0.037 ;
    END
  END io_outs_down[25]
  PIN io_outs_down[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.448 0 8.472 0.084 ;
    END
  END io_outs_down[26]
  PIN io_outs_down[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  7.776 0 7.794 0.037 ;
    END
  END io_outs_down[27]
  PIN io_outs_down[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.56 0 10.584 0.084 ;
    END
  END io_outs_down[28]
  PIN io_outs_down[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.736 0 8.76 0.084 ;
    END
  END io_outs_down[29]
  PIN io_outs_down[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.848 0 22.872 0.084 ;
    END
  END io_outs_down[2]
  PIN io_outs_down[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  10.656 0 10.674 0.037 ;
    END
  END io_outs_down[30]
  PIN io_outs_down[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  11.016 0 11.034 0.037 ;
    END
  END io_outs_down[31]
  PIN io_outs_down[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  9.36 0 9.378 0.037 ;
    END
  END io_outs_down[32]
  PIN io_outs_down[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  8.496 0 8.514 0.037 ;
    END
  END io_outs_down[33]
  PIN io_outs_down[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  10.8 0 10.818 0.037 ;
    END
  END io_outs_down[34]
  PIN io_outs_down[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  8.568 0 8.586 0.037 ;
    END
  END io_outs_down[35]
  PIN io_outs_down[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.944 0 10.968 0.084 ;
    END
  END io_outs_down[36]
  PIN io_outs_down[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  10.224 0 10.242 0.037 ;
    END
  END io_outs_down[37]
  PIN io_outs_down[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  9.216 0 9.234 0.037 ;
    END
  END io_outs_down[38]
  PIN io_outs_down[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  8.424 0 8.442 0.037 ;
    END
  END io_outs_down[39]
  PIN io_outs_down[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.696 0 21.72 0.084 ;
    END
  END io_outs_down[3]
  PIN io_outs_down[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  11.232 0 11.25 0.037 ;
    END
  END io_outs_down[40]
  PIN io_outs_down[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  9.288 0 9.306 0.037 ;
    END
  END io_outs_down[41]
  PIN io_outs_down[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  10.584 0 10.602 0.037 ;
    END
  END io_outs_down[42]
  PIN io_outs_down[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  10.152 0 10.17 0.037 ;
    END
  END io_outs_down[43]
  PIN io_outs_down[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  7.392 0 7.416 0.084 ;
    END
  END io_outs_down[44]
  PIN io_outs_down[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  9.792 0 9.81 0.037 ;
    END
  END io_outs_down[45]
  PIN io_outs_down[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.848 0 10.872 0.084 ;
    END
  END io_outs_down[46]
  PIN io_outs_down[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.176 0 10.2 0.084 ;
    END
  END io_outs_down[47]
  PIN io_outs_down[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  11.304 0 11.322 0.037 ;
    END
  END io_outs_down[48]
  PIN io_outs_down[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  9.504 0 9.522 0.037 ;
    END
  END io_outs_down[49]
  PIN io_outs_down[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.12 0 21.144 0.084 ;
    END
  END io_outs_down[4]
  PIN io_outs_down[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  10.368 0 10.386 0.037 ;
    END
  END io_outs_down[50]
  PIN io_outs_down[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  10.08 0 10.098 0.037 ;
    END
  END io_outs_down[51]
  PIN io_outs_down[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.16 0 8.184 0.084 ;
    END
  END io_outs_down[52]
  PIN io_outs_down[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.544 0 8.568 0.084 ;
    END
  END io_outs_down[53]
  PIN io_outs_down[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  8.64 0 8.658 0.037 ;
    END
  END io_outs_down[54]
  PIN io_outs_down[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  9.648 0 9.666 0.037 ;
    END
  END io_outs_down[55]
  PIN io_outs_down[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  7.416 0 7.434 0.037 ;
    END
  END io_outs_down[56]
  PIN io_outs_down[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.696 0 9.72 0.084 ;
    END
  END io_outs_down[57]
  PIN io_outs_down[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  9.072 0 9.09 0.037 ;
    END
  END io_outs_down[58]
  PIN io_outs_down[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  9.576 0 9.594 0.037 ;
    END
  END io_outs_down[59]
  PIN io_outs_down[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  23.52 0 23.544 0.084 ;
    END
  END io_outs_down[5]
  PIN io_outs_down[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  7.992 0 8.01 0.037 ;
    END
  END io_outs_down[60]
  PIN io_outs_down[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.6 0 9.624 0.084 ;
    END
  END io_outs_down[61]
  PIN io_outs_down[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.08 0 10.104 0.084 ;
    END
  END io_outs_down[62]
  PIN io_outs_down[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.888 0 9.912 0.084 ;
    END
  END io_outs_down[63]
  PIN io_outs_down[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  23.832 0 23.85 0.037 ;
    END
  END io_outs_down[6]
  PIN io_outs_down[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.752 0 22.776 0.084 ;
    END
  END io_outs_down[7]
  PIN io_outs_down[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  21.984 0 22.008 0.084 ;
    END
  END io_outs_down[8]
  PIN io_outs_down[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  21.888 0 21.906 0.037 ;
    END
  END io_outs_down[9]
  PIN io_outs_left[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 13.221 0.037 13.239 ;
    END
  END io_outs_left[0]
  PIN io_outs_left[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 16.308 0.037 16.326 ;
    END
  END io_outs_left[10]
  PIN io_outs_left[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 16.38 0.037 16.398 ;
    END
  END io_outs_left[11]
  PIN io_outs_left[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 18.504 0.037 18.522 ;
    END
  END io_outs_left[12]
  PIN io_outs_left[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 16.224 0.084 16.248 ;
    END
  END io_outs_left[13]
  PIN io_outs_left[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 19.776 0.084 19.8 ;
    END
  END io_outs_left[14]
  PIN io_outs_left[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 18.936 0.037 18.954 ;
    END
  END io_outs_left[15]
  PIN io_outs_left[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 11.448 0.037 11.466 ;
    END
  END io_outs_left[16]
  PIN io_outs_left[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 10.656 0.084 10.68 ;
    END
  END io_outs_left[17]
  PIN io_outs_left[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 29.844 0.037 29.862 ;
    END
  END io_outs_left[18]
  PIN io_outs_left[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 12.096 0.084 12.12 ;
    END
  END io_outs_left[19]
  PIN io_outs_left[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 12.288 0.084 12.312 ;
    END
  END io_outs_left[1]
  PIN io_outs_left[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 17.001 0.037 17.019 ;
    END
  END io_outs_left[20]
  PIN io_outs_left[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 25.056 0.084 25.08 ;
    END
  END io_outs_left[21]
  PIN io_outs_left[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 26.4 0.084 26.424 ;
    END
  END io_outs_left[22]
  PIN io_outs_left[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 20.352 0.084 20.376 ;
    END
  END io_outs_left[23]
  PIN io_outs_left[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 29.76 0.084 29.784 ;
    END
  END io_outs_left[24]
  PIN io_outs_left[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 18.54 0.037 18.558 ;
    END
  END io_outs_left[25]
  PIN io_outs_left[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 23.616 0.084 23.64 ;
    END
  END io_outs_left[26]
  PIN io_outs_left[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 11.412 0.037 11.43 ;
    END
  END io_outs_left[27]
  PIN io_outs_left[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 22.716 0.037 22.734 ;
    END
  END io_outs_left[28]
  PIN io_outs_left[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 11.424 0.084 11.448 ;
    END
  END io_outs_left[29]
  PIN io_outs_left[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 15.228 0.037 15.246 ;
    END
  END io_outs_left[2]
  PIN io_outs_left[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 29.568 0.084 29.592 ;
    END
  END io_outs_left[30]
  PIN io_outs_left[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 13.248 0.084 13.272 ;
    END
  END io_outs_left[31]
  PIN io_outs_left[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 21.321 0.037 21.339 ;
    END
  END io_outs_left[32]
  PIN io_outs_left[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 29.961 0.037 29.979 ;
    END
  END io_outs_left[33]
  PIN io_outs_left[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 13.92 0.084 13.944 ;
    END
  END io_outs_left[34]
  PIN io_outs_left[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 26.181 0.037 26.199 ;
    END
  END io_outs_left[35]
  PIN io_outs_left[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 26.304 0.084 26.328 ;
    END
  END io_outs_left[36]
  PIN io_outs_left[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 21.984 0.084 22.008 ;
    END
  END io_outs_left[37]
  PIN io_outs_left[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 18.912 0.084 18.936 ;
    END
  END io_outs_left[38]
  PIN io_outs_left[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 10.944 0.037 10.962 ;
    END
  END io_outs_left[39]
  PIN io_outs_left[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 13.608 0.037 13.626 ;
    END
  END io_outs_left[3]
  PIN io_outs_left[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 12.192 0.084 12.216 ;
    END
  END io_outs_left[40]
  PIN io_outs_left[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 22.788 0.037 22.806 ;
    END
  END io_outs_left[41]
  PIN io_outs_left[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 10.836 0.037 10.854 ;
    END
  END io_outs_left[42]
  PIN io_outs_left[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 22.752 0.037 22.77 ;
    END
  END io_outs_left[43]
  PIN io_outs_left[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 12.024 0.037 12.042 ;
    END
  END io_outs_left[44]
  PIN io_outs_left[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 26.208 0.084 26.232 ;
    END
  END io_outs_left[45]
  PIN io_outs_left[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 26.532 0.037 26.55 ;
    END
  END io_outs_left[46]
  PIN io_outs_left[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 16.032 0.084 16.056 ;
    END
  END io_outs_left[47]
  PIN io_outs_left[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 28.8 0.037 28.818 ;
    END
  END io_outs_left[48]
  PIN io_outs_left[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 18.624 0.084 18.648 ;
    END
  END io_outs_left[49]
  PIN io_outs_left[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 17.184 0.084 17.208 ;
    END
  END io_outs_left[4]
  PIN io_outs_left[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 24.021 0.037 24.039 ;
    END
  END io_outs_left[50]
  PIN io_outs_left[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 15.921 0.037 15.939 ;
    END
  END io_outs_left[51]
  PIN io_outs_left[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 14.148 0.037 14.166 ;
    END
  END io_outs_left[52]
  PIN io_outs_left[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 11.712 0.084 11.736 ;
    END
  END io_outs_left[53]
  PIN io_outs_left[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 15.456 0.084 15.48 ;
    END
  END io_outs_left[54]
  PIN io_outs_left[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 26.88 0.084 26.904 ;
    END
  END io_outs_left[55]
  PIN io_outs_left[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 26.064 0.037 26.082 ;
    END
  END io_outs_left[56]
  PIN io_outs_left[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 11.376 0.037 11.394 ;
    END
  END io_outs_left[57]
  PIN io_outs_left[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 27.84 0.084 27.864 ;
    END
  END io_outs_left[58]
  PIN io_outs_left[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 10.908 0.037 10.926 ;
    END
  END io_outs_left[59]
  PIN io_outs_left[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 14.301 0.037 14.319 ;
    END
  END io_outs_left[5]
  PIN io_outs_left[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 12.96 0.084 12.984 ;
    END
  END io_outs_left[60]
  PIN io_outs_left[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 10.752 0.084 10.776 ;
    END
  END io_outs_left[61]
  PIN io_outs_left[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 18.816 0.084 18.84 ;
    END
  END io_outs_left[62]
  PIN io_outs_left[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 11.988 0.037 12.006 ;
    END
  END io_outs_left[63]
  PIN io_outs_left[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 15.732 0.037 15.75 ;
    END
  END io_outs_left[6]
  PIN io_outs_left[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 15.156 0.037 15.174 ;
    END
  END io_outs_left[7]
  PIN io_outs_left[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  0 17.28 0.084 17.304 ;
    END
  END io_outs_left[8]
  PIN io_outs_left[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  0 15.381 0.037 15.399 ;
    END
  END io_outs_left[9]
  PIN io_outs_right[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 26.028 43.2 26.046 ;
    END
  END io_outs_right[0]
  PIN io_outs_right[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 28.296 43.2 28.314 ;
    END
  END io_outs_right[10]
  PIN io_outs_right[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 31.428 43.2 31.446 ;
    END
  END io_outs_right[11]
  PIN io_outs_right[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 28.152 43.2 28.17 ;
    END
  END io_outs_right[12]
  PIN io_outs_right[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 24.48 43.2 24.504 ;
    END
  END io_outs_right[13]
  PIN io_outs_right[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 24.672 43.2 24.696 ;
    END
  END io_outs_right[14]
  PIN io_outs_right[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 24.516 43.2 24.534 ;
    END
  END io_outs_right[15]
  PIN io_outs_right[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 12.141 43.2 12.159 ;
    END
  END io_outs_right[16]
  PIN io_outs_right[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 11.484 43.2 11.502 ;
    END
  END io_outs_right[17]
  PIN io_outs_right[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 19.296 43.2 19.32 ;
    END
  END io_outs_right[18]
  PIN io_outs_right[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 11.04 43.2 11.064 ;
    END
  END io_outs_right[19]
  PIN io_outs_right[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 22.248 43.2 22.266 ;
    END
  END io_outs_right[1]
  PIN io_outs_right[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 25.02 43.2 25.038 ;
    END
  END io_outs_right[20]
  PIN io_outs_right[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 12.636 43.2 12.654 ;
    END
  END io_outs_right[21]
  PIN io_outs_right[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 14.076 43.2 14.094 ;
    END
  END io_outs_right[22]
  PIN io_outs_right[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 14.112 43.2 14.13 ;
    END
  END io_outs_right[23]
  PIN io_outs_right[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 21.504 43.2 21.528 ;
    END
  END io_outs_right[24]
  PIN io_outs_right[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 17.664 43.2 17.688 ;
    END
  END io_outs_right[25]
  PIN io_outs_right[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 23.136 43.2 23.16 ;
    END
  END io_outs_right[26]
  PIN io_outs_right[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 24.864 43.2 24.888 ;
    END
  END io_outs_right[27]
  PIN io_outs_right[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 11.061 43.2 11.079 ;
    END
  END io_outs_right[28]
  PIN io_outs_right[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 19.968 43.2 19.992 ;
    END
  END io_outs_right[29]
  PIN io_outs_right[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 24.192 43.2 24.216 ;
    END
  END io_outs_right[2]
  PIN io_outs_right[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 10.872 43.2 10.89 ;
    END
  END io_outs_right[30]
  PIN io_outs_right[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 11.016 43.2 11.034 ;
    END
  END io_outs_right[31]
  PIN io_outs_right[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 29.952 43.2 29.976 ;
    END
  END io_outs_right[32]
  PIN io_outs_right[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 27.612 43.2 27.63 ;
    END
  END io_outs_right[33]
  PIN io_outs_right[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 10.848 43.2 10.872 ;
    END
  END io_outs_right[34]
  PIN io_outs_right[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 28.032 43.2 28.056 ;
    END
  END io_outs_right[35]
  PIN io_outs_right[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 20.016 43.2 20.034 ;
    END
  END io_outs_right[36]
  PIN io_outs_right[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 18.144 43.2 18.168 ;
    END
  END io_outs_right[37]
  PIN io_outs_right[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 13.68 43.2 13.698 ;
    END
  END io_outs_right[38]
  PIN io_outs_right[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 17.76 43.2 17.784 ;
    END
  END io_outs_right[39]
  PIN io_outs_right[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 25.488 43.2 25.506 ;
    END
  END io_outs_right[3]
  PIN io_outs_right[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 21.408 43.2 21.432 ;
    END
  END io_outs_right[40]
  PIN io_outs_right[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 23.436 43.2 23.454 ;
    END
  END io_outs_right[41]
  PIN io_outs_right[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 11.328 43.2 11.352 ;
    END
  END io_outs_right[42]
  PIN io_outs_right[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 29.664 43.2 29.688 ;
    END
  END io_outs_right[43]
  PIN io_outs_right[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 23.52 43.2 23.544 ;
    END
  END io_outs_right[44]
  PIN io_outs_right[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 27.108 43.2 27.126 ;
    END
  END io_outs_right[45]
  PIN io_outs_right[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 23.481 43.2 23.499 ;
    END
  END io_outs_right[46]
  PIN io_outs_right[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 15.936 43.2 15.96 ;
    END
  END io_outs_right[47]
  PIN io_outs_right[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 29.808 43.2 29.826 ;
    END
  END io_outs_right[48]
  PIN io_outs_right[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 15.876 43.2 15.894 ;
    END
  END io_outs_right[49]
  PIN io_outs_right[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 32.352 43.2 32.376 ;
    END
  END io_outs_right[4]
  PIN io_outs_right[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 10.944 43.2 10.968 ;
    END
  END io_outs_right[50]
  PIN io_outs_right[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 14.652 43.2 14.67 ;
    END
  END io_outs_right[51]
  PIN io_outs_right[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 15.552 43.2 15.576 ;
    END
  END io_outs_right[52]
  PIN io_outs_right[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 11.952 43.2 11.97 ;
    END
  END io_outs_right[53]
  PIN io_outs_right[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 11.136 43.2 11.16 ;
    END
  END io_outs_right[54]
  PIN io_outs_right[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 11.808 43.2 11.832 ;
    END
  END io_outs_right[55]
  PIN io_outs_right[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 18.048 43.2 18.072 ;
    END
  END io_outs_right[56]
  PIN io_outs_right[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 20.928 43.2 20.952 ;
    END
  END io_outs_right[57]
  PIN io_outs_right[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 11.232 43.2 11.256 ;
    END
  END io_outs_right[58]
  PIN io_outs_right[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 10.98 43.2 10.998 ;
    END
  END io_outs_right[59]
  PIN io_outs_right[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 25.92 43.2 25.944 ;
    END
  END io_outs_right[5]
  PIN io_outs_right[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 14.976 43.2 15 ;
    END
  END io_outs_right[60]
  PIN io_outs_right[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 30.144 43.2 30.168 ;
    END
  END io_outs_right[61]
  PIN io_outs_right[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 14.112 43.2 14.136 ;
    END
  END io_outs_right[62]
  PIN io_outs_right[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 29.916 43.2 29.934 ;
    END
  END io_outs_right[63]
  PIN io_outs_right[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 30.42 43.2 30.438 ;
    END
  END io_outs_right[6]
  PIN io_outs_right[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 30.348 43.2 30.366 ;
    END
  END io_outs_right[7]
  PIN io_outs_right[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT  43.116 32.448 43.2 32.472 ;
    END
  END io_outs_right[8]
  PIN io_outs_right[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT  43.163 33.084 43.2 33.102 ;
    END
  END io_outs_right[9]
  PIN io_outs_up[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  30.528 43.163 30.546 43.2 ;
    END
  END io_outs_up[0]
  PIN io_outs_up[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.264 43.116 15.288 43.2 ;
    END
  END io_outs_up[10]
  PIN io_outs_up[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  26.4 43.116 26.424 43.2 ;
    END
  END io_outs_up[11]
  PIN io_outs_up[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  15.768 43.163 15.786 43.2 ;
    END
  END io_outs_up[12]
  PIN io_outs_up[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  22.176 43.116 22.2 43.2 ;
    END
  END io_outs_up[13]
  PIN io_outs_up[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  15.36 43.116 15.384 43.2 ;
    END
  END io_outs_up[14]
  PIN io_outs_up[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  26.064 43.163 26.082 43.2 ;
    END
  END io_outs_up[15]
  PIN io_outs_up[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  10.872 43.163 10.89 43.2 ;
    END
  END io_outs_up[16]
  PIN io_outs_up[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.272 43.116 10.296 43.2 ;
    END
  END io_outs_up[17]
  PIN io_outs_up[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.464 43.116 10.488 43.2 ;
    END
  END io_outs_up[18]
  PIN io_outs_up[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  8.712 43.163 8.73 43.2 ;
    END
  END io_outs_up[19]
  PIN io_outs_up[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  20.352 43.116 20.376 43.2 ;
    END
  END io_outs_up[1]
  PIN io_outs_up[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.64 43.116 8.664 43.2 ;
    END
  END io_outs_up[20]
  PIN io_outs_up[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.216 43.116 9.24 43.2 ;
    END
  END io_outs_up[21]
  PIN io_outs_up[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  9.936 43.163 9.954 43.2 ;
    END
  END io_outs_up[22]
  PIN io_outs_up[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.256 43.116 8.28 43.2 ;
    END
  END io_outs_up[23]
  PIN io_outs_up[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.408 43.116 9.432 43.2 ;
    END
  END io_outs_up[24]
  PIN io_outs_up[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  7.848 43.163 7.866 43.2 ;
    END
  END io_outs_up[25]
  PIN io_outs_up[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  7.92 43.163 7.938 43.2 ;
    END
  END io_outs_up[26]
  PIN io_outs_up[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  8.208 43.163 8.226 43.2 ;
    END
  END io_outs_up[27]
  PIN io_outs_up[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  10.44 43.163 10.458 43.2 ;
    END
  END io_outs_up[28]
  PIN io_outs_up[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  7.872 43.116 7.896 43.2 ;
    END
  END io_outs_up[29]
  PIN io_outs_up[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  20.736 43.163 20.754 43.2 ;
    END
  END io_outs_up[2]
  PIN io_outs_up[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.928 43.116 8.952 43.2 ;
    END
  END io_outs_up[30]
  PIN io_outs_up[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.368 43.116 10.392 43.2 ;
    END
  END io_outs_up[31]
  PIN io_outs_up[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  11.04 43.116 11.064 43.2 ;
    END
  END io_outs_up[32]
  PIN io_outs_up[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.504 43.116 9.528 43.2 ;
    END
  END io_outs_up[33]
  PIN io_outs_up[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.312 43.116 9.336 43.2 ;
    END
  END io_outs_up[34]
  PIN io_outs_up[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  8.784 43.163 8.802 43.2 ;
    END
  END io_outs_up[35]
  PIN io_outs_up[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.024 43.116 9.048 43.2 ;
    END
  END io_outs_up[36]
  PIN io_outs_up[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  11.088 43.163 11.106 43.2 ;
    END
  END io_outs_up[37]
  PIN io_outs_up[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  9.432 43.163 9.45 43.2 ;
    END
  END io_outs_up[38]
  PIN io_outs_up[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  7.632 43.163 7.65 43.2 ;
    END
  END io_outs_up[39]
  PIN io_outs_up[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  20.808 43.163 20.826 43.2 ;
    END
  END io_outs_up[3]
  PIN io_outs_up[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  8.136 43.163 8.154 43.2 ;
    END
  END io_outs_up[40]
  PIN io_outs_up[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  7.68 43.116 7.704 43.2 ;
    END
  END io_outs_up[41]
  PIN io_outs_up[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.832 43.116 8.856 43.2 ;
    END
  END io_outs_up[42]
  PIN io_outs_up[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  8.352 43.116 8.376 43.2 ;
    END
  END io_outs_up[43]
  PIN io_outs_up[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  10.728 43.163 10.746 43.2 ;
    END
  END io_outs_up[44]
  PIN io_outs_up[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  9.864 43.163 9.882 43.2 ;
    END
  END io_outs_up[45]
  PIN io_outs_up[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  7.968 43.116 7.992 43.2 ;
    END
  END io_outs_up[46]
  PIN io_outs_up[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  10.512 43.163 10.53 43.2 ;
    END
  END io_outs_up[47]
  PIN io_outs_up[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  10.944 43.163 10.962 43.2 ;
    END
  END io_outs_up[48]
  PIN io_outs_up[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  10.008 43.163 10.026 43.2 ;
    END
  END io_outs_up[49]
  PIN io_outs_up[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  19.392 43.116 19.416 43.2 ;
    END
  END io_outs_up[4]
  PIN io_outs_up[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  8.856 43.163 8.874 43.2 ;
    END
  END io_outs_up[50]
  PIN io_outs_up[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  7.584 43.116 7.608 43.2 ;
    END
  END io_outs_up[51]
  PIN io_outs_up[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  8.28 43.163 8.298 43.2 ;
    END
  END io_outs_up[52]
  PIN io_outs_up[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.984 43.116 10.008 43.2 ;
    END
  END io_outs_up[53]
  PIN io_outs_up[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  7.776 43.116 7.8 43.2 ;
    END
  END io_outs_up[54]
  PIN io_outs_up[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  7.488 43.163 7.506 43.2 ;
    END
  END io_outs_up[55]
  PIN io_outs_up[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  9.792 43.116 9.816 43.2 ;
    END
  END io_outs_up[56]
  PIN io_outs_up[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  11.16 43.163 11.178 43.2 ;
    END
  END io_outs_up[57]
  PIN io_outs_up[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  8.064 43.163 8.082 43.2 ;
    END
  END io_outs_up[58]
  PIN io_outs_up[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  11.136 43.116 11.16 43.2 ;
    END
  END io_outs_up[59]
  PIN io_outs_up[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  24.672 43.116 24.696 43.2 ;
    END
  END io_outs_up[5]
  PIN io_outs_up[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  7.704 43.163 7.722 43.2 ;
    END
  END io_outs_up[60]
  PIN io_outs_up[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  10.656 43.116 10.68 43.2 ;
    END
  END io_outs_up[61]
  PIN io_outs_up[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  7.488 43.116 7.512 43.2 ;
    END
  END io_outs_up[62]
  PIN io_outs_up[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  11.232 43.116 11.256 43.2 ;
    END
  END io_outs_up[63]
  PIN io_outs_up[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  27.504 43.163 27.522 43.2 ;
    END
  END io_outs_up[6]
  PIN io_outs_up[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  19.104 43.116 19.128 43.2 ;
    END
  END io_outs_up[7]
  PIN io_outs_up[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT  18.792 43.163 18.81 43.2 ;
    END
  END io_outs_up[8]
  PIN io_outs_up[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT  19.2 43.116 19.224 43.2 ;
    END
  END io_outs_up[9]
  OBS
    LAYER M1 ;
     RECT  0 0 43.2 43.2 ;
    LAYER M2 ;
     RECT  0 0 43.2 43.2 ;
    LAYER M3 ;
     RECT  0 0 43.2 43.2 ;
    LAYER M4 ;
     RECT  0 0 43.2 43.2 ;
    LAYER M5 ;
     RECT  0 0 43.2 43.2 ;
  END
END Element
END LIBRARY
