VERSION 5.6 ;
  BUSBITCHARS "[]" ;
  DIVIDERCHAR "/" ;

MACRO LDO_COMPARATOR_LATCH
  CLASS CORE ;
  ORIGIN 0.000 0.000 ;
  FOREIGN LDO_COMPARATOR_LATCH 0 0 ;
  SIZE 18.240 BY 8.140 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      #LAYER pwell ;
      #  RECT -0.130 7.925 18.370 8.355 ;
      #  RECT 2.005 6.705 18.130 7.925 ;
      #  RECT 2.005 6.475 15.290 6.705 ;
      LAYER met1 ;
        RECT 0.000 8.025 18.240 8.255 ;
    END
    PORT
      #LAYER pwell ;
      #  RECT 2.040 1.485 15.390 1.665 ;
      #  RECT 0.485 1.435 15.390 1.485 ;
      #  RECT 0.485 0.215 18.130 1.435 ;
      #  RECT -0.130 -0.215 18.370 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 18.240 0.115 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 8.055 18.240 8.225 ;
      LAYER mcon ;
        RECT 0.155 8.055 0.325 8.225 ;
        RECT 0.635 8.055 0.805 8.225 ;
        RECT 1.115 8.055 1.285 8.225 ;
        RECT 1.595 8.055 1.765 8.225 ;
        RECT 2.075 8.055 2.245 8.225 ;
        RECT 2.555 8.055 2.725 8.225 ;
        RECT 3.035 8.055 3.205 8.225 ;
        RECT 3.515 8.055 3.685 8.225 ;
        RECT 3.995 8.055 4.165 8.225 ;
        RECT 4.475 8.055 4.645 8.225 ;
        RECT 4.955 8.055 5.125 8.225 ;
        RECT 5.435 8.055 5.605 8.225 ;
        RECT 5.915 8.055 6.085 8.225 ;
        RECT 6.395 8.055 6.565 8.225 ;
        RECT 6.875 8.055 7.045 8.225 ;
        RECT 7.355 8.055 7.525 8.225 ;
        RECT 7.835 8.055 8.005 8.225 ;
        RECT 8.315 8.055 8.485 8.225 ;
        RECT 8.795 8.055 8.965 8.225 ;
        RECT 9.275 8.055 9.445 8.225 ;
        RECT 15.995 8.055 16.165 8.225 ;
        RECT 16.475 8.055 16.645 8.225 ;
        RECT 16.955 8.055 17.125 8.225 ;
        RECT 17.435 8.055 17.605 8.225 ;
        RECT 17.915 8.055 18.085 8.225 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 18.240 0.085 ;
      LAYER mcon ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 15.995 -0.085 16.165 0.085 ;
        RECT 16.475 -0.085 16.645 0.085 ;
        RECT 16.955 -0.085 17.125 0.085 ;
        RECT 17.435 -0.085 17.605 0.085 ;
        RECT 17.915 -0.085 18.085 0.085 ;
    END
  END vnb
  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT -0.185 7.515 18.240 7.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 18.240 0.625 ;
    END
    PORT
      LAYER li1 ;
        RECT 15.930 0.365 17.240 1.345 ;
      LAYER mcon ;
        RECT 15.960 0.395 16.130 0.565 ;
        RECT 16.320 0.395 16.490 0.565 ;
        RECT 16.680 0.395 16.850 0.565 ;
        RECT 17.040 0.395 17.210 0.565 ;
    END
    PORT
      LAYER li1 ;
        RECT 15.930 6.795 17.240 7.775 ;
      LAYER mcon ;
        RECT 15.960 7.575 16.130 7.745 ;
        RECT 16.320 7.575 16.490 7.745 ;
        RECT 16.680 7.575 16.850 7.745 ;
        RECT 17.040 7.575 17.210 7.745 ;
    END
  END vgnd
  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 4.325 18.240 4.695 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 18.240 3.815 ;
    END
    PORT
      LAYER li1 ;
        RECT 15.930 4.385 16.880 5.965 ;
        RECT 17.500 4.385 18.090 5.965 ;
      LAYER mcon ;
        RECT 15.960 4.465 16.130 4.635 ;
        RECT 16.320 4.465 16.490 4.635 ;
        RECT 16.680 4.465 16.850 4.635 ;
        RECT 17.530 4.465 17.700 4.635 ;
        RECT 17.890 4.465 18.060 4.635 ;
    END
    PORT
      LAYER li1 ;
        RECT 15.930 2.175 16.880 3.755 ;
        RECT 17.500 2.175 18.090 3.755 ;
      LAYER mcon ;
        RECT 15.960 3.505 16.130 3.675 ;
        RECT 16.320 3.505 16.490 3.675 ;
        RECT 16.680 3.505 16.850 3.675 ;
        RECT 17.530 3.505 17.700 3.675 ;
        RECT 17.890 3.505 18.060 3.675 ;
    END
  END vpwr
  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      #LAYER nwell ;
      #  RECT 15.510 6.175 18.570 6.255 ;
      #  RECT -0.440 1.965 18.570 6.175 ;
      #  RECT 15.510 1.885 18.570 1.965 ;
      LAYER met1 ;
        RECT 0.000 3.955 18.240 4.185 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 3.985 18.240 4.155 ;
      LAYER mcon ;
        RECT 2.120 3.985 2.290 4.155 ;
        RECT 2.600 3.985 2.770 4.155 ;
        RECT 3.080 3.985 3.250 4.155 ;
        RECT 3.560 3.985 3.730 4.155 ;
        RECT 4.040 3.985 4.210 4.155 ;
        RECT 4.520 3.985 4.690 4.155 ;
        RECT 5.000 3.985 5.170 4.155 ;
        RECT 5.480 3.985 5.650 4.155 ;
        RECT 5.960 3.985 6.130 4.155 ;
        RECT 6.440 3.985 6.610 4.155 ;
        RECT 6.920 3.985 7.090 4.155 ;
        RECT 10.760 3.985 10.930 4.155 ;
        RECT 15.995 3.985 16.165 4.155 ;
        RECT 16.475 3.985 16.645 4.155 ;
        RECT 16.955 3.985 17.125 4.155 ;
        RECT 17.435 3.985 17.605 4.155 ;
        RECT 17.915 3.985 18.085 4.155 ;
    END
  END vpb
  PIN VREF
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 9.005 6.130 9.335 6.475 ;
    END
  END VREF
  PIN VREG
    DIRECTION INOUT ;
    USE POWER ;
    ANTENNAGATEAREA 5.000000 ;
    PORT
      LAYER li1 ;
        RECT 9.110 1.660 9.490 2.005 ;
    END
  END VREG
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.035 5.650 1.390 5.975 ;
        RECT 1.085 2.385 1.350 5.650 ;
        RECT 1.005 2.035 1.430 2.385 ;
    END
  END CLK
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.000 5.725 17.340 6.060 ;
        RECT 17.085 1.980 17.255 5.725 ;
        RECT 17.030 1.700 17.315 1.980 ;
        RECT 17.085 1.605 17.255 1.700 ;
    END
  END OUT
  OBS
      LAYER li1 ;
        RECT 3.035 7.565 15.170 7.735 ;
        RECT 2.250 6.735 2.580 7.325 ;
        RECT 3.035 7.010 3.365 7.565 ;
        RECT 3.825 6.735 4.155 7.315 ;
        RECT 4.610 6.975 4.940 7.565 ;
        RECT 5.390 6.735 5.720 7.295 ;
        RECT 6.175 6.895 6.505 7.565 ;
        RECT 6.965 6.770 7.295 7.565 ;
        RECT 7.750 6.970 8.080 7.325 ;
        RECT 8.530 7.170 8.860 7.565 ;
        RECT 9.315 6.970 9.645 7.360 ;
        RECT 10.100 7.205 10.430 7.565 ;
        RECT 10.880 6.970 11.210 7.370 ;
        RECT 11.660 7.175 11.990 7.565 ;
        RECT 12.445 6.970 12.775 7.320 ;
        RECT 13.230 7.240 13.560 7.565 ;
        RECT 14.010 6.970 14.340 7.245 ;
        RECT 7.750 6.800 14.340 6.970 ;
        RECT 1.615 6.565 5.720 6.735 ;
        RECT 1.615 6.490 1.950 6.565 ;
        RECT 6.545 6.395 7.310 6.565 ;
        RECT 1.035 5.650 1.390 5.975 ;
        RECT 5.920 5.920 6.090 6.245 ;
        RECT 6.545 6.125 6.845 6.395 ;
        RECT 3.050 5.850 7.295 5.920 ;
        RECT 14.010 5.850 14.340 6.800 ;
        RECT 14.840 6.680 15.170 7.565 ;
        RECT 17.690 6.965 18.020 7.625 ;
        RECT 17.420 6.795 18.020 6.965 ;
        RECT 17.420 6.615 17.635 6.795 ;
        RECT 15.965 6.375 16.855 6.590 ;
        RECT 15.210 6.205 16.855 6.375 ;
        RECT 17.060 6.445 17.635 6.615 ;
        RECT 15.210 5.920 15.380 6.205 ;
        RECT 15.050 5.850 15.380 5.920 ;
        RECT 3.050 5.750 15.380 5.850 ;
        RECT 2.265 4.740 2.595 5.510 ;
        RECT 3.050 4.955 3.380 5.750 ;
        RECT 3.840 4.740 4.170 5.500 ;
        RECT 4.625 4.955 4.955 5.750 ;
        RECT 5.405 4.740 5.735 5.480 ;
        RECT 6.190 4.870 6.520 5.750 ;
        RECT 6.965 5.680 15.380 5.750 ;
        RECT 6.965 4.955 7.295 5.680 ;
        RECT 2.265 4.570 5.735 4.740 ;
        RECT 7.750 4.745 8.080 5.510 ;
        RECT 8.530 5.000 8.860 5.680 ;
        RECT 9.315 4.745 9.645 5.450 ;
        RECT 10.100 4.970 10.430 5.680 ;
        RECT 10.880 4.745 11.210 5.390 ;
        RECT 11.660 4.970 11.990 5.680 ;
        RECT 12.445 4.745 12.775 5.505 ;
        RECT 13.230 4.985 13.560 5.680 ;
        RECT 14.010 4.745 14.340 5.280 ;
        RECT 15.050 4.865 15.380 5.680 ;
        RECT 7.750 4.575 14.340 4.745 ;
        RECT 9.315 4.570 9.645 4.575 ;
        RECT 12.445 4.570 12.775 4.575 ;
        RECT 2.265 4.425 2.595 4.570 ;
        RECT 14.010 4.425 14.340 4.575 ;
        RECT 17.060 4.385 17.310 6.445 ;
        RECT 17.815 6.285 18.115 6.615 ;
        RECT 2.265 3.645 2.595 3.685 ;
        RECT 14.010 3.645 14.340 3.715 ;
        RECT 2.265 3.475 5.735 3.645 ;
        RECT 2.265 2.705 2.595 3.475 ;
        RECT 3.050 2.385 3.380 3.180 ;
        RECT 3.840 2.715 4.170 3.475 ;
        RECT 4.625 2.385 4.955 3.180 ;
        RECT 5.405 2.735 5.735 3.475 ;
        RECT 7.750 3.475 14.340 3.645 ;
        RECT 6.190 2.385 6.520 3.265 ;
        RECT 6.965 2.515 7.295 3.180 ;
        RECT 7.750 2.705 8.080 3.475 ;
        RECT 8.530 2.515 8.860 3.135 ;
        RECT 9.315 2.800 9.645 3.475 ;
        RECT 10.100 2.515 10.430 3.165 ;
        RECT 10.880 2.825 11.210 3.475 ;
        RECT 11.660 2.515 11.990 3.165 ;
        RECT 12.445 2.710 12.775 3.475 ;
        RECT 13.230 2.515 13.560 3.150 ;
        RECT 14.010 2.840 14.340 3.475 ;
        RECT 15.050 2.515 15.380 3.270 ;
        RECT 6.965 2.385 15.380 2.515 ;
        RECT 1.030 2.045 1.360 2.385 ;
        RECT 3.050 2.345 15.380 2.385 ;
        RECT 3.050 2.215 7.490 2.345 ;
        RECT 6.555 1.975 6.880 2.045 ;
        RECT 0.595 1.705 0.925 1.860 ;
        RECT 6.185 1.805 6.880 1.975 ;
        RECT 7.295 1.820 7.490 2.215 ;
        RECT 6.555 1.715 6.880 1.805 ;
        RECT 0.595 1.535 5.755 1.705 ;
        RECT 0.595 0.665 0.925 1.535 ;
        RECT 1.465 0.285 1.795 1.310 ;
        RECT 2.285 0.765 2.615 1.535 ;
        RECT 3.070 0.525 3.400 1.320 ;
        RECT 3.860 0.775 4.190 1.535 ;
        RECT 4.645 0.525 4.975 1.320 ;
        RECT 5.425 0.795 5.755 1.535 ;
        RECT 6.210 0.525 6.540 1.025 ;
        RECT 6.965 0.525 7.295 1.535 ;
        RECT 14.010 1.490 14.340 2.345 ;
        RECT 15.050 2.215 15.380 2.345 ;
        RECT 15.210 1.935 15.380 2.215 ;
        RECT 15.210 1.765 16.855 1.935 ;
        RECT 15.965 1.550 16.855 1.765 ;
        RECT 17.060 1.695 17.310 3.755 ;
        RECT 17.060 1.525 17.635 1.695 ;
        RECT 17.815 1.525 18.115 1.855 ;
        RECT 7.750 1.320 14.340 1.490 ;
        RECT 7.750 0.765 8.080 1.320 ;
        RECT 8.530 0.525 8.860 1.105 ;
        RECT 9.315 0.730 9.645 1.320 ;
        RECT 10.100 0.525 10.430 1.095 ;
        RECT 10.880 0.720 11.210 1.320 ;
        RECT 11.660 0.525 11.990 1.105 ;
        RECT 12.445 0.770 12.775 1.320 ;
        RECT 13.230 0.525 13.560 1.100 ;
        RECT 14.010 0.815 14.340 1.320 ;
        RECT 14.935 0.525 15.265 1.410 ;
        RECT 17.420 1.345 17.635 1.525 ;
        RECT 17.420 1.175 18.020 1.345 ;
        RECT 3.070 0.355 15.265 0.525 ;
        RECT 17.690 0.515 18.020 1.175 ;
      LAYER mcon ;
        RECT 1.695 6.545 1.865 6.715 ;
        RECT 7.010 6.395 7.180 6.565 ;
        RECT 5.920 6.075 6.090 6.245 ;
        RECT 1.130 5.720 1.300 5.890 ;
        RECT 17.100 6.350 17.270 6.520 ;
        RECT 2.350 4.475 2.520 4.645 ;
        RECT 14.065 4.460 14.235 4.630 ;
        RECT 17.895 6.295 18.065 6.465 ;
        RECT 2.350 3.485 2.520 3.655 ;
        RECT 14.065 3.510 14.235 3.680 ;
        RECT 1.105 2.125 1.275 2.295 ;
        RECT 0.660 1.655 0.830 1.825 ;
        RECT 7.320 1.830 7.490 2.000 ;
        RECT 1.545 0.365 1.715 0.535 ;
        RECT 17.085 1.740 17.255 1.910 ;
        RECT 17.865 1.605 18.035 1.775 ;
      LAYER met1 ;
        RECT 1.580 6.300 1.950 6.850 ;
        RECT 6.115 6.300 6.420 6.320 ;
        RECT 6.935 6.300 7.270 6.650 ;
        RECT 5.765 6.025 6.420 6.300 ;
        RECT 17.055 6.175 17.695 6.625 ;
        RECT 6.115 6.020 6.420 6.025 ;
        RECT 17.865 6.005 18.100 6.535 ;
        RECT 1.045 5.650 1.365 5.955 ;
        RECT 16.950 5.715 18.100 6.005 ;
        RECT 1.010 2.030 1.350 2.360 ;
        RECT 1.640 1.860 1.960 1.945 ;
        RECT 0.595 1.580 1.960 1.860 ;
        RECT 6.040 1.740 6.425 2.310 ;
        RECT 17.475 2.270 18.110 2.620 ;
        RECT 6.875 2.080 7.540 2.145 ;
        RECT 6.875 1.745 7.575 2.080 ;
        RECT 6.875 1.685 7.540 1.745 ;
        RECT 16.985 1.635 17.410 1.985 ;
        RECT 17.815 1.535 18.110 2.270 ;
      LAYER via ;
        RECT 1.640 6.350 1.900 6.610 ;
        RECT 6.955 6.340 7.215 6.600 ;
        RECT 17.360 6.315 17.620 6.575 ;
        RECT 6.130 6.020 6.390 6.280 ;
        RECT 1.075 5.665 1.335 5.925 ;
        RECT 17.030 5.740 17.290 6.000 ;
        RECT 1.050 2.065 1.310 2.325 ;
        RECT 17.490 2.310 17.750 2.570 ;
        RECT 1.640 1.620 1.900 1.880 ;
        RECT 6.130 1.920 6.390 2.180 ;
        RECT 6.955 1.775 7.215 2.035 ;
        RECT 17.030 1.700 17.290 1.960 ;
      LAYER met2 ;
        RECT 1.615 6.350 1.950 6.660 ;
        RECT 1.680 1.900 1.880 6.350 ;
        RECT 6.100 6.020 6.435 6.330 ;
        RECT 6.935 6.300 7.270 6.650 ;
        RECT 6.185 2.200 6.355 6.020 ;
        RECT 1.615 1.590 1.950 1.900 ;
        RECT 6.100 1.890 6.435 2.200 ;
        RECT 7.010 2.055 7.180 6.300 ;
        RECT 17.285 6.250 17.715 6.640 ;
        RECT 17.545 2.590 17.715 6.250 ;
        RECT 17.460 2.280 17.805 2.590 ;
        RECT 6.920 1.745 7.265 2.055 ;
  END
END LDO_COMPARATOR_LATCH
END LIBRARY

